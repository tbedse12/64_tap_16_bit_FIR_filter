module DA_table_2(table_in_2 , table_out_2);
input unsigned [15:0]table_in_2;
output [31:0]table_out_2;
wire  [31:0]LUT_2[65535:0]; 
wire [31:0]table_out_2; 
assign table_out_2 = LUT_2[table_in_2];
assign LUT_2[0] = 32'b00000000000000000000000000000000;
assign LUT_2[1] = 32'b11111111111111111100111000011001;
assign LUT_2[2] = 32'b00000000000000000110111000111100;
assign LUT_2[3] = 32'b00000000000000000011110001010101;
assign LUT_2[4] = 32'b11111111111111111100011101101000;
assign LUT_2[5] = 32'b11111111111111111001010110000001;
assign LUT_2[6] = 32'b00000000000000000011010110100100;
assign LUT_2[7] = 32'b00000000000000000000001110111101;
assign LUT_2[8] = 32'b11111111111111111010110001011101;
assign LUT_2[9] = 32'b11111111111111110111101001110110;
assign LUT_2[10] = 32'b00000000000000000001101010011001;
assign LUT_2[11] = 32'b11111111111111111110100010110010;
assign LUT_2[12] = 32'b11111111111111110111001111000101;
assign LUT_2[13] = 32'b11111111111111110100000111011110;
assign LUT_2[14] = 32'b11111111111111111110001000000001;
assign LUT_2[15] = 32'b11111111111111111011000000011010;
assign LUT_2[16] = 32'b11111111111111111010100100001010;
assign LUT_2[17] = 32'b11111111111111110111011100100011;
assign LUT_2[18] = 32'b00000000000000000001011101000110;
assign LUT_2[19] = 32'b11111111111111111110010101011111;
assign LUT_2[20] = 32'b11111111111111110111000001110010;
assign LUT_2[21] = 32'b11111111111111110011111010001011;
assign LUT_2[22] = 32'b11111111111111111101111010101110;
assign LUT_2[23] = 32'b11111111111111111010110011000111;
assign LUT_2[24] = 32'b11111111111111110101010101100111;
assign LUT_2[25] = 32'b11111111111111110010001110000000;
assign LUT_2[26] = 32'b11111111111111111100001110100011;
assign LUT_2[27] = 32'b11111111111111111001000110111100;
assign LUT_2[28] = 32'b11111111111111110001110011001111;
assign LUT_2[29] = 32'b11111111111111101110101011101000;
assign LUT_2[30] = 32'b11111111111111111000101100001011;
assign LUT_2[31] = 32'b11111111111111110101100100100100;
assign LUT_2[32] = 32'b00000000000000000000011011101001;
assign LUT_2[33] = 32'b11111111111111111101010100000010;
assign LUT_2[34] = 32'b00000000000000000111010100100101;
assign LUT_2[35] = 32'b00000000000000000100001100111110;
assign LUT_2[36] = 32'b11111111111111111100111001010001;
assign LUT_2[37] = 32'b11111111111111111001110001101010;
assign LUT_2[38] = 32'b00000000000000000011110010001101;
assign LUT_2[39] = 32'b00000000000000000000101010100110;
assign LUT_2[40] = 32'b11111111111111111011001101000110;
assign LUT_2[41] = 32'b11111111111111111000000101011111;
assign LUT_2[42] = 32'b00000000000000000010000110000010;
assign LUT_2[43] = 32'b11111111111111111110111110011011;
assign LUT_2[44] = 32'b11111111111111110111101010101110;
assign LUT_2[45] = 32'b11111111111111110100100011000111;
assign LUT_2[46] = 32'b11111111111111111110100011101010;
assign LUT_2[47] = 32'b11111111111111111011011100000011;
assign LUT_2[48] = 32'b11111111111111111010111111110011;
assign LUT_2[49] = 32'b11111111111111110111111000001100;
assign LUT_2[50] = 32'b00000000000000000001111000101111;
assign LUT_2[51] = 32'b11111111111111111110110001001000;
assign LUT_2[52] = 32'b11111111111111110111011101011011;
assign LUT_2[53] = 32'b11111111111111110100010101110100;
assign LUT_2[54] = 32'b11111111111111111110010110010111;
assign LUT_2[55] = 32'b11111111111111111011001110110000;
assign LUT_2[56] = 32'b11111111111111110101110001010000;
assign LUT_2[57] = 32'b11111111111111110010101001101001;
assign LUT_2[58] = 32'b11111111111111111100101010001100;
assign LUT_2[59] = 32'b11111111111111111001100010100101;
assign LUT_2[60] = 32'b11111111111111110010001110111000;
assign LUT_2[61] = 32'b11111111111111101111000111010001;
assign LUT_2[62] = 32'b11111111111111111001000111110100;
assign LUT_2[63] = 32'b11111111111111110110000000001101;
assign LUT_2[64] = 32'b11111111111111111000001000100011;
assign LUT_2[65] = 32'b11111111111111110101000000111100;
assign LUT_2[66] = 32'b11111111111111111111000001011111;
assign LUT_2[67] = 32'b11111111111111111011111001111000;
assign LUT_2[68] = 32'b11111111111111110100100110001011;
assign LUT_2[69] = 32'b11111111111111110001011110100100;
assign LUT_2[70] = 32'b11111111111111111011011111000111;
assign LUT_2[71] = 32'b11111111111111111000010111100000;
assign LUT_2[72] = 32'b11111111111111110010111010000000;
assign LUT_2[73] = 32'b11111111111111101111110010011001;
assign LUT_2[74] = 32'b11111111111111111001110010111100;
assign LUT_2[75] = 32'b11111111111111110110101011010101;
assign LUT_2[76] = 32'b11111111111111101111010111101000;
assign LUT_2[77] = 32'b11111111111111101100010000000001;
assign LUT_2[78] = 32'b11111111111111110110010000100100;
assign LUT_2[79] = 32'b11111111111111110011001000111101;
assign LUT_2[80] = 32'b11111111111111110010101100101101;
assign LUT_2[81] = 32'b11111111111111101111100101000110;
assign LUT_2[82] = 32'b11111111111111111001100101101001;
assign LUT_2[83] = 32'b11111111111111110110011110000010;
assign LUT_2[84] = 32'b11111111111111101111001010010101;
assign LUT_2[85] = 32'b11111111111111101100000010101110;
assign LUT_2[86] = 32'b11111111111111110110000011010001;
assign LUT_2[87] = 32'b11111111111111110010111011101010;
assign LUT_2[88] = 32'b11111111111111101101011110001010;
assign LUT_2[89] = 32'b11111111111111101010010110100011;
assign LUT_2[90] = 32'b11111111111111110100010111000110;
assign LUT_2[91] = 32'b11111111111111110001001111011111;
assign LUT_2[92] = 32'b11111111111111101001111011110010;
assign LUT_2[93] = 32'b11111111111111100110110100001011;
assign LUT_2[94] = 32'b11111111111111110000110100101110;
assign LUT_2[95] = 32'b11111111111111101101101101000111;
assign LUT_2[96] = 32'b11111111111111111000100100001100;
assign LUT_2[97] = 32'b11111111111111110101011100100101;
assign LUT_2[98] = 32'b11111111111111111111011101001000;
assign LUT_2[99] = 32'b11111111111111111100010101100001;
assign LUT_2[100] = 32'b11111111111111110101000001110100;
assign LUT_2[101] = 32'b11111111111111110001111010001101;
assign LUT_2[102] = 32'b11111111111111111011111010110000;
assign LUT_2[103] = 32'b11111111111111111000110011001001;
assign LUT_2[104] = 32'b11111111111111110011010101101001;
assign LUT_2[105] = 32'b11111111111111110000001110000010;
assign LUT_2[106] = 32'b11111111111111111010001110100101;
assign LUT_2[107] = 32'b11111111111111110111000110111110;
assign LUT_2[108] = 32'b11111111111111101111110011010001;
assign LUT_2[109] = 32'b11111111111111101100101011101010;
assign LUT_2[110] = 32'b11111111111111110110101100001101;
assign LUT_2[111] = 32'b11111111111111110011100100100110;
assign LUT_2[112] = 32'b11111111111111110011001000010110;
assign LUT_2[113] = 32'b11111111111111110000000000101111;
assign LUT_2[114] = 32'b11111111111111111010000001010010;
assign LUT_2[115] = 32'b11111111111111110110111001101011;
assign LUT_2[116] = 32'b11111111111111101111100101111110;
assign LUT_2[117] = 32'b11111111111111101100011110010111;
assign LUT_2[118] = 32'b11111111111111110110011110111010;
assign LUT_2[119] = 32'b11111111111111110011010111010011;
assign LUT_2[120] = 32'b11111111111111101101111001110011;
assign LUT_2[121] = 32'b11111111111111101010110010001100;
assign LUT_2[122] = 32'b11111111111111110100110010101111;
assign LUT_2[123] = 32'b11111111111111110001101011001000;
assign LUT_2[124] = 32'b11111111111111101010010111011011;
assign LUT_2[125] = 32'b11111111111111100111001111110100;
assign LUT_2[126] = 32'b11111111111111110001010000010111;
assign LUT_2[127] = 32'b11111111111111101110001000110000;
assign LUT_2[128] = 32'b00000000000000000100010100001111;
assign LUT_2[129] = 32'b00000000000000000001001100101000;
assign LUT_2[130] = 32'b00000000000000001011001101001011;
assign LUT_2[131] = 32'b00000000000000001000000101100100;
assign LUT_2[132] = 32'b00000000000000000000110001110111;
assign LUT_2[133] = 32'b11111111111111111101101010010000;
assign LUT_2[134] = 32'b00000000000000000111101010110011;
assign LUT_2[135] = 32'b00000000000000000100100011001100;
assign LUT_2[136] = 32'b11111111111111111111000101101100;
assign LUT_2[137] = 32'b11111111111111111011111110000101;
assign LUT_2[138] = 32'b00000000000000000101111110101000;
assign LUT_2[139] = 32'b00000000000000000010110111000001;
assign LUT_2[140] = 32'b11111111111111111011100011010100;
assign LUT_2[141] = 32'b11111111111111111000011011101101;
assign LUT_2[142] = 32'b00000000000000000010011100010000;
assign LUT_2[143] = 32'b11111111111111111111010100101001;
assign LUT_2[144] = 32'b11111111111111111110111000011001;
assign LUT_2[145] = 32'b11111111111111111011110000110010;
assign LUT_2[146] = 32'b00000000000000000101110001010101;
assign LUT_2[147] = 32'b00000000000000000010101001101110;
assign LUT_2[148] = 32'b11111111111111111011010110000001;
assign LUT_2[149] = 32'b11111111111111111000001110011010;
assign LUT_2[150] = 32'b00000000000000000010001110111101;
assign LUT_2[151] = 32'b11111111111111111111000111010110;
assign LUT_2[152] = 32'b11111111111111111001101001110110;
assign LUT_2[153] = 32'b11111111111111110110100010001111;
assign LUT_2[154] = 32'b00000000000000000000100010110010;
assign LUT_2[155] = 32'b11111111111111111101011011001011;
assign LUT_2[156] = 32'b11111111111111110110000111011110;
assign LUT_2[157] = 32'b11111111111111110010111111110111;
assign LUT_2[158] = 32'b11111111111111111101000000011010;
assign LUT_2[159] = 32'b11111111111111111001111000110011;
assign LUT_2[160] = 32'b00000000000000000100101111111000;
assign LUT_2[161] = 32'b00000000000000000001101000010001;
assign LUT_2[162] = 32'b00000000000000001011101000110100;
assign LUT_2[163] = 32'b00000000000000001000100001001101;
assign LUT_2[164] = 32'b00000000000000000001001101100000;
assign LUT_2[165] = 32'b11111111111111111110000101111001;
assign LUT_2[166] = 32'b00000000000000001000000110011100;
assign LUT_2[167] = 32'b00000000000000000100111110110101;
assign LUT_2[168] = 32'b11111111111111111111100001010101;
assign LUT_2[169] = 32'b11111111111111111100011001101110;
assign LUT_2[170] = 32'b00000000000000000110011010010001;
assign LUT_2[171] = 32'b00000000000000000011010010101010;
assign LUT_2[172] = 32'b11111111111111111011111110111101;
assign LUT_2[173] = 32'b11111111111111111000110111010110;
assign LUT_2[174] = 32'b00000000000000000010110111111001;
assign LUT_2[175] = 32'b11111111111111111111110000010010;
assign LUT_2[176] = 32'b11111111111111111111010100000010;
assign LUT_2[177] = 32'b11111111111111111100001100011011;
assign LUT_2[178] = 32'b00000000000000000110001100111110;
assign LUT_2[179] = 32'b00000000000000000011000101010111;
assign LUT_2[180] = 32'b11111111111111111011110001101010;
assign LUT_2[181] = 32'b11111111111111111000101010000011;
assign LUT_2[182] = 32'b00000000000000000010101010100110;
assign LUT_2[183] = 32'b11111111111111111111100010111111;
assign LUT_2[184] = 32'b11111111111111111010000101011111;
assign LUT_2[185] = 32'b11111111111111110110111101111000;
assign LUT_2[186] = 32'b00000000000000000000111110011011;
assign LUT_2[187] = 32'b11111111111111111101110110110100;
assign LUT_2[188] = 32'b11111111111111110110100011000111;
assign LUT_2[189] = 32'b11111111111111110011011011100000;
assign LUT_2[190] = 32'b11111111111111111101011100000011;
assign LUT_2[191] = 32'b11111111111111111010010100011100;
assign LUT_2[192] = 32'b11111111111111111100011100110010;
assign LUT_2[193] = 32'b11111111111111111001010101001011;
assign LUT_2[194] = 32'b00000000000000000011010101101110;
assign LUT_2[195] = 32'b00000000000000000000001110000111;
assign LUT_2[196] = 32'b11111111111111111000111010011010;
assign LUT_2[197] = 32'b11111111111111110101110010110011;
assign LUT_2[198] = 32'b11111111111111111111110011010110;
assign LUT_2[199] = 32'b11111111111111111100101011101111;
assign LUT_2[200] = 32'b11111111111111110111001110001111;
assign LUT_2[201] = 32'b11111111111111110100000110101000;
assign LUT_2[202] = 32'b11111111111111111110000111001011;
assign LUT_2[203] = 32'b11111111111111111010111111100100;
assign LUT_2[204] = 32'b11111111111111110011101011110111;
assign LUT_2[205] = 32'b11111111111111110000100100010000;
assign LUT_2[206] = 32'b11111111111111111010100100110011;
assign LUT_2[207] = 32'b11111111111111110111011101001100;
assign LUT_2[208] = 32'b11111111111111110111000000111100;
assign LUT_2[209] = 32'b11111111111111110011111001010101;
assign LUT_2[210] = 32'b11111111111111111101111001111000;
assign LUT_2[211] = 32'b11111111111111111010110010010001;
assign LUT_2[212] = 32'b11111111111111110011011110100100;
assign LUT_2[213] = 32'b11111111111111110000010110111101;
assign LUT_2[214] = 32'b11111111111111111010010111100000;
assign LUT_2[215] = 32'b11111111111111110111001111111001;
assign LUT_2[216] = 32'b11111111111111110001110010011001;
assign LUT_2[217] = 32'b11111111111111101110101010110010;
assign LUT_2[218] = 32'b11111111111111111000101011010101;
assign LUT_2[219] = 32'b11111111111111110101100011101110;
assign LUT_2[220] = 32'b11111111111111101110010000000001;
assign LUT_2[221] = 32'b11111111111111101011001000011010;
assign LUT_2[222] = 32'b11111111111111110101001000111101;
assign LUT_2[223] = 32'b11111111111111110010000001010110;
assign LUT_2[224] = 32'b11111111111111111100111000011011;
assign LUT_2[225] = 32'b11111111111111111001110000110100;
assign LUT_2[226] = 32'b00000000000000000011110001010111;
assign LUT_2[227] = 32'b00000000000000000000101001110000;
assign LUT_2[228] = 32'b11111111111111111001010110000011;
assign LUT_2[229] = 32'b11111111111111110110001110011100;
assign LUT_2[230] = 32'b00000000000000000000001110111111;
assign LUT_2[231] = 32'b11111111111111111101000111011000;
assign LUT_2[232] = 32'b11111111111111110111101001111000;
assign LUT_2[233] = 32'b11111111111111110100100010010001;
assign LUT_2[234] = 32'b11111111111111111110100010110100;
assign LUT_2[235] = 32'b11111111111111111011011011001101;
assign LUT_2[236] = 32'b11111111111111110100000111100000;
assign LUT_2[237] = 32'b11111111111111110000111111111001;
assign LUT_2[238] = 32'b11111111111111111011000000011100;
assign LUT_2[239] = 32'b11111111111111110111111000110101;
assign LUT_2[240] = 32'b11111111111111110111011100100101;
assign LUT_2[241] = 32'b11111111111111110100010100111110;
assign LUT_2[242] = 32'b11111111111111111110010101100001;
assign LUT_2[243] = 32'b11111111111111111011001101111010;
assign LUT_2[244] = 32'b11111111111111110011111010001101;
assign LUT_2[245] = 32'b11111111111111110000110010100110;
assign LUT_2[246] = 32'b11111111111111111010110011001001;
assign LUT_2[247] = 32'b11111111111111110111101011100010;
assign LUT_2[248] = 32'b11111111111111110010001110000010;
assign LUT_2[249] = 32'b11111111111111101111000110011011;
assign LUT_2[250] = 32'b11111111111111111001000110111110;
assign LUT_2[251] = 32'b11111111111111110101111111010111;
assign LUT_2[252] = 32'b11111111111111101110101011101010;
assign LUT_2[253] = 32'b11111111111111101011100100000011;
assign LUT_2[254] = 32'b11111111111111110101100100100110;
assign LUT_2[255] = 32'b11111111111111110010011100111111;
assign LUT_2[256] = 32'b00000000000000000011111110100110;
assign LUT_2[257] = 32'b00000000000000000000110110111111;
assign LUT_2[258] = 32'b00000000000000001010110111100010;
assign LUT_2[259] = 32'b00000000000000000111101111111011;
assign LUT_2[260] = 32'b00000000000000000000011100001110;
assign LUT_2[261] = 32'b11111111111111111101010100100111;
assign LUT_2[262] = 32'b00000000000000000111010101001010;
assign LUT_2[263] = 32'b00000000000000000100001101100011;
assign LUT_2[264] = 32'b11111111111111111110110000000011;
assign LUT_2[265] = 32'b11111111111111111011101000011100;
assign LUT_2[266] = 32'b00000000000000000101101000111111;
assign LUT_2[267] = 32'b00000000000000000010100001011000;
assign LUT_2[268] = 32'b11111111111111111011001101101011;
assign LUT_2[269] = 32'b11111111111111111000000110000100;
assign LUT_2[270] = 32'b00000000000000000010000110100111;
assign LUT_2[271] = 32'b11111111111111111110111111000000;
assign LUT_2[272] = 32'b11111111111111111110100010110000;
assign LUT_2[273] = 32'b11111111111111111011011011001001;
assign LUT_2[274] = 32'b00000000000000000101011011101100;
assign LUT_2[275] = 32'b00000000000000000010010100000101;
assign LUT_2[276] = 32'b11111111111111111011000000011000;
assign LUT_2[277] = 32'b11111111111111110111111000110001;
assign LUT_2[278] = 32'b00000000000000000001111001010100;
assign LUT_2[279] = 32'b11111111111111111110110001101101;
assign LUT_2[280] = 32'b11111111111111111001010100001101;
assign LUT_2[281] = 32'b11111111111111110110001100100110;
assign LUT_2[282] = 32'b00000000000000000000001101001001;
assign LUT_2[283] = 32'b11111111111111111101000101100010;
assign LUT_2[284] = 32'b11111111111111110101110001110101;
assign LUT_2[285] = 32'b11111111111111110010101010001110;
assign LUT_2[286] = 32'b11111111111111111100101010110001;
assign LUT_2[287] = 32'b11111111111111111001100011001010;
assign LUT_2[288] = 32'b00000000000000000100011010001111;
assign LUT_2[289] = 32'b00000000000000000001010010101000;
assign LUT_2[290] = 32'b00000000000000001011010011001011;
assign LUT_2[291] = 32'b00000000000000001000001011100100;
assign LUT_2[292] = 32'b00000000000000000000110111110111;
assign LUT_2[293] = 32'b11111111111111111101110000010000;
assign LUT_2[294] = 32'b00000000000000000111110000110011;
assign LUT_2[295] = 32'b00000000000000000100101001001100;
assign LUT_2[296] = 32'b11111111111111111111001011101100;
assign LUT_2[297] = 32'b11111111111111111100000100000101;
assign LUT_2[298] = 32'b00000000000000000110000100101000;
assign LUT_2[299] = 32'b00000000000000000010111101000001;
assign LUT_2[300] = 32'b11111111111111111011101001010100;
assign LUT_2[301] = 32'b11111111111111111000100001101101;
assign LUT_2[302] = 32'b00000000000000000010100010010000;
assign LUT_2[303] = 32'b11111111111111111111011010101001;
assign LUT_2[304] = 32'b11111111111111111110111110011001;
assign LUT_2[305] = 32'b11111111111111111011110110110010;
assign LUT_2[306] = 32'b00000000000000000101110111010101;
assign LUT_2[307] = 32'b00000000000000000010101111101110;
assign LUT_2[308] = 32'b11111111111111111011011100000001;
assign LUT_2[309] = 32'b11111111111111111000010100011010;
assign LUT_2[310] = 32'b00000000000000000010010100111101;
assign LUT_2[311] = 32'b11111111111111111111001101010110;
assign LUT_2[312] = 32'b11111111111111111001101111110110;
assign LUT_2[313] = 32'b11111111111111110110101000001111;
assign LUT_2[314] = 32'b00000000000000000000101000110010;
assign LUT_2[315] = 32'b11111111111111111101100001001011;
assign LUT_2[316] = 32'b11111111111111110110001101011110;
assign LUT_2[317] = 32'b11111111111111110011000101110111;
assign LUT_2[318] = 32'b11111111111111111101000110011010;
assign LUT_2[319] = 32'b11111111111111111001111110110011;
assign LUT_2[320] = 32'b11111111111111111100000111001001;
assign LUT_2[321] = 32'b11111111111111111000111111100010;
assign LUT_2[322] = 32'b00000000000000000011000000000101;
assign LUT_2[323] = 32'b11111111111111111111111000011110;
assign LUT_2[324] = 32'b11111111111111111000100100110001;
assign LUT_2[325] = 32'b11111111111111110101011101001010;
assign LUT_2[326] = 32'b11111111111111111111011101101101;
assign LUT_2[327] = 32'b11111111111111111100010110000110;
assign LUT_2[328] = 32'b11111111111111110110111000100110;
assign LUT_2[329] = 32'b11111111111111110011110000111111;
assign LUT_2[330] = 32'b11111111111111111101110001100010;
assign LUT_2[331] = 32'b11111111111111111010101001111011;
assign LUT_2[332] = 32'b11111111111111110011010110001110;
assign LUT_2[333] = 32'b11111111111111110000001110100111;
assign LUT_2[334] = 32'b11111111111111111010001111001010;
assign LUT_2[335] = 32'b11111111111111110111000111100011;
assign LUT_2[336] = 32'b11111111111111110110101011010011;
assign LUT_2[337] = 32'b11111111111111110011100011101100;
assign LUT_2[338] = 32'b11111111111111111101100100001111;
assign LUT_2[339] = 32'b11111111111111111010011100101000;
assign LUT_2[340] = 32'b11111111111111110011001000111011;
assign LUT_2[341] = 32'b11111111111111110000000001010100;
assign LUT_2[342] = 32'b11111111111111111010000001110111;
assign LUT_2[343] = 32'b11111111111111110110111010010000;
assign LUT_2[344] = 32'b11111111111111110001011100110000;
assign LUT_2[345] = 32'b11111111111111101110010101001001;
assign LUT_2[346] = 32'b11111111111111111000010101101100;
assign LUT_2[347] = 32'b11111111111111110101001110000101;
assign LUT_2[348] = 32'b11111111111111101101111010011000;
assign LUT_2[349] = 32'b11111111111111101010110010110001;
assign LUT_2[350] = 32'b11111111111111110100110011010100;
assign LUT_2[351] = 32'b11111111111111110001101011101101;
assign LUT_2[352] = 32'b11111111111111111100100010110010;
assign LUT_2[353] = 32'b11111111111111111001011011001011;
assign LUT_2[354] = 32'b00000000000000000011011011101110;
assign LUT_2[355] = 32'b00000000000000000000010100000111;
assign LUT_2[356] = 32'b11111111111111111001000000011010;
assign LUT_2[357] = 32'b11111111111111110101111000110011;
assign LUT_2[358] = 32'b11111111111111111111111001010110;
assign LUT_2[359] = 32'b11111111111111111100110001101111;
assign LUT_2[360] = 32'b11111111111111110111010100001111;
assign LUT_2[361] = 32'b11111111111111110100001100101000;
assign LUT_2[362] = 32'b11111111111111111110001101001011;
assign LUT_2[363] = 32'b11111111111111111011000101100100;
assign LUT_2[364] = 32'b11111111111111110011110001110111;
assign LUT_2[365] = 32'b11111111111111110000101010010000;
assign LUT_2[366] = 32'b11111111111111111010101010110011;
assign LUT_2[367] = 32'b11111111111111110111100011001100;
assign LUT_2[368] = 32'b11111111111111110111000110111100;
assign LUT_2[369] = 32'b11111111111111110011111111010101;
assign LUT_2[370] = 32'b11111111111111111101111111111000;
assign LUT_2[371] = 32'b11111111111111111010111000010001;
assign LUT_2[372] = 32'b11111111111111110011100100100100;
assign LUT_2[373] = 32'b11111111111111110000011100111101;
assign LUT_2[374] = 32'b11111111111111111010011101100000;
assign LUT_2[375] = 32'b11111111111111110111010101111001;
assign LUT_2[376] = 32'b11111111111111110001111000011001;
assign LUT_2[377] = 32'b11111111111111101110110000110010;
assign LUT_2[378] = 32'b11111111111111111000110001010101;
assign LUT_2[379] = 32'b11111111111111110101101001101110;
assign LUT_2[380] = 32'b11111111111111101110010110000001;
assign LUT_2[381] = 32'b11111111111111101011001110011010;
assign LUT_2[382] = 32'b11111111111111110101001110111101;
assign LUT_2[383] = 32'b11111111111111110010000111010110;
assign LUT_2[384] = 32'b00000000000000001000010010110101;
assign LUT_2[385] = 32'b00000000000000000101001011001110;
assign LUT_2[386] = 32'b00000000000000001111001011110001;
assign LUT_2[387] = 32'b00000000000000001100000100001010;
assign LUT_2[388] = 32'b00000000000000000100110000011101;
assign LUT_2[389] = 32'b00000000000000000001101000110110;
assign LUT_2[390] = 32'b00000000000000001011101001011001;
assign LUT_2[391] = 32'b00000000000000001000100001110010;
assign LUT_2[392] = 32'b00000000000000000011000100010010;
assign LUT_2[393] = 32'b11111111111111111111111100101011;
assign LUT_2[394] = 32'b00000000000000001001111101001110;
assign LUT_2[395] = 32'b00000000000000000110110101100111;
assign LUT_2[396] = 32'b11111111111111111111100001111010;
assign LUT_2[397] = 32'b11111111111111111100011010010011;
assign LUT_2[398] = 32'b00000000000000000110011010110110;
assign LUT_2[399] = 32'b00000000000000000011010011001111;
assign LUT_2[400] = 32'b00000000000000000010110110111111;
assign LUT_2[401] = 32'b11111111111111111111101111011000;
assign LUT_2[402] = 32'b00000000000000001001101111111011;
assign LUT_2[403] = 32'b00000000000000000110101000010100;
assign LUT_2[404] = 32'b11111111111111111111010100100111;
assign LUT_2[405] = 32'b11111111111111111100001101000000;
assign LUT_2[406] = 32'b00000000000000000110001101100011;
assign LUT_2[407] = 32'b00000000000000000011000101111100;
assign LUT_2[408] = 32'b11111111111111111101101000011100;
assign LUT_2[409] = 32'b11111111111111111010100000110101;
assign LUT_2[410] = 32'b00000000000000000100100001011000;
assign LUT_2[411] = 32'b00000000000000000001011001110001;
assign LUT_2[412] = 32'b11111111111111111010000110000100;
assign LUT_2[413] = 32'b11111111111111110110111110011101;
assign LUT_2[414] = 32'b00000000000000000000111111000000;
assign LUT_2[415] = 32'b11111111111111111101110111011001;
assign LUT_2[416] = 32'b00000000000000001000101110011110;
assign LUT_2[417] = 32'b00000000000000000101100110110111;
assign LUT_2[418] = 32'b00000000000000001111100111011010;
assign LUT_2[419] = 32'b00000000000000001100011111110011;
assign LUT_2[420] = 32'b00000000000000000101001100000110;
assign LUT_2[421] = 32'b00000000000000000010000100011111;
assign LUT_2[422] = 32'b00000000000000001100000101000010;
assign LUT_2[423] = 32'b00000000000000001000111101011011;
assign LUT_2[424] = 32'b00000000000000000011011111111011;
assign LUT_2[425] = 32'b00000000000000000000011000010100;
assign LUT_2[426] = 32'b00000000000000001010011000110111;
assign LUT_2[427] = 32'b00000000000000000111010001010000;
assign LUT_2[428] = 32'b11111111111111111111111101100011;
assign LUT_2[429] = 32'b11111111111111111100110101111100;
assign LUT_2[430] = 32'b00000000000000000110110110011111;
assign LUT_2[431] = 32'b00000000000000000011101110111000;
assign LUT_2[432] = 32'b00000000000000000011010010101000;
assign LUT_2[433] = 32'b00000000000000000000001011000001;
assign LUT_2[434] = 32'b00000000000000001010001011100100;
assign LUT_2[435] = 32'b00000000000000000111000011111101;
assign LUT_2[436] = 32'b11111111111111111111110000010000;
assign LUT_2[437] = 32'b11111111111111111100101000101001;
assign LUT_2[438] = 32'b00000000000000000110101001001100;
assign LUT_2[439] = 32'b00000000000000000011100001100101;
assign LUT_2[440] = 32'b11111111111111111110000100000101;
assign LUT_2[441] = 32'b11111111111111111010111100011110;
assign LUT_2[442] = 32'b00000000000000000100111101000001;
assign LUT_2[443] = 32'b00000000000000000001110101011010;
assign LUT_2[444] = 32'b11111111111111111010100001101101;
assign LUT_2[445] = 32'b11111111111111110111011010000110;
assign LUT_2[446] = 32'b00000000000000000001011010101001;
assign LUT_2[447] = 32'b11111111111111111110010011000010;
assign LUT_2[448] = 32'b00000000000000000000011011011000;
assign LUT_2[449] = 32'b11111111111111111101010011110001;
assign LUT_2[450] = 32'b00000000000000000111010100010100;
assign LUT_2[451] = 32'b00000000000000000100001100101101;
assign LUT_2[452] = 32'b11111111111111111100111001000000;
assign LUT_2[453] = 32'b11111111111111111001110001011001;
assign LUT_2[454] = 32'b00000000000000000011110001111100;
assign LUT_2[455] = 32'b00000000000000000000101010010101;
assign LUT_2[456] = 32'b11111111111111111011001100110101;
assign LUT_2[457] = 32'b11111111111111111000000101001110;
assign LUT_2[458] = 32'b00000000000000000010000101110001;
assign LUT_2[459] = 32'b11111111111111111110111110001010;
assign LUT_2[460] = 32'b11111111111111110111101010011101;
assign LUT_2[461] = 32'b11111111111111110100100010110110;
assign LUT_2[462] = 32'b11111111111111111110100011011001;
assign LUT_2[463] = 32'b11111111111111111011011011110010;
assign LUT_2[464] = 32'b11111111111111111010111111100010;
assign LUT_2[465] = 32'b11111111111111110111110111111011;
assign LUT_2[466] = 32'b00000000000000000001111000011110;
assign LUT_2[467] = 32'b11111111111111111110110000110111;
assign LUT_2[468] = 32'b11111111111111110111011101001010;
assign LUT_2[469] = 32'b11111111111111110100010101100011;
assign LUT_2[470] = 32'b11111111111111111110010110000110;
assign LUT_2[471] = 32'b11111111111111111011001110011111;
assign LUT_2[472] = 32'b11111111111111110101110000111111;
assign LUT_2[473] = 32'b11111111111111110010101001011000;
assign LUT_2[474] = 32'b11111111111111111100101001111011;
assign LUT_2[475] = 32'b11111111111111111001100010010100;
assign LUT_2[476] = 32'b11111111111111110010001110100111;
assign LUT_2[477] = 32'b11111111111111101111000111000000;
assign LUT_2[478] = 32'b11111111111111111001000111100011;
assign LUT_2[479] = 32'b11111111111111110101111111111100;
assign LUT_2[480] = 32'b00000000000000000000110111000001;
assign LUT_2[481] = 32'b11111111111111111101101111011010;
assign LUT_2[482] = 32'b00000000000000000111101111111101;
assign LUT_2[483] = 32'b00000000000000000100101000010110;
assign LUT_2[484] = 32'b11111111111111111101010100101001;
assign LUT_2[485] = 32'b11111111111111111010001101000010;
assign LUT_2[486] = 32'b00000000000000000100001101100101;
assign LUT_2[487] = 32'b00000000000000000001000101111110;
assign LUT_2[488] = 32'b11111111111111111011101000011110;
assign LUT_2[489] = 32'b11111111111111111000100000110111;
assign LUT_2[490] = 32'b00000000000000000010100001011010;
assign LUT_2[491] = 32'b11111111111111111111011001110011;
assign LUT_2[492] = 32'b11111111111111111000000110000110;
assign LUT_2[493] = 32'b11111111111111110100111110011111;
assign LUT_2[494] = 32'b11111111111111111110111111000010;
assign LUT_2[495] = 32'b11111111111111111011110111011011;
assign LUT_2[496] = 32'b11111111111111111011011011001011;
assign LUT_2[497] = 32'b11111111111111111000010011100100;
assign LUT_2[498] = 32'b00000000000000000010010100000111;
assign LUT_2[499] = 32'b11111111111111111111001100100000;
assign LUT_2[500] = 32'b11111111111111110111111000110011;
assign LUT_2[501] = 32'b11111111111111110100110001001100;
assign LUT_2[502] = 32'b11111111111111111110110001101111;
assign LUT_2[503] = 32'b11111111111111111011101010001000;
assign LUT_2[504] = 32'b11111111111111110110001100101000;
assign LUT_2[505] = 32'b11111111111111110011000101000001;
assign LUT_2[506] = 32'b11111111111111111101000101100100;
assign LUT_2[507] = 32'b11111111111111111001111101111101;
assign LUT_2[508] = 32'b11111111111111110010101010010000;
assign LUT_2[509] = 32'b11111111111111101111100010101001;
assign LUT_2[510] = 32'b11111111111111111001100011001100;
assign LUT_2[511] = 32'b11111111111111110110011011100101;
assign LUT_2[512] = 32'b00000000000000000100110001110010;
assign LUT_2[513] = 32'b00000000000000000001101010001011;
assign LUT_2[514] = 32'b00000000000000001011101010101110;
assign LUT_2[515] = 32'b00000000000000001000100011000111;
assign LUT_2[516] = 32'b00000000000000000001001111011010;
assign LUT_2[517] = 32'b11111111111111111110000111110011;
assign LUT_2[518] = 32'b00000000000000001000001000010110;
assign LUT_2[519] = 32'b00000000000000000101000000101111;
assign LUT_2[520] = 32'b11111111111111111111100011001111;
assign LUT_2[521] = 32'b11111111111111111100011011101000;
assign LUT_2[522] = 32'b00000000000000000110011100001011;
assign LUT_2[523] = 32'b00000000000000000011010100100100;
assign LUT_2[524] = 32'b11111111111111111100000000110111;
assign LUT_2[525] = 32'b11111111111111111000111001010000;
assign LUT_2[526] = 32'b00000000000000000010111001110011;
assign LUT_2[527] = 32'b11111111111111111111110010001100;
assign LUT_2[528] = 32'b11111111111111111111010101111100;
assign LUT_2[529] = 32'b11111111111111111100001110010101;
assign LUT_2[530] = 32'b00000000000000000110001110111000;
assign LUT_2[531] = 32'b00000000000000000011000111010001;
assign LUT_2[532] = 32'b11111111111111111011110011100100;
assign LUT_2[533] = 32'b11111111111111111000101011111101;
assign LUT_2[534] = 32'b00000000000000000010101100100000;
assign LUT_2[535] = 32'b11111111111111111111100100111001;
assign LUT_2[536] = 32'b11111111111111111010000111011001;
assign LUT_2[537] = 32'b11111111111111110110111111110010;
assign LUT_2[538] = 32'b00000000000000000001000000010101;
assign LUT_2[539] = 32'b11111111111111111101111000101110;
assign LUT_2[540] = 32'b11111111111111110110100101000001;
assign LUT_2[541] = 32'b11111111111111110011011101011010;
assign LUT_2[542] = 32'b11111111111111111101011101111101;
assign LUT_2[543] = 32'b11111111111111111010010110010110;
assign LUT_2[544] = 32'b00000000000000000101001101011011;
assign LUT_2[545] = 32'b00000000000000000010000101110100;
assign LUT_2[546] = 32'b00000000000000001100000110010111;
assign LUT_2[547] = 32'b00000000000000001000111110110000;
assign LUT_2[548] = 32'b00000000000000000001101011000011;
assign LUT_2[549] = 32'b11111111111111111110100011011100;
assign LUT_2[550] = 32'b00000000000000001000100011111111;
assign LUT_2[551] = 32'b00000000000000000101011100011000;
assign LUT_2[552] = 32'b11111111111111111111111110111000;
assign LUT_2[553] = 32'b11111111111111111100110111010001;
assign LUT_2[554] = 32'b00000000000000000110110111110100;
assign LUT_2[555] = 32'b00000000000000000011110000001101;
assign LUT_2[556] = 32'b11111111111111111100011100100000;
assign LUT_2[557] = 32'b11111111111111111001010100111001;
assign LUT_2[558] = 32'b00000000000000000011010101011100;
assign LUT_2[559] = 32'b00000000000000000000001101110101;
assign LUT_2[560] = 32'b11111111111111111111110001100101;
assign LUT_2[561] = 32'b11111111111111111100101001111110;
assign LUT_2[562] = 32'b00000000000000000110101010100001;
assign LUT_2[563] = 32'b00000000000000000011100010111010;
assign LUT_2[564] = 32'b11111111111111111100001111001101;
assign LUT_2[565] = 32'b11111111111111111001000111100110;
assign LUT_2[566] = 32'b00000000000000000011001000001001;
assign LUT_2[567] = 32'b00000000000000000000000000100010;
assign LUT_2[568] = 32'b11111111111111111010100011000010;
assign LUT_2[569] = 32'b11111111111111110111011011011011;
assign LUT_2[570] = 32'b00000000000000000001011011111110;
assign LUT_2[571] = 32'b11111111111111111110010100010111;
assign LUT_2[572] = 32'b11111111111111110111000000101010;
assign LUT_2[573] = 32'b11111111111111110011111001000011;
assign LUT_2[574] = 32'b11111111111111111101111001100110;
assign LUT_2[575] = 32'b11111111111111111010110001111111;
assign LUT_2[576] = 32'b11111111111111111100111010010101;
assign LUT_2[577] = 32'b11111111111111111001110010101110;
assign LUT_2[578] = 32'b00000000000000000011110011010001;
assign LUT_2[579] = 32'b00000000000000000000101011101010;
assign LUT_2[580] = 32'b11111111111111111001010111111101;
assign LUT_2[581] = 32'b11111111111111110110010000010110;
assign LUT_2[582] = 32'b00000000000000000000010000111001;
assign LUT_2[583] = 32'b11111111111111111101001001010010;
assign LUT_2[584] = 32'b11111111111111110111101011110010;
assign LUT_2[585] = 32'b11111111111111110100100100001011;
assign LUT_2[586] = 32'b11111111111111111110100100101110;
assign LUT_2[587] = 32'b11111111111111111011011101000111;
assign LUT_2[588] = 32'b11111111111111110100001001011010;
assign LUT_2[589] = 32'b11111111111111110001000001110011;
assign LUT_2[590] = 32'b11111111111111111011000010010110;
assign LUT_2[591] = 32'b11111111111111110111111010101111;
assign LUT_2[592] = 32'b11111111111111110111011110011111;
assign LUT_2[593] = 32'b11111111111111110100010110111000;
assign LUT_2[594] = 32'b11111111111111111110010111011011;
assign LUT_2[595] = 32'b11111111111111111011001111110100;
assign LUT_2[596] = 32'b11111111111111110011111100000111;
assign LUT_2[597] = 32'b11111111111111110000110100100000;
assign LUT_2[598] = 32'b11111111111111111010110101000011;
assign LUT_2[599] = 32'b11111111111111110111101101011100;
assign LUT_2[600] = 32'b11111111111111110010001111111100;
assign LUT_2[601] = 32'b11111111111111101111001000010101;
assign LUT_2[602] = 32'b11111111111111111001001000111000;
assign LUT_2[603] = 32'b11111111111111110110000001010001;
assign LUT_2[604] = 32'b11111111111111101110101101100100;
assign LUT_2[605] = 32'b11111111111111101011100101111101;
assign LUT_2[606] = 32'b11111111111111110101100110100000;
assign LUT_2[607] = 32'b11111111111111110010011110111001;
assign LUT_2[608] = 32'b11111111111111111101010101111110;
assign LUT_2[609] = 32'b11111111111111111010001110010111;
assign LUT_2[610] = 32'b00000000000000000100001110111010;
assign LUT_2[611] = 32'b00000000000000000001000111010011;
assign LUT_2[612] = 32'b11111111111111111001110011100110;
assign LUT_2[613] = 32'b11111111111111110110101011111111;
assign LUT_2[614] = 32'b00000000000000000000101100100010;
assign LUT_2[615] = 32'b11111111111111111101100100111011;
assign LUT_2[616] = 32'b11111111111111111000000111011011;
assign LUT_2[617] = 32'b11111111111111110100111111110100;
assign LUT_2[618] = 32'b11111111111111111111000000010111;
assign LUT_2[619] = 32'b11111111111111111011111000110000;
assign LUT_2[620] = 32'b11111111111111110100100101000011;
assign LUT_2[621] = 32'b11111111111111110001011101011100;
assign LUT_2[622] = 32'b11111111111111111011011101111111;
assign LUT_2[623] = 32'b11111111111111111000010110011000;
assign LUT_2[624] = 32'b11111111111111110111111010001000;
assign LUT_2[625] = 32'b11111111111111110100110010100001;
assign LUT_2[626] = 32'b11111111111111111110110011000100;
assign LUT_2[627] = 32'b11111111111111111011101011011101;
assign LUT_2[628] = 32'b11111111111111110100010111110000;
assign LUT_2[629] = 32'b11111111111111110001010000001001;
assign LUT_2[630] = 32'b11111111111111111011010000101100;
assign LUT_2[631] = 32'b11111111111111111000001001000101;
assign LUT_2[632] = 32'b11111111111111110010101011100101;
assign LUT_2[633] = 32'b11111111111111101111100011111110;
assign LUT_2[634] = 32'b11111111111111111001100100100001;
assign LUT_2[635] = 32'b11111111111111110110011100111010;
assign LUT_2[636] = 32'b11111111111111101111001001001101;
assign LUT_2[637] = 32'b11111111111111101100000001100110;
assign LUT_2[638] = 32'b11111111111111110110000010001001;
assign LUT_2[639] = 32'b11111111111111110010111010100010;
assign LUT_2[640] = 32'b00000000000000001001000110000001;
assign LUT_2[641] = 32'b00000000000000000101111110011010;
assign LUT_2[642] = 32'b00000000000000001111111110111101;
assign LUT_2[643] = 32'b00000000000000001100110111010110;
assign LUT_2[644] = 32'b00000000000000000101100011101001;
assign LUT_2[645] = 32'b00000000000000000010011100000010;
assign LUT_2[646] = 32'b00000000000000001100011100100101;
assign LUT_2[647] = 32'b00000000000000001001010100111110;
assign LUT_2[648] = 32'b00000000000000000011110111011110;
assign LUT_2[649] = 32'b00000000000000000000101111110111;
assign LUT_2[650] = 32'b00000000000000001010110000011010;
assign LUT_2[651] = 32'b00000000000000000111101000110011;
assign LUT_2[652] = 32'b00000000000000000000010101000110;
assign LUT_2[653] = 32'b11111111111111111101001101011111;
assign LUT_2[654] = 32'b00000000000000000111001110000010;
assign LUT_2[655] = 32'b00000000000000000100000110011011;
assign LUT_2[656] = 32'b00000000000000000011101010001011;
assign LUT_2[657] = 32'b00000000000000000000100010100100;
assign LUT_2[658] = 32'b00000000000000001010100011000111;
assign LUT_2[659] = 32'b00000000000000000111011011100000;
assign LUT_2[660] = 32'b00000000000000000000000111110011;
assign LUT_2[661] = 32'b11111111111111111101000000001100;
assign LUT_2[662] = 32'b00000000000000000111000000101111;
assign LUT_2[663] = 32'b00000000000000000011111001001000;
assign LUT_2[664] = 32'b11111111111111111110011011101000;
assign LUT_2[665] = 32'b11111111111111111011010100000001;
assign LUT_2[666] = 32'b00000000000000000101010100100100;
assign LUT_2[667] = 32'b00000000000000000010001100111101;
assign LUT_2[668] = 32'b11111111111111111010111001010000;
assign LUT_2[669] = 32'b11111111111111110111110001101001;
assign LUT_2[670] = 32'b00000000000000000001110010001100;
assign LUT_2[671] = 32'b11111111111111111110101010100101;
assign LUT_2[672] = 32'b00000000000000001001100001101010;
assign LUT_2[673] = 32'b00000000000000000110011010000011;
assign LUT_2[674] = 32'b00000000000000010000011010100110;
assign LUT_2[675] = 32'b00000000000000001101010010111111;
assign LUT_2[676] = 32'b00000000000000000101111111010010;
assign LUT_2[677] = 32'b00000000000000000010110111101011;
assign LUT_2[678] = 32'b00000000000000001100111000001110;
assign LUT_2[679] = 32'b00000000000000001001110000100111;
assign LUT_2[680] = 32'b00000000000000000100010011000111;
assign LUT_2[681] = 32'b00000000000000000001001011100000;
assign LUT_2[682] = 32'b00000000000000001011001100000011;
assign LUT_2[683] = 32'b00000000000000001000000100011100;
assign LUT_2[684] = 32'b00000000000000000000110000101111;
assign LUT_2[685] = 32'b11111111111111111101101001001000;
assign LUT_2[686] = 32'b00000000000000000111101001101011;
assign LUT_2[687] = 32'b00000000000000000100100010000100;
assign LUT_2[688] = 32'b00000000000000000100000101110100;
assign LUT_2[689] = 32'b00000000000000000000111110001101;
assign LUT_2[690] = 32'b00000000000000001010111110110000;
assign LUT_2[691] = 32'b00000000000000000111110111001001;
assign LUT_2[692] = 32'b00000000000000000000100011011100;
assign LUT_2[693] = 32'b11111111111111111101011011110101;
assign LUT_2[694] = 32'b00000000000000000111011100011000;
assign LUT_2[695] = 32'b00000000000000000100010100110001;
assign LUT_2[696] = 32'b11111111111111111110110111010001;
assign LUT_2[697] = 32'b11111111111111111011101111101010;
assign LUT_2[698] = 32'b00000000000000000101110000001101;
assign LUT_2[699] = 32'b00000000000000000010101000100110;
assign LUT_2[700] = 32'b11111111111111111011010100111001;
assign LUT_2[701] = 32'b11111111111111111000001101010010;
assign LUT_2[702] = 32'b00000000000000000010001101110101;
assign LUT_2[703] = 32'b11111111111111111111000110001110;
assign LUT_2[704] = 32'b00000000000000000001001110100100;
assign LUT_2[705] = 32'b11111111111111111110000110111101;
assign LUT_2[706] = 32'b00000000000000001000000111100000;
assign LUT_2[707] = 32'b00000000000000000100111111111001;
assign LUT_2[708] = 32'b11111111111111111101101100001100;
assign LUT_2[709] = 32'b11111111111111111010100100100101;
assign LUT_2[710] = 32'b00000000000000000100100101001000;
assign LUT_2[711] = 32'b00000000000000000001011101100001;
assign LUT_2[712] = 32'b11111111111111111100000000000001;
assign LUT_2[713] = 32'b11111111111111111000111000011010;
assign LUT_2[714] = 32'b00000000000000000010111000111101;
assign LUT_2[715] = 32'b11111111111111111111110001010110;
assign LUT_2[716] = 32'b11111111111111111000011101101001;
assign LUT_2[717] = 32'b11111111111111110101010110000010;
assign LUT_2[718] = 32'b11111111111111111111010110100101;
assign LUT_2[719] = 32'b11111111111111111100001110111110;
assign LUT_2[720] = 32'b11111111111111111011110010101110;
assign LUT_2[721] = 32'b11111111111111111000101011000111;
assign LUT_2[722] = 32'b00000000000000000010101011101010;
assign LUT_2[723] = 32'b11111111111111111111100100000011;
assign LUT_2[724] = 32'b11111111111111111000010000010110;
assign LUT_2[725] = 32'b11111111111111110101001000101111;
assign LUT_2[726] = 32'b11111111111111111111001001010010;
assign LUT_2[727] = 32'b11111111111111111100000001101011;
assign LUT_2[728] = 32'b11111111111111110110100100001011;
assign LUT_2[729] = 32'b11111111111111110011011100100100;
assign LUT_2[730] = 32'b11111111111111111101011101000111;
assign LUT_2[731] = 32'b11111111111111111010010101100000;
assign LUT_2[732] = 32'b11111111111111110011000001110011;
assign LUT_2[733] = 32'b11111111111111101111111010001100;
assign LUT_2[734] = 32'b11111111111111111001111010101111;
assign LUT_2[735] = 32'b11111111111111110110110011001000;
assign LUT_2[736] = 32'b00000000000000000001101010001101;
assign LUT_2[737] = 32'b11111111111111111110100010100110;
assign LUT_2[738] = 32'b00000000000000001000100011001001;
assign LUT_2[739] = 32'b00000000000000000101011011100010;
assign LUT_2[740] = 32'b11111111111111111110000111110101;
assign LUT_2[741] = 32'b11111111111111111011000000001110;
assign LUT_2[742] = 32'b00000000000000000101000000110001;
assign LUT_2[743] = 32'b00000000000000000001111001001010;
assign LUT_2[744] = 32'b11111111111111111100011011101010;
assign LUT_2[745] = 32'b11111111111111111001010100000011;
assign LUT_2[746] = 32'b00000000000000000011010100100110;
assign LUT_2[747] = 32'b00000000000000000000001100111111;
assign LUT_2[748] = 32'b11111111111111111000111001010010;
assign LUT_2[749] = 32'b11111111111111110101110001101011;
assign LUT_2[750] = 32'b11111111111111111111110010001110;
assign LUT_2[751] = 32'b11111111111111111100101010100111;
assign LUT_2[752] = 32'b11111111111111111100001110010111;
assign LUT_2[753] = 32'b11111111111111111001000110110000;
assign LUT_2[754] = 32'b00000000000000000011000111010011;
assign LUT_2[755] = 32'b11111111111111111111111111101100;
assign LUT_2[756] = 32'b11111111111111111000101011111111;
assign LUT_2[757] = 32'b11111111111111110101100100011000;
assign LUT_2[758] = 32'b11111111111111111111100100111011;
assign LUT_2[759] = 32'b11111111111111111100011101010100;
assign LUT_2[760] = 32'b11111111111111110110111111110100;
assign LUT_2[761] = 32'b11111111111111110011111000001101;
assign LUT_2[762] = 32'b11111111111111111101111000110000;
assign LUT_2[763] = 32'b11111111111111111010110001001001;
assign LUT_2[764] = 32'b11111111111111110011011101011100;
assign LUT_2[765] = 32'b11111111111111110000010101110101;
assign LUT_2[766] = 32'b11111111111111111010010110011000;
assign LUT_2[767] = 32'b11111111111111110111001110110001;
assign LUT_2[768] = 32'b00000000000000001000110000011000;
assign LUT_2[769] = 32'b00000000000000000101101000110001;
assign LUT_2[770] = 32'b00000000000000001111101001010100;
assign LUT_2[771] = 32'b00000000000000001100100001101101;
assign LUT_2[772] = 32'b00000000000000000101001110000000;
assign LUT_2[773] = 32'b00000000000000000010000110011001;
assign LUT_2[774] = 32'b00000000000000001100000110111100;
assign LUT_2[775] = 32'b00000000000000001000111111010101;
assign LUT_2[776] = 32'b00000000000000000011100001110101;
assign LUT_2[777] = 32'b00000000000000000000011010001110;
assign LUT_2[778] = 32'b00000000000000001010011010110001;
assign LUT_2[779] = 32'b00000000000000000111010011001010;
assign LUT_2[780] = 32'b11111111111111111111111111011101;
assign LUT_2[781] = 32'b11111111111111111100110111110110;
assign LUT_2[782] = 32'b00000000000000000110111000011001;
assign LUT_2[783] = 32'b00000000000000000011110000110010;
assign LUT_2[784] = 32'b00000000000000000011010100100010;
assign LUT_2[785] = 32'b00000000000000000000001100111011;
assign LUT_2[786] = 32'b00000000000000001010001101011110;
assign LUT_2[787] = 32'b00000000000000000111000101110111;
assign LUT_2[788] = 32'b11111111111111111111110010001010;
assign LUT_2[789] = 32'b11111111111111111100101010100011;
assign LUT_2[790] = 32'b00000000000000000110101011000110;
assign LUT_2[791] = 32'b00000000000000000011100011011111;
assign LUT_2[792] = 32'b11111111111111111110000101111111;
assign LUT_2[793] = 32'b11111111111111111010111110011000;
assign LUT_2[794] = 32'b00000000000000000100111110111011;
assign LUT_2[795] = 32'b00000000000000000001110111010100;
assign LUT_2[796] = 32'b11111111111111111010100011100111;
assign LUT_2[797] = 32'b11111111111111110111011100000000;
assign LUT_2[798] = 32'b00000000000000000001011100100011;
assign LUT_2[799] = 32'b11111111111111111110010100111100;
assign LUT_2[800] = 32'b00000000000000001001001100000001;
assign LUT_2[801] = 32'b00000000000000000110000100011010;
assign LUT_2[802] = 32'b00000000000000010000000100111101;
assign LUT_2[803] = 32'b00000000000000001100111101010110;
assign LUT_2[804] = 32'b00000000000000000101101001101001;
assign LUT_2[805] = 32'b00000000000000000010100010000010;
assign LUT_2[806] = 32'b00000000000000001100100010100101;
assign LUT_2[807] = 32'b00000000000000001001011010111110;
assign LUT_2[808] = 32'b00000000000000000011111101011110;
assign LUT_2[809] = 32'b00000000000000000000110101110111;
assign LUT_2[810] = 32'b00000000000000001010110110011010;
assign LUT_2[811] = 32'b00000000000000000111101110110011;
assign LUT_2[812] = 32'b00000000000000000000011011000110;
assign LUT_2[813] = 32'b11111111111111111101010011011111;
assign LUT_2[814] = 32'b00000000000000000111010100000010;
assign LUT_2[815] = 32'b00000000000000000100001100011011;
assign LUT_2[816] = 32'b00000000000000000011110000001011;
assign LUT_2[817] = 32'b00000000000000000000101000100100;
assign LUT_2[818] = 32'b00000000000000001010101001000111;
assign LUT_2[819] = 32'b00000000000000000111100001100000;
assign LUT_2[820] = 32'b00000000000000000000001101110011;
assign LUT_2[821] = 32'b11111111111111111101000110001100;
assign LUT_2[822] = 32'b00000000000000000111000110101111;
assign LUT_2[823] = 32'b00000000000000000011111111001000;
assign LUT_2[824] = 32'b11111111111111111110100001101000;
assign LUT_2[825] = 32'b11111111111111111011011010000001;
assign LUT_2[826] = 32'b00000000000000000101011010100100;
assign LUT_2[827] = 32'b00000000000000000010010010111101;
assign LUT_2[828] = 32'b11111111111111111010111111010000;
assign LUT_2[829] = 32'b11111111111111110111110111101001;
assign LUT_2[830] = 32'b00000000000000000001111000001100;
assign LUT_2[831] = 32'b11111111111111111110110000100101;
assign LUT_2[832] = 32'b00000000000000000000111000111011;
assign LUT_2[833] = 32'b11111111111111111101110001010100;
assign LUT_2[834] = 32'b00000000000000000111110001110111;
assign LUT_2[835] = 32'b00000000000000000100101010010000;
assign LUT_2[836] = 32'b11111111111111111101010110100011;
assign LUT_2[837] = 32'b11111111111111111010001110111100;
assign LUT_2[838] = 32'b00000000000000000100001111011111;
assign LUT_2[839] = 32'b00000000000000000001000111111000;
assign LUT_2[840] = 32'b11111111111111111011101010011000;
assign LUT_2[841] = 32'b11111111111111111000100010110001;
assign LUT_2[842] = 32'b00000000000000000010100011010100;
assign LUT_2[843] = 32'b11111111111111111111011011101101;
assign LUT_2[844] = 32'b11111111111111111000001000000000;
assign LUT_2[845] = 32'b11111111111111110101000000011001;
assign LUT_2[846] = 32'b11111111111111111111000000111100;
assign LUT_2[847] = 32'b11111111111111111011111001010101;
assign LUT_2[848] = 32'b11111111111111111011011101000101;
assign LUT_2[849] = 32'b11111111111111111000010101011110;
assign LUT_2[850] = 32'b00000000000000000010010110000001;
assign LUT_2[851] = 32'b11111111111111111111001110011010;
assign LUT_2[852] = 32'b11111111111111110111111010101101;
assign LUT_2[853] = 32'b11111111111111110100110011000110;
assign LUT_2[854] = 32'b11111111111111111110110011101001;
assign LUT_2[855] = 32'b11111111111111111011101100000010;
assign LUT_2[856] = 32'b11111111111111110110001110100010;
assign LUT_2[857] = 32'b11111111111111110011000110111011;
assign LUT_2[858] = 32'b11111111111111111101000111011110;
assign LUT_2[859] = 32'b11111111111111111001111111110111;
assign LUT_2[860] = 32'b11111111111111110010101100001010;
assign LUT_2[861] = 32'b11111111111111101111100100100011;
assign LUT_2[862] = 32'b11111111111111111001100101000110;
assign LUT_2[863] = 32'b11111111111111110110011101011111;
assign LUT_2[864] = 32'b00000000000000000001010100100100;
assign LUT_2[865] = 32'b11111111111111111110001100111101;
assign LUT_2[866] = 32'b00000000000000001000001101100000;
assign LUT_2[867] = 32'b00000000000000000101000101111001;
assign LUT_2[868] = 32'b11111111111111111101110010001100;
assign LUT_2[869] = 32'b11111111111111111010101010100101;
assign LUT_2[870] = 32'b00000000000000000100101011001000;
assign LUT_2[871] = 32'b00000000000000000001100011100001;
assign LUT_2[872] = 32'b11111111111111111100000110000001;
assign LUT_2[873] = 32'b11111111111111111000111110011010;
assign LUT_2[874] = 32'b00000000000000000010111110111101;
assign LUT_2[875] = 32'b11111111111111111111110111010110;
assign LUT_2[876] = 32'b11111111111111111000100011101001;
assign LUT_2[877] = 32'b11111111111111110101011100000010;
assign LUT_2[878] = 32'b11111111111111111111011100100101;
assign LUT_2[879] = 32'b11111111111111111100010100111110;
assign LUT_2[880] = 32'b11111111111111111011111000101110;
assign LUT_2[881] = 32'b11111111111111111000110001000111;
assign LUT_2[882] = 32'b00000000000000000010110001101010;
assign LUT_2[883] = 32'b11111111111111111111101010000011;
assign LUT_2[884] = 32'b11111111111111111000010110010110;
assign LUT_2[885] = 32'b11111111111111110101001110101111;
assign LUT_2[886] = 32'b11111111111111111111001111010010;
assign LUT_2[887] = 32'b11111111111111111100000111101011;
assign LUT_2[888] = 32'b11111111111111110110101010001011;
assign LUT_2[889] = 32'b11111111111111110011100010100100;
assign LUT_2[890] = 32'b11111111111111111101100011000111;
assign LUT_2[891] = 32'b11111111111111111010011011100000;
assign LUT_2[892] = 32'b11111111111111110011000111110011;
assign LUT_2[893] = 32'b11111111111111110000000000001100;
assign LUT_2[894] = 32'b11111111111111111010000000101111;
assign LUT_2[895] = 32'b11111111111111110110111001001000;
assign LUT_2[896] = 32'b00000000000000001101000100100111;
assign LUT_2[897] = 32'b00000000000000001001111101000000;
assign LUT_2[898] = 32'b00000000000000010011111101100011;
assign LUT_2[899] = 32'b00000000000000010000110101111100;
assign LUT_2[900] = 32'b00000000000000001001100010001111;
assign LUT_2[901] = 32'b00000000000000000110011010101000;
assign LUT_2[902] = 32'b00000000000000010000011011001011;
assign LUT_2[903] = 32'b00000000000000001101010011100100;
assign LUT_2[904] = 32'b00000000000000000111110110000100;
assign LUT_2[905] = 32'b00000000000000000100101110011101;
assign LUT_2[906] = 32'b00000000000000001110101111000000;
assign LUT_2[907] = 32'b00000000000000001011100111011001;
assign LUT_2[908] = 32'b00000000000000000100010011101100;
assign LUT_2[909] = 32'b00000000000000000001001100000101;
assign LUT_2[910] = 32'b00000000000000001011001100101000;
assign LUT_2[911] = 32'b00000000000000001000000101000001;
assign LUT_2[912] = 32'b00000000000000000111101000110001;
assign LUT_2[913] = 32'b00000000000000000100100001001010;
assign LUT_2[914] = 32'b00000000000000001110100001101101;
assign LUT_2[915] = 32'b00000000000000001011011010000110;
assign LUT_2[916] = 32'b00000000000000000100000110011001;
assign LUT_2[917] = 32'b00000000000000000000111110110010;
assign LUT_2[918] = 32'b00000000000000001010111111010101;
assign LUT_2[919] = 32'b00000000000000000111110111101110;
assign LUT_2[920] = 32'b00000000000000000010011010001110;
assign LUT_2[921] = 32'b11111111111111111111010010100111;
assign LUT_2[922] = 32'b00000000000000001001010011001010;
assign LUT_2[923] = 32'b00000000000000000110001011100011;
assign LUT_2[924] = 32'b11111111111111111110110111110110;
assign LUT_2[925] = 32'b11111111111111111011110000001111;
assign LUT_2[926] = 32'b00000000000000000101110000110010;
assign LUT_2[927] = 32'b00000000000000000010101001001011;
assign LUT_2[928] = 32'b00000000000000001101100000010000;
assign LUT_2[929] = 32'b00000000000000001010011000101001;
assign LUT_2[930] = 32'b00000000000000010100011001001100;
assign LUT_2[931] = 32'b00000000000000010001010001100101;
assign LUT_2[932] = 32'b00000000000000001001111101111000;
assign LUT_2[933] = 32'b00000000000000000110110110010001;
assign LUT_2[934] = 32'b00000000000000010000110110110100;
assign LUT_2[935] = 32'b00000000000000001101101111001101;
assign LUT_2[936] = 32'b00000000000000001000010001101101;
assign LUT_2[937] = 32'b00000000000000000101001010000110;
assign LUT_2[938] = 32'b00000000000000001111001010101001;
assign LUT_2[939] = 32'b00000000000000001100000011000010;
assign LUT_2[940] = 32'b00000000000000000100101111010101;
assign LUT_2[941] = 32'b00000000000000000001100111101110;
assign LUT_2[942] = 32'b00000000000000001011101000010001;
assign LUT_2[943] = 32'b00000000000000001000100000101010;
assign LUT_2[944] = 32'b00000000000000001000000100011010;
assign LUT_2[945] = 32'b00000000000000000100111100110011;
assign LUT_2[946] = 32'b00000000000000001110111101010110;
assign LUT_2[947] = 32'b00000000000000001011110101101111;
assign LUT_2[948] = 32'b00000000000000000100100010000010;
assign LUT_2[949] = 32'b00000000000000000001011010011011;
assign LUT_2[950] = 32'b00000000000000001011011010111110;
assign LUT_2[951] = 32'b00000000000000001000010011010111;
assign LUT_2[952] = 32'b00000000000000000010110101110111;
assign LUT_2[953] = 32'b11111111111111111111101110010000;
assign LUT_2[954] = 32'b00000000000000001001101110110011;
assign LUT_2[955] = 32'b00000000000000000110100111001100;
assign LUT_2[956] = 32'b11111111111111111111010011011111;
assign LUT_2[957] = 32'b11111111111111111100001011111000;
assign LUT_2[958] = 32'b00000000000000000110001100011011;
assign LUT_2[959] = 32'b00000000000000000011000100110100;
assign LUT_2[960] = 32'b00000000000000000101001101001010;
assign LUT_2[961] = 32'b00000000000000000010000101100011;
assign LUT_2[962] = 32'b00000000000000001100000110000110;
assign LUT_2[963] = 32'b00000000000000001000111110011111;
assign LUT_2[964] = 32'b00000000000000000001101010110010;
assign LUT_2[965] = 32'b11111111111111111110100011001011;
assign LUT_2[966] = 32'b00000000000000001000100011101110;
assign LUT_2[967] = 32'b00000000000000000101011100000111;
assign LUT_2[968] = 32'b11111111111111111111111110100111;
assign LUT_2[969] = 32'b11111111111111111100110111000000;
assign LUT_2[970] = 32'b00000000000000000110110111100011;
assign LUT_2[971] = 32'b00000000000000000011101111111100;
assign LUT_2[972] = 32'b11111111111111111100011100001111;
assign LUT_2[973] = 32'b11111111111111111001010100101000;
assign LUT_2[974] = 32'b00000000000000000011010101001011;
assign LUT_2[975] = 32'b00000000000000000000001101100100;
assign LUT_2[976] = 32'b11111111111111111111110001010100;
assign LUT_2[977] = 32'b11111111111111111100101001101101;
assign LUT_2[978] = 32'b00000000000000000110101010010000;
assign LUT_2[979] = 32'b00000000000000000011100010101001;
assign LUT_2[980] = 32'b11111111111111111100001110111100;
assign LUT_2[981] = 32'b11111111111111111001000111010101;
assign LUT_2[982] = 32'b00000000000000000011000111111000;
assign LUT_2[983] = 32'b00000000000000000000000000010001;
assign LUT_2[984] = 32'b11111111111111111010100010110001;
assign LUT_2[985] = 32'b11111111111111110111011011001010;
assign LUT_2[986] = 32'b00000000000000000001011011101101;
assign LUT_2[987] = 32'b11111111111111111110010100000110;
assign LUT_2[988] = 32'b11111111111111110111000000011001;
assign LUT_2[989] = 32'b11111111111111110011111000110010;
assign LUT_2[990] = 32'b11111111111111111101111001010101;
assign LUT_2[991] = 32'b11111111111111111010110001101110;
assign LUT_2[992] = 32'b00000000000000000101101000110011;
assign LUT_2[993] = 32'b00000000000000000010100001001100;
assign LUT_2[994] = 32'b00000000000000001100100001101111;
assign LUT_2[995] = 32'b00000000000000001001011010001000;
assign LUT_2[996] = 32'b00000000000000000010000110011011;
assign LUT_2[997] = 32'b11111111111111111110111110110100;
assign LUT_2[998] = 32'b00000000000000001000111111010111;
assign LUT_2[999] = 32'b00000000000000000101110111110000;
assign LUT_2[1000] = 32'b00000000000000000000011010010000;
assign LUT_2[1001] = 32'b11111111111111111101010010101001;
assign LUT_2[1002] = 32'b00000000000000000111010011001100;
assign LUT_2[1003] = 32'b00000000000000000100001011100101;
assign LUT_2[1004] = 32'b11111111111111111100110111111000;
assign LUT_2[1005] = 32'b11111111111111111001110000010001;
assign LUT_2[1006] = 32'b00000000000000000011110000110100;
assign LUT_2[1007] = 32'b00000000000000000000101001001101;
assign LUT_2[1008] = 32'b00000000000000000000001100111101;
assign LUT_2[1009] = 32'b11111111111111111101000101010110;
assign LUT_2[1010] = 32'b00000000000000000111000101111001;
assign LUT_2[1011] = 32'b00000000000000000011111110010010;
assign LUT_2[1012] = 32'b11111111111111111100101010100101;
assign LUT_2[1013] = 32'b11111111111111111001100010111110;
assign LUT_2[1014] = 32'b00000000000000000011100011100001;
assign LUT_2[1015] = 32'b00000000000000000000011011111010;
assign LUT_2[1016] = 32'b11111111111111111010111110011010;
assign LUT_2[1017] = 32'b11111111111111110111110110110011;
assign LUT_2[1018] = 32'b00000000000000000001110111010110;
assign LUT_2[1019] = 32'b11111111111111111110101111101111;
assign LUT_2[1020] = 32'b11111111111111110111011100000010;
assign LUT_2[1021] = 32'b11111111111111110100010100011011;
assign LUT_2[1022] = 32'b11111111111111111110010100111110;
assign LUT_2[1023] = 32'b11111111111111111011001101010111;
assign LUT_2[1024] = 32'b00000000000000000110101100000101;
assign LUT_2[1025] = 32'b00000000000000000011100100011110;
assign LUT_2[1026] = 32'b00000000000000001101100101000001;
assign LUT_2[1027] = 32'b00000000000000001010011101011010;
assign LUT_2[1028] = 32'b00000000000000000011001001101101;
assign LUT_2[1029] = 32'b00000000000000000000000010000110;
assign LUT_2[1030] = 32'b00000000000000001010000010101001;
assign LUT_2[1031] = 32'b00000000000000000110111011000010;
assign LUT_2[1032] = 32'b00000000000000000001011101100010;
assign LUT_2[1033] = 32'b11111111111111111110010101111011;
assign LUT_2[1034] = 32'b00000000000000001000010110011110;
assign LUT_2[1035] = 32'b00000000000000000101001110110111;
assign LUT_2[1036] = 32'b11111111111111111101111011001010;
assign LUT_2[1037] = 32'b11111111111111111010110011100011;
assign LUT_2[1038] = 32'b00000000000000000100110100000110;
assign LUT_2[1039] = 32'b00000000000000000001101100011111;
assign LUT_2[1040] = 32'b00000000000000000001010000001111;
assign LUT_2[1041] = 32'b11111111111111111110001000101000;
assign LUT_2[1042] = 32'b00000000000000001000001001001011;
assign LUT_2[1043] = 32'b00000000000000000101000001100100;
assign LUT_2[1044] = 32'b11111111111111111101101101110111;
assign LUT_2[1045] = 32'b11111111111111111010100110010000;
assign LUT_2[1046] = 32'b00000000000000000100100110110011;
assign LUT_2[1047] = 32'b00000000000000000001011111001100;
assign LUT_2[1048] = 32'b11111111111111111100000001101100;
assign LUT_2[1049] = 32'b11111111111111111000111010000101;
assign LUT_2[1050] = 32'b00000000000000000010111010101000;
assign LUT_2[1051] = 32'b11111111111111111111110011000001;
assign LUT_2[1052] = 32'b11111111111111111000011111010100;
assign LUT_2[1053] = 32'b11111111111111110101010111101101;
assign LUT_2[1054] = 32'b11111111111111111111011000010000;
assign LUT_2[1055] = 32'b11111111111111111100010000101001;
assign LUT_2[1056] = 32'b00000000000000000111000111101110;
assign LUT_2[1057] = 32'b00000000000000000100000000000111;
assign LUT_2[1058] = 32'b00000000000000001110000000101010;
assign LUT_2[1059] = 32'b00000000000000001010111001000011;
assign LUT_2[1060] = 32'b00000000000000000011100101010110;
assign LUT_2[1061] = 32'b00000000000000000000011101101111;
assign LUT_2[1062] = 32'b00000000000000001010011110010010;
assign LUT_2[1063] = 32'b00000000000000000111010110101011;
assign LUT_2[1064] = 32'b00000000000000000001111001001011;
assign LUT_2[1065] = 32'b11111111111111111110110001100100;
assign LUT_2[1066] = 32'b00000000000000001000110010000111;
assign LUT_2[1067] = 32'b00000000000000000101101010100000;
assign LUT_2[1068] = 32'b11111111111111111110010110110011;
assign LUT_2[1069] = 32'b11111111111111111011001111001100;
assign LUT_2[1070] = 32'b00000000000000000101001111101111;
assign LUT_2[1071] = 32'b00000000000000000010001000001000;
assign LUT_2[1072] = 32'b00000000000000000001101011111000;
assign LUT_2[1073] = 32'b11111111111111111110100100010001;
assign LUT_2[1074] = 32'b00000000000000001000100100110100;
assign LUT_2[1075] = 32'b00000000000000000101011101001101;
assign LUT_2[1076] = 32'b11111111111111111110001001100000;
assign LUT_2[1077] = 32'b11111111111111111011000001111001;
assign LUT_2[1078] = 32'b00000000000000000101000010011100;
assign LUT_2[1079] = 32'b00000000000000000001111010110101;
assign LUT_2[1080] = 32'b11111111111111111100011101010101;
assign LUT_2[1081] = 32'b11111111111111111001010101101110;
assign LUT_2[1082] = 32'b00000000000000000011010110010001;
assign LUT_2[1083] = 32'b00000000000000000000001110101010;
assign LUT_2[1084] = 32'b11111111111111111000111010111101;
assign LUT_2[1085] = 32'b11111111111111110101110011010110;
assign LUT_2[1086] = 32'b11111111111111111111110011111001;
assign LUT_2[1087] = 32'b11111111111111111100101100010010;
assign LUT_2[1088] = 32'b11111111111111111110110100101000;
assign LUT_2[1089] = 32'b11111111111111111011101101000001;
assign LUT_2[1090] = 32'b00000000000000000101101101100100;
assign LUT_2[1091] = 32'b00000000000000000010100101111101;
assign LUT_2[1092] = 32'b11111111111111111011010010010000;
assign LUT_2[1093] = 32'b11111111111111111000001010101001;
assign LUT_2[1094] = 32'b00000000000000000010001011001100;
assign LUT_2[1095] = 32'b11111111111111111111000011100101;
assign LUT_2[1096] = 32'b11111111111111111001100110000101;
assign LUT_2[1097] = 32'b11111111111111110110011110011110;
assign LUT_2[1098] = 32'b00000000000000000000011111000001;
assign LUT_2[1099] = 32'b11111111111111111101010111011010;
assign LUT_2[1100] = 32'b11111111111111110110000011101101;
assign LUT_2[1101] = 32'b11111111111111110010111100000110;
assign LUT_2[1102] = 32'b11111111111111111100111100101001;
assign LUT_2[1103] = 32'b11111111111111111001110101000010;
assign LUT_2[1104] = 32'b11111111111111111001011000110010;
assign LUT_2[1105] = 32'b11111111111111110110010001001011;
assign LUT_2[1106] = 32'b00000000000000000000010001101110;
assign LUT_2[1107] = 32'b11111111111111111101001010000111;
assign LUT_2[1108] = 32'b11111111111111110101110110011010;
assign LUT_2[1109] = 32'b11111111111111110010101110110011;
assign LUT_2[1110] = 32'b11111111111111111100101111010110;
assign LUT_2[1111] = 32'b11111111111111111001100111101111;
assign LUT_2[1112] = 32'b11111111111111110100001010001111;
assign LUT_2[1113] = 32'b11111111111111110001000010101000;
assign LUT_2[1114] = 32'b11111111111111111011000011001011;
assign LUT_2[1115] = 32'b11111111111111110111111011100100;
assign LUT_2[1116] = 32'b11111111111111110000100111110111;
assign LUT_2[1117] = 32'b11111111111111101101100000010000;
assign LUT_2[1118] = 32'b11111111111111110111100000110011;
assign LUT_2[1119] = 32'b11111111111111110100011001001100;
assign LUT_2[1120] = 32'b11111111111111111111010000010001;
assign LUT_2[1121] = 32'b11111111111111111100001000101010;
assign LUT_2[1122] = 32'b00000000000000000110001001001101;
assign LUT_2[1123] = 32'b00000000000000000011000001100110;
assign LUT_2[1124] = 32'b11111111111111111011101101111001;
assign LUT_2[1125] = 32'b11111111111111111000100110010010;
assign LUT_2[1126] = 32'b00000000000000000010100110110101;
assign LUT_2[1127] = 32'b11111111111111111111011111001110;
assign LUT_2[1128] = 32'b11111111111111111010000001101110;
assign LUT_2[1129] = 32'b11111111111111110110111010000111;
assign LUT_2[1130] = 32'b00000000000000000000111010101010;
assign LUT_2[1131] = 32'b11111111111111111101110011000011;
assign LUT_2[1132] = 32'b11111111111111110110011111010110;
assign LUT_2[1133] = 32'b11111111111111110011010111101111;
assign LUT_2[1134] = 32'b11111111111111111101011000010010;
assign LUT_2[1135] = 32'b11111111111111111010010000101011;
assign LUT_2[1136] = 32'b11111111111111111001110100011011;
assign LUT_2[1137] = 32'b11111111111111110110101100110100;
assign LUT_2[1138] = 32'b00000000000000000000101101010111;
assign LUT_2[1139] = 32'b11111111111111111101100101110000;
assign LUT_2[1140] = 32'b11111111111111110110010010000011;
assign LUT_2[1141] = 32'b11111111111111110011001010011100;
assign LUT_2[1142] = 32'b11111111111111111101001010111111;
assign LUT_2[1143] = 32'b11111111111111111010000011011000;
assign LUT_2[1144] = 32'b11111111111111110100100101111000;
assign LUT_2[1145] = 32'b11111111111111110001011110010001;
assign LUT_2[1146] = 32'b11111111111111111011011110110100;
assign LUT_2[1147] = 32'b11111111111111111000010111001101;
assign LUT_2[1148] = 32'b11111111111111110001000011100000;
assign LUT_2[1149] = 32'b11111111111111101101111011111001;
assign LUT_2[1150] = 32'b11111111111111110111111100011100;
assign LUT_2[1151] = 32'b11111111111111110100110100110101;
assign LUT_2[1152] = 32'b00000000000000001011000000010100;
assign LUT_2[1153] = 32'b00000000000000000111111000101101;
assign LUT_2[1154] = 32'b00000000000000010001111001010000;
assign LUT_2[1155] = 32'b00000000000000001110110001101001;
assign LUT_2[1156] = 32'b00000000000000000111011101111100;
assign LUT_2[1157] = 32'b00000000000000000100010110010101;
assign LUT_2[1158] = 32'b00000000000000001110010110111000;
assign LUT_2[1159] = 32'b00000000000000001011001111010001;
assign LUT_2[1160] = 32'b00000000000000000101110001110001;
assign LUT_2[1161] = 32'b00000000000000000010101010001010;
assign LUT_2[1162] = 32'b00000000000000001100101010101101;
assign LUT_2[1163] = 32'b00000000000000001001100011000110;
assign LUT_2[1164] = 32'b00000000000000000010001111011001;
assign LUT_2[1165] = 32'b11111111111111111111000111110010;
assign LUT_2[1166] = 32'b00000000000000001001001000010101;
assign LUT_2[1167] = 32'b00000000000000000110000000101110;
assign LUT_2[1168] = 32'b00000000000000000101100100011110;
assign LUT_2[1169] = 32'b00000000000000000010011100110111;
assign LUT_2[1170] = 32'b00000000000000001100011101011010;
assign LUT_2[1171] = 32'b00000000000000001001010101110011;
assign LUT_2[1172] = 32'b00000000000000000010000010000110;
assign LUT_2[1173] = 32'b11111111111111111110111010011111;
assign LUT_2[1174] = 32'b00000000000000001000111011000010;
assign LUT_2[1175] = 32'b00000000000000000101110011011011;
assign LUT_2[1176] = 32'b00000000000000000000010101111011;
assign LUT_2[1177] = 32'b11111111111111111101001110010100;
assign LUT_2[1178] = 32'b00000000000000000111001110110111;
assign LUT_2[1179] = 32'b00000000000000000100000111010000;
assign LUT_2[1180] = 32'b11111111111111111100110011100011;
assign LUT_2[1181] = 32'b11111111111111111001101011111100;
assign LUT_2[1182] = 32'b00000000000000000011101100011111;
assign LUT_2[1183] = 32'b00000000000000000000100100111000;
assign LUT_2[1184] = 32'b00000000000000001011011011111101;
assign LUT_2[1185] = 32'b00000000000000001000010100010110;
assign LUT_2[1186] = 32'b00000000000000010010010100111001;
assign LUT_2[1187] = 32'b00000000000000001111001101010010;
assign LUT_2[1188] = 32'b00000000000000000111111001100101;
assign LUT_2[1189] = 32'b00000000000000000100110001111110;
assign LUT_2[1190] = 32'b00000000000000001110110010100001;
assign LUT_2[1191] = 32'b00000000000000001011101010111010;
assign LUT_2[1192] = 32'b00000000000000000110001101011010;
assign LUT_2[1193] = 32'b00000000000000000011000101110011;
assign LUT_2[1194] = 32'b00000000000000001101000110010110;
assign LUT_2[1195] = 32'b00000000000000001001111110101111;
assign LUT_2[1196] = 32'b00000000000000000010101011000010;
assign LUT_2[1197] = 32'b11111111111111111111100011011011;
assign LUT_2[1198] = 32'b00000000000000001001100011111110;
assign LUT_2[1199] = 32'b00000000000000000110011100010111;
assign LUT_2[1200] = 32'b00000000000000000110000000000111;
assign LUT_2[1201] = 32'b00000000000000000010111000100000;
assign LUT_2[1202] = 32'b00000000000000001100111001000011;
assign LUT_2[1203] = 32'b00000000000000001001110001011100;
assign LUT_2[1204] = 32'b00000000000000000010011101101111;
assign LUT_2[1205] = 32'b11111111111111111111010110001000;
assign LUT_2[1206] = 32'b00000000000000001001010110101011;
assign LUT_2[1207] = 32'b00000000000000000110001111000100;
assign LUT_2[1208] = 32'b00000000000000000000110001100100;
assign LUT_2[1209] = 32'b11111111111111111101101001111101;
assign LUT_2[1210] = 32'b00000000000000000111101010100000;
assign LUT_2[1211] = 32'b00000000000000000100100010111001;
assign LUT_2[1212] = 32'b11111111111111111101001111001100;
assign LUT_2[1213] = 32'b11111111111111111010000111100101;
assign LUT_2[1214] = 32'b00000000000000000100001000001000;
assign LUT_2[1215] = 32'b00000000000000000001000000100001;
assign LUT_2[1216] = 32'b00000000000000000011001000110111;
assign LUT_2[1217] = 32'b00000000000000000000000001010000;
assign LUT_2[1218] = 32'b00000000000000001010000001110011;
assign LUT_2[1219] = 32'b00000000000000000110111010001100;
assign LUT_2[1220] = 32'b11111111111111111111100110011111;
assign LUT_2[1221] = 32'b11111111111111111100011110111000;
assign LUT_2[1222] = 32'b00000000000000000110011111011011;
assign LUT_2[1223] = 32'b00000000000000000011010111110100;
assign LUT_2[1224] = 32'b11111111111111111101111010010100;
assign LUT_2[1225] = 32'b11111111111111111010110010101101;
assign LUT_2[1226] = 32'b00000000000000000100110011010000;
assign LUT_2[1227] = 32'b00000000000000000001101011101001;
assign LUT_2[1228] = 32'b11111111111111111010010111111100;
assign LUT_2[1229] = 32'b11111111111111110111010000010101;
assign LUT_2[1230] = 32'b00000000000000000001010000111000;
assign LUT_2[1231] = 32'b11111111111111111110001001010001;
assign LUT_2[1232] = 32'b11111111111111111101101101000001;
assign LUT_2[1233] = 32'b11111111111111111010100101011010;
assign LUT_2[1234] = 32'b00000000000000000100100101111101;
assign LUT_2[1235] = 32'b00000000000000000001011110010110;
assign LUT_2[1236] = 32'b11111111111111111010001010101001;
assign LUT_2[1237] = 32'b11111111111111110111000011000010;
assign LUT_2[1238] = 32'b00000000000000000001000011100101;
assign LUT_2[1239] = 32'b11111111111111111101111011111110;
assign LUT_2[1240] = 32'b11111111111111111000011110011110;
assign LUT_2[1241] = 32'b11111111111111110101010110110111;
assign LUT_2[1242] = 32'b11111111111111111111010111011010;
assign LUT_2[1243] = 32'b11111111111111111100001111110011;
assign LUT_2[1244] = 32'b11111111111111110100111100000110;
assign LUT_2[1245] = 32'b11111111111111110001110100011111;
assign LUT_2[1246] = 32'b11111111111111111011110101000010;
assign LUT_2[1247] = 32'b11111111111111111000101101011011;
assign LUT_2[1248] = 32'b00000000000000000011100100100000;
assign LUT_2[1249] = 32'b00000000000000000000011100111001;
assign LUT_2[1250] = 32'b00000000000000001010011101011100;
assign LUT_2[1251] = 32'b00000000000000000111010101110101;
assign LUT_2[1252] = 32'b00000000000000000000000010001000;
assign LUT_2[1253] = 32'b11111111111111111100111010100001;
assign LUT_2[1254] = 32'b00000000000000000110111011000100;
assign LUT_2[1255] = 32'b00000000000000000011110011011101;
assign LUT_2[1256] = 32'b11111111111111111110010101111101;
assign LUT_2[1257] = 32'b11111111111111111011001110010110;
assign LUT_2[1258] = 32'b00000000000000000101001110111001;
assign LUT_2[1259] = 32'b00000000000000000010000111010010;
assign LUT_2[1260] = 32'b11111111111111111010110011100101;
assign LUT_2[1261] = 32'b11111111111111110111101011111110;
assign LUT_2[1262] = 32'b00000000000000000001101100100001;
assign LUT_2[1263] = 32'b11111111111111111110100100111010;
assign LUT_2[1264] = 32'b11111111111111111110001000101010;
assign LUT_2[1265] = 32'b11111111111111111011000001000011;
assign LUT_2[1266] = 32'b00000000000000000101000001100110;
assign LUT_2[1267] = 32'b00000000000000000001111001111111;
assign LUT_2[1268] = 32'b11111111111111111010100110010010;
assign LUT_2[1269] = 32'b11111111111111110111011110101011;
assign LUT_2[1270] = 32'b00000000000000000001011111001110;
assign LUT_2[1271] = 32'b11111111111111111110010111100111;
assign LUT_2[1272] = 32'b11111111111111111000111010000111;
assign LUT_2[1273] = 32'b11111111111111110101110010100000;
assign LUT_2[1274] = 32'b11111111111111111111110011000011;
assign LUT_2[1275] = 32'b11111111111111111100101011011100;
assign LUT_2[1276] = 32'b11111111111111110101010111101111;
assign LUT_2[1277] = 32'b11111111111111110010010000001000;
assign LUT_2[1278] = 32'b11111111111111111100010000101011;
assign LUT_2[1279] = 32'b11111111111111111001001001000100;
assign LUT_2[1280] = 32'b00000000000000001010101010101011;
assign LUT_2[1281] = 32'b00000000000000000111100011000100;
assign LUT_2[1282] = 32'b00000000000000010001100011100111;
assign LUT_2[1283] = 32'b00000000000000001110011100000000;
assign LUT_2[1284] = 32'b00000000000000000111001000010011;
assign LUT_2[1285] = 32'b00000000000000000100000000101100;
assign LUT_2[1286] = 32'b00000000000000001110000001001111;
assign LUT_2[1287] = 32'b00000000000000001010111001101000;
assign LUT_2[1288] = 32'b00000000000000000101011100001000;
assign LUT_2[1289] = 32'b00000000000000000010010100100001;
assign LUT_2[1290] = 32'b00000000000000001100010101000100;
assign LUT_2[1291] = 32'b00000000000000001001001101011101;
assign LUT_2[1292] = 32'b00000000000000000001111001110000;
assign LUT_2[1293] = 32'b11111111111111111110110010001001;
assign LUT_2[1294] = 32'b00000000000000001000110010101100;
assign LUT_2[1295] = 32'b00000000000000000101101011000101;
assign LUT_2[1296] = 32'b00000000000000000101001110110101;
assign LUT_2[1297] = 32'b00000000000000000010000111001110;
assign LUT_2[1298] = 32'b00000000000000001100000111110001;
assign LUT_2[1299] = 32'b00000000000000001001000000001010;
assign LUT_2[1300] = 32'b00000000000000000001101100011101;
assign LUT_2[1301] = 32'b11111111111111111110100100110110;
assign LUT_2[1302] = 32'b00000000000000001000100101011001;
assign LUT_2[1303] = 32'b00000000000000000101011101110010;
assign LUT_2[1304] = 32'b00000000000000000000000000010010;
assign LUT_2[1305] = 32'b11111111111111111100111000101011;
assign LUT_2[1306] = 32'b00000000000000000110111001001110;
assign LUT_2[1307] = 32'b00000000000000000011110001100111;
assign LUT_2[1308] = 32'b11111111111111111100011101111010;
assign LUT_2[1309] = 32'b11111111111111111001010110010011;
assign LUT_2[1310] = 32'b00000000000000000011010110110110;
assign LUT_2[1311] = 32'b00000000000000000000001111001111;
assign LUT_2[1312] = 32'b00000000000000001011000110010100;
assign LUT_2[1313] = 32'b00000000000000000111111110101101;
assign LUT_2[1314] = 32'b00000000000000010001111111010000;
assign LUT_2[1315] = 32'b00000000000000001110110111101001;
assign LUT_2[1316] = 32'b00000000000000000111100011111100;
assign LUT_2[1317] = 32'b00000000000000000100011100010101;
assign LUT_2[1318] = 32'b00000000000000001110011100111000;
assign LUT_2[1319] = 32'b00000000000000001011010101010001;
assign LUT_2[1320] = 32'b00000000000000000101110111110001;
assign LUT_2[1321] = 32'b00000000000000000010110000001010;
assign LUT_2[1322] = 32'b00000000000000001100110000101101;
assign LUT_2[1323] = 32'b00000000000000001001101001000110;
assign LUT_2[1324] = 32'b00000000000000000010010101011001;
assign LUT_2[1325] = 32'b11111111111111111111001101110010;
assign LUT_2[1326] = 32'b00000000000000001001001110010101;
assign LUT_2[1327] = 32'b00000000000000000110000110101110;
assign LUT_2[1328] = 32'b00000000000000000101101010011110;
assign LUT_2[1329] = 32'b00000000000000000010100010110111;
assign LUT_2[1330] = 32'b00000000000000001100100011011010;
assign LUT_2[1331] = 32'b00000000000000001001011011110011;
assign LUT_2[1332] = 32'b00000000000000000010001000000110;
assign LUT_2[1333] = 32'b11111111111111111111000000011111;
assign LUT_2[1334] = 32'b00000000000000001001000001000010;
assign LUT_2[1335] = 32'b00000000000000000101111001011011;
assign LUT_2[1336] = 32'b00000000000000000000011011111011;
assign LUT_2[1337] = 32'b11111111111111111101010100010100;
assign LUT_2[1338] = 32'b00000000000000000111010100110111;
assign LUT_2[1339] = 32'b00000000000000000100001101010000;
assign LUT_2[1340] = 32'b11111111111111111100111001100011;
assign LUT_2[1341] = 32'b11111111111111111001110001111100;
assign LUT_2[1342] = 32'b00000000000000000011110010011111;
assign LUT_2[1343] = 32'b00000000000000000000101010111000;
assign LUT_2[1344] = 32'b00000000000000000010110011001110;
assign LUT_2[1345] = 32'b11111111111111111111101011100111;
assign LUT_2[1346] = 32'b00000000000000001001101100001010;
assign LUT_2[1347] = 32'b00000000000000000110100100100011;
assign LUT_2[1348] = 32'b11111111111111111111010000110110;
assign LUT_2[1349] = 32'b11111111111111111100001001001111;
assign LUT_2[1350] = 32'b00000000000000000110001001110010;
assign LUT_2[1351] = 32'b00000000000000000011000010001011;
assign LUT_2[1352] = 32'b11111111111111111101100100101011;
assign LUT_2[1353] = 32'b11111111111111111010011101000100;
assign LUT_2[1354] = 32'b00000000000000000100011101100111;
assign LUT_2[1355] = 32'b00000000000000000001010110000000;
assign LUT_2[1356] = 32'b11111111111111111010000010010011;
assign LUT_2[1357] = 32'b11111111111111110110111010101100;
assign LUT_2[1358] = 32'b00000000000000000000111011001111;
assign LUT_2[1359] = 32'b11111111111111111101110011101000;
assign LUT_2[1360] = 32'b11111111111111111101010111011000;
assign LUT_2[1361] = 32'b11111111111111111010001111110001;
assign LUT_2[1362] = 32'b00000000000000000100010000010100;
assign LUT_2[1363] = 32'b00000000000000000001001000101101;
assign LUT_2[1364] = 32'b11111111111111111001110101000000;
assign LUT_2[1365] = 32'b11111111111111110110101101011001;
assign LUT_2[1366] = 32'b00000000000000000000101101111100;
assign LUT_2[1367] = 32'b11111111111111111101100110010101;
assign LUT_2[1368] = 32'b11111111111111111000001000110101;
assign LUT_2[1369] = 32'b11111111111111110101000001001110;
assign LUT_2[1370] = 32'b11111111111111111111000001110001;
assign LUT_2[1371] = 32'b11111111111111111011111010001010;
assign LUT_2[1372] = 32'b11111111111111110100100110011101;
assign LUT_2[1373] = 32'b11111111111111110001011110110110;
assign LUT_2[1374] = 32'b11111111111111111011011111011001;
assign LUT_2[1375] = 32'b11111111111111111000010111110010;
assign LUT_2[1376] = 32'b00000000000000000011001110110111;
assign LUT_2[1377] = 32'b00000000000000000000000111010000;
assign LUT_2[1378] = 32'b00000000000000001010000111110011;
assign LUT_2[1379] = 32'b00000000000000000111000000001100;
assign LUT_2[1380] = 32'b11111111111111111111101100011111;
assign LUT_2[1381] = 32'b11111111111111111100100100111000;
assign LUT_2[1382] = 32'b00000000000000000110100101011011;
assign LUT_2[1383] = 32'b00000000000000000011011101110100;
assign LUT_2[1384] = 32'b11111111111111111110000000010100;
assign LUT_2[1385] = 32'b11111111111111111010111000101101;
assign LUT_2[1386] = 32'b00000000000000000100111001010000;
assign LUT_2[1387] = 32'b00000000000000000001110001101001;
assign LUT_2[1388] = 32'b11111111111111111010011101111100;
assign LUT_2[1389] = 32'b11111111111111110111010110010101;
assign LUT_2[1390] = 32'b00000000000000000001010110111000;
assign LUT_2[1391] = 32'b11111111111111111110001111010001;
assign LUT_2[1392] = 32'b11111111111111111101110011000001;
assign LUT_2[1393] = 32'b11111111111111111010101011011010;
assign LUT_2[1394] = 32'b00000000000000000100101011111101;
assign LUT_2[1395] = 32'b00000000000000000001100100010110;
assign LUT_2[1396] = 32'b11111111111111111010010000101001;
assign LUT_2[1397] = 32'b11111111111111110111001001000010;
assign LUT_2[1398] = 32'b00000000000000000001001001100101;
assign LUT_2[1399] = 32'b11111111111111111110000001111110;
assign LUT_2[1400] = 32'b11111111111111111000100100011110;
assign LUT_2[1401] = 32'b11111111111111110101011100110111;
assign LUT_2[1402] = 32'b11111111111111111111011101011010;
assign LUT_2[1403] = 32'b11111111111111111100010101110011;
assign LUT_2[1404] = 32'b11111111111111110101000010000110;
assign LUT_2[1405] = 32'b11111111111111110001111010011111;
assign LUT_2[1406] = 32'b11111111111111111011111011000010;
assign LUT_2[1407] = 32'b11111111111111111000110011011011;
assign LUT_2[1408] = 32'b00000000000000001110111110111010;
assign LUT_2[1409] = 32'b00000000000000001011110111010011;
assign LUT_2[1410] = 32'b00000000000000010101110111110110;
assign LUT_2[1411] = 32'b00000000000000010010110000001111;
assign LUT_2[1412] = 32'b00000000000000001011011100100010;
assign LUT_2[1413] = 32'b00000000000000001000010100111011;
assign LUT_2[1414] = 32'b00000000000000010010010101011110;
assign LUT_2[1415] = 32'b00000000000000001111001101110111;
assign LUT_2[1416] = 32'b00000000000000001001110000010111;
assign LUT_2[1417] = 32'b00000000000000000110101000110000;
assign LUT_2[1418] = 32'b00000000000000010000101001010011;
assign LUT_2[1419] = 32'b00000000000000001101100001101100;
assign LUT_2[1420] = 32'b00000000000000000110001101111111;
assign LUT_2[1421] = 32'b00000000000000000011000110011000;
assign LUT_2[1422] = 32'b00000000000000001101000110111011;
assign LUT_2[1423] = 32'b00000000000000001001111111010100;
assign LUT_2[1424] = 32'b00000000000000001001100011000100;
assign LUT_2[1425] = 32'b00000000000000000110011011011101;
assign LUT_2[1426] = 32'b00000000000000010000011100000000;
assign LUT_2[1427] = 32'b00000000000000001101010100011001;
assign LUT_2[1428] = 32'b00000000000000000110000000101100;
assign LUT_2[1429] = 32'b00000000000000000010111001000101;
assign LUT_2[1430] = 32'b00000000000000001100111001101000;
assign LUT_2[1431] = 32'b00000000000000001001110010000001;
assign LUT_2[1432] = 32'b00000000000000000100010100100001;
assign LUT_2[1433] = 32'b00000000000000000001001100111010;
assign LUT_2[1434] = 32'b00000000000000001011001101011101;
assign LUT_2[1435] = 32'b00000000000000001000000101110110;
assign LUT_2[1436] = 32'b00000000000000000000110010001001;
assign LUT_2[1437] = 32'b11111111111111111101101010100010;
assign LUT_2[1438] = 32'b00000000000000000111101011000101;
assign LUT_2[1439] = 32'b00000000000000000100100011011110;
assign LUT_2[1440] = 32'b00000000000000001111011010100011;
assign LUT_2[1441] = 32'b00000000000000001100010010111100;
assign LUT_2[1442] = 32'b00000000000000010110010011011111;
assign LUT_2[1443] = 32'b00000000000000010011001011111000;
assign LUT_2[1444] = 32'b00000000000000001011111000001011;
assign LUT_2[1445] = 32'b00000000000000001000110000100100;
assign LUT_2[1446] = 32'b00000000000000010010110001000111;
assign LUT_2[1447] = 32'b00000000000000001111101001100000;
assign LUT_2[1448] = 32'b00000000000000001010001100000000;
assign LUT_2[1449] = 32'b00000000000000000111000100011001;
assign LUT_2[1450] = 32'b00000000000000010001000100111100;
assign LUT_2[1451] = 32'b00000000000000001101111101010101;
assign LUT_2[1452] = 32'b00000000000000000110101001101000;
assign LUT_2[1453] = 32'b00000000000000000011100010000001;
assign LUT_2[1454] = 32'b00000000000000001101100010100100;
assign LUT_2[1455] = 32'b00000000000000001010011010111101;
assign LUT_2[1456] = 32'b00000000000000001001111110101101;
assign LUT_2[1457] = 32'b00000000000000000110110111000110;
assign LUT_2[1458] = 32'b00000000000000010000110111101001;
assign LUT_2[1459] = 32'b00000000000000001101110000000010;
assign LUT_2[1460] = 32'b00000000000000000110011100010101;
assign LUT_2[1461] = 32'b00000000000000000011010100101110;
assign LUT_2[1462] = 32'b00000000000000001101010101010001;
assign LUT_2[1463] = 32'b00000000000000001010001101101010;
assign LUT_2[1464] = 32'b00000000000000000100110000001010;
assign LUT_2[1465] = 32'b00000000000000000001101000100011;
assign LUT_2[1466] = 32'b00000000000000001011101001000110;
assign LUT_2[1467] = 32'b00000000000000001000100001011111;
assign LUT_2[1468] = 32'b00000000000000000001001101110010;
assign LUT_2[1469] = 32'b11111111111111111110000110001011;
assign LUT_2[1470] = 32'b00000000000000001000000110101110;
assign LUT_2[1471] = 32'b00000000000000000100111111000111;
assign LUT_2[1472] = 32'b00000000000000000111000111011101;
assign LUT_2[1473] = 32'b00000000000000000011111111110110;
assign LUT_2[1474] = 32'b00000000000000001110000000011001;
assign LUT_2[1475] = 32'b00000000000000001010111000110010;
assign LUT_2[1476] = 32'b00000000000000000011100101000101;
assign LUT_2[1477] = 32'b00000000000000000000011101011110;
assign LUT_2[1478] = 32'b00000000000000001010011110000001;
assign LUT_2[1479] = 32'b00000000000000000111010110011010;
assign LUT_2[1480] = 32'b00000000000000000001111000111010;
assign LUT_2[1481] = 32'b11111111111111111110110001010011;
assign LUT_2[1482] = 32'b00000000000000001000110001110110;
assign LUT_2[1483] = 32'b00000000000000000101101010001111;
assign LUT_2[1484] = 32'b11111111111111111110010110100010;
assign LUT_2[1485] = 32'b11111111111111111011001110111011;
assign LUT_2[1486] = 32'b00000000000000000101001111011110;
assign LUT_2[1487] = 32'b00000000000000000010000111110111;
assign LUT_2[1488] = 32'b00000000000000000001101011100111;
assign LUT_2[1489] = 32'b11111111111111111110100100000000;
assign LUT_2[1490] = 32'b00000000000000001000100100100011;
assign LUT_2[1491] = 32'b00000000000000000101011100111100;
assign LUT_2[1492] = 32'b11111111111111111110001001001111;
assign LUT_2[1493] = 32'b11111111111111111011000001101000;
assign LUT_2[1494] = 32'b00000000000000000101000010001011;
assign LUT_2[1495] = 32'b00000000000000000001111010100100;
assign LUT_2[1496] = 32'b11111111111111111100011101000100;
assign LUT_2[1497] = 32'b11111111111111111001010101011101;
assign LUT_2[1498] = 32'b00000000000000000011010110000000;
assign LUT_2[1499] = 32'b00000000000000000000001110011001;
assign LUT_2[1500] = 32'b11111111111111111000111010101100;
assign LUT_2[1501] = 32'b11111111111111110101110011000101;
assign LUT_2[1502] = 32'b11111111111111111111110011101000;
assign LUT_2[1503] = 32'b11111111111111111100101100000001;
assign LUT_2[1504] = 32'b00000000000000000111100011000110;
assign LUT_2[1505] = 32'b00000000000000000100011011011111;
assign LUT_2[1506] = 32'b00000000000000001110011100000010;
assign LUT_2[1507] = 32'b00000000000000001011010100011011;
assign LUT_2[1508] = 32'b00000000000000000100000000101110;
assign LUT_2[1509] = 32'b00000000000000000000111001000111;
assign LUT_2[1510] = 32'b00000000000000001010111001101010;
assign LUT_2[1511] = 32'b00000000000000000111110010000011;
assign LUT_2[1512] = 32'b00000000000000000010010100100011;
assign LUT_2[1513] = 32'b11111111111111111111001100111100;
assign LUT_2[1514] = 32'b00000000000000001001001101011111;
assign LUT_2[1515] = 32'b00000000000000000110000101111000;
assign LUT_2[1516] = 32'b11111111111111111110110010001011;
assign LUT_2[1517] = 32'b11111111111111111011101010100100;
assign LUT_2[1518] = 32'b00000000000000000101101011000111;
assign LUT_2[1519] = 32'b00000000000000000010100011100000;
assign LUT_2[1520] = 32'b00000000000000000010000111010000;
assign LUT_2[1521] = 32'b11111111111111111110111111101001;
assign LUT_2[1522] = 32'b00000000000000001001000000001100;
assign LUT_2[1523] = 32'b00000000000000000101111000100101;
assign LUT_2[1524] = 32'b11111111111111111110100100111000;
assign LUT_2[1525] = 32'b11111111111111111011011101010001;
assign LUT_2[1526] = 32'b00000000000000000101011101110100;
assign LUT_2[1527] = 32'b00000000000000000010010110001101;
assign LUT_2[1528] = 32'b11111111111111111100111000101101;
assign LUT_2[1529] = 32'b11111111111111111001110001000110;
assign LUT_2[1530] = 32'b00000000000000000011110001101001;
assign LUT_2[1531] = 32'b00000000000000000000101010000010;
assign LUT_2[1532] = 32'b11111111111111111001010110010101;
assign LUT_2[1533] = 32'b11111111111111110110001110101110;
assign LUT_2[1534] = 32'b00000000000000000000001111010001;
assign LUT_2[1535] = 32'b11111111111111111101000111101010;
assign LUT_2[1536] = 32'b00000000000000001011011101110111;
assign LUT_2[1537] = 32'b00000000000000001000010110010000;
assign LUT_2[1538] = 32'b00000000000000010010010110110011;
assign LUT_2[1539] = 32'b00000000000000001111001111001100;
assign LUT_2[1540] = 32'b00000000000000000111111011011111;
assign LUT_2[1541] = 32'b00000000000000000100110011111000;
assign LUT_2[1542] = 32'b00000000000000001110110100011011;
assign LUT_2[1543] = 32'b00000000000000001011101100110100;
assign LUT_2[1544] = 32'b00000000000000000110001111010100;
assign LUT_2[1545] = 32'b00000000000000000011000111101101;
assign LUT_2[1546] = 32'b00000000000000001101001000010000;
assign LUT_2[1547] = 32'b00000000000000001010000000101001;
assign LUT_2[1548] = 32'b00000000000000000010101100111100;
assign LUT_2[1549] = 32'b11111111111111111111100101010101;
assign LUT_2[1550] = 32'b00000000000000001001100101111000;
assign LUT_2[1551] = 32'b00000000000000000110011110010001;
assign LUT_2[1552] = 32'b00000000000000000110000010000001;
assign LUT_2[1553] = 32'b00000000000000000010111010011010;
assign LUT_2[1554] = 32'b00000000000000001100111010111101;
assign LUT_2[1555] = 32'b00000000000000001001110011010110;
assign LUT_2[1556] = 32'b00000000000000000010011111101001;
assign LUT_2[1557] = 32'b11111111111111111111011000000010;
assign LUT_2[1558] = 32'b00000000000000001001011000100101;
assign LUT_2[1559] = 32'b00000000000000000110010000111110;
assign LUT_2[1560] = 32'b00000000000000000000110011011110;
assign LUT_2[1561] = 32'b11111111111111111101101011110111;
assign LUT_2[1562] = 32'b00000000000000000111101100011010;
assign LUT_2[1563] = 32'b00000000000000000100100100110011;
assign LUT_2[1564] = 32'b11111111111111111101010001000110;
assign LUT_2[1565] = 32'b11111111111111111010001001011111;
assign LUT_2[1566] = 32'b00000000000000000100001010000010;
assign LUT_2[1567] = 32'b00000000000000000001000010011011;
assign LUT_2[1568] = 32'b00000000000000001011111001100000;
assign LUT_2[1569] = 32'b00000000000000001000110001111001;
assign LUT_2[1570] = 32'b00000000000000010010110010011100;
assign LUT_2[1571] = 32'b00000000000000001111101010110101;
assign LUT_2[1572] = 32'b00000000000000001000010111001000;
assign LUT_2[1573] = 32'b00000000000000000101001111100001;
assign LUT_2[1574] = 32'b00000000000000001111010000000100;
assign LUT_2[1575] = 32'b00000000000000001100001000011101;
assign LUT_2[1576] = 32'b00000000000000000110101010111101;
assign LUT_2[1577] = 32'b00000000000000000011100011010110;
assign LUT_2[1578] = 32'b00000000000000001101100011111001;
assign LUT_2[1579] = 32'b00000000000000001010011100010010;
assign LUT_2[1580] = 32'b00000000000000000011001000100101;
assign LUT_2[1581] = 32'b00000000000000000000000000111110;
assign LUT_2[1582] = 32'b00000000000000001010000001100001;
assign LUT_2[1583] = 32'b00000000000000000110111001111010;
assign LUT_2[1584] = 32'b00000000000000000110011101101010;
assign LUT_2[1585] = 32'b00000000000000000011010110000011;
assign LUT_2[1586] = 32'b00000000000000001101010110100110;
assign LUT_2[1587] = 32'b00000000000000001010001110111111;
assign LUT_2[1588] = 32'b00000000000000000010111011010010;
assign LUT_2[1589] = 32'b11111111111111111111110011101011;
assign LUT_2[1590] = 32'b00000000000000001001110100001110;
assign LUT_2[1591] = 32'b00000000000000000110101100100111;
assign LUT_2[1592] = 32'b00000000000000000001001111000111;
assign LUT_2[1593] = 32'b11111111111111111110000111100000;
assign LUT_2[1594] = 32'b00000000000000001000001000000011;
assign LUT_2[1595] = 32'b00000000000000000101000000011100;
assign LUT_2[1596] = 32'b11111111111111111101101100101111;
assign LUT_2[1597] = 32'b11111111111111111010100101001000;
assign LUT_2[1598] = 32'b00000000000000000100100101101011;
assign LUT_2[1599] = 32'b00000000000000000001011110000100;
assign LUT_2[1600] = 32'b00000000000000000011100110011010;
assign LUT_2[1601] = 32'b00000000000000000000011110110011;
assign LUT_2[1602] = 32'b00000000000000001010011111010110;
assign LUT_2[1603] = 32'b00000000000000000111010111101111;
assign LUT_2[1604] = 32'b00000000000000000000000100000010;
assign LUT_2[1605] = 32'b11111111111111111100111100011011;
assign LUT_2[1606] = 32'b00000000000000000110111100111110;
assign LUT_2[1607] = 32'b00000000000000000011110101010111;
assign LUT_2[1608] = 32'b11111111111111111110010111110111;
assign LUT_2[1609] = 32'b11111111111111111011010000010000;
assign LUT_2[1610] = 32'b00000000000000000101010000110011;
assign LUT_2[1611] = 32'b00000000000000000010001001001100;
assign LUT_2[1612] = 32'b11111111111111111010110101011111;
assign LUT_2[1613] = 32'b11111111111111110111101101111000;
assign LUT_2[1614] = 32'b00000000000000000001101110011011;
assign LUT_2[1615] = 32'b11111111111111111110100110110100;
assign LUT_2[1616] = 32'b11111111111111111110001010100100;
assign LUT_2[1617] = 32'b11111111111111111011000010111101;
assign LUT_2[1618] = 32'b00000000000000000101000011100000;
assign LUT_2[1619] = 32'b00000000000000000001111011111001;
assign LUT_2[1620] = 32'b11111111111111111010101000001100;
assign LUT_2[1621] = 32'b11111111111111110111100000100101;
assign LUT_2[1622] = 32'b00000000000000000001100001001000;
assign LUT_2[1623] = 32'b11111111111111111110011001100001;
assign LUT_2[1624] = 32'b11111111111111111000111100000001;
assign LUT_2[1625] = 32'b11111111111111110101110100011010;
assign LUT_2[1626] = 32'b11111111111111111111110100111101;
assign LUT_2[1627] = 32'b11111111111111111100101101010110;
assign LUT_2[1628] = 32'b11111111111111110101011001101001;
assign LUT_2[1629] = 32'b11111111111111110010010010000010;
assign LUT_2[1630] = 32'b11111111111111111100010010100101;
assign LUT_2[1631] = 32'b11111111111111111001001010111110;
assign LUT_2[1632] = 32'b00000000000000000100000010000011;
assign LUT_2[1633] = 32'b00000000000000000000111010011100;
assign LUT_2[1634] = 32'b00000000000000001010111010111111;
assign LUT_2[1635] = 32'b00000000000000000111110011011000;
assign LUT_2[1636] = 32'b00000000000000000000011111101011;
assign LUT_2[1637] = 32'b11111111111111111101011000000100;
assign LUT_2[1638] = 32'b00000000000000000111011000100111;
assign LUT_2[1639] = 32'b00000000000000000100010001000000;
assign LUT_2[1640] = 32'b11111111111111111110110011100000;
assign LUT_2[1641] = 32'b11111111111111111011101011111001;
assign LUT_2[1642] = 32'b00000000000000000101101100011100;
assign LUT_2[1643] = 32'b00000000000000000010100100110101;
assign LUT_2[1644] = 32'b11111111111111111011010001001000;
assign LUT_2[1645] = 32'b11111111111111111000001001100001;
assign LUT_2[1646] = 32'b00000000000000000010001010000100;
assign LUT_2[1647] = 32'b11111111111111111111000010011101;
assign LUT_2[1648] = 32'b11111111111111111110100110001101;
assign LUT_2[1649] = 32'b11111111111111111011011110100110;
assign LUT_2[1650] = 32'b00000000000000000101011111001001;
assign LUT_2[1651] = 32'b00000000000000000010010111100010;
assign LUT_2[1652] = 32'b11111111111111111011000011110101;
assign LUT_2[1653] = 32'b11111111111111110111111100001110;
assign LUT_2[1654] = 32'b00000000000000000001111100110001;
assign LUT_2[1655] = 32'b11111111111111111110110101001010;
assign LUT_2[1656] = 32'b11111111111111111001010111101010;
assign LUT_2[1657] = 32'b11111111111111110110010000000011;
assign LUT_2[1658] = 32'b00000000000000000000010000100110;
assign LUT_2[1659] = 32'b11111111111111111101001000111111;
assign LUT_2[1660] = 32'b11111111111111110101110101010010;
assign LUT_2[1661] = 32'b11111111111111110010101101101011;
assign LUT_2[1662] = 32'b11111111111111111100101110001110;
assign LUT_2[1663] = 32'b11111111111111111001100110100111;
assign LUT_2[1664] = 32'b00000000000000001111110010000110;
assign LUT_2[1665] = 32'b00000000000000001100101010011111;
assign LUT_2[1666] = 32'b00000000000000010110101011000010;
assign LUT_2[1667] = 32'b00000000000000010011100011011011;
assign LUT_2[1668] = 32'b00000000000000001100001111101110;
assign LUT_2[1669] = 32'b00000000000000001001001000000111;
assign LUT_2[1670] = 32'b00000000000000010011001000101010;
assign LUT_2[1671] = 32'b00000000000000010000000001000011;
assign LUT_2[1672] = 32'b00000000000000001010100011100011;
assign LUT_2[1673] = 32'b00000000000000000111011011111100;
assign LUT_2[1674] = 32'b00000000000000010001011100011111;
assign LUT_2[1675] = 32'b00000000000000001110010100111000;
assign LUT_2[1676] = 32'b00000000000000000111000001001011;
assign LUT_2[1677] = 32'b00000000000000000011111001100100;
assign LUT_2[1678] = 32'b00000000000000001101111010000111;
assign LUT_2[1679] = 32'b00000000000000001010110010100000;
assign LUT_2[1680] = 32'b00000000000000001010010110010000;
assign LUT_2[1681] = 32'b00000000000000000111001110101001;
assign LUT_2[1682] = 32'b00000000000000010001001111001100;
assign LUT_2[1683] = 32'b00000000000000001110000111100101;
assign LUT_2[1684] = 32'b00000000000000000110110011111000;
assign LUT_2[1685] = 32'b00000000000000000011101100010001;
assign LUT_2[1686] = 32'b00000000000000001101101100110100;
assign LUT_2[1687] = 32'b00000000000000001010100101001101;
assign LUT_2[1688] = 32'b00000000000000000101000111101101;
assign LUT_2[1689] = 32'b00000000000000000010000000000110;
assign LUT_2[1690] = 32'b00000000000000001100000000101001;
assign LUT_2[1691] = 32'b00000000000000001000111001000010;
assign LUT_2[1692] = 32'b00000000000000000001100101010101;
assign LUT_2[1693] = 32'b11111111111111111110011101101110;
assign LUT_2[1694] = 32'b00000000000000001000011110010001;
assign LUT_2[1695] = 32'b00000000000000000101010110101010;
assign LUT_2[1696] = 32'b00000000000000010000001101101111;
assign LUT_2[1697] = 32'b00000000000000001101000110001000;
assign LUT_2[1698] = 32'b00000000000000010111000110101011;
assign LUT_2[1699] = 32'b00000000000000010011111111000100;
assign LUT_2[1700] = 32'b00000000000000001100101011010111;
assign LUT_2[1701] = 32'b00000000000000001001100011110000;
assign LUT_2[1702] = 32'b00000000000000010011100100010011;
assign LUT_2[1703] = 32'b00000000000000010000011100101100;
assign LUT_2[1704] = 32'b00000000000000001010111111001100;
assign LUT_2[1705] = 32'b00000000000000000111110111100101;
assign LUT_2[1706] = 32'b00000000000000010001111000001000;
assign LUT_2[1707] = 32'b00000000000000001110110000100001;
assign LUT_2[1708] = 32'b00000000000000000111011100110100;
assign LUT_2[1709] = 32'b00000000000000000100010101001101;
assign LUT_2[1710] = 32'b00000000000000001110010101110000;
assign LUT_2[1711] = 32'b00000000000000001011001110001001;
assign LUT_2[1712] = 32'b00000000000000001010110001111001;
assign LUT_2[1713] = 32'b00000000000000000111101010010010;
assign LUT_2[1714] = 32'b00000000000000010001101010110101;
assign LUT_2[1715] = 32'b00000000000000001110100011001110;
assign LUT_2[1716] = 32'b00000000000000000111001111100001;
assign LUT_2[1717] = 32'b00000000000000000100000111111010;
assign LUT_2[1718] = 32'b00000000000000001110001000011101;
assign LUT_2[1719] = 32'b00000000000000001011000000110110;
assign LUT_2[1720] = 32'b00000000000000000101100011010110;
assign LUT_2[1721] = 32'b00000000000000000010011011101111;
assign LUT_2[1722] = 32'b00000000000000001100011100010010;
assign LUT_2[1723] = 32'b00000000000000001001010100101011;
assign LUT_2[1724] = 32'b00000000000000000010000000111110;
assign LUT_2[1725] = 32'b11111111111111111110111001010111;
assign LUT_2[1726] = 32'b00000000000000001000111001111010;
assign LUT_2[1727] = 32'b00000000000000000101110010010011;
assign LUT_2[1728] = 32'b00000000000000000111111010101001;
assign LUT_2[1729] = 32'b00000000000000000100110011000010;
assign LUT_2[1730] = 32'b00000000000000001110110011100101;
assign LUT_2[1731] = 32'b00000000000000001011101011111110;
assign LUT_2[1732] = 32'b00000000000000000100011000010001;
assign LUT_2[1733] = 32'b00000000000000000001010000101010;
assign LUT_2[1734] = 32'b00000000000000001011010001001101;
assign LUT_2[1735] = 32'b00000000000000001000001001100110;
assign LUT_2[1736] = 32'b00000000000000000010101100000110;
assign LUT_2[1737] = 32'b11111111111111111111100100011111;
assign LUT_2[1738] = 32'b00000000000000001001100101000010;
assign LUT_2[1739] = 32'b00000000000000000110011101011011;
assign LUT_2[1740] = 32'b11111111111111111111001001101110;
assign LUT_2[1741] = 32'b11111111111111111100000010000111;
assign LUT_2[1742] = 32'b00000000000000000110000010101010;
assign LUT_2[1743] = 32'b00000000000000000010111011000011;
assign LUT_2[1744] = 32'b00000000000000000010011110110011;
assign LUT_2[1745] = 32'b11111111111111111111010111001100;
assign LUT_2[1746] = 32'b00000000000000001001010111101111;
assign LUT_2[1747] = 32'b00000000000000000110010000001000;
assign LUT_2[1748] = 32'b11111111111111111110111100011011;
assign LUT_2[1749] = 32'b11111111111111111011110100110100;
assign LUT_2[1750] = 32'b00000000000000000101110101010111;
assign LUT_2[1751] = 32'b00000000000000000010101101110000;
assign LUT_2[1752] = 32'b11111111111111111101010000010000;
assign LUT_2[1753] = 32'b11111111111111111010001000101001;
assign LUT_2[1754] = 32'b00000000000000000100001001001100;
assign LUT_2[1755] = 32'b00000000000000000001000001100101;
assign LUT_2[1756] = 32'b11111111111111111001101101111000;
assign LUT_2[1757] = 32'b11111111111111110110100110010001;
assign LUT_2[1758] = 32'b00000000000000000000100110110100;
assign LUT_2[1759] = 32'b11111111111111111101011111001101;
assign LUT_2[1760] = 32'b00000000000000001000010110010010;
assign LUT_2[1761] = 32'b00000000000000000101001110101011;
assign LUT_2[1762] = 32'b00000000000000001111001111001110;
assign LUT_2[1763] = 32'b00000000000000001100000111100111;
assign LUT_2[1764] = 32'b00000000000000000100110011111010;
assign LUT_2[1765] = 32'b00000000000000000001101100010011;
assign LUT_2[1766] = 32'b00000000000000001011101100110110;
assign LUT_2[1767] = 32'b00000000000000001000100101001111;
assign LUT_2[1768] = 32'b00000000000000000011000111101111;
assign LUT_2[1769] = 32'b00000000000000000000000000001000;
assign LUT_2[1770] = 32'b00000000000000001010000000101011;
assign LUT_2[1771] = 32'b00000000000000000110111001000100;
assign LUT_2[1772] = 32'b11111111111111111111100101010111;
assign LUT_2[1773] = 32'b11111111111111111100011101110000;
assign LUT_2[1774] = 32'b00000000000000000110011110010011;
assign LUT_2[1775] = 32'b00000000000000000011010110101100;
assign LUT_2[1776] = 32'b00000000000000000010111010011100;
assign LUT_2[1777] = 32'b11111111111111111111110010110101;
assign LUT_2[1778] = 32'b00000000000000001001110011011000;
assign LUT_2[1779] = 32'b00000000000000000110101011110001;
assign LUT_2[1780] = 32'b11111111111111111111011000000100;
assign LUT_2[1781] = 32'b11111111111111111100010000011101;
assign LUT_2[1782] = 32'b00000000000000000110010001000000;
assign LUT_2[1783] = 32'b00000000000000000011001001011001;
assign LUT_2[1784] = 32'b11111111111111111101101011111001;
assign LUT_2[1785] = 32'b11111111111111111010100100010010;
assign LUT_2[1786] = 32'b00000000000000000100100100110101;
assign LUT_2[1787] = 32'b00000000000000000001011101001110;
assign LUT_2[1788] = 32'b11111111111111111010001001100001;
assign LUT_2[1789] = 32'b11111111111111110111000001111010;
assign LUT_2[1790] = 32'b00000000000000000001000010011101;
assign LUT_2[1791] = 32'b11111111111111111101111010110110;
assign LUT_2[1792] = 32'b00000000000000001111011100011101;
assign LUT_2[1793] = 32'b00000000000000001100010100110110;
assign LUT_2[1794] = 32'b00000000000000010110010101011001;
assign LUT_2[1795] = 32'b00000000000000010011001101110010;
assign LUT_2[1796] = 32'b00000000000000001011111010000101;
assign LUT_2[1797] = 32'b00000000000000001000110010011110;
assign LUT_2[1798] = 32'b00000000000000010010110011000001;
assign LUT_2[1799] = 32'b00000000000000001111101011011010;
assign LUT_2[1800] = 32'b00000000000000001010001101111010;
assign LUT_2[1801] = 32'b00000000000000000111000110010011;
assign LUT_2[1802] = 32'b00000000000000010001000110110110;
assign LUT_2[1803] = 32'b00000000000000001101111111001111;
assign LUT_2[1804] = 32'b00000000000000000110101011100010;
assign LUT_2[1805] = 32'b00000000000000000011100011111011;
assign LUT_2[1806] = 32'b00000000000000001101100100011110;
assign LUT_2[1807] = 32'b00000000000000001010011100110111;
assign LUT_2[1808] = 32'b00000000000000001010000000100111;
assign LUT_2[1809] = 32'b00000000000000000110111001000000;
assign LUT_2[1810] = 32'b00000000000000010000111001100011;
assign LUT_2[1811] = 32'b00000000000000001101110001111100;
assign LUT_2[1812] = 32'b00000000000000000110011110001111;
assign LUT_2[1813] = 32'b00000000000000000011010110101000;
assign LUT_2[1814] = 32'b00000000000000001101010111001011;
assign LUT_2[1815] = 32'b00000000000000001010001111100100;
assign LUT_2[1816] = 32'b00000000000000000100110010000100;
assign LUT_2[1817] = 32'b00000000000000000001101010011101;
assign LUT_2[1818] = 32'b00000000000000001011101011000000;
assign LUT_2[1819] = 32'b00000000000000001000100011011001;
assign LUT_2[1820] = 32'b00000000000000000001001111101100;
assign LUT_2[1821] = 32'b11111111111111111110001000000101;
assign LUT_2[1822] = 32'b00000000000000001000001000101000;
assign LUT_2[1823] = 32'b00000000000000000101000001000001;
assign LUT_2[1824] = 32'b00000000000000001111111000000110;
assign LUT_2[1825] = 32'b00000000000000001100110000011111;
assign LUT_2[1826] = 32'b00000000000000010110110001000010;
assign LUT_2[1827] = 32'b00000000000000010011101001011011;
assign LUT_2[1828] = 32'b00000000000000001100010101101110;
assign LUT_2[1829] = 32'b00000000000000001001001110000111;
assign LUT_2[1830] = 32'b00000000000000010011001110101010;
assign LUT_2[1831] = 32'b00000000000000010000000111000011;
assign LUT_2[1832] = 32'b00000000000000001010101001100011;
assign LUT_2[1833] = 32'b00000000000000000111100001111100;
assign LUT_2[1834] = 32'b00000000000000010001100010011111;
assign LUT_2[1835] = 32'b00000000000000001110011010111000;
assign LUT_2[1836] = 32'b00000000000000000111000111001011;
assign LUT_2[1837] = 32'b00000000000000000011111111100100;
assign LUT_2[1838] = 32'b00000000000000001110000000000111;
assign LUT_2[1839] = 32'b00000000000000001010111000100000;
assign LUT_2[1840] = 32'b00000000000000001010011100010000;
assign LUT_2[1841] = 32'b00000000000000000111010100101001;
assign LUT_2[1842] = 32'b00000000000000010001010101001100;
assign LUT_2[1843] = 32'b00000000000000001110001101100101;
assign LUT_2[1844] = 32'b00000000000000000110111001111000;
assign LUT_2[1845] = 32'b00000000000000000011110010010001;
assign LUT_2[1846] = 32'b00000000000000001101110010110100;
assign LUT_2[1847] = 32'b00000000000000001010101011001101;
assign LUT_2[1848] = 32'b00000000000000000101001101101101;
assign LUT_2[1849] = 32'b00000000000000000010000110000110;
assign LUT_2[1850] = 32'b00000000000000001100000110101001;
assign LUT_2[1851] = 32'b00000000000000001000111111000010;
assign LUT_2[1852] = 32'b00000000000000000001101011010101;
assign LUT_2[1853] = 32'b11111111111111111110100011101110;
assign LUT_2[1854] = 32'b00000000000000001000100100010001;
assign LUT_2[1855] = 32'b00000000000000000101011100101010;
assign LUT_2[1856] = 32'b00000000000000000111100101000000;
assign LUT_2[1857] = 32'b00000000000000000100011101011001;
assign LUT_2[1858] = 32'b00000000000000001110011101111100;
assign LUT_2[1859] = 32'b00000000000000001011010110010101;
assign LUT_2[1860] = 32'b00000000000000000100000010101000;
assign LUT_2[1861] = 32'b00000000000000000000111011000001;
assign LUT_2[1862] = 32'b00000000000000001010111011100100;
assign LUT_2[1863] = 32'b00000000000000000111110011111101;
assign LUT_2[1864] = 32'b00000000000000000010010110011101;
assign LUT_2[1865] = 32'b11111111111111111111001110110110;
assign LUT_2[1866] = 32'b00000000000000001001001111011001;
assign LUT_2[1867] = 32'b00000000000000000110000111110010;
assign LUT_2[1868] = 32'b11111111111111111110110100000101;
assign LUT_2[1869] = 32'b11111111111111111011101100011110;
assign LUT_2[1870] = 32'b00000000000000000101101101000001;
assign LUT_2[1871] = 32'b00000000000000000010100101011010;
assign LUT_2[1872] = 32'b00000000000000000010001001001010;
assign LUT_2[1873] = 32'b11111111111111111111000001100011;
assign LUT_2[1874] = 32'b00000000000000001001000010000110;
assign LUT_2[1875] = 32'b00000000000000000101111010011111;
assign LUT_2[1876] = 32'b11111111111111111110100110110010;
assign LUT_2[1877] = 32'b11111111111111111011011111001011;
assign LUT_2[1878] = 32'b00000000000000000101011111101110;
assign LUT_2[1879] = 32'b00000000000000000010011000000111;
assign LUT_2[1880] = 32'b11111111111111111100111010100111;
assign LUT_2[1881] = 32'b11111111111111111001110011000000;
assign LUT_2[1882] = 32'b00000000000000000011110011100011;
assign LUT_2[1883] = 32'b00000000000000000000101011111100;
assign LUT_2[1884] = 32'b11111111111111111001011000001111;
assign LUT_2[1885] = 32'b11111111111111110110010000101000;
assign LUT_2[1886] = 32'b00000000000000000000010001001011;
assign LUT_2[1887] = 32'b11111111111111111101001001100100;
assign LUT_2[1888] = 32'b00000000000000001000000000101001;
assign LUT_2[1889] = 32'b00000000000000000100111001000010;
assign LUT_2[1890] = 32'b00000000000000001110111001100101;
assign LUT_2[1891] = 32'b00000000000000001011110001111110;
assign LUT_2[1892] = 32'b00000000000000000100011110010001;
assign LUT_2[1893] = 32'b00000000000000000001010110101010;
assign LUT_2[1894] = 32'b00000000000000001011010111001101;
assign LUT_2[1895] = 32'b00000000000000001000001111100110;
assign LUT_2[1896] = 32'b00000000000000000010110010000110;
assign LUT_2[1897] = 32'b11111111111111111111101010011111;
assign LUT_2[1898] = 32'b00000000000000001001101011000010;
assign LUT_2[1899] = 32'b00000000000000000110100011011011;
assign LUT_2[1900] = 32'b11111111111111111111001111101110;
assign LUT_2[1901] = 32'b11111111111111111100001000000111;
assign LUT_2[1902] = 32'b00000000000000000110001000101010;
assign LUT_2[1903] = 32'b00000000000000000011000001000011;
assign LUT_2[1904] = 32'b00000000000000000010100100110011;
assign LUT_2[1905] = 32'b11111111111111111111011101001100;
assign LUT_2[1906] = 32'b00000000000000001001011101101111;
assign LUT_2[1907] = 32'b00000000000000000110010110001000;
assign LUT_2[1908] = 32'b11111111111111111111000010011011;
assign LUT_2[1909] = 32'b11111111111111111011111010110100;
assign LUT_2[1910] = 32'b00000000000000000101111011010111;
assign LUT_2[1911] = 32'b00000000000000000010110011110000;
assign LUT_2[1912] = 32'b11111111111111111101010110010000;
assign LUT_2[1913] = 32'b11111111111111111010001110101001;
assign LUT_2[1914] = 32'b00000000000000000100001111001100;
assign LUT_2[1915] = 32'b00000000000000000001000111100101;
assign LUT_2[1916] = 32'b11111111111111111001110011111000;
assign LUT_2[1917] = 32'b11111111111111110110101100010001;
assign LUT_2[1918] = 32'b00000000000000000000101100110100;
assign LUT_2[1919] = 32'b11111111111111111101100101001101;
assign LUT_2[1920] = 32'b00000000000000010011110000101100;
assign LUT_2[1921] = 32'b00000000000000010000101001000101;
assign LUT_2[1922] = 32'b00000000000000011010101001101000;
assign LUT_2[1923] = 32'b00000000000000010111100010000001;
assign LUT_2[1924] = 32'b00000000000000010000001110010100;
assign LUT_2[1925] = 32'b00000000000000001101000110101101;
assign LUT_2[1926] = 32'b00000000000000010111000111010000;
assign LUT_2[1927] = 32'b00000000000000010011111111101001;
assign LUT_2[1928] = 32'b00000000000000001110100010001001;
assign LUT_2[1929] = 32'b00000000000000001011011010100010;
assign LUT_2[1930] = 32'b00000000000000010101011011000101;
assign LUT_2[1931] = 32'b00000000000000010010010011011110;
assign LUT_2[1932] = 32'b00000000000000001010111111110001;
assign LUT_2[1933] = 32'b00000000000000000111111000001010;
assign LUT_2[1934] = 32'b00000000000000010001111000101101;
assign LUT_2[1935] = 32'b00000000000000001110110001000110;
assign LUT_2[1936] = 32'b00000000000000001110010100110110;
assign LUT_2[1937] = 32'b00000000000000001011001101001111;
assign LUT_2[1938] = 32'b00000000000000010101001101110010;
assign LUT_2[1939] = 32'b00000000000000010010000110001011;
assign LUT_2[1940] = 32'b00000000000000001010110010011110;
assign LUT_2[1941] = 32'b00000000000000000111101010110111;
assign LUT_2[1942] = 32'b00000000000000010001101011011010;
assign LUT_2[1943] = 32'b00000000000000001110100011110011;
assign LUT_2[1944] = 32'b00000000000000001001000110010011;
assign LUT_2[1945] = 32'b00000000000000000101111110101100;
assign LUT_2[1946] = 32'b00000000000000001111111111001111;
assign LUT_2[1947] = 32'b00000000000000001100110111101000;
assign LUT_2[1948] = 32'b00000000000000000101100011111011;
assign LUT_2[1949] = 32'b00000000000000000010011100010100;
assign LUT_2[1950] = 32'b00000000000000001100011100110111;
assign LUT_2[1951] = 32'b00000000000000001001010101010000;
assign LUT_2[1952] = 32'b00000000000000010100001100010101;
assign LUT_2[1953] = 32'b00000000000000010001000100101110;
assign LUT_2[1954] = 32'b00000000000000011011000101010001;
assign LUT_2[1955] = 32'b00000000000000010111111101101010;
assign LUT_2[1956] = 32'b00000000000000010000101001111101;
assign LUT_2[1957] = 32'b00000000000000001101100010010110;
assign LUT_2[1958] = 32'b00000000000000010111100010111001;
assign LUT_2[1959] = 32'b00000000000000010100011011010010;
assign LUT_2[1960] = 32'b00000000000000001110111101110010;
assign LUT_2[1961] = 32'b00000000000000001011110110001011;
assign LUT_2[1962] = 32'b00000000000000010101110110101110;
assign LUT_2[1963] = 32'b00000000000000010010101111000111;
assign LUT_2[1964] = 32'b00000000000000001011011011011010;
assign LUT_2[1965] = 32'b00000000000000001000010011110011;
assign LUT_2[1966] = 32'b00000000000000010010010100010110;
assign LUT_2[1967] = 32'b00000000000000001111001100101111;
assign LUT_2[1968] = 32'b00000000000000001110110000011111;
assign LUT_2[1969] = 32'b00000000000000001011101000111000;
assign LUT_2[1970] = 32'b00000000000000010101101001011011;
assign LUT_2[1971] = 32'b00000000000000010010100001110100;
assign LUT_2[1972] = 32'b00000000000000001011001110000111;
assign LUT_2[1973] = 32'b00000000000000001000000110100000;
assign LUT_2[1974] = 32'b00000000000000010010000111000011;
assign LUT_2[1975] = 32'b00000000000000001110111111011100;
assign LUT_2[1976] = 32'b00000000000000001001100001111100;
assign LUT_2[1977] = 32'b00000000000000000110011010010101;
assign LUT_2[1978] = 32'b00000000000000010000011010111000;
assign LUT_2[1979] = 32'b00000000000000001101010011010001;
assign LUT_2[1980] = 32'b00000000000000000101111111100100;
assign LUT_2[1981] = 32'b00000000000000000010110111111101;
assign LUT_2[1982] = 32'b00000000000000001100111000100000;
assign LUT_2[1983] = 32'b00000000000000001001110000111001;
assign LUT_2[1984] = 32'b00000000000000001011111001001111;
assign LUT_2[1985] = 32'b00000000000000001000110001101000;
assign LUT_2[1986] = 32'b00000000000000010010110010001011;
assign LUT_2[1987] = 32'b00000000000000001111101010100100;
assign LUT_2[1988] = 32'b00000000000000001000010110110111;
assign LUT_2[1989] = 32'b00000000000000000101001111010000;
assign LUT_2[1990] = 32'b00000000000000001111001111110011;
assign LUT_2[1991] = 32'b00000000000000001100001000001100;
assign LUT_2[1992] = 32'b00000000000000000110101010101100;
assign LUT_2[1993] = 32'b00000000000000000011100011000101;
assign LUT_2[1994] = 32'b00000000000000001101100011101000;
assign LUT_2[1995] = 32'b00000000000000001010011100000001;
assign LUT_2[1996] = 32'b00000000000000000011001000010100;
assign LUT_2[1997] = 32'b00000000000000000000000000101101;
assign LUT_2[1998] = 32'b00000000000000001010000001010000;
assign LUT_2[1999] = 32'b00000000000000000110111001101001;
assign LUT_2[2000] = 32'b00000000000000000110011101011001;
assign LUT_2[2001] = 32'b00000000000000000011010101110010;
assign LUT_2[2002] = 32'b00000000000000001101010110010101;
assign LUT_2[2003] = 32'b00000000000000001010001110101110;
assign LUT_2[2004] = 32'b00000000000000000010111011000001;
assign LUT_2[2005] = 32'b11111111111111111111110011011010;
assign LUT_2[2006] = 32'b00000000000000001001110011111101;
assign LUT_2[2007] = 32'b00000000000000000110101100010110;
assign LUT_2[2008] = 32'b00000000000000000001001110110110;
assign LUT_2[2009] = 32'b11111111111111111110000111001111;
assign LUT_2[2010] = 32'b00000000000000001000000111110010;
assign LUT_2[2011] = 32'b00000000000000000101000000001011;
assign LUT_2[2012] = 32'b11111111111111111101101100011110;
assign LUT_2[2013] = 32'b11111111111111111010100100110111;
assign LUT_2[2014] = 32'b00000000000000000100100101011010;
assign LUT_2[2015] = 32'b00000000000000000001011101110011;
assign LUT_2[2016] = 32'b00000000000000001100010100111000;
assign LUT_2[2017] = 32'b00000000000000001001001101010001;
assign LUT_2[2018] = 32'b00000000000000010011001101110100;
assign LUT_2[2019] = 32'b00000000000000010000000110001101;
assign LUT_2[2020] = 32'b00000000000000001000110010100000;
assign LUT_2[2021] = 32'b00000000000000000101101010111001;
assign LUT_2[2022] = 32'b00000000000000001111101011011100;
assign LUT_2[2023] = 32'b00000000000000001100100011110101;
assign LUT_2[2024] = 32'b00000000000000000111000110010101;
assign LUT_2[2025] = 32'b00000000000000000011111110101110;
assign LUT_2[2026] = 32'b00000000000000001101111111010001;
assign LUT_2[2027] = 32'b00000000000000001010110111101010;
assign LUT_2[2028] = 32'b00000000000000000011100011111101;
assign LUT_2[2029] = 32'b00000000000000000000011100010110;
assign LUT_2[2030] = 32'b00000000000000001010011100111001;
assign LUT_2[2031] = 32'b00000000000000000111010101010010;
assign LUT_2[2032] = 32'b00000000000000000110111001000010;
assign LUT_2[2033] = 32'b00000000000000000011110001011011;
assign LUT_2[2034] = 32'b00000000000000001101110001111110;
assign LUT_2[2035] = 32'b00000000000000001010101010010111;
assign LUT_2[2036] = 32'b00000000000000000011010110101010;
assign LUT_2[2037] = 32'b00000000000000000000001111000011;
assign LUT_2[2038] = 32'b00000000000000001010001111100110;
assign LUT_2[2039] = 32'b00000000000000000111000111111111;
assign LUT_2[2040] = 32'b00000000000000000001101010011111;
assign LUT_2[2041] = 32'b11111111111111111110100010111000;
assign LUT_2[2042] = 32'b00000000000000001000100011011011;
assign LUT_2[2043] = 32'b00000000000000000101011011110100;
assign LUT_2[2044] = 32'b11111111111111111110001000000111;
assign LUT_2[2045] = 32'b11111111111111111011000000100000;
assign LUT_2[2046] = 32'b00000000000000000101000001000011;
assign LUT_2[2047] = 32'b00000000000000000001111001011100;
assign LUT_2[2048] = 32'b11111111111111111011110101111100;
assign LUT_2[2049] = 32'b11111111111111111000101110010101;
assign LUT_2[2050] = 32'b00000000000000000010101110111000;
assign LUT_2[2051] = 32'b11111111111111111111100111010001;
assign LUT_2[2052] = 32'b11111111111111111000010011100100;
assign LUT_2[2053] = 32'b11111111111111110101001011111101;
assign LUT_2[2054] = 32'b11111111111111111111001100100000;
assign LUT_2[2055] = 32'b11111111111111111100000100111001;
assign LUT_2[2056] = 32'b11111111111111110110100111011001;
assign LUT_2[2057] = 32'b11111111111111110011011111110010;
assign LUT_2[2058] = 32'b11111111111111111101100000010101;
assign LUT_2[2059] = 32'b11111111111111111010011000101110;
assign LUT_2[2060] = 32'b11111111111111110011000101000001;
assign LUT_2[2061] = 32'b11111111111111101111111101011010;
assign LUT_2[2062] = 32'b11111111111111111001111101111101;
assign LUT_2[2063] = 32'b11111111111111110110110110010110;
assign LUT_2[2064] = 32'b11111111111111110110011010000110;
assign LUT_2[2065] = 32'b11111111111111110011010010011111;
assign LUT_2[2066] = 32'b11111111111111111101010011000010;
assign LUT_2[2067] = 32'b11111111111111111010001011011011;
assign LUT_2[2068] = 32'b11111111111111110010110111101110;
assign LUT_2[2069] = 32'b11111111111111101111110000000111;
assign LUT_2[2070] = 32'b11111111111111111001110000101010;
assign LUT_2[2071] = 32'b11111111111111110110101001000011;
assign LUT_2[2072] = 32'b11111111111111110001001011100011;
assign LUT_2[2073] = 32'b11111111111111101110000011111100;
assign LUT_2[2074] = 32'b11111111111111111000000100011111;
assign LUT_2[2075] = 32'b11111111111111110100111100111000;
assign LUT_2[2076] = 32'b11111111111111101101101001001011;
assign LUT_2[2077] = 32'b11111111111111101010100001100100;
assign LUT_2[2078] = 32'b11111111111111110100100010000111;
assign LUT_2[2079] = 32'b11111111111111110001011010100000;
assign LUT_2[2080] = 32'b11111111111111111100010001100101;
assign LUT_2[2081] = 32'b11111111111111111001001001111110;
assign LUT_2[2082] = 32'b00000000000000000011001010100001;
assign LUT_2[2083] = 32'b00000000000000000000000010111010;
assign LUT_2[2084] = 32'b11111111111111111000101111001101;
assign LUT_2[2085] = 32'b11111111111111110101100111100110;
assign LUT_2[2086] = 32'b11111111111111111111101000001001;
assign LUT_2[2087] = 32'b11111111111111111100100000100010;
assign LUT_2[2088] = 32'b11111111111111110111000011000010;
assign LUT_2[2089] = 32'b11111111111111110011111011011011;
assign LUT_2[2090] = 32'b11111111111111111101111011111110;
assign LUT_2[2091] = 32'b11111111111111111010110100010111;
assign LUT_2[2092] = 32'b11111111111111110011100000101010;
assign LUT_2[2093] = 32'b11111111111111110000011001000011;
assign LUT_2[2094] = 32'b11111111111111111010011001100110;
assign LUT_2[2095] = 32'b11111111111111110111010001111111;
assign LUT_2[2096] = 32'b11111111111111110110110101101111;
assign LUT_2[2097] = 32'b11111111111111110011101110001000;
assign LUT_2[2098] = 32'b11111111111111111101101110101011;
assign LUT_2[2099] = 32'b11111111111111111010100111000100;
assign LUT_2[2100] = 32'b11111111111111110011010011010111;
assign LUT_2[2101] = 32'b11111111111111110000001011110000;
assign LUT_2[2102] = 32'b11111111111111111010001100010011;
assign LUT_2[2103] = 32'b11111111111111110111000100101100;
assign LUT_2[2104] = 32'b11111111111111110001100111001100;
assign LUT_2[2105] = 32'b11111111111111101110011111100101;
assign LUT_2[2106] = 32'b11111111111111111000100000001000;
assign LUT_2[2107] = 32'b11111111111111110101011000100001;
assign LUT_2[2108] = 32'b11111111111111101110000100110100;
assign LUT_2[2109] = 32'b11111111111111101010111101001101;
assign LUT_2[2110] = 32'b11111111111111110100111101110000;
assign LUT_2[2111] = 32'b11111111111111110001110110001001;
assign LUT_2[2112] = 32'b11111111111111110011111110011111;
assign LUT_2[2113] = 32'b11111111111111110000110110111000;
assign LUT_2[2114] = 32'b11111111111111111010110111011011;
assign LUT_2[2115] = 32'b11111111111111110111101111110100;
assign LUT_2[2116] = 32'b11111111111111110000011100000111;
assign LUT_2[2117] = 32'b11111111111111101101010100100000;
assign LUT_2[2118] = 32'b11111111111111110111010101000011;
assign LUT_2[2119] = 32'b11111111111111110100001101011100;
assign LUT_2[2120] = 32'b11111111111111101110101111111100;
assign LUT_2[2121] = 32'b11111111111111101011101000010101;
assign LUT_2[2122] = 32'b11111111111111110101101000111000;
assign LUT_2[2123] = 32'b11111111111111110010100001010001;
assign LUT_2[2124] = 32'b11111111111111101011001101100100;
assign LUT_2[2125] = 32'b11111111111111101000000101111101;
assign LUT_2[2126] = 32'b11111111111111110010000110100000;
assign LUT_2[2127] = 32'b11111111111111101110111110111001;
assign LUT_2[2128] = 32'b11111111111111101110100010101001;
assign LUT_2[2129] = 32'b11111111111111101011011011000010;
assign LUT_2[2130] = 32'b11111111111111110101011011100101;
assign LUT_2[2131] = 32'b11111111111111110010010011111110;
assign LUT_2[2132] = 32'b11111111111111101011000000010001;
assign LUT_2[2133] = 32'b11111111111111100111111000101010;
assign LUT_2[2134] = 32'b11111111111111110001111001001101;
assign LUT_2[2135] = 32'b11111111111111101110110001100110;
assign LUT_2[2136] = 32'b11111111111111101001010100000110;
assign LUT_2[2137] = 32'b11111111111111100110001100011111;
assign LUT_2[2138] = 32'b11111111111111110000001101000010;
assign LUT_2[2139] = 32'b11111111111111101101000101011011;
assign LUT_2[2140] = 32'b11111111111111100101110001101110;
assign LUT_2[2141] = 32'b11111111111111100010101010000111;
assign LUT_2[2142] = 32'b11111111111111101100101010101010;
assign LUT_2[2143] = 32'b11111111111111101001100011000011;
assign LUT_2[2144] = 32'b11111111111111110100011010001000;
assign LUT_2[2145] = 32'b11111111111111110001010010100001;
assign LUT_2[2146] = 32'b11111111111111111011010011000100;
assign LUT_2[2147] = 32'b11111111111111111000001011011101;
assign LUT_2[2148] = 32'b11111111111111110000110111110000;
assign LUT_2[2149] = 32'b11111111111111101101110000001001;
assign LUT_2[2150] = 32'b11111111111111110111110000101100;
assign LUT_2[2151] = 32'b11111111111111110100101001000101;
assign LUT_2[2152] = 32'b11111111111111101111001011100101;
assign LUT_2[2153] = 32'b11111111111111101100000011111110;
assign LUT_2[2154] = 32'b11111111111111110110000100100001;
assign LUT_2[2155] = 32'b11111111111111110010111100111010;
assign LUT_2[2156] = 32'b11111111111111101011101001001101;
assign LUT_2[2157] = 32'b11111111111111101000100001100110;
assign LUT_2[2158] = 32'b11111111111111110010100010001001;
assign LUT_2[2159] = 32'b11111111111111101111011010100010;
assign LUT_2[2160] = 32'b11111111111111101110111110010010;
assign LUT_2[2161] = 32'b11111111111111101011110110101011;
assign LUT_2[2162] = 32'b11111111111111110101110111001110;
assign LUT_2[2163] = 32'b11111111111111110010101111100111;
assign LUT_2[2164] = 32'b11111111111111101011011011111010;
assign LUT_2[2165] = 32'b11111111111111101000010100010011;
assign LUT_2[2166] = 32'b11111111111111110010010100110110;
assign LUT_2[2167] = 32'b11111111111111101111001101001111;
assign LUT_2[2168] = 32'b11111111111111101001101111101111;
assign LUT_2[2169] = 32'b11111111111111100110101000001000;
assign LUT_2[2170] = 32'b11111111111111110000101000101011;
assign LUT_2[2171] = 32'b11111111111111101101100001000100;
assign LUT_2[2172] = 32'b11111111111111100110001101010111;
assign LUT_2[2173] = 32'b11111111111111100011000101110000;
assign LUT_2[2174] = 32'b11111111111111101101000110010011;
assign LUT_2[2175] = 32'b11111111111111101001111110101100;
assign LUT_2[2176] = 32'b00000000000000000000001010001011;
assign LUT_2[2177] = 32'b11111111111111111101000010100100;
assign LUT_2[2178] = 32'b00000000000000000111000011000111;
assign LUT_2[2179] = 32'b00000000000000000011111011100000;
assign LUT_2[2180] = 32'b11111111111111111100100111110011;
assign LUT_2[2181] = 32'b11111111111111111001100000001100;
assign LUT_2[2182] = 32'b00000000000000000011100000101111;
assign LUT_2[2183] = 32'b00000000000000000000011001001000;
assign LUT_2[2184] = 32'b11111111111111111010111011101000;
assign LUT_2[2185] = 32'b11111111111111110111110100000001;
assign LUT_2[2186] = 32'b00000000000000000001110100100100;
assign LUT_2[2187] = 32'b11111111111111111110101100111101;
assign LUT_2[2188] = 32'b11111111111111110111011001010000;
assign LUT_2[2189] = 32'b11111111111111110100010001101001;
assign LUT_2[2190] = 32'b11111111111111111110010010001100;
assign LUT_2[2191] = 32'b11111111111111111011001010100101;
assign LUT_2[2192] = 32'b11111111111111111010101110010101;
assign LUT_2[2193] = 32'b11111111111111110111100110101110;
assign LUT_2[2194] = 32'b00000000000000000001100111010001;
assign LUT_2[2195] = 32'b11111111111111111110011111101010;
assign LUT_2[2196] = 32'b11111111111111110111001011111101;
assign LUT_2[2197] = 32'b11111111111111110100000100010110;
assign LUT_2[2198] = 32'b11111111111111111110000100111001;
assign LUT_2[2199] = 32'b11111111111111111010111101010010;
assign LUT_2[2200] = 32'b11111111111111110101011111110010;
assign LUT_2[2201] = 32'b11111111111111110010011000001011;
assign LUT_2[2202] = 32'b11111111111111111100011000101110;
assign LUT_2[2203] = 32'b11111111111111111001010001000111;
assign LUT_2[2204] = 32'b11111111111111110001111101011010;
assign LUT_2[2205] = 32'b11111111111111101110110101110011;
assign LUT_2[2206] = 32'b11111111111111111000110110010110;
assign LUT_2[2207] = 32'b11111111111111110101101110101111;
assign LUT_2[2208] = 32'b00000000000000000000100101110100;
assign LUT_2[2209] = 32'b11111111111111111101011110001101;
assign LUT_2[2210] = 32'b00000000000000000111011110110000;
assign LUT_2[2211] = 32'b00000000000000000100010111001001;
assign LUT_2[2212] = 32'b11111111111111111101000011011100;
assign LUT_2[2213] = 32'b11111111111111111001111011110101;
assign LUT_2[2214] = 32'b00000000000000000011111100011000;
assign LUT_2[2215] = 32'b00000000000000000000110100110001;
assign LUT_2[2216] = 32'b11111111111111111011010111010001;
assign LUT_2[2217] = 32'b11111111111111111000001111101010;
assign LUT_2[2218] = 32'b00000000000000000010010000001101;
assign LUT_2[2219] = 32'b11111111111111111111001000100110;
assign LUT_2[2220] = 32'b11111111111111110111110100111001;
assign LUT_2[2221] = 32'b11111111111111110100101101010010;
assign LUT_2[2222] = 32'b11111111111111111110101101110101;
assign LUT_2[2223] = 32'b11111111111111111011100110001110;
assign LUT_2[2224] = 32'b11111111111111111011001001111110;
assign LUT_2[2225] = 32'b11111111111111111000000010010111;
assign LUT_2[2226] = 32'b00000000000000000010000010111010;
assign LUT_2[2227] = 32'b11111111111111111110111011010011;
assign LUT_2[2228] = 32'b11111111111111110111100111100110;
assign LUT_2[2229] = 32'b11111111111111110100011111111111;
assign LUT_2[2230] = 32'b11111111111111111110100000100010;
assign LUT_2[2231] = 32'b11111111111111111011011000111011;
assign LUT_2[2232] = 32'b11111111111111110101111011011011;
assign LUT_2[2233] = 32'b11111111111111110010110011110100;
assign LUT_2[2234] = 32'b11111111111111111100110100010111;
assign LUT_2[2235] = 32'b11111111111111111001101100110000;
assign LUT_2[2236] = 32'b11111111111111110010011001000011;
assign LUT_2[2237] = 32'b11111111111111101111010001011100;
assign LUT_2[2238] = 32'b11111111111111111001010001111111;
assign LUT_2[2239] = 32'b11111111111111110110001010011000;
assign LUT_2[2240] = 32'b11111111111111111000010010101110;
assign LUT_2[2241] = 32'b11111111111111110101001011000111;
assign LUT_2[2242] = 32'b11111111111111111111001011101010;
assign LUT_2[2243] = 32'b11111111111111111100000100000011;
assign LUT_2[2244] = 32'b11111111111111110100110000010110;
assign LUT_2[2245] = 32'b11111111111111110001101000101111;
assign LUT_2[2246] = 32'b11111111111111111011101001010010;
assign LUT_2[2247] = 32'b11111111111111111000100001101011;
assign LUT_2[2248] = 32'b11111111111111110011000100001011;
assign LUT_2[2249] = 32'b11111111111111101111111100100100;
assign LUT_2[2250] = 32'b11111111111111111001111101000111;
assign LUT_2[2251] = 32'b11111111111111110110110101100000;
assign LUT_2[2252] = 32'b11111111111111101111100001110011;
assign LUT_2[2253] = 32'b11111111111111101100011010001100;
assign LUT_2[2254] = 32'b11111111111111110110011010101111;
assign LUT_2[2255] = 32'b11111111111111110011010011001000;
assign LUT_2[2256] = 32'b11111111111111110010110110111000;
assign LUT_2[2257] = 32'b11111111111111101111101111010001;
assign LUT_2[2258] = 32'b11111111111111111001101111110100;
assign LUT_2[2259] = 32'b11111111111111110110101000001101;
assign LUT_2[2260] = 32'b11111111111111101111010100100000;
assign LUT_2[2261] = 32'b11111111111111101100001100111001;
assign LUT_2[2262] = 32'b11111111111111110110001101011100;
assign LUT_2[2263] = 32'b11111111111111110011000101110101;
assign LUT_2[2264] = 32'b11111111111111101101101000010101;
assign LUT_2[2265] = 32'b11111111111111101010100000101110;
assign LUT_2[2266] = 32'b11111111111111110100100001010001;
assign LUT_2[2267] = 32'b11111111111111110001011001101010;
assign LUT_2[2268] = 32'b11111111111111101010000101111101;
assign LUT_2[2269] = 32'b11111111111111100110111110010110;
assign LUT_2[2270] = 32'b11111111111111110000111110111001;
assign LUT_2[2271] = 32'b11111111111111101101110111010010;
assign LUT_2[2272] = 32'b11111111111111111000101110010111;
assign LUT_2[2273] = 32'b11111111111111110101100110110000;
assign LUT_2[2274] = 32'b11111111111111111111100111010011;
assign LUT_2[2275] = 32'b11111111111111111100011111101100;
assign LUT_2[2276] = 32'b11111111111111110101001011111111;
assign LUT_2[2277] = 32'b11111111111111110010000100011000;
assign LUT_2[2278] = 32'b11111111111111111100000100111011;
assign LUT_2[2279] = 32'b11111111111111111000111101010100;
assign LUT_2[2280] = 32'b11111111111111110011011111110100;
assign LUT_2[2281] = 32'b11111111111111110000011000001101;
assign LUT_2[2282] = 32'b11111111111111111010011000110000;
assign LUT_2[2283] = 32'b11111111111111110111010001001001;
assign LUT_2[2284] = 32'b11111111111111101111111101011100;
assign LUT_2[2285] = 32'b11111111111111101100110101110101;
assign LUT_2[2286] = 32'b11111111111111110110110110011000;
assign LUT_2[2287] = 32'b11111111111111110011101110110001;
assign LUT_2[2288] = 32'b11111111111111110011010010100001;
assign LUT_2[2289] = 32'b11111111111111110000001010111010;
assign LUT_2[2290] = 32'b11111111111111111010001011011101;
assign LUT_2[2291] = 32'b11111111111111110111000011110110;
assign LUT_2[2292] = 32'b11111111111111101111110000001001;
assign LUT_2[2293] = 32'b11111111111111101100101000100010;
assign LUT_2[2294] = 32'b11111111111111110110101001000101;
assign LUT_2[2295] = 32'b11111111111111110011100001011110;
assign LUT_2[2296] = 32'b11111111111111101110000011111110;
assign LUT_2[2297] = 32'b11111111111111101010111100010111;
assign LUT_2[2298] = 32'b11111111111111110100111100111010;
assign LUT_2[2299] = 32'b11111111111111110001110101010011;
assign LUT_2[2300] = 32'b11111111111111101010100001100110;
assign LUT_2[2301] = 32'b11111111111111100111011001111111;
assign LUT_2[2302] = 32'b11111111111111110001011010100010;
assign LUT_2[2303] = 32'b11111111111111101110010010111011;
assign LUT_2[2304] = 32'b11111111111111111111110100100010;
assign LUT_2[2305] = 32'b11111111111111111100101100111011;
assign LUT_2[2306] = 32'b00000000000000000110101101011110;
assign LUT_2[2307] = 32'b00000000000000000011100101110111;
assign LUT_2[2308] = 32'b11111111111111111100010010001010;
assign LUT_2[2309] = 32'b11111111111111111001001010100011;
assign LUT_2[2310] = 32'b00000000000000000011001011000110;
assign LUT_2[2311] = 32'b00000000000000000000000011011111;
assign LUT_2[2312] = 32'b11111111111111111010100101111111;
assign LUT_2[2313] = 32'b11111111111111110111011110011000;
assign LUT_2[2314] = 32'b00000000000000000001011110111011;
assign LUT_2[2315] = 32'b11111111111111111110010111010100;
assign LUT_2[2316] = 32'b11111111111111110111000011100111;
assign LUT_2[2317] = 32'b11111111111111110011111100000000;
assign LUT_2[2318] = 32'b11111111111111111101111100100011;
assign LUT_2[2319] = 32'b11111111111111111010110100111100;
assign LUT_2[2320] = 32'b11111111111111111010011000101100;
assign LUT_2[2321] = 32'b11111111111111110111010001000101;
assign LUT_2[2322] = 32'b00000000000000000001010001101000;
assign LUT_2[2323] = 32'b11111111111111111110001010000001;
assign LUT_2[2324] = 32'b11111111111111110110110110010100;
assign LUT_2[2325] = 32'b11111111111111110011101110101101;
assign LUT_2[2326] = 32'b11111111111111111101101111010000;
assign LUT_2[2327] = 32'b11111111111111111010100111101001;
assign LUT_2[2328] = 32'b11111111111111110101001010001001;
assign LUT_2[2329] = 32'b11111111111111110010000010100010;
assign LUT_2[2330] = 32'b11111111111111111100000011000101;
assign LUT_2[2331] = 32'b11111111111111111000111011011110;
assign LUT_2[2332] = 32'b11111111111111110001100111110001;
assign LUT_2[2333] = 32'b11111111111111101110100000001010;
assign LUT_2[2334] = 32'b11111111111111111000100000101101;
assign LUT_2[2335] = 32'b11111111111111110101011001000110;
assign LUT_2[2336] = 32'b00000000000000000000010000001011;
assign LUT_2[2337] = 32'b11111111111111111101001000100100;
assign LUT_2[2338] = 32'b00000000000000000111001001000111;
assign LUT_2[2339] = 32'b00000000000000000100000001100000;
assign LUT_2[2340] = 32'b11111111111111111100101101110011;
assign LUT_2[2341] = 32'b11111111111111111001100110001100;
assign LUT_2[2342] = 32'b00000000000000000011100110101111;
assign LUT_2[2343] = 32'b00000000000000000000011111001000;
assign LUT_2[2344] = 32'b11111111111111111011000001101000;
assign LUT_2[2345] = 32'b11111111111111110111111010000001;
assign LUT_2[2346] = 32'b00000000000000000001111010100100;
assign LUT_2[2347] = 32'b11111111111111111110110010111101;
assign LUT_2[2348] = 32'b11111111111111110111011111010000;
assign LUT_2[2349] = 32'b11111111111111110100010111101001;
assign LUT_2[2350] = 32'b11111111111111111110011000001100;
assign LUT_2[2351] = 32'b11111111111111111011010000100101;
assign LUT_2[2352] = 32'b11111111111111111010110100010101;
assign LUT_2[2353] = 32'b11111111111111110111101100101110;
assign LUT_2[2354] = 32'b00000000000000000001101101010001;
assign LUT_2[2355] = 32'b11111111111111111110100101101010;
assign LUT_2[2356] = 32'b11111111111111110111010001111101;
assign LUT_2[2357] = 32'b11111111111111110100001010010110;
assign LUT_2[2358] = 32'b11111111111111111110001010111001;
assign LUT_2[2359] = 32'b11111111111111111011000011010010;
assign LUT_2[2360] = 32'b11111111111111110101100101110010;
assign LUT_2[2361] = 32'b11111111111111110010011110001011;
assign LUT_2[2362] = 32'b11111111111111111100011110101110;
assign LUT_2[2363] = 32'b11111111111111111001010111000111;
assign LUT_2[2364] = 32'b11111111111111110010000011011010;
assign LUT_2[2365] = 32'b11111111111111101110111011110011;
assign LUT_2[2366] = 32'b11111111111111111000111100010110;
assign LUT_2[2367] = 32'b11111111111111110101110100101111;
assign LUT_2[2368] = 32'b11111111111111110111111101000101;
assign LUT_2[2369] = 32'b11111111111111110100110101011110;
assign LUT_2[2370] = 32'b11111111111111111110110110000001;
assign LUT_2[2371] = 32'b11111111111111111011101110011010;
assign LUT_2[2372] = 32'b11111111111111110100011010101101;
assign LUT_2[2373] = 32'b11111111111111110001010011000110;
assign LUT_2[2374] = 32'b11111111111111111011010011101001;
assign LUT_2[2375] = 32'b11111111111111111000001100000010;
assign LUT_2[2376] = 32'b11111111111111110010101110100010;
assign LUT_2[2377] = 32'b11111111111111101111100110111011;
assign LUT_2[2378] = 32'b11111111111111111001100111011110;
assign LUT_2[2379] = 32'b11111111111111110110011111110111;
assign LUT_2[2380] = 32'b11111111111111101111001100001010;
assign LUT_2[2381] = 32'b11111111111111101100000100100011;
assign LUT_2[2382] = 32'b11111111111111110110000101000110;
assign LUT_2[2383] = 32'b11111111111111110010111101011111;
assign LUT_2[2384] = 32'b11111111111111110010100001001111;
assign LUT_2[2385] = 32'b11111111111111101111011001101000;
assign LUT_2[2386] = 32'b11111111111111111001011010001011;
assign LUT_2[2387] = 32'b11111111111111110110010010100100;
assign LUT_2[2388] = 32'b11111111111111101110111110110111;
assign LUT_2[2389] = 32'b11111111111111101011110111010000;
assign LUT_2[2390] = 32'b11111111111111110101110111110011;
assign LUT_2[2391] = 32'b11111111111111110010110000001100;
assign LUT_2[2392] = 32'b11111111111111101101010010101100;
assign LUT_2[2393] = 32'b11111111111111101010001011000101;
assign LUT_2[2394] = 32'b11111111111111110100001011101000;
assign LUT_2[2395] = 32'b11111111111111110001000100000001;
assign LUT_2[2396] = 32'b11111111111111101001110000010100;
assign LUT_2[2397] = 32'b11111111111111100110101000101101;
assign LUT_2[2398] = 32'b11111111111111110000101001010000;
assign LUT_2[2399] = 32'b11111111111111101101100001101001;
assign LUT_2[2400] = 32'b11111111111111111000011000101110;
assign LUT_2[2401] = 32'b11111111111111110101010001000111;
assign LUT_2[2402] = 32'b11111111111111111111010001101010;
assign LUT_2[2403] = 32'b11111111111111111100001010000011;
assign LUT_2[2404] = 32'b11111111111111110100110110010110;
assign LUT_2[2405] = 32'b11111111111111110001101110101111;
assign LUT_2[2406] = 32'b11111111111111111011101111010010;
assign LUT_2[2407] = 32'b11111111111111111000100111101011;
assign LUT_2[2408] = 32'b11111111111111110011001010001011;
assign LUT_2[2409] = 32'b11111111111111110000000010100100;
assign LUT_2[2410] = 32'b11111111111111111010000011000111;
assign LUT_2[2411] = 32'b11111111111111110110111011100000;
assign LUT_2[2412] = 32'b11111111111111101111100111110011;
assign LUT_2[2413] = 32'b11111111111111101100100000001100;
assign LUT_2[2414] = 32'b11111111111111110110100000101111;
assign LUT_2[2415] = 32'b11111111111111110011011001001000;
assign LUT_2[2416] = 32'b11111111111111110010111100111000;
assign LUT_2[2417] = 32'b11111111111111101111110101010001;
assign LUT_2[2418] = 32'b11111111111111111001110101110100;
assign LUT_2[2419] = 32'b11111111111111110110101110001101;
assign LUT_2[2420] = 32'b11111111111111101111011010100000;
assign LUT_2[2421] = 32'b11111111111111101100010010111001;
assign LUT_2[2422] = 32'b11111111111111110110010011011100;
assign LUT_2[2423] = 32'b11111111111111110011001011110101;
assign LUT_2[2424] = 32'b11111111111111101101101110010101;
assign LUT_2[2425] = 32'b11111111111111101010100110101110;
assign LUT_2[2426] = 32'b11111111111111110100100111010001;
assign LUT_2[2427] = 32'b11111111111111110001011111101010;
assign LUT_2[2428] = 32'b11111111111111101010001011111101;
assign LUT_2[2429] = 32'b11111111111111100111000100010110;
assign LUT_2[2430] = 32'b11111111111111110001000100111001;
assign LUT_2[2431] = 32'b11111111111111101101111101010010;
assign LUT_2[2432] = 32'b00000000000000000100001000110001;
assign LUT_2[2433] = 32'b00000000000000000001000001001010;
assign LUT_2[2434] = 32'b00000000000000001011000001101101;
assign LUT_2[2435] = 32'b00000000000000000111111010000110;
assign LUT_2[2436] = 32'b00000000000000000000100110011001;
assign LUT_2[2437] = 32'b11111111111111111101011110110010;
assign LUT_2[2438] = 32'b00000000000000000111011111010101;
assign LUT_2[2439] = 32'b00000000000000000100010111101110;
assign LUT_2[2440] = 32'b11111111111111111110111010001110;
assign LUT_2[2441] = 32'b11111111111111111011110010100111;
assign LUT_2[2442] = 32'b00000000000000000101110011001010;
assign LUT_2[2443] = 32'b00000000000000000010101011100011;
assign LUT_2[2444] = 32'b11111111111111111011010111110110;
assign LUT_2[2445] = 32'b11111111111111111000010000001111;
assign LUT_2[2446] = 32'b00000000000000000010010000110010;
assign LUT_2[2447] = 32'b11111111111111111111001001001011;
assign LUT_2[2448] = 32'b11111111111111111110101100111011;
assign LUT_2[2449] = 32'b11111111111111111011100101010100;
assign LUT_2[2450] = 32'b00000000000000000101100101110111;
assign LUT_2[2451] = 32'b00000000000000000010011110010000;
assign LUT_2[2452] = 32'b11111111111111111011001010100011;
assign LUT_2[2453] = 32'b11111111111111111000000010111100;
assign LUT_2[2454] = 32'b00000000000000000010000011011111;
assign LUT_2[2455] = 32'b11111111111111111110111011111000;
assign LUT_2[2456] = 32'b11111111111111111001011110011000;
assign LUT_2[2457] = 32'b11111111111111110110010110110001;
assign LUT_2[2458] = 32'b00000000000000000000010111010100;
assign LUT_2[2459] = 32'b11111111111111111101001111101101;
assign LUT_2[2460] = 32'b11111111111111110101111100000000;
assign LUT_2[2461] = 32'b11111111111111110010110100011001;
assign LUT_2[2462] = 32'b11111111111111111100110100111100;
assign LUT_2[2463] = 32'b11111111111111111001101101010101;
assign LUT_2[2464] = 32'b00000000000000000100100100011010;
assign LUT_2[2465] = 32'b00000000000000000001011100110011;
assign LUT_2[2466] = 32'b00000000000000001011011101010110;
assign LUT_2[2467] = 32'b00000000000000001000010101101111;
assign LUT_2[2468] = 32'b00000000000000000001000010000010;
assign LUT_2[2469] = 32'b11111111111111111101111010011011;
assign LUT_2[2470] = 32'b00000000000000000111111010111110;
assign LUT_2[2471] = 32'b00000000000000000100110011010111;
assign LUT_2[2472] = 32'b11111111111111111111010101110111;
assign LUT_2[2473] = 32'b11111111111111111100001110010000;
assign LUT_2[2474] = 32'b00000000000000000110001110110011;
assign LUT_2[2475] = 32'b00000000000000000011000111001100;
assign LUT_2[2476] = 32'b11111111111111111011110011011111;
assign LUT_2[2477] = 32'b11111111111111111000101011111000;
assign LUT_2[2478] = 32'b00000000000000000010101100011011;
assign LUT_2[2479] = 32'b11111111111111111111100100110100;
assign LUT_2[2480] = 32'b11111111111111111111001000100100;
assign LUT_2[2481] = 32'b11111111111111111100000000111101;
assign LUT_2[2482] = 32'b00000000000000000110000001100000;
assign LUT_2[2483] = 32'b00000000000000000010111001111001;
assign LUT_2[2484] = 32'b11111111111111111011100110001100;
assign LUT_2[2485] = 32'b11111111111111111000011110100101;
assign LUT_2[2486] = 32'b00000000000000000010011111001000;
assign LUT_2[2487] = 32'b11111111111111111111010111100001;
assign LUT_2[2488] = 32'b11111111111111111001111010000001;
assign LUT_2[2489] = 32'b11111111111111110110110010011010;
assign LUT_2[2490] = 32'b00000000000000000000110010111101;
assign LUT_2[2491] = 32'b11111111111111111101101011010110;
assign LUT_2[2492] = 32'b11111111111111110110010111101001;
assign LUT_2[2493] = 32'b11111111111111110011010000000010;
assign LUT_2[2494] = 32'b11111111111111111101010000100101;
assign LUT_2[2495] = 32'b11111111111111111010001000111110;
assign LUT_2[2496] = 32'b11111111111111111100010001010100;
assign LUT_2[2497] = 32'b11111111111111111001001001101101;
assign LUT_2[2498] = 32'b00000000000000000011001010010000;
assign LUT_2[2499] = 32'b00000000000000000000000010101001;
assign LUT_2[2500] = 32'b11111111111111111000101110111100;
assign LUT_2[2501] = 32'b11111111111111110101100111010101;
assign LUT_2[2502] = 32'b11111111111111111111100111111000;
assign LUT_2[2503] = 32'b11111111111111111100100000010001;
assign LUT_2[2504] = 32'b11111111111111110111000010110001;
assign LUT_2[2505] = 32'b11111111111111110011111011001010;
assign LUT_2[2506] = 32'b11111111111111111101111011101101;
assign LUT_2[2507] = 32'b11111111111111111010110100000110;
assign LUT_2[2508] = 32'b11111111111111110011100000011001;
assign LUT_2[2509] = 32'b11111111111111110000011000110010;
assign LUT_2[2510] = 32'b11111111111111111010011001010101;
assign LUT_2[2511] = 32'b11111111111111110111010001101110;
assign LUT_2[2512] = 32'b11111111111111110110110101011110;
assign LUT_2[2513] = 32'b11111111111111110011101101110111;
assign LUT_2[2514] = 32'b11111111111111111101101110011010;
assign LUT_2[2515] = 32'b11111111111111111010100110110011;
assign LUT_2[2516] = 32'b11111111111111110011010011000110;
assign LUT_2[2517] = 32'b11111111111111110000001011011111;
assign LUT_2[2518] = 32'b11111111111111111010001100000010;
assign LUT_2[2519] = 32'b11111111111111110111000100011011;
assign LUT_2[2520] = 32'b11111111111111110001100110111011;
assign LUT_2[2521] = 32'b11111111111111101110011111010100;
assign LUT_2[2522] = 32'b11111111111111111000011111110111;
assign LUT_2[2523] = 32'b11111111111111110101011000010000;
assign LUT_2[2524] = 32'b11111111111111101110000100100011;
assign LUT_2[2525] = 32'b11111111111111101010111100111100;
assign LUT_2[2526] = 32'b11111111111111110100111101011111;
assign LUT_2[2527] = 32'b11111111111111110001110101111000;
assign LUT_2[2528] = 32'b11111111111111111100101100111101;
assign LUT_2[2529] = 32'b11111111111111111001100101010110;
assign LUT_2[2530] = 32'b00000000000000000011100101111001;
assign LUT_2[2531] = 32'b00000000000000000000011110010010;
assign LUT_2[2532] = 32'b11111111111111111001001010100101;
assign LUT_2[2533] = 32'b11111111111111110110000010111110;
assign LUT_2[2534] = 32'b00000000000000000000000011100001;
assign LUT_2[2535] = 32'b11111111111111111100111011111010;
assign LUT_2[2536] = 32'b11111111111111110111011110011010;
assign LUT_2[2537] = 32'b11111111111111110100010110110011;
assign LUT_2[2538] = 32'b11111111111111111110010111010110;
assign LUT_2[2539] = 32'b11111111111111111011001111101111;
assign LUT_2[2540] = 32'b11111111111111110011111100000010;
assign LUT_2[2541] = 32'b11111111111111110000110100011011;
assign LUT_2[2542] = 32'b11111111111111111010110100111110;
assign LUT_2[2543] = 32'b11111111111111110111101101010111;
assign LUT_2[2544] = 32'b11111111111111110111010001000111;
assign LUT_2[2545] = 32'b11111111111111110100001001100000;
assign LUT_2[2546] = 32'b11111111111111111110001010000011;
assign LUT_2[2547] = 32'b11111111111111111011000010011100;
assign LUT_2[2548] = 32'b11111111111111110011101110101111;
assign LUT_2[2549] = 32'b11111111111111110000100111001000;
assign LUT_2[2550] = 32'b11111111111111111010100111101011;
assign LUT_2[2551] = 32'b11111111111111110111100000000100;
assign LUT_2[2552] = 32'b11111111111111110010000010100100;
assign LUT_2[2553] = 32'b11111111111111101110111010111101;
assign LUT_2[2554] = 32'b11111111111111111000111011100000;
assign LUT_2[2555] = 32'b11111111111111110101110011111001;
assign LUT_2[2556] = 32'b11111111111111101110100000001100;
assign LUT_2[2557] = 32'b11111111111111101011011000100101;
assign LUT_2[2558] = 32'b11111111111111110101011001001000;
assign LUT_2[2559] = 32'b11111111111111110010010001100001;
assign LUT_2[2560] = 32'b00000000000000000000100111101110;
assign LUT_2[2561] = 32'b11111111111111111101100000000111;
assign LUT_2[2562] = 32'b00000000000000000111100000101010;
assign LUT_2[2563] = 32'b00000000000000000100011001000011;
assign LUT_2[2564] = 32'b11111111111111111101000101010110;
assign LUT_2[2565] = 32'b11111111111111111001111101101111;
assign LUT_2[2566] = 32'b00000000000000000011111110010010;
assign LUT_2[2567] = 32'b00000000000000000000110110101011;
assign LUT_2[2568] = 32'b11111111111111111011011001001011;
assign LUT_2[2569] = 32'b11111111111111111000010001100100;
assign LUT_2[2570] = 32'b00000000000000000010010010000111;
assign LUT_2[2571] = 32'b11111111111111111111001010100000;
assign LUT_2[2572] = 32'b11111111111111110111110110110011;
assign LUT_2[2573] = 32'b11111111111111110100101111001100;
assign LUT_2[2574] = 32'b11111111111111111110101111101111;
assign LUT_2[2575] = 32'b11111111111111111011101000001000;
assign LUT_2[2576] = 32'b11111111111111111011001011111000;
assign LUT_2[2577] = 32'b11111111111111111000000100010001;
assign LUT_2[2578] = 32'b00000000000000000010000100110100;
assign LUT_2[2579] = 32'b11111111111111111110111101001101;
assign LUT_2[2580] = 32'b11111111111111110111101001100000;
assign LUT_2[2581] = 32'b11111111111111110100100001111001;
assign LUT_2[2582] = 32'b11111111111111111110100010011100;
assign LUT_2[2583] = 32'b11111111111111111011011010110101;
assign LUT_2[2584] = 32'b11111111111111110101111101010101;
assign LUT_2[2585] = 32'b11111111111111110010110101101110;
assign LUT_2[2586] = 32'b11111111111111111100110110010001;
assign LUT_2[2587] = 32'b11111111111111111001101110101010;
assign LUT_2[2588] = 32'b11111111111111110010011010111101;
assign LUT_2[2589] = 32'b11111111111111101111010011010110;
assign LUT_2[2590] = 32'b11111111111111111001010011111001;
assign LUT_2[2591] = 32'b11111111111111110110001100010010;
assign LUT_2[2592] = 32'b00000000000000000001000011010111;
assign LUT_2[2593] = 32'b11111111111111111101111011110000;
assign LUT_2[2594] = 32'b00000000000000000111111100010011;
assign LUT_2[2595] = 32'b00000000000000000100110100101100;
assign LUT_2[2596] = 32'b11111111111111111101100000111111;
assign LUT_2[2597] = 32'b11111111111111111010011001011000;
assign LUT_2[2598] = 32'b00000000000000000100011001111011;
assign LUT_2[2599] = 32'b00000000000000000001010010010100;
assign LUT_2[2600] = 32'b11111111111111111011110100110100;
assign LUT_2[2601] = 32'b11111111111111111000101101001101;
assign LUT_2[2602] = 32'b00000000000000000010101101110000;
assign LUT_2[2603] = 32'b11111111111111111111100110001001;
assign LUT_2[2604] = 32'b11111111111111111000010010011100;
assign LUT_2[2605] = 32'b11111111111111110101001010110101;
assign LUT_2[2606] = 32'b11111111111111111111001011011000;
assign LUT_2[2607] = 32'b11111111111111111100000011110001;
assign LUT_2[2608] = 32'b11111111111111111011100111100001;
assign LUT_2[2609] = 32'b11111111111111111000011111111010;
assign LUT_2[2610] = 32'b00000000000000000010100000011101;
assign LUT_2[2611] = 32'b11111111111111111111011000110110;
assign LUT_2[2612] = 32'b11111111111111111000000101001001;
assign LUT_2[2613] = 32'b11111111111111110100111101100010;
assign LUT_2[2614] = 32'b11111111111111111110111110000101;
assign LUT_2[2615] = 32'b11111111111111111011110110011110;
assign LUT_2[2616] = 32'b11111111111111110110011000111110;
assign LUT_2[2617] = 32'b11111111111111110011010001010111;
assign LUT_2[2618] = 32'b11111111111111111101010001111010;
assign LUT_2[2619] = 32'b11111111111111111010001010010011;
assign LUT_2[2620] = 32'b11111111111111110010110110100110;
assign LUT_2[2621] = 32'b11111111111111101111101110111111;
assign LUT_2[2622] = 32'b11111111111111111001101111100010;
assign LUT_2[2623] = 32'b11111111111111110110100111111011;
assign LUT_2[2624] = 32'b11111111111111111000110000010001;
assign LUT_2[2625] = 32'b11111111111111110101101000101010;
assign LUT_2[2626] = 32'b11111111111111111111101001001101;
assign LUT_2[2627] = 32'b11111111111111111100100001100110;
assign LUT_2[2628] = 32'b11111111111111110101001101111001;
assign LUT_2[2629] = 32'b11111111111111110010000110010010;
assign LUT_2[2630] = 32'b11111111111111111100000110110101;
assign LUT_2[2631] = 32'b11111111111111111000111111001110;
assign LUT_2[2632] = 32'b11111111111111110011100001101110;
assign LUT_2[2633] = 32'b11111111111111110000011010000111;
assign LUT_2[2634] = 32'b11111111111111111010011010101010;
assign LUT_2[2635] = 32'b11111111111111110111010011000011;
assign LUT_2[2636] = 32'b11111111111111101111111111010110;
assign LUT_2[2637] = 32'b11111111111111101100110111101111;
assign LUT_2[2638] = 32'b11111111111111110110111000010010;
assign LUT_2[2639] = 32'b11111111111111110011110000101011;
assign LUT_2[2640] = 32'b11111111111111110011010100011011;
assign LUT_2[2641] = 32'b11111111111111110000001100110100;
assign LUT_2[2642] = 32'b11111111111111111010001101010111;
assign LUT_2[2643] = 32'b11111111111111110111000101110000;
assign LUT_2[2644] = 32'b11111111111111101111110010000011;
assign LUT_2[2645] = 32'b11111111111111101100101010011100;
assign LUT_2[2646] = 32'b11111111111111110110101010111111;
assign LUT_2[2647] = 32'b11111111111111110011100011011000;
assign LUT_2[2648] = 32'b11111111111111101110000101111000;
assign LUT_2[2649] = 32'b11111111111111101010111110010001;
assign LUT_2[2650] = 32'b11111111111111110100111110110100;
assign LUT_2[2651] = 32'b11111111111111110001110111001101;
assign LUT_2[2652] = 32'b11111111111111101010100011100000;
assign LUT_2[2653] = 32'b11111111111111100111011011111001;
assign LUT_2[2654] = 32'b11111111111111110001011100011100;
assign LUT_2[2655] = 32'b11111111111111101110010100110101;
assign LUT_2[2656] = 32'b11111111111111111001001011111010;
assign LUT_2[2657] = 32'b11111111111111110110000100010011;
assign LUT_2[2658] = 32'b00000000000000000000000100110110;
assign LUT_2[2659] = 32'b11111111111111111100111101001111;
assign LUT_2[2660] = 32'b11111111111111110101101001100010;
assign LUT_2[2661] = 32'b11111111111111110010100001111011;
assign LUT_2[2662] = 32'b11111111111111111100100010011110;
assign LUT_2[2663] = 32'b11111111111111111001011010110111;
assign LUT_2[2664] = 32'b11111111111111110011111101010111;
assign LUT_2[2665] = 32'b11111111111111110000110101110000;
assign LUT_2[2666] = 32'b11111111111111111010110110010011;
assign LUT_2[2667] = 32'b11111111111111110111101110101100;
assign LUT_2[2668] = 32'b11111111111111110000011010111111;
assign LUT_2[2669] = 32'b11111111111111101101010011011000;
assign LUT_2[2670] = 32'b11111111111111110111010011111011;
assign LUT_2[2671] = 32'b11111111111111110100001100010100;
assign LUT_2[2672] = 32'b11111111111111110011110000000100;
assign LUT_2[2673] = 32'b11111111111111110000101000011101;
assign LUT_2[2674] = 32'b11111111111111111010101001000000;
assign LUT_2[2675] = 32'b11111111111111110111100001011001;
assign LUT_2[2676] = 32'b11111111111111110000001101101100;
assign LUT_2[2677] = 32'b11111111111111101101000110000101;
assign LUT_2[2678] = 32'b11111111111111110111000110101000;
assign LUT_2[2679] = 32'b11111111111111110011111111000001;
assign LUT_2[2680] = 32'b11111111111111101110100001100001;
assign LUT_2[2681] = 32'b11111111111111101011011001111010;
assign LUT_2[2682] = 32'b11111111111111110101011010011101;
assign LUT_2[2683] = 32'b11111111111111110010010010110110;
assign LUT_2[2684] = 32'b11111111111111101010111111001001;
assign LUT_2[2685] = 32'b11111111111111100111110111100010;
assign LUT_2[2686] = 32'b11111111111111110001111000000101;
assign LUT_2[2687] = 32'b11111111111111101110110000011110;
assign LUT_2[2688] = 32'b00000000000000000100111011111101;
assign LUT_2[2689] = 32'b00000000000000000001110100010110;
assign LUT_2[2690] = 32'b00000000000000001011110100111001;
assign LUT_2[2691] = 32'b00000000000000001000101101010010;
assign LUT_2[2692] = 32'b00000000000000000001011001100101;
assign LUT_2[2693] = 32'b11111111111111111110010001111110;
assign LUT_2[2694] = 32'b00000000000000001000010010100001;
assign LUT_2[2695] = 32'b00000000000000000101001010111010;
assign LUT_2[2696] = 32'b11111111111111111111101101011010;
assign LUT_2[2697] = 32'b11111111111111111100100101110011;
assign LUT_2[2698] = 32'b00000000000000000110100110010110;
assign LUT_2[2699] = 32'b00000000000000000011011110101111;
assign LUT_2[2700] = 32'b11111111111111111100001011000010;
assign LUT_2[2701] = 32'b11111111111111111001000011011011;
assign LUT_2[2702] = 32'b00000000000000000011000011111110;
assign LUT_2[2703] = 32'b11111111111111111111111100010111;
assign LUT_2[2704] = 32'b11111111111111111111100000000111;
assign LUT_2[2705] = 32'b11111111111111111100011000100000;
assign LUT_2[2706] = 32'b00000000000000000110011001000011;
assign LUT_2[2707] = 32'b00000000000000000011010001011100;
assign LUT_2[2708] = 32'b11111111111111111011111101101111;
assign LUT_2[2709] = 32'b11111111111111111000110110001000;
assign LUT_2[2710] = 32'b00000000000000000010110110101011;
assign LUT_2[2711] = 32'b11111111111111111111101111000100;
assign LUT_2[2712] = 32'b11111111111111111010010001100100;
assign LUT_2[2713] = 32'b11111111111111110111001001111101;
assign LUT_2[2714] = 32'b00000000000000000001001010100000;
assign LUT_2[2715] = 32'b11111111111111111110000010111001;
assign LUT_2[2716] = 32'b11111111111111110110101111001100;
assign LUT_2[2717] = 32'b11111111111111110011100111100101;
assign LUT_2[2718] = 32'b11111111111111111101101000001000;
assign LUT_2[2719] = 32'b11111111111111111010100000100001;
assign LUT_2[2720] = 32'b00000000000000000101010111100110;
assign LUT_2[2721] = 32'b00000000000000000010001111111111;
assign LUT_2[2722] = 32'b00000000000000001100010000100010;
assign LUT_2[2723] = 32'b00000000000000001001001000111011;
assign LUT_2[2724] = 32'b00000000000000000001110101001110;
assign LUT_2[2725] = 32'b11111111111111111110101101100111;
assign LUT_2[2726] = 32'b00000000000000001000101110001010;
assign LUT_2[2727] = 32'b00000000000000000101100110100011;
assign LUT_2[2728] = 32'b00000000000000000000001001000011;
assign LUT_2[2729] = 32'b11111111111111111101000001011100;
assign LUT_2[2730] = 32'b00000000000000000111000001111111;
assign LUT_2[2731] = 32'b00000000000000000011111010011000;
assign LUT_2[2732] = 32'b11111111111111111100100110101011;
assign LUT_2[2733] = 32'b11111111111111111001011111000100;
assign LUT_2[2734] = 32'b00000000000000000011011111100111;
assign LUT_2[2735] = 32'b00000000000000000000011000000000;
assign LUT_2[2736] = 32'b11111111111111111111111011110000;
assign LUT_2[2737] = 32'b11111111111111111100110100001001;
assign LUT_2[2738] = 32'b00000000000000000110110100101100;
assign LUT_2[2739] = 32'b00000000000000000011101101000101;
assign LUT_2[2740] = 32'b11111111111111111100011001011000;
assign LUT_2[2741] = 32'b11111111111111111001010001110001;
assign LUT_2[2742] = 32'b00000000000000000011010010010100;
assign LUT_2[2743] = 32'b00000000000000000000001010101101;
assign LUT_2[2744] = 32'b11111111111111111010101101001101;
assign LUT_2[2745] = 32'b11111111111111110111100101100110;
assign LUT_2[2746] = 32'b00000000000000000001100110001001;
assign LUT_2[2747] = 32'b11111111111111111110011110100010;
assign LUT_2[2748] = 32'b11111111111111110111001010110101;
assign LUT_2[2749] = 32'b11111111111111110100000011001110;
assign LUT_2[2750] = 32'b11111111111111111110000011110001;
assign LUT_2[2751] = 32'b11111111111111111010111100001010;
assign LUT_2[2752] = 32'b11111111111111111101000100100000;
assign LUT_2[2753] = 32'b11111111111111111001111100111001;
assign LUT_2[2754] = 32'b00000000000000000011111101011100;
assign LUT_2[2755] = 32'b00000000000000000000110101110101;
assign LUT_2[2756] = 32'b11111111111111111001100010001000;
assign LUT_2[2757] = 32'b11111111111111110110011010100001;
assign LUT_2[2758] = 32'b00000000000000000000011011000100;
assign LUT_2[2759] = 32'b11111111111111111101010011011101;
assign LUT_2[2760] = 32'b11111111111111110111110101111101;
assign LUT_2[2761] = 32'b11111111111111110100101110010110;
assign LUT_2[2762] = 32'b11111111111111111110101110111001;
assign LUT_2[2763] = 32'b11111111111111111011100111010010;
assign LUT_2[2764] = 32'b11111111111111110100010011100101;
assign LUT_2[2765] = 32'b11111111111111110001001011111110;
assign LUT_2[2766] = 32'b11111111111111111011001100100001;
assign LUT_2[2767] = 32'b11111111111111111000000100111010;
assign LUT_2[2768] = 32'b11111111111111110111101000101010;
assign LUT_2[2769] = 32'b11111111111111110100100001000011;
assign LUT_2[2770] = 32'b11111111111111111110100001100110;
assign LUT_2[2771] = 32'b11111111111111111011011001111111;
assign LUT_2[2772] = 32'b11111111111111110100000110010010;
assign LUT_2[2773] = 32'b11111111111111110000111110101011;
assign LUT_2[2774] = 32'b11111111111111111010111111001110;
assign LUT_2[2775] = 32'b11111111111111110111110111100111;
assign LUT_2[2776] = 32'b11111111111111110010011010000111;
assign LUT_2[2777] = 32'b11111111111111101111010010100000;
assign LUT_2[2778] = 32'b11111111111111111001010011000011;
assign LUT_2[2779] = 32'b11111111111111110110001011011100;
assign LUT_2[2780] = 32'b11111111111111101110110111101111;
assign LUT_2[2781] = 32'b11111111111111101011110000001000;
assign LUT_2[2782] = 32'b11111111111111110101110000101011;
assign LUT_2[2783] = 32'b11111111111111110010101001000100;
assign LUT_2[2784] = 32'b11111111111111111101100000001001;
assign LUT_2[2785] = 32'b11111111111111111010011000100010;
assign LUT_2[2786] = 32'b00000000000000000100011001000101;
assign LUT_2[2787] = 32'b00000000000000000001010001011110;
assign LUT_2[2788] = 32'b11111111111111111001111101110001;
assign LUT_2[2789] = 32'b11111111111111110110110110001010;
assign LUT_2[2790] = 32'b00000000000000000000110110101101;
assign LUT_2[2791] = 32'b11111111111111111101101111000110;
assign LUT_2[2792] = 32'b11111111111111111000010001100110;
assign LUT_2[2793] = 32'b11111111111111110101001001111111;
assign LUT_2[2794] = 32'b11111111111111111111001010100010;
assign LUT_2[2795] = 32'b11111111111111111100000010111011;
assign LUT_2[2796] = 32'b11111111111111110100101111001110;
assign LUT_2[2797] = 32'b11111111111111110001100111100111;
assign LUT_2[2798] = 32'b11111111111111111011101000001010;
assign LUT_2[2799] = 32'b11111111111111111000100000100011;
assign LUT_2[2800] = 32'b11111111111111111000000100010011;
assign LUT_2[2801] = 32'b11111111111111110100111100101100;
assign LUT_2[2802] = 32'b11111111111111111110111101001111;
assign LUT_2[2803] = 32'b11111111111111111011110101101000;
assign LUT_2[2804] = 32'b11111111111111110100100001111011;
assign LUT_2[2805] = 32'b11111111111111110001011010010100;
assign LUT_2[2806] = 32'b11111111111111111011011010110111;
assign LUT_2[2807] = 32'b11111111111111111000010011010000;
assign LUT_2[2808] = 32'b11111111111111110010110101110000;
assign LUT_2[2809] = 32'b11111111111111101111101110001001;
assign LUT_2[2810] = 32'b11111111111111111001101110101100;
assign LUT_2[2811] = 32'b11111111111111110110100111000101;
assign LUT_2[2812] = 32'b11111111111111101111010011011000;
assign LUT_2[2813] = 32'b11111111111111101100001011110001;
assign LUT_2[2814] = 32'b11111111111111110110001100010100;
assign LUT_2[2815] = 32'b11111111111111110011000100101101;
assign LUT_2[2816] = 32'b00000000000000000100100110010100;
assign LUT_2[2817] = 32'b00000000000000000001011110101101;
assign LUT_2[2818] = 32'b00000000000000001011011111010000;
assign LUT_2[2819] = 32'b00000000000000001000010111101001;
assign LUT_2[2820] = 32'b00000000000000000001000011111100;
assign LUT_2[2821] = 32'b11111111111111111101111100010101;
assign LUT_2[2822] = 32'b00000000000000000111111100111000;
assign LUT_2[2823] = 32'b00000000000000000100110101010001;
assign LUT_2[2824] = 32'b11111111111111111111010111110001;
assign LUT_2[2825] = 32'b11111111111111111100010000001010;
assign LUT_2[2826] = 32'b00000000000000000110010000101101;
assign LUT_2[2827] = 32'b00000000000000000011001001000110;
assign LUT_2[2828] = 32'b11111111111111111011110101011001;
assign LUT_2[2829] = 32'b11111111111111111000101101110010;
assign LUT_2[2830] = 32'b00000000000000000010101110010101;
assign LUT_2[2831] = 32'b11111111111111111111100110101110;
assign LUT_2[2832] = 32'b11111111111111111111001010011110;
assign LUT_2[2833] = 32'b11111111111111111100000010110111;
assign LUT_2[2834] = 32'b00000000000000000110000011011010;
assign LUT_2[2835] = 32'b00000000000000000010111011110011;
assign LUT_2[2836] = 32'b11111111111111111011101000000110;
assign LUT_2[2837] = 32'b11111111111111111000100000011111;
assign LUT_2[2838] = 32'b00000000000000000010100001000010;
assign LUT_2[2839] = 32'b11111111111111111111011001011011;
assign LUT_2[2840] = 32'b11111111111111111001111011111011;
assign LUT_2[2841] = 32'b11111111111111110110110100010100;
assign LUT_2[2842] = 32'b00000000000000000000110100110111;
assign LUT_2[2843] = 32'b11111111111111111101101101010000;
assign LUT_2[2844] = 32'b11111111111111110110011001100011;
assign LUT_2[2845] = 32'b11111111111111110011010001111100;
assign LUT_2[2846] = 32'b11111111111111111101010010011111;
assign LUT_2[2847] = 32'b11111111111111111010001010111000;
assign LUT_2[2848] = 32'b00000000000000000101000001111101;
assign LUT_2[2849] = 32'b00000000000000000001111010010110;
assign LUT_2[2850] = 32'b00000000000000001011111010111001;
assign LUT_2[2851] = 32'b00000000000000001000110011010010;
assign LUT_2[2852] = 32'b00000000000000000001011111100101;
assign LUT_2[2853] = 32'b11111111111111111110010111111110;
assign LUT_2[2854] = 32'b00000000000000001000011000100001;
assign LUT_2[2855] = 32'b00000000000000000101010000111010;
assign LUT_2[2856] = 32'b11111111111111111111110011011010;
assign LUT_2[2857] = 32'b11111111111111111100101011110011;
assign LUT_2[2858] = 32'b00000000000000000110101100010110;
assign LUT_2[2859] = 32'b00000000000000000011100100101111;
assign LUT_2[2860] = 32'b11111111111111111100010001000010;
assign LUT_2[2861] = 32'b11111111111111111001001001011011;
assign LUT_2[2862] = 32'b00000000000000000011001001111110;
assign LUT_2[2863] = 32'b00000000000000000000000010010111;
assign LUT_2[2864] = 32'b11111111111111111111100110000111;
assign LUT_2[2865] = 32'b11111111111111111100011110100000;
assign LUT_2[2866] = 32'b00000000000000000110011111000011;
assign LUT_2[2867] = 32'b00000000000000000011010111011100;
assign LUT_2[2868] = 32'b11111111111111111100000011101111;
assign LUT_2[2869] = 32'b11111111111111111000111100001000;
assign LUT_2[2870] = 32'b00000000000000000010111100101011;
assign LUT_2[2871] = 32'b11111111111111111111110101000100;
assign LUT_2[2872] = 32'b11111111111111111010010111100100;
assign LUT_2[2873] = 32'b11111111111111110111001111111101;
assign LUT_2[2874] = 32'b00000000000000000001010000100000;
assign LUT_2[2875] = 32'b11111111111111111110001000111001;
assign LUT_2[2876] = 32'b11111111111111110110110101001100;
assign LUT_2[2877] = 32'b11111111111111110011101101100101;
assign LUT_2[2878] = 32'b11111111111111111101101110001000;
assign LUT_2[2879] = 32'b11111111111111111010100110100001;
assign LUT_2[2880] = 32'b11111111111111111100101110110111;
assign LUT_2[2881] = 32'b11111111111111111001100111010000;
assign LUT_2[2882] = 32'b00000000000000000011100111110011;
assign LUT_2[2883] = 32'b00000000000000000000100000001100;
assign LUT_2[2884] = 32'b11111111111111111001001100011111;
assign LUT_2[2885] = 32'b11111111111111110110000100111000;
assign LUT_2[2886] = 32'b00000000000000000000000101011011;
assign LUT_2[2887] = 32'b11111111111111111100111101110100;
assign LUT_2[2888] = 32'b11111111111111110111100000010100;
assign LUT_2[2889] = 32'b11111111111111110100011000101101;
assign LUT_2[2890] = 32'b11111111111111111110011001010000;
assign LUT_2[2891] = 32'b11111111111111111011010001101001;
assign LUT_2[2892] = 32'b11111111111111110011111101111100;
assign LUT_2[2893] = 32'b11111111111111110000110110010101;
assign LUT_2[2894] = 32'b11111111111111111010110110111000;
assign LUT_2[2895] = 32'b11111111111111110111101111010001;
assign LUT_2[2896] = 32'b11111111111111110111010011000001;
assign LUT_2[2897] = 32'b11111111111111110100001011011010;
assign LUT_2[2898] = 32'b11111111111111111110001011111101;
assign LUT_2[2899] = 32'b11111111111111111011000100010110;
assign LUT_2[2900] = 32'b11111111111111110011110000101001;
assign LUT_2[2901] = 32'b11111111111111110000101001000010;
assign LUT_2[2902] = 32'b11111111111111111010101001100101;
assign LUT_2[2903] = 32'b11111111111111110111100001111110;
assign LUT_2[2904] = 32'b11111111111111110010000100011110;
assign LUT_2[2905] = 32'b11111111111111101110111100110111;
assign LUT_2[2906] = 32'b11111111111111111000111101011010;
assign LUT_2[2907] = 32'b11111111111111110101110101110011;
assign LUT_2[2908] = 32'b11111111111111101110100010000110;
assign LUT_2[2909] = 32'b11111111111111101011011010011111;
assign LUT_2[2910] = 32'b11111111111111110101011011000010;
assign LUT_2[2911] = 32'b11111111111111110010010011011011;
assign LUT_2[2912] = 32'b11111111111111111101001010100000;
assign LUT_2[2913] = 32'b11111111111111111010000010111001;
assign LUT_2[2914] = 32'b00000000000000000100000011011100;
assign LUT_2[2915] = 32'b00000000000000000000111011110101;
assign LUT_2[2916] = 32'b11111111111111111001101000001000;
assign LUT_2[2917] = 32'b11111111111111110110100000100001;
assign LUT_2[2918] = 32'b00000000000000000000100001000100;
assign LUT_2[2919] = 32'b11111111111111111101011001011101;
assign LUT_2[2920] = 32'b11111111111111110111111011111101;
assign LUT_2[2921] = 32'b11111111111111110100110100010110;
assign LUT_2[2922] = 32'b11111111111111111110110100111001;
assign LUT_2[2923] = 32'b11111111111111111011101101010010;
assign LUT_2[2924] = 32'b11111111111111110100011001100101;
assign LUT_2[2925] = 32'b11111111111111110001010001111110;
assign LUT_2[2926] = 32'b11111111111111111011010010100001;
assign LUT_2[2927] = 32'b11111111111111111000001010111010;
assign LUT_2[2928] = 32'b11111111111111110111101110101010;
assign LUT_2[2929] = 32'b11111111111111110100100111000011;
assign LUT_2[2930] = 32'b11111111111111111110100111100110;
assign LUT_2[2931] = 32'b11111111111111111011011111111111;
assign LUT_2[2932] = 32'b11111111111111110100001100010010;
assign LUT_2[2933] = 32'b11111111111111110001000100101011;
assign LUT_2[2934] = 32'b11111111111111111011000101001110;
assign LUT_2[2935] = 32'b11111111111111110111111101100111;
assign LUT_2[2936] = 32'b11111111111111110010100000000111;
assign LUT_2[2937] = 32'b11111111111111101111011000100000;
assign LUT_2[2938] = 32'b11111111111111111001011001000011;
assign LUT_2[2939] = 32'b11111111111111110110010001011100;
assign LUT_2[2940] = 32'b11111111111111101110111101101111;
assign LUT_2[2941] = 32'b11111111111111101011110110001000;
assign LUT_2[2942] = 32'b11111111111111110101110110101011;
assign LUT_2[2943] = 32'b11111111111111110010101111000100;
assign LUT_2[2944] = 32'b00000000000000001000111010100011;
assign LUT_2[2945] = 32'b00000000000000000101110010111100;
assign LUT_2[2946] = 32'b00000000000000001111110011011111;
assign LUT_2[2947] = 32'b00000000000000001100101011111000;
assign LUT_2[2948] = 32'b00000000000000000101011000001011;
assign LUT_2[2949] = 32'b00000000000000000010010000100100;
assign LUT_2[2950] = 32'b00000000000000001100010001000111;
assign LUT_2[2951] = 32'b00000000000000001001001001100000;
assign LUT_2[2952] = 32'b00000000000000000011101100000000;
assign LUT_2[2953] = 32'b00000000000000000000100100011001;
assign LUT_2[2954] = 32'b00000000000000001010100100111100;
assign LUT_2[2955] = 32'b00000000000000000111011101010101;
assign LUT_2[2956] = 32'b00000000000000000000001001101000;
assign LUT_2[2957] = 32'b11111111111111111101000010000001;
assign LUT_2[2958] = 32'b00000000000000000111000010100100;
assign LUT_2[2959] = 32'b00000000000000000011111010111101;
assign LUT_2[2960] = 32'b00000000000000000011011110101101;
assign LUT_2[2961] = 32'b00000000000000000000010111000110;
assign LUT_2[2962] = 32'b00000000000000001010010111101001;
assign LUT_2[2963] = 32'b00000000000000000111010000000010;
assign LUT_2[2964] = 32'b11111111111111111111111100010101;
assign LUT_2[2965] = 32'b11111111111111111100110100101110;
assign LUT_2[2966] = 32'b00000000000000000110110101010001;
assign LUT_2[2967] = 32'b00000000000000000011101101101010;
assign LUT_2[2968] = 32'b11111111111111111110010000001010;
assign LUT_2[2969] = 32'b11111111111111111011001000100011;
assign LUT_2[2970] = 32'b00000000000000000101001001000110;
assign LUT_2[2971] = 32'b00000000000000000010000001011111;
assign LUT_2[2972] = 32'b11111111111111111010101101110010;
assign LUT_2[2973] = 32'b11111111111111110111100110001011;
assign LUT_2[2974] = 32'b00000000000000000001100110101110;
assign LUT_2[2975] = 32'b11111111111111111110011111000111;
assign LUT_2[2976] = 32'b00000000000000001001010110001100;
assign LUT_2[2977] = 32'b00000000000000000110001110100101;
assign LUT_2[2978] = 32'b00000000000000010000001111001000;
assign LUT_2[2979] = 32'b00000000000000001101000111100001;
assign LUT_2[2980] = 32'b00000000000000000101110011110100;
assign LUT_2[2981] = 32'b00000000000000000010101100001101;
assign LUT_2[2982] = 32'b00000000000000001100101100110000;
assign LUT_2[2983] = 32'b00000000000000001001100101001001;
assign LUT_2[2984] = 32'b00000000000000000100000111101001;
assign LUT_2[2985] = 32'b00000000000000000001000000000010;
assign LUT_2[2986] = 32'b00000000000000001011000000100101;
assign LUT_2[2987] = 32'b00000000000000000111111000111110;
assign LUT_2[2988] = 32'b00000000000000000000100101010001;
assign LUT_2[2989] = 32'b11111111111111111101011101101010;
assign LUT_2[2990] = 32'b00000000000000000111011110001101;
assign LUT_2[2991] = 32'b00000000000000000100010110100110;
assign LUT_2[2992] = 32'b00000000000000000011111010010110;
assign LUT_2[2993] = 32'b00000000000000000000110010101111;
assign LUT_2[2994] = 32'b00000000000000001010110011010010;
assign LUT_2[2995] = 32'b00000000000000000111101011101011;
assign LUT_2[2996] = 32'b00000000000000000000010111111110;
assign LUT_2[2997] = 32'b11111111111111111101010000010111;
assign LUT_2[2998] = 32'b00000000000000000111010000111010;
assign LUT_2[2999] = 32'b00000000000000000100001001010011;
assign LUT_2[3000] = 32'b11111111111111111110101011110011;
assign LUT_2[3001] = 32'b11111111111111111011100100001100;
assign LUT_2[3002] = 32'b00000000000000000101100100101111;
assign LUT_2[3003] = 32'b00000000000000000010011101001000;
assign LUT_2[3004] = 32'b11111111111111111011001001011011;
assign LUT_2[3005] = 32'b11111111111111111000000001110100;
assign LUT_2[3006] = 32'b00000000000000000010000010010111;
assign LUT_2[3007] = 32'b11111111111111111110111010110000;
assign LUT_2[3008] = 32'b00000000000000000001000011000110;
assign LUT_2[3009] = 32'b11111111111111111101111011011111;
assign LUT_2[3010] = 32'b00000000000000000111111100000010;
assign LUT_2[3011] = 32'b00000000000000000100110100011011;
assign LUT_2[3012] = 32'b11111111111111111101100000101110;
assign LUT_2[3013] = 32'b11111111111111111010011001000111;
assign LUT_2[3014] = 32'b00000000000000000100011001101010;
assign LUT_2[3015] = 32'b00000000000000000001010010000011;
assign LUT_2[3016] = 32'b11111111111111111011110100100011;
assign LUT_2[3017] = 32'b11111111111111111000101100111100;
assign LUT_2[3018] = 32'b00000000000000000010101101011111;
assign LUT_2[3019] = 32'b11111111111111111111100101111000;
assign LUT_2[3020] = 32'b11111111111111111000010010001011;
assign LUT_2[3021] = 32'b11111111111111110101001010100100;
assign LUT_2[3022] = 32'b11111111111111111111001011000111;
assign LUT_2[3023] = 32'b11111111111111111100000011100000;
assign LUT_2[3024] = 32'b11111111111111111011100111010000;
assign LUT_2[3025] = 32'b11111111111111111000011111101001;
assign LUT_2[3026] = 32'b00000000000000000010100000001100;
assign LUT_2[3027] = 32'b11111111111111111111011000100101;
assign LUT_2[3028] = 32'b11111111111111111000000100111000;
assign LUT_2[3029] = 32'b11111111111111110100111101010001;
assign LUT_2[3030] = 32'b11111111111111111110111101110100;
assign LUT_2[3031] = 32'b11111111111111111011110110001101;
assign LUT_2[3032] = 32'b11111111111111110110011000101101;
assign LUT_2[3033] = 32'b11111111111111110011010001000110;
assign LUT_2[3034] = 32'b11111111111111111101010001101001;
assign LUT_2[3035] = 32'b11111111111111111010001010000010;
assign LUT_2[3036] = 32'b11111111111111110010110110010101;
assign LUT_2[3037] = 32'b11111111111111101111101110101110;
assign LUT_2[3038] = 32'b11111111111111111001101111010001;
assign LUT_2[3039] = 32'b11111111111111110110100111101010;
assign LUT_2[3040] = 32'b00000000000000000001011110101111;
assign LUT_2[3041] = 32'b11111111111111111110010111001000;
assign LUT_2[3042] = 32'b00000000000000001000010111101011;
assign LUT_2[3043] = 32'b00000000000000000101010000000100;
assign LUT_2[3044] = 32'b11111111111111111101111100010111;
assign LUT_2[3045] = 32'b11111111111111111010110100110000;
assign LUT_2[3046] = 32'b00000000000000000100110101010011;
assign LUT_2[3047] = 32'b00000000000000000001101101101100;
assign LUT_2[3048] = 32'b11111111111111111100010000001100;
assign LUT_2[3049] = 32'b11111111111111111001001000100101;
assign LUT_2[3050] = 32'b00000000000000000011001001001000;
assign LUT_2[3051] = 32'b00000000000000000000000001100001;
assign LUT_2[3052] = 32'b11111111111111111000101101110100;
assign LUT_2[3053] = 32'b11111111111111110101100110001101;
assign LUT_2[3054] = 32'b11111111111111111111100110110000;
assign LUT_2[3055] = 32'b11111111111111111100011111001001;
assign LUT_2[3056] = 32'b11111111111111111100000010111001;
assign LUT_2[3057] = 32'b11111111111111111000111011010010;
assign LUT_2[3058] = 32'b00000000000000000010111011110101;
assign LUT_2[3059] = 32'b11111111111111111111110100001110;
assign LUT_2[3060] = 32'b11111111111111111000100000100001;
assign LUT_2[3061] = 32'b11111111111111110101011000111010;
assign LUT_2[3062] = 32'b11111111111111111111011001011101;
assign LUT_2[3063] = 32'b11111111111111111100010001110110;
assign LUT_2[3064] = 32'b11111111111111110110110100010110;
assign LUT_2[3065] = 32'b11111111111111110011101100101111;
assign LUT_2[3066] = 32'b11111111111111111101101101010010;
assign LUT_2[3067] = 32'b11111111111111111010100101101011;
assign LUT_2[3068] = 32'b11111111111111110011010001111110;
assign LUT_2[3069] = 32'b11111111111111110000001010010111;
assign LUT_2[3070] = 32'b11111111111111111010001010111010;
assign LUT_2[3071] = 32'b11111111111111110111000011010011;
assign LUT_2[3072] = 32'b00000000000000000010100010000001;
assign LUT_2[3073] = 32'b11111111111111111111011010011010;
assign LUT_2[3074] = 32'b00000000000000001001011010111101;
assign LUT_2[3075] = 32'b00000000000000000110010011010110;
assign LUT_2[3076] = 32'b11111111111111111110111111101001;
assign LUT_2[3077] = 32'b11111111111111111011111000000010;
assign LUT_2[3078] = 32'b00000000000000000101111000100101;
assign LUT_2[3079] = 32'b00000000000000000010110000111110;
assign LUT_2[3080] = 32'b11111111111111111101010011011110;
assign LUT_2[3081] = 32'b11111111111111111010001011110111;
assign LUT_2[3082] = 32'b00000000000000000100001100011010;
assign LUT_2[3083] = 32'b00000000000000000001000100110011;
assign LUT_2[3084] = 32'b11111111111111111001110001000110;
assign LUT_2[3085] = 32'b11111111111111110110101001011111;
assign LUT_2[3086] = 32'b00000000000000000000101010000010;
assign LUT_2[3087] = 32'b11111111111111111101100010011011;
assign LUT_2[3088] = 32'b11111111111111111101000110001011;
assign LUT_2[3089] = 32'b11111111111111111001111110100100;
assign LUT_2[3090] = 32'b00000000000000000011111111000111;
assign LUT_2[3091] = 32'b00000000000000000000110111100000;
assign LUT_2[3092] = 32'b11111111111111111001100011110011;
assign LUT_2[3093] = 32'b11111111111111110110011100001100;
assign LUT_2[3094] = 32'b00000000000000000000011100101111;
assign LUT_2[3095] = 32'b11111111111111111101010101001000;
assign LUT_2[3096] = 32'b11111111111111110111110111101000;
assign LUT_2[3097] = 32'b11111111111111110100110000000001;
assign LUT_2[3098] = 32'b11111111111111111110110000100100;
assign LUT_2[3099] = 32'b11111111111111111011101000111101;
assign LUT_2[3100] = 32'b11111111111111110100010101010000;
assign LUT_2[3101] = 32'b11111111111111110001001101101001;
assign LUT_2[3102] = 32'b11111111111111111011001110001100;
assign LUT_2[3103] = 32'b11111111111111111000000110100101;
assign LUT_2[3104] = 32'b00000000000000000010111101101010;
assign LUT_2[3105] = 32'b11111111111111111111110110000011;
assign LUT_2[3106] = 32'b00000000000000001001110110100110;
assign LUT_2[3107] = 32'b00000000000000000110101110111111;
assign LUT_2[3108] = 32'b11111111111111111111011011010010;
assign LUT_2[3109] = 32'b11111111111111111100010011101011;
assign LUT_2[3110] = 32'b00000000000000000110010100001110;
assign LUT_2[3111] = 32'b00000000000000000011001100100111;
assign LUT_2[3112] = 32'b11111111111111111101101111000111;
assign LUT_2[3113] = 32'b11111111111111111010100111100000;
assign LUT_2[3114] = 32'b00000000000000000100101000000011;
assign LUT_2[3115] = 32'b00000000000000000001100000011100;
assign LUT_2[3116] = 32'b11111111111111111010001100101111;
assign LUT_2[3117] = 32'b11111111111111110111000101001000;
assign LUT_2[3118] = 32'b00000000000000000001000101101011;
assign LUT_2[3119] = 32'b11111111111111111101111110000100;
assign LUT_2[3120] = 32'b11111111111111111101100001110100;
assign LUT_2[3121] = 32'b11111111111111111010011010001101;
assign LUT_2[3122] = 32'b00000000000000000100011010110000;
assign LUT_2[3123] = 32'b00000000000000000001010011001001;
assign LUT_2[3124] = 32'b11111111111111111001111111011100;
assign LUT_2[3125] = 32'b11111111111111110110110111110101;
assign LUT_2[3126] = 32'b00000000000000000000111000011000;
assign LUT_2[3127] = 32'b11111111111111111101110000110001;
assign LUT_2[3128] = 32'b11111111111111111000010011010001;
assign LUT_2[3129] = 32'b11111111111111110101001011101010;
assign LUT_2[3130] = 32'b11111111111111111111001100001101;
assign LUT_2[3131] = 32'b11111111111111111100000100100110;
assign LUT_2[3132] = 32'b11111111111111110100110000111001;
assign LUT_2[3133] = 32'b11111111111111110001101001010010;
assign LUT_2[3134] = 32'b11111111111111111011101001110101;
assign LUT_2[3135] = 32'b11111111111111111000100010001110;
assign LUT_2[3136] = 32'b11111111111111111010101010100100;
assign LUT_2[3137] = 32'b11111111111111110111100010111101;
assign LUT_2[3138] = 32'b00000000000000000001100011100000;
assign LUT_2[3139] = 32'b11111111111111111110011011111001;
assign LUT_2[3140] = 32'b11111111111111110111001000001100;
assign LUT_2[3141] = 32'b11111111111111110100000000100101;
assign LUT_2[3142] = 32'b11111111111111111110000001001000;
assign LUT_2[3143] = 32'b11111111111111111010111001100001;
assign LUT_2[3144] = 32'b11111111111111110101011100000001;
assign LUT_2[3145] = 32'b11111111111111110010010100011010;
assign LUT_2[3146] = 32'b11111111111111111100010100111101;
assign LUT_2[3147] = 32'b11111111111111111001001101010110;
assign LUT_2[3148] = 32'b11111111111111110001111001101001;
assign LUT_2[3149] = 32'b11111111111111101110110010000010;
assign LUT_2[3150] = 32'b11111111111111111000110010100101;
assign LUT_2[3151] = 32'b11111111111111110101101010111110;
assign LUT_2[3152] = 32'b11111111111111110101001110101110;
assign LUT_2[3153] = 32'b11111111111111110010000111000111;
assign LUT_2[3154] = 32'b11111111111111111100000111101010;
assign LUT_2[3155] = 32'b11111111111111111001000000000011;
assign LUT_2[3156] = 32'b11111111111111110001101100010110;
assign LUT_2[3157] = 32'b11111111111111101110100100101111;
assign LUT_2[3158] = 32'b11111111111111111000100101010010;
assign LUT_2[3159] = 32'b11111111111111110101011101101011;
assign LUT_2[3160] = 32'b11111111111111110000000000001011;
assign LUT_2[3161] = 32'b11111111111111101100111000100100;
assign LUT_2[3162] = 32'b11111111111111110110111001000111;
assign LUT_2[3163] = 32'b11111111111111110011110001100000;
assign LUT_2[3164] = 32'b11111111111111101100011101110011;
assign LUT_2[3165] = 32'b11111111111111101001010110001100;
assign LUT_2[3166] = 32'b11111111111111110011010110101111;
assign LUT_2[3167] = 32'b11111111111111110000001111001000;
assign LUT_2[3168] = 32'b11111111111111111011000110001101;
assign LUT_2[3169] = 32'b11111111111111110111111110100110;
assign LUT_2[3170] = 32'b00000000000000000001111111001001;
assign LUT_2[3171] = 32'b11111111111111111110110111100010;
assign LUT_2[3172] = 32'b11111111111111110111100011110101;
assign LUT_2[3173] = 32'b11111111111111110100011100001110;
assign LUT_2[3174] = 32'b11111111111111111110011100110001;
assign LUT_2[3175] = 32'b11111111111111111011010101001010;
assign LUT_2[3176] = 32'b11111111111111110101110111101010;
assign LUT_2[3177] = 32'b11111111111111110010110000000011;
assign LUT_2[3178] = 32'b11111111111111111100110000100110;
assign LUT_2[3179] = 32'b11111111111111111001101000111111;
assign LUT_2[3180] = 32'b11111111111111110010010101010010;
assign LUT_2[3181] = 32'b11111111111111101111001101101011;
assign LUT_2[3182] = 32'b11111111111111111001001110001110;
assign LUT_2[3183] = 32'b11111111111111110110000110100111;
assign LUT_2[3184] = 32'b11111111111111110101101010010111;
assign LUT_2[3185] = 32'b11111111111111110010100010110000;
assign LUT_2[3186] = 32'b11111111111111111100100011010011;
assign LUT_2[3187] = 32'b11111111111111111001011011101100;
assign LUT_2[3188] = 32'b11111111111111110010000111111111;
assign LUT_2[3189] = 32'b11111111111111101111000000011000;
assign LUT_2[3190] = 32'b11111111111111111001000000111011;
assign LUT_2[3191] = 32'b11111111111111110101111001010100;
assign LUT_2[3192] = 32'b11111111111111110000011011110100;
assign LUT_2[3193] = 32'b11111111111111101101010100001101;
assign LUT_2[3194] = 32'b11111111111111110111010100110000;
assign LUT_2[3195] = 32'b11111111111111110100001101001001;
assign LUT_2[3196] = 32'b11111111111111101100111001011100;
assign LUT_2[3197] = 32'b11111111111111101001110001110101;
assign LUT_2[3198] = 32'b11111111111111110011110010011000;
assign LUT_2[3199] = 32'b11111111111111110000101010110001;
assign LUT_2[3200] = 32'b00000000000000000110110110010000;
assign LUT_2[3201] = 32'b00000000000000000011101110101001;
assign LUT_2[3202] = 32'b00000000000000001101101111001100;
assign LUT_2[3203] = 32'b00000000000000001010100111100101;
assign LUT_2[3204] = 32'b00000000000000000011010011111000;
assign LUT_2[3205] = 32'b00000000000000000000001100010001;
assign LUT_2[3206] = 32'b00000000000000001010001100110100;
assign LUT_2[3207] = 32'b00000000000000000111000101001101;
assign LUT_2[3208] = 32'b00000000000000000001100111101101;
assign LUT_2[3209] = 32'b11111111111111111110100000000110;
assign LUT_2[3210] = 32'b00000000000000001000100000101001;
assign LUT_2[3211] = 32'b00000000000000000101011001000010;
assign LUT_2[3212] = 32'b11111111111111111110000101010101;
assign LUT_2[3213] = 32'b11111111111111111010111101101110;
assign LUT_2[3214] = 32'b00000000000000000100111110010001;
assign LUT_2[3215] = 32'b00000000000000000001110110101010;
assign LUT_2[3216] = 32'b00000000000000000001011010011010;
assign LUT_2[3217] = 32'b11111111111111111110010010110011;
assign LUT_2[3218] = 32'b00000000000000001000010011010110;
assign LUT_2[3219] = 32'b00000000000000000101001011101111;
assign LUT_2[3220] = 32'b11111111111111111101111000000010;
assign LUT_2[3221] = 32'b11111111111111111010110000011011;
assign LUT_2[3222] = 32'b00000000000000000100110000111110;
assign LUT_2[3223] = 32'b00000000000000000001101001010111;
assign LUT_2[3224] = 32'b11111111111111111100001011110111;
assign LUT_2[3225] = 32'b11111111111111111001000100010000;
assign LUT_2[3226] = 32'b00000000000000000011000100110011;
assign LUT_2[3227] = 32'b11111111111111111111111101001100;
assign LUT_2[3228] = 32'b11111111111111111000101001011111;
assign LUT_2[3229] = 32'b11111111111111110101100001111000;
assign LUT_2[3230] = 32'b11111111111111111111100010011011;
assign LUT_2[3231] = 32'b11111111111111111100011010110100;
assign LUT_2[3232] = 32'b00000000000000000111010001111001;
assign LUT_2[3233] = 32'b00000000000000000100001010010010;
assign LUT_2[3234] = 32'b00000000000000001110001010110101;
assign LUT_2[3235] = 32'b00000000000000001011000011001110;
assign LUT_2[3236] = 32'b00000000000000000011101111100001;
assign LUT_2[3237] = 32'b00000000000000000000100111111010;
assign LUT_2[3238] = 32'b00000000000000001010101000011101;
assign LUT_2[3239] = 32'b00000000000000000111100000110110;
assign LUT_2[3240] = 32'b00000000000000000010000011010110;
assign LUT_2[3241] = 32'b11111111111111111110111011101111;
assign LUT_2[3242] = 32'b00000000000000001000111100010010;
assign LUT_2[3243] = 32'b00000000000000000101110100101011;
assign LUT_2[3244] = 32'b11111111111111111110100000111110;
assign LUT_2[3245] = 32'b11111111111111111011011001010111;
assign LUT_2[3246] = 32'b00000000000000000101011001111010;
assign LUT_2[3247] = 32'b00000000000000000010010010010011;
assign LUT_2[3248] = 32'b00000000000000000001110110000011;
assign LUT_2[3249] = 32'b11111111111111111110101110011100;
assign LUT_2[3250] = 32'b00000000000000001000101110111111;
assign LUT_2[3251] = 32'b00000000000000000101100111011000;
assign LUT_2[3252] = 32'b11111111111111111110010011101011;
assign LUT_2[3253] = 32'b11111111111111111011001100000100;
assign LUT_2[3254] = 32'b00000000000000000101001100100111;
assign LUT_2[3255] = 32'b00000000000000000010000101000000;
assign LUT_2[3256] = 32'b11111111111111111100100111100000;
assign LUT_2[3257] = 32'b11111111111111111001011111111001;
assign LUT_2[3258] = 32'b00000000000000000011100000011100;
assign LUT_2[3259] = 32'b00000000000000000000011000110101;
assign LUT_2[3260] = 32'b11111111111111111001000101001000;
assign LUT_2[3261] = 32'b11111111111111110101111101100001;
assign LUT_2[3262] = 32'b11111111111111111111111110000100;
assign LUT_2[3263] = 32'b11111111111111111100110110011101;
assign LUT_2[3264] = 32'b11111111111111111110111110110011;
assign LUT_2[3265] = 32'b11111111111111111011110111001100;
assign LUT_2[3266] = 32'b00000000000000000101110111101111;
assign LUT_2[3267] = 32'b00000000000000000010110000001000;
assign LUT_2[3268] = 32'b11111111111111111011011100011011;
assign LUT_2[3269] = 32'b11111111111111111000010100110100;
assign LUT_2[3270] = 32'b00000000000000000010010101010111;
assign LUT_2[3271] = 32'b11111111111111111111001101110000;
assign LUT_2[3272] = 32'b11111111111111111001110000010000;
assign LUT_2[3273] = 32'b11111111111111110110101000101001;
assign LUT_2[3274] = 32'b00000000000000000000101001001100;
assign LUT_2[3275] = 32'b11111111111111111101100001100101;
assign LUT_2[3276] = 32'b11111111111111110110001101111000;
assign LUT_2[3277] = 32'b11111111111111110011000110010001;
assign LUT_2[3278] = 32'b11111111111111111101000110110100;
assign LUT_2[3279] = 32'b11111111111111111001111111001101;
assign LUT_2[3280] = 32'b11111111111111111001100010111101;
assign LUT_2[3281] = 32'b11111111111111110110011011010110;
assign LUT_2[3282] = 32'b00000000000000000000011011111001;
assign LUT_2[3283] = 32'b11111111111111111101010100010010;
assign LUT_2[3284] = 32'b11111111111111110110000000100101;
assign LUT_2[3285] = 32'b11111111111111110010111000111110;
assign LUT_2[3286] = 32'b11111111111111111100111001100001;
assign LUT_2[3287] = 32'b11111111111111111001110001111010;
assign LUT_2[3288] = 32'b11111111111111110100010100011010;
assign LUT_2[3289] = 32'b11111111111111110001001100110011;
assign LUT_2[3290] = 32'b11111111111111111011001101010110;
assign LUT_2[3291] = 32'b11111111111111111000000101101111;
assign LUT_2[3292] = 32'b11111111111111110000110010000010;
assign LUT_2[3293] = 32'b11111111111111101101101010011011;
assign LUT_2[3294] = 32'b11111111111111110111101010111110;
assign LUT_2[3295] = 32'b11111111111111110100100011010111;
assign LUT_2[3296] = 32'b11111111111111111111011010011100;
assign LUT_2[3297] = 32'b11111111111111111100010010110101;
assign LUT_2[3298] = 32'b00000000000000000110010011011000;
assign LUT_2[3299] = 32'b00000000000000000011001011110001;
assign LUT_2[3300] = 32'b11111111111111111011111000000100;
assign LUT_2[3301] = 32'b11111111111111111000110000011101;
assign LUT_2[3302] = 32'b00000000000000000010110001000000;
assign LUT_2[3303] = 32'b11111111111111111111101001011001;
assign LUT_2[3304] = 32'b11111111111111111010001011111001;
assign LUT_2[3305] = 32'b11111111111111110111000100010010;
assign LUT_2[3306] = 32'b00000000000000000001000100110101;
assign LUT_2[3307] = 32'b11111111111111111101111101001110;
assign LUT_2[3308] = 32'b11111111111111110110101001100001;
assign LUT_2[3309] = 32'b11111111111111110011100001111010;
assign LUT_2[3310] = 32'b11111111111111111101100010011101;
assign LUT_2[3311] = 32'b11111111111111111010011010110110;
assign LUT_2[3312] = 32'b11111111111111111001111110100110;
assign LUT_2[3313] = 32'b11111111111111110110110110111111;
assign LUT_2[3314] = 32'b00000000000000000000110111100010;
assign LUT_2[3315] = 32'b11111111111111111101101111111011;
assign LUT_2[3316] = 32'b11111111111111110110011100001110;
assign LUT_2[3317] = 32'b11111111111111110011010100100111;
assign LUT_2[3318] = 32'b11111111111111111101010101001010;
assign LUT_2[3319] = 32'b11111111111111111010001101100011;
assign LUT_2[3320] = 32'b11111111111111110100110000000011;
assign LUT_2[3321] = 32'b11111111111111110001101000011100;
assign LUT_2[3322] = 32'b11111111111111111011101000111111;
assign LUT_2[3323] = 32'b11111111111111111000100001011000;
assign LUT_2[3324] = 32'b11111111111111110001001101101011;
assign LUT_2[3325] = 32'b11111111111111101110000110000100;
assign LUT_2[3326] = 32'b11111111111111111000000110100111;
assign LUT_2[3327] = 32'b11111111111111110100111111000000;
assign LUT_2[3328] = 32'b00000000000000000110100000100111;
assign LUT_2[3329] = 32'b00000000000000000011011001000000;
assign LUT_2[3330] = 32'b00000000000000001101011001100011;
assign LUT_2[3331] = 32'b00000000000000001010010001111100;
assign LUT_2[3332] = 32'b00000000000000000010111110001111;
assign LUT_2[3333] = 32'b11111111111111111111110110101000;
assign LUT_2[3334] = 32'b00000000000000001001110111001011;
assign LUT_2[3335] = 32'b00000000000000000110101111100100;
assign LUT_2[3336] = 32'b00000000000000000001010010000100;
assign LUT_2[3337] = 32'b11111111111111111110001010011101;
assign LUT_2[3338] = 32'b00000000000000001000001011000000;
assign LUT_2[3339] = 32'b00000000000000000101000011011001;
assign LUT_2[3340] = 32'b11111111111111111101101111101100;
assign LUT_2[3341] = 32'b11111111111111111010101000000101;
assign LUT_2[3342] = 32'b00000000000000000100101000101000;
assign LUT_2[3343] = 32'b00000000000000000001100001000001;
assign LUT_2[3344] = 32'b00000000000000000001000100110001;
assign LUT_2[3345] = 32'b11111111111111111101111101001010;
assign LUT_2[3346] = 32'b00000000000000000111111101101101;
assign LUT_2[3347] = 32'b00000000000000000100110110000110;
assign LUT_2[3348] = 32'b11111111111111111101100010011001;
assign LUT_2[3349] = 32'b11111111111111111010011010110010;
assign LUT_2[3350] = 32'b00000000000000000100011011010101;
assign LUT_2[3351] = 32'b00000000000000000001010011101110;
assign LUT_2[3352] = 32'b11111111111111111011110110001110;
assign LUT_2[3353] = 32'b11111111111111111000101110100111;
assign LUT_2[3354] = 32'b00000000000000000010101111001010;
assign LUT_2[3355] = 32'b11111111111111111111100111100011;
assign LUT_2[3356] = 32'b11111111111111111000010011110110;
assign LUT_2[3357] = 32'b11111111111111110101001100001111;
assign LUT_2[3358] = 32'b11111111111111111111001100110010;
assign LUT_2[3359] = 32'b11111111111111111100000101001011;
assign LUT_2[3360] = 32'b00000000000000000110111100010000;
assign LUT_2[3361] = 32'b00000000000000000011110100101001;
assign LUT_2[3362] = 32'b00000000000000001101110101001100;
assign LUT_2[3363] = 32'b00000000000000001010101101100101;
assign LUT_2[3364] = 32'b00000000000000000011011001111000;
assign LUT_2[3365] = 32'b00000000000000000000010010010001;
assign LUT_2[3366] = 32'b00000000000000001010010010110100;
assign LUT_2[3367] = 32'b00000000000000000111001011001101;
assign LUT_2[3368] = 32'b00000000000000000001101101101101;
assign LUT_2[3369] = 32'b11111111111111111110100110000110;
assign LUT_2[3370] = 32'b00000000000000001000100110101001;
assign LUT_2[3371] = 32'b00000000000000000101011111000010;
assign LUT_2[3372] = 32'b11111111111111111110001011010101;
assign LUT_2[3373] = 32'b11111111111111111011000011101110;
assign LUT_2[3374] = 32'b00000000000000000101000100010001;
assign LUT_2[3375] = 32'b00000000000000000001111100101010;
assign LUT_2[3376] = 32'b00000000000000000001100000011010;
assign LUT_2[3377] = 32'b11111111111111111110011000110011;
assign LUT_2[3378] = 32'b00000000000000001000011001010110;
assign LUT_2[3379] = 32'b00000000000000000101010001101111;
assign LUT_2[3380] = 32'b11111111111111111101111110000010;
assign LUT_2[3381] = 32'b11111111111111111010110110011011;
assign LUT_2[3382] = 32'b00000000000000000100110110111110;
assign LUT_2[3383] = 32'b00000000000000000001101111010111;
assign LUT_2[3384] = 32'b11111111111111111100010001110111;
assign LUT_2[3385] = 32'b11111111111111111001001010010000;
assign LUT_2[3386] = 32'b00000000000000000011001010110011;
assign LUT_2[3387] = 32'b00000000000000000000000011001100;
assign LUT_2[3388] = 32'b11111111111111111000101111011111;
assign LUT_2[3389] = 32'b11111111111111110101100111111000;
assign LUT_2[3390] = 32'b11111111111111111111101000011011;
assign LUT_2[3391] = 32'b11111111111111111100100000110100;
assign LUT_2[3392] = 32'b11111111111111111110101001001010;
assign LUT_2[3393] = 32'b11111111111111111011100001100011;
assign LUT_2[3394] = 32'b00000000000000000101100010000110;
assign LUT_2[3395] = 32'b00000000000000000010011010011111;
assign LUT_2[3396] = 32'b11111111111111111011000110110010;
assign LUT_2[3397] = 32'b11111111111111110111111111001011;
assign LUT_2[3398] = 32'b00000000000000000001111111101110;
assign LUT_2[3399] = 32'b11111111111111111110111000000111;
assign LUT_2[3400] = 32'b11111111111111111001011010100111;
assign LUT_2[3401] = 32'b11111111111111110110010011000000;
assign LUT_2[3402] = 32'b00000000000000000000010011100011;
assign LUT_2[3403] = 32'b11111111111111111101001011111100;
assign LUT_2[3404] = 32'b11111111111111110101111000001111;
assign LUT_2[3405] = 32'b11111111111111110010110000101000;
assign LUT_2[3406] = 32'b11111111111111111100110001001011;
assign LUT_2[3407] = 32'b11111111111111111001101001100100;
assign LUT_2[3408] = 32'b11111111111111111001001101010100;
assign LUT_2[3409] = 32'b11111111111111110110000101101101;
assign LUT_2[3410] = 32'b00000000000000000000000110010000;
assign LUT_2[3411] = 32'b11111111111111111100111110101001;
assign LUT_2[3412] = 32'b11111111111111110101101010111100;
assign LUT_2[3413] = 32'b11111111111111110010100011010101;
assign LUT_2[3414] = 32'b11111111111111111100100011111000;
assign LUT_2[3415] = 32'b11111111111111111001011100010001;
assign LUT_2[3416] = 32'b11111111111111110011111110110001;
assign LUT_2[3417] = 32'b11111111111111110000110111001010;
assign LUT_2[3418] = 32'b11111111111111111010110111101101;
assign LUT_2[3419] = 32'b11111111111111110111110000000110;
assign LUT_2[3420] = 32'b11111111111111110000011100011001;
assign LUT_2[3421] = 32'b11111111111111101101010100110010;
assign LUT_2[3422] = 32'b11111111111111110111010101010101;
assign LUT_2[3423] = 32'b11111111111111110100001101101110;
assign LUT_2[3424] = 32'b11111111111111111111000100110011;
assign LUT_2[3425] = 32'b11111111111111111011111101001100;
assign LUT_2[3426] = 32'b00000000000000000101111101101111;
assign LUT_2[3427] = 32'b00000000000000000010110110001000;
assign LUT_2[3428] = 32'b11111111111111111011100010011011;
assign LUT_2[3429] = 32'b11111111111111111000011010110100;
assign LUT_2[3430] = 32'b00000000000000000010011011010111;
assign LUT_2[3431] = 32'b11111111111111111111010011110000;
assign LUT_2[3432] = 32'b11111111111111111001110110010000;
assign LUT_2[3433] = 32'b11111111111111110110101110101001;
assign LUT_2[3434] = 32'b00000000000000000000101111001100;
assign LUT_2[3435] = 32'b11111111111111111101100111100101;
assign LUT_2[3436] = 32'b11111111111111110110010011111000;
assign LUT_2[3437] = 32'b11111111111111110011001100010001;
assign LUT_2[3438] = 32'b11111111111111111101001100110100;
assign LUT_2[3439] = 32'b11111111111111111010000101001101;
assign LUT_2[3440] = 32'b11111111111111111001101000111101;
assign LUT_2[3441] = 32'b11111111111111110110100001010110;
assign LUT_2[3442] = 32'b00000000000000000000100001111001;
assign LUT_2[3443] = 32'b11111111111111111101011010010010;
assign LUT_2[3444] = 32'b11111111111111110110000110100101;
assign LUT_2[3445] = 32'b11111111111111110010111110111110;
assign LUT_2[3446] = 32'b11111111111111111100111111100001;
assign LUT_2[3447] = 32'b11111111111111111001110111111010;
assign LUT_2[3448] = 32'b11111111111111110100011010011010;
assign LUT_2[3449] = 32'b11111111111111110001010010110011;
assign LUT_2[3450] = 32'b11111111111111111011010011010110;
assign LUT_2[3451] = 32'b11111111111111111000001011101111;
assign LUT_2[3452] = 32'b11111111111111110000111000000010;
assign LUT_2[3453] = 32'b11111111111111101101110000011011;
assign LUT_2[3454] = 32'b11111111111111110111110000111110;
assign LUT_2[3455] = 32'b11111111111111110100101001010111;
assign LUT_2[3456] = 32'b00000000000000001010110100110110;
assign LUT_2[3457] = 32'b00000000000000000111101101001111;
assign LUT_2[3458] = 32'b00000000000000010001101101110010;
assign LUT_2[3459] = 32'b00000000000000001110100110001011;
assign LUT_2[3460] = 32'b00000000000000000111010010011110;
assign LUT_2[3461] = 32'b00000000000000000100001010110111;
assign LUT_2[3462] = 32'b00000000000000001110001011011010;
assign LUT_2[3463] = 32'b00000000000000001011000011110011;
assign LUT_2[3464] = 32'b00000000000000000101100110010011;
assign LUT_2[3465] = 32'b00000000000000000010011110101100;
assign LUT_2[3466] = 32'b00000000000000001100011111001111;
assign LUT_2[3467] = 32'b00000000000000001001010111101000;
assign LUT_2[3468] = 32'b00000000000000000010000011111011;
assign LUT_2[3469] = 32'b11111111111111111110111100010100;
assign LUT_2[3470] = 32'b00000000000000001000111100110111;
assign LUT_2[3471] = 32'b00000000000000000101110101010000;
assign LUT_2[3472] = 32'b00000000000000000101011001000000;
assign LUT_2[3473] = 32'b00000000000000000010010001011001;
assign LUT_2[3474] = 32'b00000000000000001100010001111100;
assign LUT_2[3475] = 32'b00000000000000001001001010010101;
assign LUT_2[3476] = 32'b00000000000000000001110110101000;
assign LUT_2[3477] = 32'b11111111111111111110101111000001;
assign LUT_2[3478] = 32'b00000000000000001000101111100100;
assign LUT_2[3479] = 32'b00000000000000000101100111111101;
assign LUT_2[3480] = 32'b00000000000000000000001010011101;
assign LUT_2[3481] = 32'b11111111111111111101000010110110;
assign LUT_2[3482] = 32'b00000000000000000111000011011001;
assign LUT_2[3483] = 32'b00000000000000000011111011110010;
assign LUT_2[3484] = 32'b11111111111111111100101000000101;
assign LUT_2[3485] = 32'b11111111111111111001100000011110;
assign LUT_2[3486] = 32'b00000000000000000011100001000001;
assign LUT_2[3487] = 32'b00000000000000000000011001011010;
assign LUT_2[3488] = 32'b00000000000000001011010000011111;
assign LUT_2[3489] = 32'b00000000000000001000001000111000;
assign LUT_2[3490] = 32'b00000000000000010010001001011011;
assign LUT_2[3491] = 32'b00000000000000001111000001110100;
assign LUT_2[3492] = 32'b00000000000000000111101110000111;
assign LUT_2[3493] = 32'b00000000000000000100100110100000;
assign LUT_2[3494] = 32'b00000000000000001110100111000011;
assign LUT_2[3495] = 32'b00000000000000001011011111011100;
assign LUT_2[3496] = 32'b00000000000000000110000001111100;
assign LUT_2[3497] = 32'b00000000000000000010111010010101;
assign LUT_2[3498] = 32'b00000000000000001100111010111000;
assign LUT_2[3499] = 32'b00000000000000001001110011010001;
assign LUT_2[3500] = 32'b00000000000000000010011111100100;
assign LUT_2[3501] = 32'b11111111111111111111010111111101;
assign LUT_2[3502] = 32'b00000000000000001001011000100000;
assign LUT_2[3503] = 32'b00000000000000000110010000111001;
assign LUT_2[3504] = 32'b00000000000000000101110100101001;
assign LUT_2[3505] = 32'b00000000000000000010101101000010;
assign LUT_2[3506] = 32'b00000000000000001100101101100101;
assign LUT_2[3507] = 32'b00000000000000001001100101111110;
assign LUT_2[3508] = 32'b00000000000000000010010010010001;
assign LUT_2[3509] = 32'b11111111111111111111001010101010;
assign LUT_2[3510] = 32'b00000000000000001001001011001101;
assign LUT_2[3511] = 32'b00000000000000000110000011100110;
assign LUT_2[3512] = 32'b00000000000000000000100110000110;
assign LUT_2[3513] = 32'b11111111111111111101011110011111;
assign LUT_2[3514] = 32'b00000000000000000111011111000010;
assign LUT_2[3515] = 32'b00000000000000000100010111011011;
assign LUT_2[3516] = 32'b11111111111111111101000011101110;
assign LUT_2[3517] = 32'b11111111111111111001111100000111;
assign LUT_2[3518] = 32'b00000000000000000011111100101010;
assign LUT_2[3519] = 32'b00000000000000000000110101000011;
assign LUT_2[3520] = 32'b00000000000000000010111101011001;
assign LUT_2[3521] = 32'b11111111111111111111110101110010;
assign LUT_2[3522] = 32'b00000000000000001001110110010101;
assign LUT_2[3523] = 32'b00000000000000000110101110101110;
assign LUT_2[3524] = 32'b11111111111111111111011011000001;
assign LUT_2[3525] = 32'b11111111111111111100010011011010;
assign LUT_2[3526] = 32'b00000000000000000110010011111101;
assign LUT_2[3527] = 32'b00000000000000000011001100010110;
assign LUT_2[3528] = 32'b11111111111111111101101110110110;
assign LUT_2[3529] = 32'b11111111111111111010100111001111;
assign LUT_2[3530] = 32'b00000000000000000100100111110010;
assign LUT_2[3531] = 32'b00000000000000000001100000001011;
assign LUT_2[3532] = 32'b11111111111111111010001100011110;
assign LUT_2[3533] = 32'b11111111111111110111000100110111;
assign LUT_2[3534] = 32'b00000000000000000001000101011010;
assign LUT_2[3535] = 32'b11111111111111111101111101110011;
assign LUT_2[3536] = 32'b11111111111111111101100001100011;
assign LUT_2[3537] = 32'b11111111111111111010011001111100;
assign LUT_2[3538] = 32'b00000000000000000100011010011111;
assign LUT_2[3539] = 32'b00000000000000000001010010111000;
assign LUT_2[3540] = 32'b11111111111111111001111111001011;
assign LUT_2[3541] = 32'b11111111111111110110110111100100;
assign LUT_2[3542] = 32'b00000000000000000000111000000111;
assign LUT_2[3543] = 32'b11111111111111111101110000100000;
assign LUT_2[3544] = 32'b11111111111111111000010011000000;
assign LUT_2[3545] = 32'b11111111111111110101001011011001;
assign LUT_2[3546] = 32'b11111111111111111111001011111100;
assign LUT_2[3547] = 32'b11111111111111111100000100010101;
assign LUT_2[3548] = 32'b11111111111111110100110000101000;
assign LUT_2[3549] = 32'b11111111111111110001101001000001;
assign LUT_2[3550] = 32'b11111111111111111011101001100100;
assign LUT_2[3551] = 32'b11111111111111111000100001111101;
assign LUT_2[3552] = 32'b00000000000000000011011001000010;
assign LUT_2[3553] = 32'b00000000000000000000010001011011;
assign LUT_2[3554] = 32'b00000000000000001010010001111110;
assign LUT_2[3555] = 32'b00000000000000000111001010010111;
assign LUT_2[3556] = 32'b11111111111111111111110110101010;
assign LUT_2[3557] = 32'b11111111111111111100101111000011;
assign LUT_2[3558] = 32'b00000000000000000110101111100110;
assign LUT_2[3559] = 32'b00000000000000000011100111111111;
assign LUT_2[3560] = 32'b11111111111111111110001010011111;
assign LUT_2[3561] = 32'b11111111111111111011000010111000;
assign LUT_2[3562] = 32'b00000000000000000101000011011011;
assign LUT_2[3563] = 32'b00000000000000000001111011110100;
assign LUT_2[3564] = 32'b11111111111111111010101000000111;
assign LUT_2[3565] = 32'b11111111111111110111100000100000;
assign LUT_2[3566] = 32'b00000000000000000001100001000011;
assign LUT_2[3567] = 32'b11111111111111111110011001011100;
assign LUT_2[3568] = 32'b11111111111111111101111101001100;
assign LUT_2[3569] = 32'b11111111111111111010110101100101;
assign LUT_2[3570] = 32'b00000000000000000100110110001000;
assign LUT_2[3571] = 32'b00000000000000000001101110100001;
assign LUT_2[3572] = 32'b11111111111111111010011010110100;
assign LUT_2[3573] = 32'b11111111111111110111010011001101;
assign LUT_2[3574] = 32'b00000000000000000001010011110000;
assign LUT_2[3575] = 32'b11111111111111111110001100001001;
assign LUT_2[3576] = 32'b11111111111111111000101110101001;
assign LUT_2[3577] = 32'b11111111111111110101100111000010;
assign LUT_2[3578] = 32'b11111111111111111111100111100101;
assign LUT_2[3579] = 32'b11111111111111111100011111111110;
assign LUT_2[3580] = 32'b11111111111111110101001100010001;
assign LUT_2[3581] = 32'b11111111111111110010000100101010;
assign LUT_2[3582] = 32'b11111111111111111100000101001101;
assign LUT_2[3583] = 32'b11111111111111111000111101100110;
assign LUT_2[3584] = 32'b00000000000000000111010011110011;
assign LUT_2[3585] = 32'b00000000000000000100001100001100;
assign LUT_2[3586] = 32'b00000000000000001110001100101111;
assign LUT_2[3587] = 32'b00000000000000001011000101001000;
assign LUT_2[3588] = 32'b00000000000000000011110001011011;
assign LUT_2[3589] = 32'b00000000000000000000101001110100;
assign LUT_2[3590] = 32'b00000000000000001010101010010111;
assign LUT_2[3591] = 32'b00000000000000000111100010110000;
assign LUT_2[3592] = 32'b00000000000000000010000101010000;
assign LUT_2[3593] = 32'b11111111111111111110111101101001;
assign LUT_2[3594] = 32'b00000000000000001000111110001100;
assign LUT_2[3595] = 32'b00000000000000000101110110100101;
assign LUT_2[3596] = 32'b11111111111111111110100010111000;
assign LUT_2[3597] = 32'b11111111111111111011011011010001;
assign LUT_2[3598] = 32'b00000000000000000101011011110100;
assign LUT_2[3599] = 32'b00000000000000000010010100001101;
assign LUT_2[3600] = 32'b00000000000000000001110111111101;
assign LUT_2[3601] = 32'b11111111111111111110110000010110;
assign LUT_2[3602] = 32'b00000000000000001000110000111001;
assign LUT_2[3603] = 32'b00000000000000000101101001010010;
assign LUT_2[3604] = 32'b11111111111111111110010101100101;
assign LUT_2[3605] = 32'b11111111111111111011001101111110;
assign LUT_2[3606] = 32'b00000000000000000101001110100001;
assign LUT_2[3607] = 32'b00000000000000000010000110111010;
assign LUT_2[3608] = 32'b11111111111111111100101001011010;
assign LUT_2[3609] = 32'b11111111111111111001100001110011;
assign LUT_2[3610] = 32'b00000000000000000011100010010110;
assign LUT_2[3611] = 32'b00000000000000000000011010101111;
assign LUT_2[3612] = 32'b11111111111111111001000111000010;
assign LUT_2[3613] = 32'b11111111111111110101111111011011;
assign LUT_2[3614] = 32'b11111111111111111111111111111110;
assign LUT_2[3615] = 32'b11111111111111111100111000010111;
assign LUT_2[3616] = 32'b00000000000000000111101111011100;
assign LUT_2[3617] = 32'b00000000000000000100100111110101;
assign LUT_2[3618] = 32'b00000000000000001110101000011000;
assign LUT_2[3619] = 32'b00000000000000001011100000110001;
assign LUT_2[3620] = 32'b00000000000000000100001101000100;
assign LUT_2[3621] = 32'b00000000000000000001000101011101;
assign LUT_2[3622] = 32'b00000000000000001011000110000000;
assign LUT_2[3623] = 32'b00000000000000000111111110011001;
assign LUT_2[3624] = 32'b00000000000000000010100000111001;
assign LUT_2[3625] = 32'b11111111111111111111011001010010;
assign LUT_2[3626] = 32'b00000000000000001001011001110101;
assign LUT_2[3627] = 32'b00000000000000000110010010001110;
assign LUT_2[3628] = 32'b11111111111111111110111110100001;
assign LUT_2[3629] = 32'b11111111111111111011110110111010;
assign LUT_2[3630] = 32'b00000000000000000101110111011101;
assign LUT_2[3631] = 32'b00000000000000000010101111110110;
assign LUT_2[3632] = 32'b00000000000000000010010011100110;
assign LUT_2[3633] = 32'b11111111111111111111001011111111;
assign LUT_2[3634] = 32'b00000000000000001001001100100010;
assign LUT_2[3635] = 32'b00000000000000000110000100111011;
assign LUT_2[3636] = 32'b11111111111111111110110001001110;
assign LUT_2[3637] = 32'b11111111111111111011101001100111;
assign LUT_2[3638] = 32'b00000000000000000101101010001010;
assign LUT_2[3639] = 32'b00000000000000000010100010100011;
assign LUT_2[3640] = 32'b11111111111111111101000101000011;
assign LUT_2[3641] = 32'b11111111111111111001111101011100;
assign LUT_2[3642] = 32'b00000000000000000011111101111111;
assign LUT_2[3643] = 32'b00000000000000000000110110011000;
assign LUT_2[3644] = 32'b11111111111111111001100010101011;
assign LUT_2[3645] = 32'b11111111111111110110011011000100;
assign LUT_2[3646] = 32'b00000000000000000000011011100111;
assign LUT_2[3647] = 32'b11111111111111111101010100000000;
assign LUT_2[3648] = 32'b11111111111111111111011100010110;
assign LUT_2[3649] = 32'b11111111111111111100010100101111;
assign LUT_2[3650] = 32'b00000000000000000110010101010010;
assign LUT_2[3651] = 32'b00000000000000000011001101101011;
assign LUT_2[3652] = 32'b11111111111111111011111001111110;
assign LUT_2[3653] = 32'b11111111111111111000110010010111;
assign LUT_2[3654] = 32'b00000000000000000010110010111010;
assign LUT_2[3655] = 32'b11111111111111111111101011010011;
assign LUT_2[3656] = 32'b11111111111111111010001101110011;
assign LUT_2[3657] = 32'b11111111111111110111000110001100;
assign LUT_2[3658] = 32'b00000000000000000001000110101111;
assign LUT_2[3659] = 32'b11111111111111111101111111001000;
assign LUT_2[3660] = 32'b11111111111111110110101011011011;
assign LUT_2[3661] = 32'b11111111111111110011100011110100;
assign LUT_2[3662] = 32'b11111111111111111101100100010111;
assign LUT_2[3663] = 32'b11111111111111111010011100110000;
assign LUT_2[3664] = 32'b11111111111111111010000000100000;
assign LUT_2[3665] = 32'b11111111111111110110111000111001;
assign LUT_2[3666] = 32'b00000000000000000000111001011100;
assign LUT_2[3667] = 32'b11111111111111111101110001110101;
assign LUT_2[3668] = 32'b11111111111111110110011110001000;
assign LUT_2[3669] = 32'b11111111111111110011010110100001;
assign LUT_2[3670] = 32'b11111111111111111101010111000100;
assign LUT_2[3671] = 32'b11111111111111111010001111011101;
assign LUT_2[3672] = 32'b11111111111111110100110001111101;
assign LUT_2[3673] = 32'b11111111111111110001101010010110;
assign LUT_2[3674] = 32'b11111111111111111011101010111001;
assign LUT_2[3675] = 32'b11111111111111111000100011010010;
assign LUT_2[3676] = 32'b11111111111111110001001111100101;
assign LUT_2[3677] = 32'b11111111111111101110000111111110;
assign LUT_2[3678] = 32'b11111111111111111000001000100001;
assign LUT_2[3679] = 32'b11111111111111110101000000111010;
assign LUT_2[3680] = 32'b11111111111111111111110111111111;
assign LUT_2[3681] = 32'b11111111111111111100110000011000;
assign LUT_2[3682] = 32'b00000000000000000110110000111011;
assign LUT_2[3683] = 32'b00000000000000000011101001010100;
assign LUT_2[3684] = 32'b11111111111111111100010101100111;
assign LUT_2[3685] = 32'b11111111111111111001001110000000;
assign LUT_2[3686] = 32'b00000000000000000011001110100011;
assign LUT_2[3687] = 32'b00000000000000000000000110111100;
assign LUT_2[3688] = 32'b11111111111111111010101001011100;
assign LUT_2[3689] = 32'b11111111111111110111100001110101;
assign LUT_2[3690] = 32'b00000000000000000001100010011000;
assign LUT_2[3691] = 32'b11111111111111111110011010110001;
assign LUT_2[3692] = 32'b11111111111111110111000111000100;
assign LUT_2[3693] = 32'b11111111111111110011111111011101;
assign LUT_2[3694] = 32'b11111111111111111110000000000000;
assign LUT_2[3695] = 32'b11111111111111111010111000011001;
assign LUT_2[3696] = 32'b11111111111111111010011100001001;
assign LUT_2[3697] = 32'b11111111111111110111010100100010;
assign LUT_2[3698] = 32'b00000000000000000001010101000101;
assign LUT_2[3699] = 32'b11111111111111111110001101011110;
assign LUT_2[3700] = 32'b11111111111111110110111001110001;
assign LUT_2[3701] = 32'b11111111111111110011110010001010;
assign LUT_2[3702] = 32'b11111111111111111101110010101101;
assign LUT_2[3703] = 32'b11111111111111111010101011000110;
assign LUT_2[3704] = 32'b11111111111111110101001101100110;
assign LUT_2[3705] = 32'b11111111111111110010000101111111;
assign LUT_2[3706] = 32'b11111111111111111100000110100010;
assign LUT_2[3707] = 32'b11111111111111111000111110111011;
assign LUT_2[3708] = 32'b11111111111111110001101011001110;
assign LUT_2[3709] = 32'b11111111111111101110100011100111;
assign LUT_2[3710] = 32'b11111111111111111000100100001010;
assign LUT_2[3711] = 32'b11111111111111110101011100100011;
assign LUT_2[3712] = 32'b00000000000000001011101000000010;
assign LUT_2[3713] = 32'b00000000000000001000100000011011;
assign LUT_2[3714] = 32'b00000000000000010010100000111110;
assign LUT_2[3715] = 32'b00000000000000001111011001010111;
assign LUT_2[3716] = 32'b00000000000000001000000101101010;
assign LUT_2[3717] = 32'b00000000000000000100111110000011;
assign LUT_2[3718] = 32'b00000000000000001110111110100110;
assign LUT_2[3719] = 32'b00000000000000001011110110111111;
assign LUT_2[3720] = 32'b00000000000000000110011001011111;
assign LUT_2[3721] = 32'b00000000000000000011010001111000;
assign LUT_2[3722] = 32'b00000000000000001101010010011011;
assign LUT_2[3723] = 32'b00000000000000001010001010110100;
assign LUT_2[3724] = 32'b00000000000000000010110111000111;
assign LUT_2[3725] = 32'b11111111111111111111101111100000;
assign LUT_2[3726] = 32'b00000000000000001001110000000011;
assign LUT_2[3727] = 32'b00000000000000000110101000011100;
assign LUT_2[3728] = 32'b00000000000000000110001100001100;
assign LUT_2[3729] = 32'b00000000000000000011000100100101;
assign LUT_2[3730] = 32'b00000000000000001101000101001000;
assign LUT_2[3731] = 32'b00000000000000001001111101100001;
assign LUT_2[3732] = 32'b00000000000000000010101001110100;
assign LUT_2[3733] = 32'b11111111111111111111100010001101;
assign LUT_2[3734] = 32'b00000000000000001001100010110000;
assign LUT_2[3735] = 32'b00000000000000000110011011001001;
assign LUT_2[3736] = 32'b00000000000000000000111101101001;
assign LUT_2[3737] = 32'b11111111111111111101110110000010;
assign LUT_2[3738] = 32'b00000000000000000111110110100101;
assign LUT_2[3739] = 32'b00000000000000000100101110111110;
assign LUT_2[3740] = 32'b11111111111111111101011011010001;
assign LUT_2[3741] = 32'b11111111111111111010010011101010;
assign LUT_2[3742] = 32'b00000000000000000100010100001101;
assign LUT_2[3743] = 32'b00000000000000000001001100100110;
assign LUT_2[3744] = 32'b00000000000000001100000011101011;
assign LUT_2[3745] = 32'b00000000000000001000111100000100;
assign LUT_2[3746] = 32'b00000000000000010010111100100111;
assign LUT_2[3747] = 32'b00000000000000001111110101000000;
assign LUT_2[3748] = 32'b00000000000000001000100001010011;
assign LUT_2[3749] = 32'b00000000000000000101011001101100;
assign LUT_2[3750] = 32'b00000000000000001111011010001111;
assign LUT_2[3751] = 32'b00000000000000001100010010101000;
assign LUT_2[3752] = 32'b00000000000000000110110101001000;
assign LUT_2[3753] = 32'b00000000000000000011101101100001;
assign LUT_2[3754] = 32'b00000000000000001101101110000100;
assign LUT_2[3755] = 32'b00000000000000001010100110011101;
assign LUT_2[3756] = 32'b00000000000000000011010010110000;
assign LUT_2[3757] = 32'b00000000000000000000001011001001;
assign LUT_2[3758] = 32'b00000000000000001010001011101100;
assign LUT_2[3759] = 32'b00000000000000000111000100000101;
assign LUT_2[3760] = 32'b00000000000000000110100111110101;
assign LUT_2[3761] = 32'b00000000000000000011100000001110;
assign LUT_2[3762] = 32'b00000000000000001101100000110001;
assign LUT_2[3763] = 32'b00000000000000001010011001001010;
assign LUT_2[3764] = 32'b00000000000000000011000101011101;
assign LUT_2[3765] = 32'b11111111111111111111111101110110;
assign LUT_2[3766] = 32'b00000000000000001001111110011001;
assign LUT_2[3767] = 32'b00000000000000000110110110110010;
assign LUT_2[3768] = 32'b00000000000000000001011001010010;
assign LUT_2[3769] = 32'b11111111111111111110010001101011;
assign LUT_2[3770] = 32'b00000000000000001000010010001110;
assign LUT_2[3771] = 32'b00000000000000000101001010100111;
assign LUT_2[3772] = 32'b11111111111111111101110110111010;
assign LUT_2[3773] = 32'b11111111111111111010101111010011;
assign LUT_2[3774] = 32'b00000000000000000100101111110110;
assign LUT_2[3775] = 32'b00000000000000000001101000001111;
assign LUT_2[3776] = 32'b00000000000000000011110000100101;
assign LUT_2[3777] = 32'b00000000000000000000101000111110;
assign LUT_2[3778] = 32'b00000000000000001010101001100001;
assign LUT_2[3779] = 32'b00000000000000000111100001111010;
assign LUT_2[3780] = 32'b00000000000000000000001110001101;
assign LUT_2[3781] = 32'b11111111111111111101000110100110;
assign LUT_2[3782] = 32'b00000000000000000111000111001001;
assign LUT_2[3783] = 32'b00000000000000000011111111100010;
assign LUT_2[3784] = 32'b11111111111111111110100010000010;
assign LUT_2[3785] = 32'b11111111111111111011011010011011;
assign LUT_2[3786] = 32'b00000000000000000101011010111110;
assign LUT_2[3787] = 32'b00000000000000000010010011010111;
assign LUT_2[3788] = 32'b11111111111111111010111111101010;
assign LUT_2[3789] = 32'b11111111111111110111111000000011;
assign LUT_2[3790] = 32'b00000000000000000001111000100110;
assign LUT_2[3791] = 32'b11111111111111111110110000111111;
assign LUT_2[3792] = 32'b11111111111111111110010100101111;
assign LUT_2[3793] = 32'b11111111111111111011001101001000;
assign LUT_2[3794] = 32'b00000000000000000101001101101011;
assign LUT_2[3795] = 32'b00000000000000000010000110000100;
assign LUT_2[3796] = 32'b11111111111111111010110010010111;
assign LUT_2[3797] = 32'b11111111111111110111101010110000;
assign LUT_2[3798] = 32'b00000000000000000001101011010011;
assign LUT_2[3799] = 32'b11111111111111111110100011101100;
assign LUT_2[3800] = 32'b11111111111111111001000110001100;
assign LUT_2[3801] = 32'b11111111111111110101111110100101;
assign LUT_2[3802] = 32'b11111111111111111111111111001000;
assign LUT_2[3803] = 32'b11111111111111111100110111100001;
assign LUT_2[3804] = 32'b11111111111111110101100011110100;
assign LUT_2[3805] = 32'b11111111111111110010011100001101;
assign LUT_2[3806] = 32'b11111111111111111100011100110000;
assign LUT_2[3807] = 32'b11111111111111111001010101001001;
assign LUT_2[3808] = 32'b00000000000000000100001100001110;
assign LUT_2[3809] = 32'b00000000000000000001000100100111;
assign LUT_2[3810] = 32'b00000000000000001011000101001010;
assign LUT_2[3811] = 32'b00000000000000000111111101100011;
assign LUT_2[3812] = 32'b00000000000000000000101001110110;
assign LUT_2[3813] = 32'b11111111111111111101100010001111;
assign LUT_2[3814] = 32'b00000000000000000111100010110010;
assign LUT_2[3815] = 32'b00000000000000000100011011001011;
assign LUT_2[3816] = 32'b11111111111111111110111101101011;
assign LUT_2[3817] = 32'b11111111111111111011110110000100;
assign LUT_2[3818] = 32'b00000000000000000101110110100111;
assign LUT_2[3819] = 32'b00000000000000000010101111000000;
assign LUT_2[3820] = 32'b11111111111111111011011011010011;
assign LUT_2[3821] = 32'b11111111111111111000010011101100;
assign LUT_2[3822] = 32'b00000000000000000010010100001111;
assign LUT_2[3823] = 32'b11111111111111111111001100101000;
assign LUT_2[3824] = 32'b11111111111111111110110000011000;
assign LUT_2[3825] = 32'b11111111111111111011101000110001;
assign LUT_2[3826] = 32'b00000000000000000101101001010100;
assign LUT_2[3827] = 32'b00000000000000000010100001101101;
assign LUT_2[3828] = 32'b11111111111111111011001110000000;
assign LUT_2[3829] = 32'b11111111111111111000000110011001;
assign LUT_2[3830] = 32'b00000000000000000010000110111100;
assign LUT_2[3831] = 32'b11111111111111111110111111010101;
assign LUT_2[3832] = 32'b11111111111111111001100001110101;
assign LUT_2[3833] = 32'b11111111111111110110011010001110;
assign LUT_2[3834] = 32'b00000000000000000000011010110001;
assign LUT_2[3835] = 32'b11111111111111111101010011001010;
assign LUT_2[3836] = 32'b11111111111111110101111111011101;
assign LUT_2[3837] = 32'b11111111111111110010110111110110;
assign LUT_2[3838] = 32'b11111111111111111100111000011001;
assign LUT_2[3839] = 32'b11111111111111111001110000110010;
assign LUT_2[3840] = 32'b00000000000000001011010010011001;
assign LUT_2[3841] = 32'b00000000000000001000001010110010;
assign LUT_2[3842] = 32'b00000000000000010010001011010101;
assign LUT_2[3843] = 32'b00000000000000001111000011101110;
assign LUT_2[3844] = 32'b00000000000000000111110000000001;
assign LUT_2[3845] = 32'b00000000000000000100101000011010;
assign LUT_2[3846] = 32'b00000000000000001110101000111101;
assign LUT_2[3847] = 32'b00000000000000001011100001010110;
assign LUT_2[3848] = 32'b00000000000000000110000011110110;
assign LUT_2[3849] = 32'b00000000000000000010111100001111;
assign LUT_2[3850] = 32'b00000000000000001100111100110010;
assign LUT_2[3851] = 32'b00000000000000001001110101001011;
assign LUT_2[3852] = 32'b00000000000000000010100001011110;
assign LUT_2[3853] = 32'b11111111111111111111011001110111;
assign LUT_2[3854] = 32'b00000000000000001001011010011010;
assign LUT_2[3855] = 32'b00000000000000000110010010110011;
assign LUT_2[3856] = 32'b00000000000000000101110110100011;
assign LUT_2[3857] = 32'b00000000000000000010101110111100;
assign LUT_2[3858] = 32'b00000000000000001100101111011111;
assign LUT_2[3859] = 32'b00000000000000001001100111111000;
assign LUT_2[3860] = 32'b00000000000000000010010100001011;
assign LUT_2[3861] = 32'b11111111111111111111001100100100;
assign LUT_2[3862] = 32'b00000000000000001001001101000111;
assign LUT_2[3863] = 32'b00000000000000000110000101100000;
assign LUT_2[3864] = 32'b00000000000000000000101000000000;
assign LUT_2[3865] = 32'b11111111111111111101100000011001;
assign LUT_2[3866] = 32'b00000000000000000111100000111100;
assign LUT_2[3867] = 32'b00000000000000000100011001010101;
assign LUT_2[3868] = 32'b11111111111111111101000101101000;
assign LUT_2[3869] = 32'b11111111111111111001111110000001;
assign LUT_2[3870] = 32'b00000000000000000011111110100100;
assign LUT_2[3871] = 32'b00000000000000000000110110111101;
assign LUT_2[3872] = 32'b00000000000000001011101110000010;
assign LUT_2[3873] = 32'b00000000000000001000100110011011;
assign LUT_2[3874] = 32'b00000000000000010010100110111110;
assign LUT_2[3875] = 32'b00000000000000001111011111010111;
assign LUT_2[3876] = 32'b00000000000000001000001011101010;
assign LUT_2[3877] = 32'b00000000000000000101000100000011;
assign LUT_2[3878] = 32'b00000000000000001111000100100110;
assign LUT_2[3879] = 32'b00000000000000001011111100111111;
assign LUT_2[3880] = 32'b00000000000000000110011111011111;
assign LUT_2[3881] = 32'b00000000000000000011010111111000;
assign LUT_2[3882] = 32'b00000000000000001101011000011011;
assign LUT_2[3883] = 32'b00000000000000001010010000110100;
assign LUT_2[3884] = 32'b00000000000000000010111101000111;
assign LUT_2[3885] = 32'b11111111111111111111110101100000;
assign LUT_2[3886] = 32'b00000000000000001001110110000011;
assign LUT_2[3887] = 32'b00000000000000000110101110011100;
assign LUT_2[3888] = 32'b00000000000000000110010010001100;
assign LUT_2[3889] = 32'b00000000000000000011001010100101;
assign LUT_2[3890] = 32'b00000000000000001101001011001000;
assign LUT_2[3891] = 32'b00000000000000001010000011100001;
assign LUT_2[3892] = 32'b00000000000000000010101111110100;
assign LUT_2[3893] = 32'b11111111111111111111101000001101;
assign LUT_2[3894] = 32'b00000000000000001001101000110000;
assign LUT_2[3895] = 32'b00000000000000000110100001001001;
assign LUT_2[3896] = 32'b00000000000000000001000011101001;
assign LUT_2[3897] = 32'b11111111111111111101111100000010;
assign LUT_2[3898] = 32'b00000000000000000111111100100101;
assign LUT_2[3899] = 32'b00000000000000000100110100111110;
assign LUT_2[3900] = 32'b11111111111111111101100001010001;
assign LUT_2[3901] = 32'b11111111111111111010011001101010;
assign LUT_2[3902] = 32'b00000000000000000100011010001101;
assign LUT_2[3903] = 32'b00000000000000000001010010100110;
assign LUT_2[3904] = 32'b00000000000000000011011010111100;
assign LUT_2[3905] = 32'b00000000000000000000010011010101;
assign LUT_2[3906] = 32'b00000000000000001010010011111000;
assign LUT_2[3907] = 32'b00000000000000000111001100010001;
assign LUT_2[3908] = 32'b11111111111111111111111000100100;
assign LUT_2[3909] = 32'b11111111111111111100110000111101;
assign LUT_2[3910] = 32'b00000000000000000110110001100000;
assign LUT_2[3911] = 32'b00000000000000000011101001111001;
assign LUT_2[3912] = 32'b11111111111111111110001100011001;
assign LUT_2[3913] = 32'b11111111111111111011000100110010;
assign LUT_2[3914] = 32'b00000000000000000101000101010101;
assign LUT_2[3915] = 32'b00000000000000000001111101101110;
assign LUT_2[3916] = 32'b11111111111111111010101010000001;
assign LUT_2[3917] = 32'b11111111111111110111100010011010;
assign LUT_2[3918] = 32'b00000000000000000001100010111101;
assign LUT_2[3919] = 32'b11111111111111111110011011010110;
assign LUT_2[3920] = 32'b11111111111111111101111111000110;
assign LUT_2[3921] = 32'b11111111111111111010110111011111;
assign LUT_2[3922] = 32'b00000000000000000100111000000010;
assign LUT_2[3923] = 32'b00000000000000000001110000011011;
assign LUT_2[3924] = 32'b11111111111111111010011100101110;
assign LUT_2[3925] = 32'b11111111111111110111010101000111;
assign LUT_2[3926] = 32'b00000000000000000001010101101010;
assign LUT_2[3927] = 32'b11111111111111111110001110000011;
assign LUT_2[3928] = 32'b11111111111111111000110000100011;
assign LUT_2[3929] = 32'b11111111111111110101101000111100;
assign LUT_2[3930] = 32'b11111111111111111111101001011111;
assign LUT_2[3931] = 32'b11111111111111111100100001111000;
assign LUT_2[3932] = 32'b11111111111111110101001110001011;
assign LUT_2[3933] = 32'b11111111111111110010000110100100;
assign LUT_2[3934] = 32'b11111111111111111100000111000111;
assign LUT_2[3935] = 32'b11111111111111111000111111100000;
assign LUT_2[3936] = 32'b00000000000000000011110110100101;
assign LUT_2[3937] = 32'b00000000000000000000101110111110;
assign LUT_2[3938] = 32'b00000000000000001010101111100001;
assign LUT_2[3939] = 32'b00000000000000000111100111111010;
assign LUT_2[3940] = 32'b00000000000000000000010100001101;
assign LUT_2[3941] = 32'b11111111111111111101001100100110;
assign LUT_2[3942] = 32'b00000000000000000111001101001001;
assign LUT_2[3943] = 32'b00000000000000000100000101100010;
assign LUT_2[3944] = 32'b11111111111111111110101000000010;
assign LUT_2[3945] = 32'b11111111111111111011100000011011;
assign LUT_2[3946] = 32'b00000000000000000101100000111110;
assign LUT_2[3947] = 32'b00000000000000000010011001010111;
assign LUT_2[3948] = 32'b11111111111111111011000101101010;
assign LUT_2[3949] = 32'b11111111111111110111111110000011;
assign LUT_2[3950] = 32'b00000000000000000001111110100110;
assign LUT_2[3951] = 32'b11111111111111111110110110111111;
assign LUT_2[3952] = 32'b11111111111111111110011010101111;
assign LUT_2[3953] = 32'b11111111111111111011010011001000;
assign LUT_2[3954] = 32'b00000000000000000101010011101011;
assign LUT_2[3955] = 32'b00000000000000000010001100000100;
assign LUT_2[3956] = 32'b11111111111111111010111000010111;
assign LUT_2[3957] = 32'b11111111111111110111110000110000;
assign LUT_2[3958] = 32'b00000000000000000001110001010011;
assign LUT_2[3959] = 32'b11111111111111111110101001101100;
assign LUT_2[3960] = 32'b11111111111111111001001100001100;
assign LUT_2[3961] = 32'b11111111111111110110000100100101;
assign LUT_2[3962] = 32'b00000000000000000000000101001000;
assign LUT_2[3963] = 32'b11111111111111111100111101100001;
assign LUT_2[3964] = 32'b11111111111111110101101001110100;
assign LUT_2[3965] = 32'b11111111111111110010100010001101;
assign LUT_2[3966] = 32'b11111111111111111100100010110000;
assign LUT_2[3967] = 32'b11111111111111111001011011001001;
assign LUT_2[3968] = 32'b00000000000000001111100110101000;
assign LUT_2[3969] = 32'b00000000000000001100011111000001;
assign LUT_2[3970] = 32'b00000000000000010110011111100100;
assign LUT_2[3971] = 32'b00000000000000010011010111111101;
assign LUT_2[3972] = 32'b00000000000000001100000100010000;
assign LUT_2[3973] = 32'b00000000000000001000111100101001;
assign LUT_2[3974] = 32'b00000000000000010010111101001100;
assign LUT_2[3975] = 32'b00000000000000001111110101100101;
assign LUT_2[3976] = 32'b00000000000000001010011000000101;
assign LUT_2[3977] = 32'b00000000000000000111010000011110;
assign LUT_2[3978] = 32'b00000000000000010001010001000001;
assign LUT_2[3979] = 32'b00000000000000001110001001011010;
assign LUT_2[3980] = 32'b00000000000000000110110101101101;
assign LUT_2[3981] = 32'b00000000000000000011101110000110;
assign LUT_2[3982] = 32'b00000000000000001101101110101001;
assign LUT_2[3983] = 32'b00000000000000001010100111000010;
assign LUT_2[3984] = 32'b00000000000000001010001010110010;
assign LUT_2[3985] = 32'b00000000000000000111000011001011;
assign LUT_2[3986] = 32'b00000000000000010001000011101110;
assign LUT_2[3987] = 32'b00000000000000001101111100000111;
assign LUT_2[3988] = 32'b00000000000000000110101000011010;
assign LUT_2[3989] = 32'b00000000000000000011100000110011;
assign LUT_2[3990] = 32'b00000000000000001101100001010110;
assign LUT_2[3991] = 32'b00000000000000001010011001101111;
assign LUT_2[3992] = 32'b00000000000000000100111100001111;
assign LUT_2[3993] = 32'b00000000000000000001110100101000;
assign LUT_2[3994] = 32'b00000000000000001011110101001011;
assign LUT_2[3995] = 32'b00000000000000001000101101100100;
assign LUT_2[3996] = 32'b00000000000000000001011001110111;
assign LUT_2[3997] = 32'b11111111111111111110010010010000;
assign LUT_2[3998] = 32'b00000000000000001000010010110011;
assign LUT_2[3999] = 32'b00000000000000000101001011001100;
assign LUT_2[4000] = 32'b00000000000000010000000010010001;
assign LUT_2[4001] = 32'b00000000000000001100111010101010;
assign LUT_2[4002] = 32'b00000000000000010110111011001101;
assign LUT_2[4003] = 32'b00000000000000010011110011100110;
assign LUT_2[4004] = 32'b00000000000000001100011111111001;
assign LUT_2[4005] = 32'b00000000000000001001011000010010;
assign LUT_2[4006] = 32'b00000000000000010011011000110101;
assign LUT_2[4007] = 32'b00000000000000010000010001001110;
assign LUT_2[4008] = 32'b00000000000000001010110011101110;
assign LUT_2[4009] = 32'b00000000000000000111101100000111;
assign LUT_2[4010] = 32'b00000000000000010001101100101010;
assign LUT_2[4011] = 32'b00000000000000001110100101000011;
assign LUT_2[4012] = 32'b00000000000000000111010001010110;
assign LUT_2[4013] = 32'b00000000000000000100001001101111;
assign LUT_2[4014] = 32'b00000000000000001110001010010010;
assign LUT_2[4015] = 32'b00000000000000001011000010101011;
assign LUT_2[4016] = 32'b00000000000000001010100110011011;
assign LUT_2[4017] = 32'b00000000000000000111011110110100;
assign LUT_2[4018] = 32'b00000000000000010001011111010111;
assign LUT_2[4019] = 32'b00000000000000001110010111110000;
assign LUT_2[4020] = 32'b00000000000000000111000100000011;
assign LUT_2[4021] = 32'b00000000000000000011111100011100;
assign LUT_2[4022] = 32'b00000000000000001101111100111111;
assign LUT_2[4023] = 32'b00000000000000001010110101011000;
assign LUT_2[4024] = 32'b00000000000000000101010111111000;
assign LUT_2[4025] = 32'b00000000000000000010010000010001;
assign LUT_2[4026] = 32'b00000000000000001100010000110100;
assign LUT_2[4027] = 32'b00000000000000001001001001001101;
assign LUT_2[4028] = 32'b00000000000000000001110101100000;
assign LUT_2[4029] = 32'b11111111111111111110101101111001;
assign LUT_2[4030] = 32'b00000000000000001000101110011100;
assign LUT_2[4031] = 32'b00000000000000000101100110110101;
assign LUT_2[4032] = 32'b00000000000000000111101111001011;
assign LUT_2[4033] = 32'b00000000000000000100100111100100;
assign LUT_2[4034] = 32'b00000000000000001110101000000111;
assign LUT_2[4035] = 32'b00000000000000001011100000100000;
assign LUT_2[4036] = 32'b00000000000000000100001100110011;
assign LUT_2[4037] = 32'b00000000000000000001000101001100;
assign LUT_2[4038] = 32'b00000000000000001011000101101111;
assign LUT_2[4039] = 32'b00000000000000000111111110001000;
assign LUT_2[4040] = 32'b00000000000000000010100000101000;
assign LUT_2[4041] = 32'b11111111111111111111011001000001;
assign LUT_2[4042] = 32'b00000000000000001001011001100100;
assign LUT_2[4043] = 32'b00000000000000000110010001111101;
assign LUT_2[4044] = 32'b11111111111111111110111110010000;
assign LUT_2[4045] = 32'b11111111111111111011110110101001;
assign LUT_2[4046] = 32'b00000000000000000101110111001100;
assign LUT_2[4047] = 32'b00000000000000000010101111100101;
assign LUT_2[4048] = 32'b00000000000000000010010011010101;
assign LUT_2[4049] = 32'b11111111111111111111001011101110;
assign LUT_2[4050] = 32'b00000000000000001001001100010001;
assign LUT_2[4051] = 32'b00000000000000000110000100101010;
assign LUT_2[4052] = 32'b11111111111111111110110000111101;
assign LUT_2[4053] = 32'b11111111111111111011101001010110;
assign LUT_2[4054] = 32'b00000000000000000101101001111001;
assign LUT_2[4055] = 32'b00000000000000000010100010010010;
assign LUT_2[4056] = 32'b11111111111111111101000100110010;
assign LUT_2[4057] = 32'b11111111111111111001111101001011;
assign LUT_2[4058] = 32'b00000000000000000011111101101110;
assign LUT_2[4059] = 32'b00000000000000000000110110000111;
assign LUT_2[4060] = 32'b11111111111111111001100010011010;
assign LUT_2[4061] = 32'b11111111111111110110011010110011;
assign LUT_2[4062] = 32'b00000000000000000000011011010110;
assign LUT_2[4063] = 32'b11111111111111111101010011101111;
assign LUT_2[4064] = 32'b00000000000000001000001010110100;
assign LUT_2[4065] = 32'b00000000000000000101000011001101;
assign LUT_2[4066] = 32'b00000000000000001111000011110000;
assign LUT_2[4067] = 32'b00000000000000001011111100001001;
assign LUT_2[4068] = 32'b00000000000000000100101000011100;
assign LUT_2[4069] = 32'b00000000000000000001100000110101;
assign LUT_2[4070] = 32'b00000000000000001011100001011000;
assign LUT_2[4071] = 32'b00000000000000001000011001110001;
assign LUT_2[4072] = 32'b00000000000000000010111100010001;
assign LUT_2[4073] = 32'b11111111111111111111110100101010;
assign LUT_2[4074] = 32'b00000000000000001001110101001101;
assign LUT_2[4075] = 32'b00000000000000000110101101100110;
assign LUT_2[4076] = 32'b11111111111111111111011001111001;
assign LUT_2[4077] = 32'b11111111111111111100010010010010;
assign LUT_2[4078] = 32'b00000000000000000110010010110101;
assign LUT_2[4079] = 32'b00000000000000000011001011001110;
assign LUT_2[4080] = 32'b00000000000000000010101110111110;
assign LUT_2[4081] = 32'b11111111111111111111100111010111;
assign LUT_2[4082] = 32'b00000000000000001001100111111010;
assign LUT_2[4083] = 32'b00000000000000000110100000010011;
assign LUT_2[4084] = 32'b11111111111111111111001100100110;
assign LUT_2[4085] = 32'b11111111111111111100000100111111;
assign LUT_2[4086] = 32'b00000000000000000110000101100010;
assign LUT_2[4087] = 32'b00000000000000000010111101111011;
assign LUT_2[4088] = 32'b11111111111111111101100000011011;
assign LUT_2[4089] = 32'b11111111111111111010011000110100;
assign LUT_2[4090] = 32'b00000000000000000100011001010111;
assign LUT_2[4091] = 32'b00000000000000000001010001110000;
assign LUT_2[4092] = 32'b11111111111111111001111110000011;
assign LUT_2[4093] = 32'b11111111111111110110110110011100;
assign LUT_2[4094] = 32'b00000000000000000000110110111111;
assign LUT_2[4095] = 32'b11111111111111111101101111011000;
assign LUT_2[4096] = 32'b11111111111111111111000100001011;
assign LUT_2[4097] = 32'b11111111111111111011111100100100;
assign LUT_2[4098] = 32'b00000000000000000101111101000111;
assign LUT_2[4099] = 32'b00000000000000000010110101100000;
assign LUT_2[4100] = 32'b11111111111111111011100001110011;
assign LUT_2[4101] = 32'b11111111111111111000011010001100;
assign LUT_2[4102] = 32'b00000000000000000010011010101111;
assign LUT_2[4103] = 32'b11111111111111111111010011001000;
assign LUT_2[4104] = 32'b11111111111111111001110101101000;
assign LUT_2[4105] = 32'b11111111111111110110101110000001;
assign LUT_2[4106] = 32'b00000000000000000000101110100100;
assign LUT_2[4107] = 32'b11111111111111111101100110111101;
assign LUT_2[4108] = 32'b11111111111111110110010011010000;
assign LUT_2[4109] = 32'b11111111111111110011001011101001;
assign LUT_2[4110] = 32'b11111111111111111101001100001100;
assign LUT_2[4111] = 32'b11111111111111111010000100100101;
assign LUT_2[4112] = 32'b11111111111111111001101000010101;
assign LUT_2[4113] = 32'b11111111111111110110100000101110;
assign LUT_2[4114] = 32'b00000000000000000000100001010001;
assign LUT_2[4115] = 32'b11111111111111111101011001101010;
assign LUT_2[4116] = 32'b11111111111111110110000101111101;
assign LUT_2[4117] = 32'b11111111111111110010111110010110;
assign LUT_2[4118] = 32'b11111111111111111100111110111001;
assign LUT_2[4119] = 32'b11111111111111111001110111010010;
assign LUT_2[4120] = 32'b11111111111111110100011001110010;
assign LUT_2[4121] = 32'b11111111111111110001010010001011;
assign LUT_2[4122] = 32'b11111111111111111011010010101110;
assign LUT_2[4123] = 32'b11111111111111111000001011000111;
assign LUT_2[4124] = 32'b11111111111111110000110111011010;
assign LUT_2[4125] = 32'b11111111111111101101101111110011;
assign LUT_2[4126] = 32'b11111111111111110111110000010110;
assign LUT_2[4127] = 32'b11111111111111110100101000101111;
assign LUT_2[4128] = 32'b11111111111111111111011111110100;
assign LUT_2[4129] = 32'b11111111111111111100011000001101;
assign LUT_2[4130] = 32'b00000000000000000110011000110000;
assign LUT_2[4131] = 32'b00000000000000000011010001001001;
assign LUT_2[4132] = 32'b11111111111111111011111101011100;
assign LUT_2[4133] = 32'b11111111111111111000110101110101;
assign LUT_2[4134] = 32'b00000000000000000010110110011000;
assign LUT_2[4135] = 32'b11111111111111111111101110110001;
assign LUT_2[4136] = 32'b11111111111111111010010001010001;
assign LUT_2[4137] = 32'b11111111111111110111001001101010;
assign LUT_2[4138] = 32'b00000000000000000001001010001101;
assign LUT_2[4139] = 32'b11111111111111111110000010100110;
assign LUT_2[4140] = 32'b11111111111111110110101110111001;
assign LUT_2[4141] = 32'b11111111111111110011100111010010;
assign LUT_2[4142] = 32'b11111111111111111101100111110101;
assign LUT_2[4143] = 32'b11111111111111111010100000001110;
assign LUT_2[4144] = 32'b11111111111111111010000011111110;
assign LUT_2[4145] = 32'b11111111111111110110111100010111;
assign LUT_2[4146] = 32'b00000000000000000000111100111010;
assign LUT_2[4147] = 32'b11111111111111111101110101010011;
assign LUT_2[4148] = 32'b11111111111111110110100001100110;
assign LUT_2[4149] = 32'b11111111111111110011011001111111;
assign LUT_2[4150] = 32'b11111111111111111101011010100010;
assign LUT_2[4151] = 32'b11111111111111111010010010111011;
assign LUT_2[4152] = 32'b11111111111111110100110101011011;
assign LUT_2[4153] = 32'b11111111111111110001101101110100;
assign LUT_2[4154] = 32'b11111111111111111011101110010111;
assign LUT_2[4155] = 32'b11111111111111111000100110110000;
assign LUT_2[4156] = 32'b11111111111111110001010011000011;
assign LUT_2[4157] = 32'b11111111111111101110001011011100;
assign LUT_2[4158] = 32'b11111111111111111000001011111111;
assign LUT_2[4159] = 32'b11111111111111110101000100011000;
assign LUT_2[4160] = 32'b11111111111111110111001100101110;
assign LUT_2[4161] = 32'b11111111111111110100000101000111;
assign LUT_2[4162] = 32'b11111111111111111110000101101010;
assign LUT_2[4163] = 32'b11111111111111111010111110000011;
assign LUT_2[4164] = 32'b11111111111111110011101010010110;
assign LUT_2[4165] = 32'b11111111111111110000100010101111;
assign LUT_2[4166] = 32'b11111111111111111010100011010010;
assign LUT_2[4167] = 32'b11111111111111110111011011101011;
assign LUT_2[4168] = 32'b11111111111111110001111110001011;
assign LUT_2[4169] = 32'b11111111111111101110110110100100;
assign LUT_2[4170] = 32'b11111111111111111000110111000111;
assign LUT_2[4171] = 32'b11111111111111110101101111100000;
assign LUT_2[4172] = 32'b11111111111111101110011011110011;
assign LUT_2[4173] = 32'b11111111111111101011010100001100;
assign LUT_2[4174] = 32'b11111111111111110101010100101111;
assign LUT_2[4175] = 32'b11111111111111110010001101001000;
assign LUT_2[4176] = 32'b11111111111111110001110000111000;
assign LUT_2[4177] = 32'b11111111111111101110101001010001;
assign LUT_2[4178] = 32'b11111111111111111000101001110100;
assign LUT_2[4179] = 32'b11111111111111110101100010001101;
assign LUT_2[4180] = 32'b11111111111111101110001110100000;
assign LUT_2[4181] = 32'b11111111111111101011000110111001;
assign LUT_2[4182] = 32'b11111111111111110101000111011100;
assign LUT_2[4183] = 32'b11111111111111110001111111110101;
assign LUT_2[4184] = 32'b11111111111111101100100010010101;
assign LUT_2[4185] = 32'b11111111111111101001011010101110;
assign LUT_2[4186] = 32'b11111111111111110011011011010001;
assign LUT_2[4187] = 32'b11111111111111110000010011101010;
assign LUT_2[4188] = 32'b11111111111111101000111111111101;
assign LUT_2[4189] = 32'b11111111111111100101111000010110;
assign LUT_2[4190] = 32'b11111111111111101111111000111001;
assign LUT_2[4191] = 32'b11111111111111101100110001010010;
assign LUT_2[4192] = 32'b11111111111111110111101000010111;
assign LUT_2[4193] = 32'b11111111111111110100100000110000;
assign LUT_2[4194] = 32'b11111111111111111110100001010011;
assign LUT_2[4195] = 32'b11111111111111111011011001101100;
assign LUT_2[4196] = 32'b11111111111111110100000101111111;
assign LUT_2[4197] = 32'b11111111111111110000111110011000;
assign LUT_2[4198] = 32'b11111111111111111010111110111011;
assign LUT_2[4199] = 32'b11111111111111110111110111010100;
assign LUT_2[4200] = 32'b11111111111111110010011001110100;
assign LUT_2[4201] = 32'b11111111111111101111010010001101;
assign LUT_2[4202] = 32'b11111111111111111001010010110000;
assign LUT_2[4203] = 32'b11111111111111110110001011001001;
assign LUT_2[4204] = 32'b11111111111111101110110111011100;
assign LUT_2[4205] = 32'b11111111111111101011101111110101;
assign LUT_2[4206] = 32'b11111111111111110101110000011000;
assign LUT_2[4207] = 32'b11111111111111110010101000110001;
assign LUT_2[4208] = 32'b11111111111111110010001100100001;
assign LUT_2[4209] = 32'b11111111111111101111000100111010;
assign LUT_2[4210] = 32'b11111111111111111001000101011101;
assign LUT_2[4211] = 32'b11111111111111110101111101110110;
assign LUT_2[4212] = 32'b11111111111111101110101010001001;
assign LUT_2[4213] = 32'b11111111111111101011100010100010;
assign LUT_2[4214] = 32'b11111111111111110101100011000101;
assign LUT_2[4215] = 32'b11111111111111110010011011011110;
assign LUT_2[4216] = 32'b11111111111111101100111101111110;
assign LUT_2[4217] = 32'b11111111111111101001110110010111;
assign LUT_2[4218] = 32'b11111111111111110011110110111010;
assign LUT_2[4219] = 32'b11111111111111110000101111010011;
assign LUT_2[4220] = 32'b11111111111111101001011011100110;
assign LUT_2[4221] = 32'b11111111111111100110010011111111;
assign LUT_2[4222] = 32'b11111111111111110000010100100010;
assign LUT_2[4223] = 32'b11111111111111101101001100111011;
assign LUT_2[4224] = 32'b00000000000000000011011000011010;
assign LUT_2[4225] = 32'b00000000000000000000010000110011;
assign LUT_2[4226] = 32'b00000000000000001010010001010110;
assign LUT_2[4227] = 32'b00000000000000000111001001101111;
assign LUT_2[4228] = 32'b11111111111111111111110110000010;
assign LUT_2[4229] = 32'b11111111111111111100101110011011;
assign LUT_2[4230] = 32'b00000000000000000110101110111110;
assign LUT_2[4231] = 32'b00000000000000000011100111010111;
assign LUT_2[4232] = 32'b11111111111111111110001001110111;
assign LUT_2[4233] = 32'b11111111111111111011000010010000;
assign LUT_2[4234] = 32'b00000000000000000101000010110011;
assign LUT_2[4235] = 32'b00000000000000000001111011001100;
assign LUT_2[4236] = 32'b11111111111111111010100111011111;
assign LUT_2[4237] = 32'b11111111111111110111011111111000;
assign LUT_2[4238] = 32'b00000000000000000001100000011011;
assign LUT_2[4239] = 32'b11111111111111111110011000110100;
assign LUT_2[4240] = 32'b11111111111111111101111100100100;
assign LUT_2[4241] = 32'b11111111111111111010110100111101;
assign LUT_2[4242] = 32'b00000000000000000100110101100000;
assign LUT_2[4243] = 32'b00000000000000000001101101111001;
assign LUT_2[4244] = 32'b11111111111111111010011010001100;
assign LUT_2[4245] = 32'b11111111111111110111010010100101;
assign LUT_2[4246] = 32'b00000000000000000001010011001000;
assign LUT_2[4247] = 32'b11111111111111111110001011100001;
assign LUT_2[4248] = 32'b11111111111111111000101110000001;
assign LUT_2[4249] = 32'b11111111111111110101100110011010;
assign LUT_2[4250] = 32'b11111111111111111111100110111101;
assign LUT_2[4251] = 32'b11111111111111111100011111010110;
assign LUT_2[4252] = 32'b11111111111111110101001011101001;
assign LUT_2[4253] = 32'b11111111111111110010000100000010;
assign LUT_2[4254] = 32'b11111111111111111100000100100101;
assign LUT_2[4255] = 32'b11111111111111111000111100111110;
assign LUT_2[4256] = 32'b00000000000000000011110100000011;
assign LUT_2[4257] = 32'b00000000000000000000101100011100;
assign LUT_2[4258] = 32'b00000000000000001010101100111111;
assign LUT_2[4259] = 32'b00000000000000000111100101011000;
assign LUT_2[4260] = 32'b00000000000000000000010001101011;
assign LUT_2[4261] = 32'b11111111111111111101001010000100;
assign LUT_2[4262] = 32'b00000000000000000111001010100111;
assign LUT_2[4263] = 32'b00000000000000000100000011000000;
assign LUT_2[4264] = 32'b11111111111111111110100101100000;
assign LUT_2[4265] = 32'b11111111111111111011011101111001;
assign LUT_2[4266] = 32'b00000000000000000101011110011100;
assign LUT_2[4267] = 32'b00000000000000000010010110110101;
assign LUT_2[4268] = 32'b11111111111111111011000011001000;
assign LUT_2[4269] = 32'b11111111111111110111111011100001;
assign LUT_2[4270] = 32'b00000000000000000001111100000100;
assign LUT_2[4271] = 32'b11111111111111111110110100011101;
assign LUT_2[4272] = 32'b11111111111111111110011000001101;
assign LUT_2[4273] = 32'b11111111111111111011010000100110;
assign LUT_2[4274] = 32'b00000000000000000101010001001001;
assign LUT_2[4275] = 32'b00000000000000000010001001100010;
assign LUT_2[4276] = 32'b11111111111111111010110101110101;
assign LUT_2[4277] = 32'b11111111111111110111101110001110;
assign LUT_2[4278] = 32'b00000000000000000001101110110001;
assign LUT_2[4279] = 32'b11111111111111111110100111001010;
assign LUT_2[4280] = 32'b11111111111111111001001001101010;
assign LUT_2[4281] = 32'b11111111111111110110000010000011;
assign LUT_2[4282] = 32'b00000000000000000000000010100110;
assign LUT_2[4283] = 32'b11111111111111111100111010111111;
assign LUT_2[4284] = 32'b11111111111111110101100111010010;
assign LUT_2[4285] = 32'b11111111111111110010011111101011;
assign LUT_2[4286] = 32'b11111111111111111100100000001110;
assign LUT_2[4287] = 32'b11111111111111111001011000100111;
assign LUT_2[4288] = 32'b11111111111111111011100000111101;
assign LUT_2[4289] = 32'b11111111111111111000011001010110;
assign LUT_2[4290] = 32'b00000000000000000010011001111001;
assign LUT_2[4291] = 32'b11111111111111111111010010010010;
assign LUT_2[4292] = 32'b11111111111111110111111110100101;
assign LUT_2[4293] = 32'b11111111111111110100110110111110;
assign LUT_2[4294] = 32'b11111111111111111110110111100001;
assign LUT_2[4295] = 32'b11111111111111111011101111111010;
assign LUT_2[4296] = 32'b11111111111111110110010010011010;
assign LUT_2[4297] = 32'b11111111111111110011001010110011;
assign LUT_2[4298] = 32'b11111111111111111101001011010110;
assign LUT_2[4299] = 32'b11111111111111111010000011101111;
assign LUT_2[4300] = 32'b11111111111111110010110000000010;
assign LUT_2[4301] = 32'b11111111111111101111101000011011;
assign LUT_2[4302] = 32'b11111111111111111001101000111110;
assign LUT_2[4303] = 32'b11111111111111110110100001010111;
assign LUT_2[4304] = 32'b11111111111111110110000101000111;
assign LUT_2[4305] = 32'b11111111111111110010111101100000;
assign LUT_2[4306] = 32'b11111111111111111100111110000011;
assign LUT_2[4307] = 32'b11111111111111111001110110011100;
assign LUT_2[4308] = 32'b11111111111111110010100010101111;
assign LUT_2[4309] = 32'b11111111111111101111011011001000;
assign LUT_2[4310] = 32'b11111111111111111001011011101011;
assign LUT_2[4311] = 32'b11111111111111110110010100000100;
assign LUT_2[4312] = 32'b11111111111111110000110110100100;
assign LUT_2[4313] = 32'b11111111111111101101101110111101;
assign LUT_2[4314] = 32'b11111111111111110111101111100000;
assign LUT_2[4315] = 32'b11111111111111110100100111111001;
assign LUT_2[4316] = 32'b11111111111111101101010100001100;
assign LUT_2[4317] = 32'b11111111111111101010001100100101;
assign LUT_2[4318] = 32'b11111111111111110100001101001000;
assign LUT_2[4319] = 32'b11111111111111110001000101100001;
assign LUT_2[4320] = 32'b11111111111111111011111100100110;
assign LUT_2[4321] = 32'b11111111111111111000110100111111;
assign LUT_2[4322] = 32'b00000000000000000010110101100010;
assign LUT_2[4323] = 32'b11111111111111111111101101111011;
assign LUT_2[4324] = 32'b11111111111111111000011010001110;
assign LUT_2[4325] = 32'b11111111111111110101010010100111;
assign LUT_2[4326] = 32'b11111111111111111111010011001010;
assign LUT_2[4327] = 32'b11111111111111111100001011100011;
assign LUT_2[4328] = 32'b11111111111111110110101110000011;
assign LUT_2[4329] = 32'b11111111111111110011100110011100;
assign LUT_2[4330] = 32'b11111111111111111101100110111111;
assign LUT_2[4331] = 32'b11111111111111111010011111011000;
assign LUT_2[4332] = 32'b11111111111111110011001011101011;
assign LUT_2[4333] = 32'b11111111111111110000000100000100;
assign LUT_2[4334] = 32'b11111111111111111010000100100111;
assign LUT_2[4335] = 32'b11111111111111110110111101000000;
assign LUT_2[4336] = 32'b11111111111111110110100000110000;
assign LUT_2[4337] = 32'b11111111111111110011011001001001;
assign LUT_2[4338] = 32'b11111111111111111101011001101100;
assign LUT_2[4339] = 32'b11111111111111111010010010000101;
assign LUT_2[4340] = 32'b11111111111111110010111110011000;
assign LUT_2[4341] = 32'b11111111111111101111110110110001;
assign LUT_2[4342] = 32'b11111111111111111001110111010100;
assign LUT_2[4343] = 32'b11111111111111110110101111101101;
assign LUT_2[4344] = 32'b11111111111111110001010010001101;
assign LUT_2[4345] = 32'b11111111111111101110001010100110;
assign LUT_2[4346] = 32'b11111111111111111000001011001001;
assign LUT_2[4347] = 32'b11111111111111110101000011100010;
assign LUT_2[4348] = 32'b11111111111111101101101111110101;
assign LUT_2[4349] = 32'b11111111111111101010101000001110;
assign LUT_2[4350] = 32'b11111111111111110100101000110001;
assign LUT_2[4351] = 32'b11111111111111110001100001001010;
assign LUT_2[4352] = 32'b00000000000000000011000010110001;
assign LUT_2[4353] = 32'b11111111111111111111111011001010;
assign LUT_2[4354] = 32'b00000000000000001001111011101101;
assign LUT_2[4355] = 32'b00000000000000000110110100000110;
assign LUT_2[4356] = 32'b11111111111111111111100000011001;
assign LUT_2[4357] = 32'b11111111111111111100011000110010;
assign LUT_2[4358] = 32'b00000000000000000110011001010101;
assign LUT_2[4359] = 32'b00000000000000000011010001101110;
assign LUT_2[4360] = 32'b11111111111111111101110100001110;
assign LUT_2[4361] = 32'b11111111111111111010101100100111;
assign LUT_2[4362] = 32'b00000000000000000100101101001010;
assign LUT_2[4363] = 32'b00000000000000000001100101100011;
assign LUT_2[4364] = 32'b11111111111111111010010001110110;
assign LUT_2[4365] = 32'b11111111111111110111001010001111;
assign LUT_2[4366] = 32'b00000000000000000001001010110010;
assign LUT_2[4367] = 32'b11111111111111111110000011001011;
assign LUT_2[4368] = 32'b11111111111111111101100110111011;
assign LUT_2[4369] = 32'b11111111111111111010011111010100;
assign LUT_2[4370] = 32'b00000000000000000100011111110111;
assign LUT_2[4371] = 32'b00000000000000000001011000010000;
assign LUT_2[4372] = 32'b11111111111111111010000100100011;
assign LUT_2[4373] = 32'b11111111111111110110111100111100;
assign LUT_2[4374] = 32'b00000000000000000000111101011111;
assign LUT_2[4375] = 32'b11111111111111111101110101111000;
assign LUT_2[4376] = 32'b11111111111111111000011000011000;
assign LUT_2[4377] = 32'b11111111111111110101010000110001;
assign LUT_2[4378] = 32'b11111111111111111111010001010100;
assign LUT_2[4379] = 32'b11111111111111111100001001101101;
assign LUT_2[4380] = 32'b11111111111111110100110110000000;
assign LUT_2[4381] = 32'b11111111111111110001101110011001;
assign LUT_2[4382] = 32'b11111111111111111011101110111100;
assign LUT_2[4383] = 32'b11111111111111111000100111010101;
assign LUT_2[4384] = 32'b00000000000000000011011110011010;
assign LUT_2[4385] = 32'b00000000000000000000010110110011;
assign LUT_2[4386] = 32'b00000000000000001010010111010110;
assign LUT_2[4387] = 32'b00000000000000000111001111101111;
assign LUT_2[4388] = 32'b11111111111111111111111100000010;
assign LUT_2[4389] = 32'b11111111111111111100110100011011;
assign LUT_2[4390] = 32'b00000000000000000110110100111110;
assign LUT_2[4391] = 32'b00000000000000000011101101010111;
assign LUT_2[4392] = 32'b11111111111111111110001111110111;
assign LUT_2[4393] = 32'b11111111111111111011001000010000;
assign LUT_2[4394] = 32'b00000000000000000101001000110011;
assign LUT_2[4395] = 32'b00000000000000000010000001001100;
assign LUT_2[4396] = 32'b11111111111111111010101101011111;
assign LUT_2[4397] = 32'b11111111111111110111100101111000;
assign LUT_2[4398] = 32'b00000000000000000001100110011011;
assign LUT_2[4399] = 32'b11111111111111111110011110110100;
assign LUT_2[4400] = 32'b11111111111111111110000010100100;
assign LUT_2[4401] = 32'b11111111111111111010111010111101;
assign LUT_2[4402] = 32'b00000000000000000100111011100000;
assign LUT_2[4403] = 32'b00000000000000000001110011111001;
assign LUT_2[4404] = 32'b11111111111111111010100000001100;
assign LUT_2[4405] = 32'b11111111111111110111011000100101;
assign LUT_2[4406] = 32'b00000000000000000001011001001000;
assign LUT_2[4407] = 32'b11111111111111111110010001100001;
assign LUT_2[4408] = 32'b11111111111111111000110100000001;
assign LUT_2[4409] = 32'b11111111111111110101101100011010;
assign LUT_2[4410] = 32'b11111111111111111111101100111101;
assign LUT_2[4411] = 32'b11111111111111111100100101010110;
assign LUT_2[4412] = 32'b11111111111111110101010001101001;
assign LUT_2[4413] = 32'b11111111111111110010001010000010;
assign LUT_2[4414] = 32'b11111111111111111100001010100101;
assign LUT_2[4415] = 32'b11111111111111111001000010111110;
assign LUT_2[4416] = 32'b11111111111111111011001011010100;
assign LUT_2[4417] = 32'b11111111111111111000000011101101;
assign LUT_2[4418] = 32'b00000000000000000010000100010000;
assign LUT_2[4419] = 32'b11111111111111111110111100101001;
assign LUT_2[4420] = 32'b11111111111111110111101000111100;
assign LUT_2[4421] = 32'b11111111111111110100100001010101;
assign LUT_2[4422] = 32'b11111111111111111110100001111000;
assign LUT_2[4423] = 32'b11111111111111111011011010010001;
assign LUT_2[4424] = 32'b11111111111111110101111100110001;
assign LUT_2[4425] = 32'b11111111111111110010110101001010;
assign LUT_2[4426] = 32'b11111111111111111100110101101101;
assign LUT_2[4427] = 32'b11111111111111111001101110000110;
assign LUT_2[4428] = 32'b11111111111111110010011010011001;
assign LUT_2[4429] = 32'b11111111111111101111010010110010;
assign LUT_2[4430] = 32'b11111111111111111001010011010101;
assign LUT_2[4431] = 32'b11111111111111110110001011101110;
assign LUT_2[4432] = 32'b11111111111111110101101111011110;
assign LUT_2[4433] = 32'b11111111111111110010100111110111;
assign LUT_2[4434] = 32'b11111111111111111100101000011010;
assign LUT_2[4435] = 32'b11111111111111111001100000110011;
assign LUT_2[4436] = 32'b11111111111111110010001101000110;
assign LUT_2[4437] = 32'b11111111111111101111000101011111;
assign LUT_2[4438] = 32'b11111111111111111001000110000010;
assign LUT_2[4439] = 32'b11111111111111110101111110011011;
assign LUT_2[4440] = 32'b11111111111111110000100000111011;
assign LUT_2[4441] = 32'b11111111111111101101011001010100;
assign LUT_2[4442] = 32'b11111111111111110111011001110111;
assign LUT_2[4443] = 32'b11111111111111110100010010010000;
assign LUT_2[4444] = 32'b11111111111111101100111110100011;
assign LUT_2[4445] = 32'b11111111111111101001110110111100;
assign LUT_2[4446] = 32'b11111111111111110011110111011111;
assign LUT_2[4447] = 32'b11111111111111110000101111111000;
assign LUT_2[4448] = 32'b11111111111111111011100110111101;
assign LUT_2[4449] = 32'b11111111111111111000011111010110;
assign LUT_2[4450] = 32'b00000000000000000010011111111001;
assign LUT_2[4451] = 32'b11111111111111111111011000010010;
assign LUT_2[4452] = 32'b11111111111111111000000100100101;
assign LUT_2[4453] = 32'b11111111111111110100111100111110;
assign LUT_2[4454] = 32'b11111111111111111110111101100001;
assign LUT_2[4455] = 32'b11111111111111111011110101111010;
assign LUT_2[4456] = 32'b11111111111111110110011000011010;
assign LUT_2[4457] = 32'b11111111111111110011010000110011;
assign LUT_2[4458] = 32'b11111111111111111101010001010110;
assign LUT_2[4459] = 32'b11111111111111111010001001101111;
assign LUT_2[4460] = 32'b11111111111111110010110110000010;
assign LUT_2[4461] = 32'b11111111111111101111101110011011;
assign LUT_2[4462] = 32'b11111111111111111001101110111110;
assign LUT_2[4463] = 32'b11111111111111110110100111010111;
assign LUT_2[4464] = 32'b11111111111111110110001011000111;
assign LUT_2[4465] = 32'b11111111111111110011000011100000;
assign LUT_2[4466] = 32'b11111111111111111101000100000011;
assign LUT_2[4467] = 32'b11111111111111111001111100011100;
assign LUT_2[4468] = 32'b11111111111111110010101000101111;
assign LUT_2[4469] = 32'b11111111111111101111100001001000;
assign LUT_2[4470] = 32'b11111111111111111001100001101011;
assign LUT_2[4471] = 32'b11111111111111110110011010000100;
assign LUT_2[4472] = 32'b11111111111111110000111100100100;
assign LUT_2[4473] = 32'b11111111111111101101110100111101;
assign LUT_2[4474] = 32'b11111111111111110111110101100000;
assign LUT_2[4475] = 32'b11111111111111110100101101111001;
assign LUT_2[4476] = 32'b11111111111111101101011010001100;
assign LUT_2[4477] = 32'b11111111111111101010010010100101;
assign LUT_2[4478] = 32'b11111111111111110100010011001000;
assign LUT_2[4479] = 32'b11111111111111110001001011100001;
assign LUT_2[4480] = 32'b00000000000000000111010111000000;
assign LUT_2[4481] = 32'b00000000000000000100001111011001;
assign LUT_2[4482] = 32'b00000000000000001110001111111100;
assign LUT_2[4483] = 32'b00000000000000001011001000010101;
assign LUT_2[4484] = 32'b00000000000000000011110100101000;
assign LUT_2[4485] = 32'b00000000000000000000101101000001;
assign LUT_2[4486] = 32'b00000000000000001010101101100100;
assign LUT_2[4487] = 32'b00000000000000000111100101111101;
assign LUT_2[4488] = 32'b00000000000000000010001000011101;
assign LUT_2[4489] = 32'b11111111111111111111000000110110;
assign LUT_2[4490] = 32'b00000000000000001001000001011001;
assign LUT_2[4491] = 32'b00000000000000000101111001110010;
assign LUT_2[4492] = 32'b11111111111111111110100110000101;
assign LUT_2[4493] = 32'b11111111111111111011011110011110;
assign LUT_2[4494] = 32'b00000000000000000101011111000001;
assign LUT_2[4495] = 32'b00000000000000000010010111011010;
assign LUT_2[4496] = 32'b00000000000000000001111011001010;
assign LUT_2[4497] = 32'b11111111111111111110110011100011;
assign LUT_2[4498] = 32'b00000000000000001000110100000110;
assign LUT_2[4499] = 32'b00000000000000000101101100011111;
assign LUT_2[4500] = 32'b11111111111111111110011000110010;
assign LUT_2[4501] = 32'b11111111111111111011010001001011;
assign LUT_2[4502] = 32'b00000000000000000101010001101110;
assign LUT_2[4503] = 32'b00000000000000000010001010000111;
assign LUT_2[4504] = 32'b11111111111111111100101100100111;
assign LUT_2[4505] = 32'b11111111111111111001100101000000;
assign LUT_2[4506] = 32'b00000000000000000011100101100011;
assign LUT_2[4507] = 32'b00000000000000000000011101111100;
assign LUT_2[4508] = 32'b11111111111111111001001010001111;
assign LUT_2[4509] = 32'b11111111111111110110000010101000;
assign LUT_2[4510] = 32'b00000000000000000000000011001011;
assign LUT_2[4511] = 32'b11111111111111111100111011100100;
assign LUT_2[4512] = 32'b00000000000000000111110010101001;
assign LUT_2[4513] = 32'b00000000000000000100101011000010;
assign LUT_2[4514] = 32'b00000000000000001110101011100101;
assign LUT_2[4515] = 32'b00000000000000001011100011111110;
assign LUT_2[4516] = 32'b00000000000000000100010000010001;
assign LUT_2[4517] = 32'b00000000000000000001001000101010;
assign LUT_2[4518] = 32'b00000000000000001011001001001101;
assign LUT_2[4519] = 32'b00000000000000001000000001100110;
assign LUT_2[4520] = 32'b00000000000000000010100100000110;
assign LUT_2[4521] = 32'b11111111111111111111011100011111;
assign LUT_2[4522] = 32'b00000000000000001001011101000010;
assign LUT_2[4523] = 32'b00000000000000000110010101011011;
assign LUT_2[4524] = 32'b11111111111111111111000001101110;
assign LUT_2[4525] = 32'b11111111111111111011111010000111;
assign LUT_2[4526] = 32'b00000000000000000101111010101010;
assign LUT_2[4527] = 32'b00000000000000000010110011000011;
assign LUT_2[4528] = 32'b00000000000000000010010110110011;
assign LUT_2[4529] = 32'b11111111111111111111001111001100;
assign LUT_2[4530] = 32'b00000000000000001001001111101111;
assign LUT_2[4531] = 32'b00000000000000000110001000001000;
assign LUT_2[4532] = 32'b11111111111111111110110100011011;
assign LUT_2[4533] = 32'b11111111111111111011101100110100;
assign LUT_2[4534] = 32'b00000000000000000101101101010111;
assign LUT_2[4535] = 32'b00000000000000000010100101110000;
assign LUT_2[4536] = 32'b11111111111111111101001000010000;
assign LUT_2[4537] = 32'b11111111111111111010000000101001;
assign LUT_2[4538] = 32'b00000000000000000100000001001100;
assign LUT_2[4539] = 32'b00000000000000000000111001100101;
assign LUT_2[4540] = 32'b11111111111111111001100101111000;
assign LUT_2[4541] = 32'b11111111111111110110011110010001;
assign LUT_2[4542] = 32'b00000000000000000000011110110100;
assign LUT_2[4543] = 32'b11111111111111111101010111001101;
assign LUT_2[4544] = 32'b11111111111111111111011111100011;
assign LUT_2[4545] = 32'b11111111111111111100010111111100;
assign LUT_2[4546] = 32'b00000000000000000110011000011111;
assign LUT_2[4547] = 32'b00000000000000000011010000111000;
assign LUT_2[4548] = 32'b11111111111111111011111101001011;
assign LUT_2[4549] = 32'b11111111111111111000110101100100;
assign LUT_2[4550] = 32'b00000000000000000010110110000111;
assign LUT_2[4551] = 32'b11111111111111111111101110100000;
assign LUT_2[4552] = 32'b11111111111111111010010001000000;
assign LUT_2[4553] = 32'b11111111111111110111001001011001;
assign LUT_2[4554] = 32'b00000000000000000001001001111100;
assign LUT_2[4555] = 32'b11111111111111111110000010010101;
assign LUT_2[4556] = 32'b11111111111111110110101110101000;
assign LUT_2[4557] = 32'b11111111111111110011100111000001;
assign LUT_2[4558] = 32'b11111111111111111101100111100100;
assign LUT_2[4559] = 32'b11111111111111111010011111111101;
assign LUT_2[4560] = 32'b11111111111111111010000011101101;
assign LUT_2[4561] = 32'b11111111111111110110111100000110;
assign LUT_2[4562] = 32'b00000000000000000000111100101001;
assign LUT_2[4563] = 32'b11111111111111111101110101000010;
assign LUT_2[4564] = 32'b11111111111111110110100001010101;
assign LUT_2[4565] = 32'b11111111111111110011011001101110;
assign LUT_2[4566] = 32'b11111111111111111101011010010001;
assign LUT_2[4567] = 32'b11111111111111111010010010101010;
assign LUT_2[4568] = 32'b11111111111111110100110101001010;
assign LUT_2[4569] = 32'b11111111111111110001101101100011;
assign LUT_2[4570] = 32'b11111111111111111011101110000110;
assign LUT_2[4571] = 32'b11111111111111111000100110011111;
assign LUT_2[4572] = 32'b11111111111111110001010010110010;
assign LUT_2[4573] = 32'b11111111111111101110001011001011;
assign LUT_2[4574] = 32'b11111111111111111000001011101110;
assign LUT_2[4575] = 32'b11111111111111110101000100000111;
assign LUT_2[4576] = 32'b11111111111111111111111011001100;
assign LUT_2[4577] = 32'b11111111111111111100110011100101;
assign LUT_2[4578] = 32'b00000000000000000110110100001000;
assign LUT_2[4579] = 32'b00000000000000000011101100100001;
assign LUT_2[4580] = 32'b11111111111111111100011000110100;
assign LUT_2[4581] = 32'b11111111111111111001010001001101;
assign LUT_2[4582] = 32'b00000000000000000011010001110000;
assign LUT_2[4583] = 32'b00000000000000000000001010001001;
assign LUT_2[4584] = 32'b11111111111111111010101100101001;
assign LUT_2[4585] = 32'b11111111111111110111100101000010;
assign LUT_2[4586] = 32'b00000000000000000001100101100101;
assign LUT_2[4587] = 32'b11111111111111111110011101111110;
assign LUT_2[4588] = 32'b11111111111111110111001010010001;
assign LUT_2[4589] = 32'b11111111111111110100000010101010;
assign LUT_2[4590] = 32'b11111111111111111110000011001101;
assign LUT_2[4591] = 32'b11111111111111111010111011100110;
assign LUT_2[4592] = 32'b11111111111111111010011111010110;
assign LUT_2[4593] = 32'b11111111111111110111010111101111;
assign LUT_2[4594] = 32'b00000000000000000001011000010010;
assign LUT_2[4595] = 32'b11111111111111111110010000101011;
assign LUT_2[4596] = 32'b11111111111111110110111100111110;
assign LUT_2[4597] = 32'b11111111111111110011110101010111;
assign LUT_2[4598] = 32'b11111111111111111101110101111010;
assign LUT_2[4599] = 32'b11111111111111111010101110010011;
assign LUT_2[4600] = 32'b11111111111111110101010000110011;
assign LUT_2[4601] = 32'b11111111111111110010001001001100;
assign LUT_2[4602] = 32'b11111111111111111100001001101111;
assign LUT_2[4603] = 32'b11111111111111111001000010001000;
assign LUT_2[4604] = 32'b11111111111111110001101110011011;
assign LUT_2[4605] = 32'b11111111111111101110100110110100;
assign LUT_2[4606] = 32'b11111111111111111000100111010111;
assign LUT_2[4607] = 32'b11111111111111110101011111110000;
assign LUT_2[4608] = 32'b00000000000000000011110101111101;
assign LUT_2[4609] = 32'b00000000000000000000101110010110;
assign LUT_2[4610] = 32'b00000000000000001010101110111001;
assign LUT_2[4611] = 32'b00000000000000000111100111010010;
assign LUT_2[4612] = 32'b00000000000000000000010011100101;
assign LUT_2[4613] = 32'b11111111111111111101001011111110;
assign LUT_2[4614] = 32'b00000000000000000111001100100001;
assign LUT_2[4615] = 32'b00000000000000000100000100111010;
assign LUT_2[4616] = 32'b11111111111111111110100111011010;
assign LUT_2[4617] = 32'b11111111111111111011011111110011;
assign LUT_2[4618] = 32'b00000000000000000101100000010110;
assign LUT_2[4619] = 32'b00000000000000000010011000101111;
assign LUT_2[4620] = 32'b11111111111111111011000101000010;
assign LUT_2[4621] = 32'b11111111111111110111111101011011;
assign LUT_2[4622] = 32'b00000000000000000001111101111110;
assign LUT_2[4623] = 32'b11111111111111111110110110010111;
assign LUT_2[4624] = 32'b11111111111111111110011010000111;
assign LUT_2[4625] = 32'b11111111111111111011010010100000;
assign LUT_2[4626] = 32'b00000000000000000101010011000011;
assign LUT_2[4627] = 32'b00000000000000000010001011011100;
assign LUT_2[4628] = 32'b11111111111111111010110111101111;
assign LUT_2[4629] = 32'b11111111111111110111110000001000;
assign LUT_2[4630] = 32'b00000000000000000001110000101011;
assign LUT_2[4631] = 32'b11111111111111111110101001000100;
assign LUT_2[4632] = 32'b11111111111111111001001011100100;
assign LUT_2[4633] = 32'b11111111111111110110000011111101;
assign LUT_2[4634] = 32'b00000000000000000000000100100000;
assign LUT_2[4635] = 32'b11111111111111111100111100111001;
assign LUT_2[4636] = 32'b11111111111111110101101001001100;
assign LUT_2[4637] = 32'b11111111111111110010100001100101;
assign LUT_2[4638] = 32'b11111111111111111100100010001000;
assign LUT_2[4639] = 32'b11111111111111111001011010100001;
assign LUT_2[4640] = 32'b00000000000000000100010001100110;
assign LUT_2[4641] = 32'b00000000000000000001001001111111;
assign LUT_2[4642] = 32'b00000000000000001011001010100010;
assign LUT_2[4643] = 32'b00000000000000001000000010111011;
assign LUT_2[4644] = 32'b00000000000000000000101111001110;
assign LUT_2[4645] = 32'b11111111111111111101100111100111;
assign LUT_2[4646] = 32'b00000000000000000111101000001010;
assign LUT_2[4647] = 32'b00000000000000000100100000100011;
assign LUT_2[4648] = 32'b11111111111111111111000011000011;
assign LUT_2[4649] = 32'b11111111111111111011111011011100;
assign LUT_2[4650] = 32'b00000000000000000101111011111111;
assign LUT_2[4651] = 32'b00000000000000000010110100011000;
assign LUT_2[4652] = 32'b11111111111111111011100000101011;
assign LUT_2[4653] = 32'b11111111111111111000011001000100;
assign LUT_2[4654] = 32'b00000000000000000010011001100111;
assign LUT_2[4655] = 32'b11111111111111111111010010000000;
assign LUT_2[4656] = 32'b11111111111111111110110101110000;
assign LUT_2[4657] = 32'b11111111111111111011101110001001;
assign LUT_2[4658] = 32'b00000000000000000101101110101100;
assign LUT_2[4659] = 32'b00000000000000000010100111000101;
assign LUT_2[4660] = 32'b11111111111111111011010011011000;
assign LUT_2[4661] = 32'b11111111111111111000001011110001;
assign LUT_2[4662] = 32'b00000000000000000010001100010100;
assign LUT_2[4663] = 32'b11111111111111111111000100101101;
assign LUT_2[4664] = 32'b11111111111111111001100111001101;
assign LUT_2[4665] = 32'b11111111111111110110011111100110;
assign LUT_2[4666] = 32'b00000000000000000000100000001001;
assign LUT_2[4667] = 32'b11111111111111111101011000100010;
assign LUT_2[4668] = 32'b11111111111111110110000100110101;
assign LUT_2[4669] = 32'b11111111111111110010111101001110;
assign LUT_2[4670] = 32'b11111111111111111100111101110001;
assign LUT_2[4671] = 32'b11111111111111111001110110001010;
assign LUT_2[4672] = 32'b11111111111111111011111110100000;
assign LUT_2[4673] = 32'b11111111111111111000110110111001;
assign LUT_2[4674] = 32'b00000000000000000010110111011100;
assign LUT_2[4675] = 32'b11111111111111111111101111110101;
assign LUT_2[4676] = 32'b11111111111111111000011100001000;
assign LUT_2[4677] = 32'b11111111111111110101010100100001;
assign LUT_2[4678] = 32'b11111111111111111111010101000100;
assign LUT_2[4679] = 32'b11111111111111111100001101011101;
assign LUT_2[4680] = 32'b11111111111111110110101111111101;
assign LUT_2[4681] = 32'b11111111111111110011101000010110;
assign LUT_2[4682] = 32'b11111111111111111101101000111001;
assign LUT_2[4683] = 32'b11111111111111111010100001010010;
assign LUT_2[4684] = 32'b11111111111111110011001101100101;
assign LUT_2[4685] = 32'b11111111111111110000000101111110;
assign LUT_2[4686] = 32'b11111111111111111010000110100001;
assign LUT_2[4687] = 32'b11111111111111110110111110111010;
assign LUT_2[4688] = 32'b11111111111111110110100010101010;
assign LUT_2[4689] = 32'b11111111111111110011011011000011;
assign LUT_2[4690] = 32'b11111111111111111101011011100110;
assign LUT_2[4691] = 32'b11111111111111111010010011111111;
assign LUT_2[4692] = 32'b11111111111111110011000000010010;
assign LUT_2[4693] = 32'b11111111111111101111111000101011;
assign LUT_2[4694] = 32'b11111111111111111001111001001110;
assign LUT_2[4695] = 32'b11111111111111110110110001100111;
assign LUT_2[4696] = 32'b11111111111111110001010100000111;
assign LUT_2[4697] = 32'b11111111111111101110001100100000;
assign LUT_2[4698] = 32'b11111111111111111000001101000011;
assign LUT_2[4699] = 32'b11111111111111110101000101011100;
assign LUT_2[4700] = 32'b11111111111111101101110001101111;
assign LUT_2[4701] = 32'b11111111111111101010101010001000;
assign LUT_2[4702] = 32'b11111111111111110100101010101011;
assign LUT_2[4703] = 32'b11111111111111110001100011000100;
assign LUT_2[4704] = 32'b11111111111111111100011010001001;
assign LUT_2[4705] = 32'b11111111111111111001010010100010;
assign LUT_2[4706] = 32'b00000000000000000011010011000101;
assign LUT_2[4707] = 32'b00000000000000000000001011011110;
assign LUT_2[4708] = 32'b11111111111111111000110111110001;
assign LUT_2[4709] = 32'b11111111111111110101110000001010;
assign LUT_2[4710] = 32'b11111111111111111111110000101101;
assign LUT_2[4711] = 32'b11111111111111111100101001000110;
assign LUT_2[4712] = 32'b11111111111111110111001011100110;
assign LUT_2[4713] = 32'b11111111111111110100000011111111;
assign LUT_2[4714] = 32'b11111111111111111110000100100010;
assign LUT_2[4715] = 32'b11111111111111111010111100111011;
assign LUT_2[4716] = 32'b11111111111111110011101001001110;
assign LUT_2[4717] = 32'b11111111111111110000100001100111;
assign LUT_2[4718] = 32'b11111111111111111010100010001010;
assign LUT_2[4719] = 32'b11111111111111110111011010100011;
assign LUT_2[4720] = 32'b11111111111111110110111110010011;
assign LUT_2[4721] = 32'b11111111111111110011110110101100;
assign LUT_2[4722] = 32'b11111111111111111101110111001111;
assign LUT_2[4723] = 32'b11111111111111111010101111101000;
assign LUT_2[4724] = 32'b11111111111111110011011011111011;
assign LUT_2[4725] = 32'b11111111111111110000010100010100;
assign LUT_2[4726] = 32'b11111111111111111010010100110111;
assign LUT_2[4727] = 32'b11111111111111110111001101010000;
assign LUT_2[4728] = 32'b11111111111111110001101111110000;
assign LUT_2[4729] = 32'b11111111111111101110101000001001;
assign LUT_2[4730] = 32'b11111111111111111000101000101100;
assign LUT_2[4731] = 32'b11111111111111110101100001000101;
assign LUT_2[4732] = 32'b11111111111111101110001101011000;
assign LUT_2[4733] = 32'b11111111111111101011000101110001;
assign LUT_2[4734] = 32'b11111111111111110101000110010100;
assign LUT_2[4735] = 32'b11111111111111110001111110101101;
assign LUT_2[4736] = 32'b00000000000000001000001010001100;
assign LUT_2[4737] = 32'b00000000000000000101000010100101;
assign LUT_2[4738] = 32'b00000000000000001111000011001000;
assign LUT_2[4739] = 32'b00000000000000001011111011100001;
assign LUT_2[4740] = 32'b00000000000000000100100111110100;
assign LUT_2[4741] = 32'b00000000000000000001100000001101;
assign LUT_2[4742] = 32'b00000000000000001011100000110000;
assign LUT_2[4743] = 32'b00000000000000001000011001001001;
assign LUT_2[4744] = 32'b00000000000000000010111011101001;
assign LUT_2[4745] = 32'b11111111111111111111110100000010;
assign LUT_2[4746] = 32'b00000000000000001001110100100101;
assign LUT_2[4747] = 32'b00000000000000000110101100111110;
assign LUT_2[4748] = 32'b11111111111111111111011001010001;
assign LUT_2[4749] = 32'b11111111111111111100010001101010;
assign LUT_2[4750] = 32'b00000000000000000110010010001101;
assign LUT_2[4751] = 32'b00000000000000000011001010100110;
assign LUT_2[4752] = 32'b00000000000000000010101110010110;
assign LUT_2[4753] = 32'b11111111111111111111100110101111;
assign LUT_2[4754] = 32'b00000000000000001001100111010010;
assign LUT_2[4755] = 32'b00000000000000000110011111101011;
assign LUT_2[4756] = 32'b11111111111111111111001011111110;
assign LUT_2[4757] = 32'b11111111111111111100000100010111;
assign LUT_2[4758] = 32'b00000000000000000110000100111010;
assign LUT_2[4759] = 32'b00000000000000000010111101010011;
assign LUT_2[4760] = 32'b11111111111111111101011111110011;
assign LUT_2[4761] = 32'b11111111111111111010011000001100;
assign LUT_2[4762] = 32'b00000000000000000100011000101111;
assign LUT_2[4763] = 32'b00000000000000000001010001001000;
assign LUT_2[4764] = 32'b11111111111111111001111101011011;
assign LUT_2[4765] = 32'b11111111111111110110110101110100;
assign LUT_2[4766] = 32'b00000000000000000000110110010111;
assign LUT_2[4767] = 32'b11111111111111111101101110110000;
assign LUT_2[4768] = 32'b00000000000000001000100101110101;
assign LUT_2[4769] = 32'b00000000000000000101011110001110;
assign LUT_2[4770] = 32'b00000000000000001111011110110001;
assign LUT_2[4771] = 32'b00000000000000001100010111001010;
assign LUT_2[4772] = 32'b00000000000000000101000011011101;
assign LUT_2[4773] = 32'b00000000000000000001111011110110;
assign LUT_2[4774] = 32'b00000000000000001011111100011001;
assign LUT_2[4775] = 32'b00000000000000001000110100110010;
assign LUT_2[4776] = 32'b00000000000000000011010111010010;
assign LUT_2[4777] = 32'b00000000000000000000001111101011;
assign LUT_2[4778] = 32'b00000000000000001010010000001110;
assign LUT_2[4779] = 32'b00000000000000000111001000100111;
assign LUT_2[4780] = 32'b11111111111111111111110100111010;
assign LUT_2[4781] = 32'b11111111111111111100101101010011;
assign LUT_2[4782] = 32'b00000000000000000110101101110110;
assign LUT_2[4783] = 32'b00000000000000000011100110001111;
assign LUT_2[4784] = 32'b00000000000000000011001001111111;
assign LUT_2[4785] = 32'b00000000000000000000000010011000;
assign LUT_2[4786] = 32'b00000000000000001010000010111011;
assign LUT_2[4787] = 32'b00000000000000000110111011010100;
assign LUT_2[4788] = 32'b11111111111111111111100111100111;
assign LUT_2[4789] = 32'b11111111111111111100100000000000;
assign LUT_2[4790] = 32'b00000000000000000110100000100011;
assign LUT_2[4791] = 32'b00000000000000000011011000111100;
assign LUT_2[4792] = 32'b11111111111111111101111011011100;
assign LUT_2[4793] = 32'b11111111111111111010110011110101;
assign LUT_2[4794] = 32'b00000000000000000100110100011000;
assign LUT_2[4795] = 32'b00000000000000000001101100110001;
assign LUT_2[4796] = 32'b11111111111111111010011001000100;
assign LUT_2[4797] = 32'b11111111111111110111010001011101;
assign LUT_2[4798] = 32'b00000000000000000001010010000000;
assign LUT_2[4799] = 32'b11111111111111111110001010011001;
assign LUT_2[4800] = 32'b00000000000000000000010010101111;
assign LUT_2[4801] = 32'b11111111111111111101001011001000;
assign LUT_2[4802] = 32'b00000000000000000111001011101011;
assign LUT_2[4803] = 32'b00000000000000000100000100000100;
assign LUT_2[4804] = 32'b11111111111111111100110000010111;
assign LUT_2[4805] = 32'b11111111111111111001101000110000;
assign LUT_2[4806] = 32'b00000000000000000011101001010011;
assign LUT_2[4807] = 32'b00000000000000000000100001101100;
assign LUT_2[4808] = 32'b11111111111111111011000100001100;
assign LUT_2[4809] = 32'b11111111111111110111111100100101;
assign LUT_2[4810] = 32'b00000000000000000001111101001000;
assign LUT_2[4811] = 32'b11111111111111111110110101100001;
assign LUT_2[4812] = 32'b11111111111111110111100001110100;
assign LUT_2[4813] = 32'b11111111111111110100011010001101;
assign LUT_2[4814] = 32'b11111111111111111110011010110000;
assign LUT_2[4815] = 32'b11111111111111111011010011001001;
assign LUT_2[4816] = 32'b11111111111111111010110110111001;
assign LUT_2[4817] = 32'b11111111111111110111101111010010;
assign LUT_2[4818] = 32'b00000000000000000001101111110101;
assign LUT_2[4819] = 32'b11111111111111111110101000001110;
assign LUT_2[4820] = 32'b11111111111111110111010100100001;
assign LUT_2[4821] = 32'b11111111111111110100001100111010;
assign LUT_2[4822] = 32'b11111111111111111110001101011101;
assign LUT_2[4823] = 32'b11111111111111111011000101110110;
assign LUT_2[4824] = 32'b11111111111111110101101000010110;
assign LUT_2[4825] = 32'b11111111111111110010100000101111;
assign LUT_2[4826] = 32'b11111111111111111100100001010010;
assign LUT_2[4827] = 32'b11111111111111111001011001101011;
assign LUT_2[4828] = 32'b11111111111111110010000101111110;
assign LUT_2[4829] = 32'b11111111111111101110111110010111;
assign LUT_2[4830] = 32'b11111111111111111000111110111010;
assign LUT_2[4831] = 32'b11111111111111110101110111010011;
assign LUT_2[4832] = 32'b00000000000000000000101110011000;
assign LUT_2[4833] = 32'b11111111111111111101100110110001;
assign LUT_2[4834] = 32'b00000000000000000111100111010100;
assign LUT_2[4835] = 32'b00000000000000000100011111101101;
assign LUT_2[4836] = 32'b11111111111111111101001100000000;
assign LUT_2[4837] = 32'b11111111111111111010000100011001;
assign LUT_2[4838] = 32'b00000000000000000100000100111100;
assign LUT_2[4839] = 32'b00000000000000000000111101010101;
assign LUT_2[4840] = 32'b11111111111111111011011111110101;
assign LUT_2[4841] = 32'b11111111111111111000011000001110;
assign LUT_2[4842] = 32'b00000000000000000010011000110001;
assign LUT_2[4843] = 32'b11111111111111111111010001001010;
assign LUT_2[4844] = 32'b11111111111111110111111101011101;
assign LUT_2[4845] = 32'b11111111111111110100110101110110;
assign LUT_2[4846] = 32'b11111111111111111110110110011001;
assign LUT_2[4847] = 32'b11111111111111111011101110110010;
assign LUT_2[4848] = 32'b11111111111111111011010010100010;
assign LUT_2[4849] = 32'b11111111111111111000001010111011;
assign LUT_2[4850] = 32'b00000000000000000010001011011110;
assign LUT_2[4851] = 32'b11111111111111111111000011110111;
assign LUT_2[4852] = 32'b11111111111111110111110000001010;
assign LUT_2[4853] = 32'b11111111111111110100101000100011;
assign LUT_2[4854] = 32'b11111111111111111110101001000110;
assign LUT_2[4855] = 32'b11111111111111111011100001011111;
assign LUT_2[4856] = 32'b11111111111111110110000011111111;
assign LUT_2[4857] = 32'b11111111111111110010111100011000;
assign LUT_2[4858] = 32'b11111111111111111100111100111011;
assign LUT_2[4859] = 32'b11111111111111111001110101010100;
assign LUT_2[4860] = 32'b11111111111111110010100001100111;
assign LUT_2[4861] = 32'b11111111111111101111011010000000;
assign LUT_2[4862] = 32'b11111111111111111001011010100011;
assign LUT_2[4863] = 32'b11111111111111110110010010111100;
assign LUT_2[4864] = 32'b00000000000000000111110100100011;
assign LUT_2[4865] = 32'b00000000000000000100101100111100;
assign LUT_2[4866] = 32'b00000000000000001110101101011111;
assign LUT_2[4867] = 32'b00000000000000001011100101111000;
assign LUT_2[4868] = 32'b00000000000000000100010010001011;
assign LUT_2[4869] = 32'b00000000000000000001001010100100;
assign LUT_2[4870] = 32'b00000000000000001011001011000111;
assign LUT_2[4871] = 32'b00000000000000001000000011100000;
assign LUT_2[4872] = 32'b00000000000000000010100110000000;
assign LUT_2[4873] = 32'b11111111111111111111011110011001;
assign LUT_2[4874] = 32'b00000000000000001001011110111100;
assign LUT_2[4875] = 32'b00000000000000000110010111010101;
assign LUT_2[4876] = 32'b11111111111111111111000011101000;
assign LUT_2[4877] = 32'b11111111111111111011111100000001;
assign LUT_2[4878] = 32'b00000000000000000101111100100100;
assign LUT_2[4879] = 32'b00000000000000000010110100111101;
assign LUT_2[4880] = 32'b00000000000000000010011000101101;
assign LUT_2[4881] = 32'b11111111111111111111010001000110;
assign LUT_2[4882] = 32'b00000000000000001001010001101001;
assign LUT_2[4883] = 32'b00000000000000000110001010000010;
assign LUT_2[4884] = 32'b11111111111111111110110110010101;
assign LUT_2[4885] = 32'b11111111111111111011101110101110;
assign LUT_2[4886] = 32'b00000000000000000101101111010001;
assign LUT_2[4887] = 32'b00000000000000000010100111101010;
assign LUT_2[4888] = 32'b11111111111111111101001010001010;
assign LUT_2[4889] = 32'b11111111111111111010000010100011;
assign LUT_2[4890] = 32'b00000000000000000100000011000110;
assign LUT_2[4891] = 32'b00000000000000000000111011011111;
assign LUT_2[4892] = 32'b11111111111111111001100111110010;
assign LUT_2[4893] = 32'b11111111111111110110100000001011;
assign LUT_2[4894] = 32'b00000000000000000000100000101110;
assign LUT_2[4895] = 32'b11111111111111111101011001000111;
assign LUT_2[4896] = 32'b00000000000000001000010000001100;
assign LUT_2[4897] = 32'b00000000000000000101001000100101;
assign LUT_2[4898] = 32'b00000000000000001111001001001000;
assign LUT_2[4899] = 32'b00000000000000001100000001100001;
assign LUT_2[4900] = 32'b00000000000000000100101101110100;
assign LUT_2[4901] = 32'b00000000000000000001100110001101;
assign LUT_2[4902] = 32'b00000000000000001011100110110000;
assign LUT_2[4903] = 32'b00000000000000001000011111001001;
assign LUT_2[4904] = 32'b00000000000000000011000001101001;
assign LUT_2[4905] = 32'b11111111111111111111111010000010;
assign LUT_2[4906] = 32'b00000000000000001001111010100101;
assign LUT_2[4907] = 32'b00000000000000000110110010111110;
assign LUT_2[4908] = 32'b11111111111111111111011111010001;
assign LUT_2[4909] = 32'b11111111111111111100010111101010;
assign LUT_2[4910] = 32'b00000000000000000110011000001101;
assign LUT_2[4911] = 32'b00000000000000000011010000100110;
assign LUT_2[4912] = 32'b00000000000000000010110100010110;
assign LUT_2[4913] = 32'b11111111111111111111101100101111;
assign LUT_2[4914] = 32'b00000000000000001001101101010010;
assign LUT_2[4915] = 32'b00000000000000000110100101101011;
assign LUT_2[4916] = 32'b11111111111111111111010001111110;
assign LUT_2[4917] = 32'b11111111111111111100001010010111;
assign LUT_2[4918] = 32'b00000000000000000110001010111010;
assign LUT_2[4919] = 32'b00000000000000000011000011010011;
assign LUT_2[4920] = 32'b11111111111111111101100101110011;
assign LUT_2[4921] = 32'b11111111111111111010011110001100;
assign LUT_2[4922] = 32'b00000000000000000100011110101111;
assign LUT_2[4923] = 32'b00000000000000000001010111001000;
assign LUT_2[4924] = 32'b11111111111111111010000011011011;
assign LUT_2[4925] = 32'b11111111111111110110111011110100;
assign LUT_2[4926] = 32'b00000000000000000000111100010111;
assign LUT_2[4927] = 32'b11111111111111111101110100110000;
assign LUT_2[4928] = 32'b11111111111111111111111101000110;
assign LUT_2[4929] = 32'b11111111111111111100110101011111;
assign LUT_2[4930] = 32'b00000000000000000110110110000010;
assign LUT_2[4931] = 32'b00000000000000000011101110011011;
assign LUT_2[4932] = 32'b11111111111111111100011010101110;
assign LUT_2[4933] = 32'b11111111111111111001010011000111;
assign LUT_2[4934] = 32'b00000000000000000011010011101010;
assign LUT_2[4935] = 32'b00000000000000000000001100000011;
assign LUT_2[4936] = 32'b11111111111111111010101110100011;
assign LUT_2[4937] = 32'b11111111111111110111100110111100;
assign LUT_2[4938] = 32'b00000000000000000001100111011111;
assign LUT_2[4939] = 32'b11111111111111111110011111111000;
assign LUT_2[4940] = 32'b11111111111111110111001100001011;
assign LUT_2[4941] = 32'b11111111111111110100000100100100;
assign LUT_2[4942] = 32'b11111111111111111110000101000111;
assign LUT_2[4943] = 32'b11111111111111111010111101100000;
assign LUT_2[4944] = 32'b11111111111111111010100001010000;
assign LUT_2[4945] = 32'b11111111111111110111011001101001;
assign LUT_2[4946] = 32'b00000000000000000001011010001100;
assign LUT_2[4947] = 32'b11111111111111111110010010100101;
assign LUT_2[4948] = 32'b11111111111111110110111110111000;
assign LUT_2[4949] = 32'b11111111111111110011110111010001;
assign LUT_2[4950] = 32'b11111111111111111101110111110100;
assign LUT_2[4951] = 32'b11111111111111111010110000001101;
assign LUT_2[4952] = 32'b11111111111111110101010010101101;
assign LUT_2[4953] = 32'b11111111111111110010001011000110;
assign LUT_2[4954] = 32'b11111111111111111100001011101001;
assign LUT_2[4955] = 32'b11111111111111111001000100000010;
assign LUT_2[4956] = 32'b11111111111111110001110000010101;
assign LUT_2[4957] = 32'b11111111111111101110101000101110;
assign LUT_2[4958] = 32'b11111111111111111000101001010001;
assign LUT_2[4959] = 32'b11111111111111110101100001101010;
assign LUT_2[4960] = 32'b00000000000000000000011000101111;
assign LUT_2[4961] = 32'b11111111111111111101010001001000;
assign LUT_2[4962] = 32'b00000000000000000111010001101011;
assign LUT_2[4963] = 32'b00000000000000000100001010000100;
assign LUT_2[4964] = 32'b11111111111111111100110110010111;
assign LUT_2[4965] = 32'b11111111111111111001101110110000;
assign LUT_2[4966] = 32'b00000000000000000011101111010011;
assign LUT_2[4967] = 32'b00000000000000000000100111101100;
assign LUT_2[4968] = 32'b11111111111111111011001010001100;
assign LUT_2[4969] = 32'b11111111111111111000000010100101;
assign LUT_2[4970] = 32'b00000000000000000010000011001000;
assign LUT_2[4971] = 32'b11111111111111111110111011100001;
assign LUT_2[4972] = 32'b11111111111111110111100111110100;
assign LUT_2[4973] = 32'b11111111111111110100100000001101;
assign LUT_2[4974] = 32'b11111111111111111110100000110000;
assign LUT_2[4975] = 32'b11111111111111111011011001001001;
assign LUT_2[4976] = 32'b11111111111111111010111100111001;
assign LUT_2[4977] = 32'b11111111111111110111110101010010;
assign LUT_2[4978] = 32'b00000000000000000001110101110101;
assign LUT_2[4979] = 32'b11111111111111111110101110001110;
assign LUT_2[4980] = 32'b11111111111111110111011010100001;
assign LUT_2[4981] = 32'b11111111111111110100010010111010;
assign LUT_2[4982] = 32'b11111111111111111110010011011101;
assign LUT_2[4983] = 32'b11111111111111111011001011110110;
assign LUT_2[4984] = 32'b11111111111111110101101110010110;
assign LUT_2[4985] = 32'b11111111111111110010100110101111;
assign LUT_2[4986] = 32'b11111111111111111100100111010010;
assign LUT_2[4987] = 32'b11111111111111111001011111101011;
assign LUT_2[4988] = 32'b11111111111111110010001011111110;
assign LUT_2[4989] = 32'b11111111111111101111000100010111;
assign LUT_2[4990] = 32'b11111111111111111001000100111010;
assign LUT_2[4991] = 32'b11111111111111110101111101010011;
assign LUT_2[4992] = 32'b00000000000000001100001000110010;
assign LUT_2[4993] = 32'b00000000000000001001000001001011;
assign LUT_2[4994] = 32'b00000000000000010011000001101110;
assign LUT_2[4995] = 32'b00000000000000001111111010000111;
assign LUT_2[4996] = 32'b00000000000000001000100110011010;
assign LUT_2[4997] = 32'b00000000000000000101011110110011;
assign LUT_2[4998] = 32'b00000000000000001111011111010110;
assign LUT_2[4999] = 32'b00000000000000001100010111101111;
assign LUT_2[5000] = 32'b00000000000000000110111010001111;
assign LUT_2[5001] = 32'b00000000000000000011110010101000;
assign LUT_2[5002] = 32'b00000000000000001101110011001011;
assign LUT_2[5003] = 32'b00000000000000001010101011100100;
assign LUT_2[5004] = 32'b00000000000000000011010111110111;
assign LUT_2[5005] = 32'b00000000000000000000010000010000;
assign LUT_2[5006] = 32'b00000000000000001010010000110011;
assign LUT_2[5007] = 32'b00000000000000000111001001001100;
assign LUT_2[5008] = 32'b00000000000000000110101100111100;
assign LUT_2[5009] = 32'b00000000000000000011100101010101;
assign LUT_2[5010] = 32'b00000000000000001101100101111000;
assign LUT_2[5011] = 32'b00000000000000001010011110010001;
assign LUT_2[5012] = 32'b00000000000000000011001010100100;
assign LUT_2[5013] = 32'b00000000000000000000000010111101;
assign LUT_2[5014] = 32'b00000000000000001010000011100000;
assign LUT_2[5015] = 32'b00000000000000000110111011111001;
assign LUT_2[5016] = 32'b00000000000000000001011110011001;
assign LUT_2[5017] = 32'b11111111111111111110010110110010;
assign LUT_2[5018] = 32'b00000000000000001000010111010101;
assign LUT_2[5019] = 32'b00000000000000000101001111101110;
assign LUT_2[5020] = 32'b11111111111111111101111100000001;
assign LUT_2[5021] = 32'b11111111111111111010110100011010;
assign LUT_2[5022] = 32'b00000000000000000100110100111101;
assign LUT_2[5023] = 32'b00000000000000000001101101010110;
assign LUT_2[5024] = 32'b00000000000000001100100100011011;
assign LUT_2[5025] = 32'b00000000000000001001011100110100;
assign LUT_2[5026] = 32'b00000000000000010011011101010111;
assign LUT_2[5027] = 32'b00000000000000010000010101110000;
assign LUT_2[5028] = 32'b00000000000000001001000010000011;
assign LUT_2[5029] = 32'b00000000000000000101111010011100;
assign LUT_2[5030] = 32'b00000000000000001111111010111111;
assign LUT_2[5031] = 32'b00000000000000001100110011011000;
assign LUT_2[5032] = 32'b00000000000000000111010101111000;
assign LUT_2[5033] = 32'b00000000000000000100001110010001;
assign LUT_2[5034] = 32'b00000000000000001110001110110100;
assign LUT_2[5035] = 32'b00000000000000001011000111001101;
assign LUT_2[5036] = 32'b00000000000000000011110011100000;
assign LUT_2[5037] = 32'b00000000000000000000101011111001;
assign LUT_2[5038] = 32'b00000000000000001010101100011100;
assign LUT_2[5039] = 32'b00000000000000000111100100110101;
assign LUT_2[5040] = 32'b00000000000000000111001000100101;
assign LUT_2[5041] = 32'b00000000000000000100000000111110;
assign LUT_2[5042] = 32'b00000000000000001110000001100001;
assign LUT_2[5043] = 32'b00000000000000001010111001111010;
assign LUT_2[5044] = 32'b00000000000000000011100110001101;
assign LUT_2[5045] = 32'b00000000000000000000011110100110;
assign LUT_2[5046] = 32'b00000000000000001010011111001001;
assign LUT_2[5047] = 32'b00000000000000000111010111100010;
assign LUT_2[5048] = 32'b00000000000000000001111010000010;
assign LUT_2[5049] = 32'b11111111111111111110110010011011;
assign LUT_2[5050] = 32'b00000000000000001000110010111110;
assign LUT_2[5051] = 32'b00000000000000000101101011010111;
assign LUT_2[5052] = 32'b11111111111111111110010111101010;
assign LUT_2[5053] = 32'b11111111111111111011010000000011;
assign LUT_2[5054] = 32'b00000000000000000101010000100110;
assign LUT_2[5055] = 32'b00000000000000000010001000111111;
assign LUT_2[5056] = 32'b00000000000000000100010001010101;
assign LUT_2[5057] = 32'b00000000000000000001001001101110;
assign LUT_2[5058] = 32'b00000000000000001011001010010001;
assign LUT_2[5059] = 32'b00000000000000001000000010101010;
assign LUT_2[5060] = 32'b00000000000000000000101110111101;
assign LUT_2[5061] = 32'b11111111111111111101100111010110;
assign LUT_2[5062] = 32'b00000000000000000111100111111001;
assign LUT_2[5063] = 32'b00000000000000000100100000010010;
assign LUT_2[5064] = 32'b11111111111111111111000010110010;
assign LUT_2[5065] = 32'b11111111111111111011111011001011;
assign LUT_2[5066] = 32'b00000000000000000101111011101110;
assign LUT_2[5067] = 32'b00000000000000000010110100000111;
assign LUT_2[5068] = 32'b11111111111111111011100000011010;
assign LUT_2[5069] = 32'b11111111111111111000011000110011;
assign LUT_2[5070] = 32'b00000000000000000010011001010110;
assign LUT_2[5071] = 32'b11111111111111111111010001101111;
assign LUT_2[5072] = 32'b11111111111111111110110101011111;
assign LUT_2[5073] = 32'b11111111111111111011101101111000;
assign LUT_2[5074] = 32'b00000000000000000101101110011011;
assign LUT_2[5075] = 32'b00000000000000000010100110110100;
assign LUT_2[5076] = 32'b11111111111111111011010011000111;
assign LUT_2[5077] = 32'b11111111111111111000001011100000;
assign LUT_2[5078] = 32'b00000000000000000010001100000011;
assign LUT_2[5079] = 32'b11111111111111111111000100011100;
assign LUT_2[5080] = 32'b11111111111111111001100110111100;
assign LUT_2[5081] = 32'b11111111111111110110011111010101;
assign LUT_2[5082] = 32'b00000000000000000000011111111000;
assign LUT_2[5083] = 32'b11111111111111111101011000010001;
assign LUT_2[5084] = 32'b11111111111111110110000100100100;
assign LUT_2[5085] = 32'b11111111111111110010111100111101;
assign LUT_2[5086] = 32'b11111111111111111100111101100000;
assign LUT_2[5087] = 32'b11111111111111111001110101111001;
assign LUT_2[5088] = 32'b00000000000000000100101100111110;
assign LUT_2[5089] = 32'b00000000000000000001100101010111;
assign LUT_2[5090] = 32'b00000000000000001011100101111010;
assign LUT_2[5091] = 32'b00000000000000001000011110010011;
assign LUT_2[5092] = 32'b00000000000000000001001010100110;
assign LUT_2[5093] = 32'b11111111111111111110000010111111;
assign LUT_2[5094] = 32'b00000000000000001000000011100010;
assign LUT_2[5095] = 32'b00000000000000000100111011111011;
assign LUT_2[5096] = 32'b11111111111111111111011110011011;
assign LUT_2[5097] = 32'b11111111111111111100010110110100;
assign LUT_2[5098] = 32'b00000000000000000110010111010111;
assign LUT_2[5099] = 32'b00000000000000000011001111110000;
assign LUT_2[5100] = 32'b11111111111111111011111100000011;
assign LUT_2[5101] = 32'b11111111111111111000110100011100;
assign LUT_2[5102] = 32'b00000000000000000010110100111111;
assign LUT_2[5103] = 32'b11111111111111111111101101011000;
assign LUT_2[5104] = 32'b11111111111111111111010001001000;
assign LUT_2[5105] = 32'b11111111111111111100001001100001;
assign LUT_2[5106] = 32'b00000000000000000110001010000100;
assign LUT_2[5107] = 32'b00000000000000000011000010011101;
assign LUT_2[5108] = 32'b11111111111111111011101110110000;
assign LUT_2[5109] = 32'b11111111111111111000100111001001;
assign LUT_2[5110] = 32'b00000000000000000010100111101100;
assign LUT_2[5111] = 32'b11111111111111111111100000000101;
assign LUT_2[5112] = 32'b11111111111111111010000010100101;
assign LUT_2[5113] = 32'b11111111111111110110111010111110;
assign LUT_2[5114] = 32'b00000000000000000000111011100001;
assign LUT_2[5115] = 32'b11111111111111111101110011111010;
assign LUT_2[5116] = 32'b11111111111111110110100000001101;
assign LUT_2[5117] = 32'b11111111111111110011011000100110;
assign LUT_2[5118] = 32'b11111111111111111101011001001001;
assign LUT_2[5119] = 32'b11111111111111111010010001100010;
assign LUT_2[5120] = 32'b00000000000000000101110000010000;
assign LUT_2[5121] = 32'b00000000000000000010101000101001;
assign LUT_2[5122] = 32'b00000000000000001100101001001100;
assign LUT_2[5123] = 32'b00000000000000001001100001100101;
assign LUT_2[5124] = 32'b00000000000000000010001101111000;
assign LUT_2[5125] = 32'b11111111111111111111000110010001;
assign LUT_2[5126] = 32'b00000000000000001001000110110100;
assign LUT_2[5127] = 32'b00000000000000000101111111001101;
assign LUT_2[5128] = 32'b00000000000000000000100001101101;
assign LUT_2[5129] = 32'b11111111111111111101011010000110;
assign LUT_2[5130] = 32'b00000000000000000111011010101001;
assign LUT_2[5131] = 32'b00000000000000000100010011000010;
assign LUT_2[5132] = 32'b11111111111111111100111111010101;
assign LUT_2[5133] = 32'b11111111111111111001110111101110;
assign LUT_2[5134] = 32'b00000000000000000011111000010001;
assign LUT_2[5135] = 32'b00000000000000000000110000101010;
assign LUT_2[5136] = 32'b00000000000000000000010100011010;
assign LUT_2[5137] = 32'b11111111111111111101001100110011;
assign LUT_2[5138] = 32'b00000000000000000111001101010110;
assign LUT_2[5139] = 32'b00000000000000000100000101101111;
assign LUT_2[5140] = 32'b11111111111111111100110010000010;
assign LUT_2[5141] = 32'b11111111111111111001101010011011;
assign LUT_2[5142] = 32'b00000000000000000011101010111110;
assign LUT_2[5143] = 32'b00000000000000000000100011010111;
assign LUT_2[5144] = 32'b11111111111111111011000101110111;
assign LUT_2[5145] = 32'b11111111111111110111111110010000;
assign LUT_2[5146] = 32'b00000000000000000001111110110011;
assign LUT_2[5147] = 32'b11111111111111111110110111001100;
assign LUT_2[5148] = 32'b11111111111111110111100011011111;
assign LUT_2[5149] = 32'b11111111111111110100011011111000;
assign LUT_2[5150] = 32'b11111111111111111110011100011011;
assign LUT_2[5151] = 32'b11111111111111111011010100110100;
assign LUT_2[5152] = 32'b00000000000000000110001011111001;
assign LUT_2[5153] = 32'b00000000000000000011000100010010;
assign LUT_2[5154] = 32'b00000000000000001101000100110101;
assign LUT_2[5155] = 32'b00000000000000001001111101001110;
assign LUT_2[5156] = 32'b00000000000000000010101001100001;
assign LUT_2[5157] = 32'b11111111111111111111100001111010;
assign LUT_2[5158] = 32'b00000000000000001001100010011101;
assign LUT_2[5159] = 32'b00000000000000000110011010110110;
assign LUT_2[5160] = 32'b00000000000000000000111101010110;
assign LUT_2[5161] = 32'b11111111111111111101110101101111;
assign LUT_2[5162] = 32'b00000000000000000111110110010010;
assign LUT_2[5163] = 32'b00000000000000000100101110101011;
assign LUT_2[5164] = 32'b11111111111111111101011010111110;
assign LUT_2[5165] = 32'b11111111111111111010010011010111;
assign LUT_2[5166] = 32'b00000000000000000100010011111010;
assign LUT_2[5167] = 32'b00000000000000000001001100010011;
assign LUT_2[5168] = 32'b00000000000000000000110000000011;
assign LUT_2[5169] = 32'b11111111111111111101101000011100;
assign LUT_2[5170] = 32'b00000000000000000111101000111111;
assign LUT_2[5171] = 32'b00000000000000000100100001011000;
assign LUT_2[5172] = 32'b11111111111111111101001101101011;
assign LUT_2[5173] = 32'b11111111111111111010000110000100;
assign LUT_2[5174] = 32'b00000000000000000100000110100111;
assign LUT_2[5175] = 32'b00000000000000000000111111000000;
assign LUT_2[5176] = 32'b11111111111111111011100001100000;
assign LUT_2[5177] = 32'b11111111111111111000011001111001;
assign LUT_2[5178] = 32'b00000000000000000010011010011100;
assign LUT_2[5179] = 32'b11111111111111111111010010110101;
assign LUT_2[5180] = 32'b11111111111111110111111111001000;
assign LUT_2[5181] = 32'b11111111111111110100110111100001;
assign LUT_2[5182] = 32'b11111111111111111110111000000100;
assign LUT_2[5183] = 32'b11111111111111111011110000011101;
assign LUT_2[5184] = 32'b11111111111111111101111000110011;
assign LUT_2[5185] = 32'b11111111111111111010110001001100;
assign LUT_2[5186] = 32'b00000000000000000100110001101111;
assign LUT_2[5187] = 32'b00000000000000000001101010001000;
assign LUT_2[5188] = 32'b11111111111111111010010110011011;
assign LUT_2[5189] = 32'b11111111111111110111001110110100;
assign LUT_2[5190] = 32'b00000000000000000001001111010111;
assign LUT_2[5191] = 32'b11111111111111111110000111110000;
assign LUT_2[5192] = 32'b11111111111111111000101010010000;
assign LUT_2[5193] = 32'b11111111111111110101100010101001;
assign LUT_2[5194] = 32'b11111111111111111111100011001100;
assign LUT_2[5195] = 32'b11111111111111111100011011100101;
assign LUT_2[5196] = 32'b11111111111111110101000111111000;
assign LUT_2[5197] = 32'b11111111111111110010000000010001;
assign LUT_2[5198] = 32'b11111111111111111100000000110100;
assign LUT_2[5199] = 32'b11111111111111111000111001001101;
assign LUT_2[5200] = 32'b11111111111111111000011100111101;
assign LUT_2[5201] = 32'b11111111111111110101010101010110;
assign LUT_2[5202] = 32'b11111111111111111111010101111001;
assign LUT_2[5203] = 32'b11111111111111111100001110010010;
assign LUT_2[5204] = 32'b11111111111111110100111010100101;
assign LUT_2[5205] = 32'b11111111111111110001110010111110;
assign LUT_2[5206] = 32'b11111111111111111011110011100001;
assign LUT_2[5207] = 32'b11111111111111111000101011111010;
assign LUT_2[5208] = 32'b11111111111111110011001110011010;
assign LUT_2[5209] = 32'b11111111111111110000000110110011;
assign LUT_2[5210] = 32'b11111111111111111010000111010110;
assign LUT_2[5211] = 32'b11111111111111110110111111101111;
assign LUT_2[5212] = 32'b11111111111111101111101100000010;
assign LUT_2[5213] = 32'b11111111111111101100100100011011;
assign LUT_2[5214] = 32'b11111111111111110110100100111110;
assign LUT_2[5215] = 32'b11111111111111110011011101010111;
assign LUT_2[5216] = 32'b11111111111111111110010100011100;
assign LUT_2[5217] = 32'b11111111111111111011001100110101;
assign LUT_2[5218] = 32'b00000000000000000101001101011000;
assign LUT_2[5219] = 32'b00000000000000000010000101110001;
assign LUT_2[5220] = 32'b11111111111111111010110010000100;
assign LUT_2[5221] = 32'b11111111111111110111101010011101;
assign LUT_2[5222] = 32'b00000000000000000001101011000000;
assign LUT_2[5223] = 32'b11111111111111111110100011011001;
assign LUT_2[5224] = 32'b11111111111111111001000101111001;
assign LUT_2[5225] = 32'b11111111111111110101111110010010;
assign LUT_2[5226] = 32'b11111111111111111111111110110101;
assign LUT_2[5227] = 32'b11111111111111111100110111001110;
assign LUT_2[5228] = 32'b11111111111111110101100011100001;
assign LUT_2[5229] = 32'b11111111111111110010011011111010;
assign LUT_2[5230] = 32'b11111111111111111100011100011101;
assign LUT_2[5231] = 32'b11111111111111111001010100110110;
assign LUT_2[5232] = 32'b11111111111111111000111000100110;
assign LUT_2[5233] = 32'b11111111111111110101110000111111;
assign LUT_2[5234] = 32'b11111111111111111111110001100010;
assign LUT_2[5235] = 32'b11111111111111111100101001111011;
assign LUT_2[5236] = 32'b11111111111111110101010110001110;
assign LUT_2[5237] = 32'b11111111111111110010001110100111;
assign LUT_2[5238] = 32'b11111111111111111100001111001010;
assign LUT_2[5239] = 32'b11111111111111111001000111100011;
assign LUT_2[5240] = 32'b11111111111111110011101010000011;
assign LUT_2[5241] = 32'b11111111111111110000100010011100;
assign LUT_2[5242] = 32'b11111111111111111010100010111111;
assign LUT_2[5243] = 32'b11111111111111110111011011011000;
assign LUT_2[5244] = 32'b11111111111111110000000111101011;
assign LUT_2[5245] = 32'b11111111111111101101000000000100;
assign LUT_2[5246] = 32'b11111111111111110111000000100111;
assign LUT_2[5247] = 32'b11111111111111110011111001000000;
assign LUT_2[5248] = 32'b00000000000000001010000100011111;
assign LUT_2[5249] = 32'b00000000000000000110111100111000;
assign LUT_2[5250] = 32'b00000000000000010000111101011011;
assign LUT_2[5251] = 32'b00000000000000001101110101110100;
assign LUT_2[5252] = 32'b00000000000000000110100010000111;
assign LUT_2[5253] = 32'b00000000000000000011011010100000;
assign LUT_2[5254] = 32'b00000000000000001101011011000011;
assign LUT_2[5255] = 32'b00000000000000001010010011011100;
assign LUT_2[5256] = 32'b00000000000000000100110101111100;
assign LUT_2[5257] = 32'b00000000000000000001101110010101;
assign LUT_2[5258] = 32'b00000000000000001011101110111000;
assign LUT_2[5259] = 32'b00000000000000001000100111010001;
assign LUT_2[5260] = 32'b00000000000000000001010011100100;
assign LUT_2[5261] = 32'b11111111111111111110001011111101;
assign LUT_2[5262] = 32'b00000000000000001000001100100000;
assign LUT_2[5263] = 32'b00000000000000000101000100111001;
assign LUT_2[5264] = 32'b00000000000000000100101000101001;
assign LUT_2[5265] = 32'b00000000000000000001100001000010;
assign LUT_2[5266] = 32'b00000000000000001011100001100101;
assign LUT_2[5267] = 32'b00000000000000001000011001111110;
assign LUT_2[5268] = 32'b00000000000000000001000110010001;
assign LUT_2[5269] = 32'b11111111111111111101111110101010;
assign LUT_2[5270] = 32'b00000000000000000111111111001101;
assign LUT_2[5271] = 32'b00000000000000000100110111100110;
assign LUT_2[5272] = 32'b11111111111111111111011010000110;
assign LUT_2[5273] = 32'b11111111111111111100010010011111;
assign LUT_2[5274] = 32'b00000000000000000110010011000010;
assign LUT_2[5275] = 32'b00000000000000000011001011011011;
assign LUT_2[5276] = 32'b11111111111111111011110111101110;
assign LUT_2[5277] = 32'b11111111111111111000110000000111;
assign LUT_2[5278] = 32'b00000000000000000010110000101010;
assign LUT_2[5279] = 32'b11111111111111111111101001000011;
assign LUT_2[5280] = 32'b00000000000000001010100000001000;
assign LUT_2[5281] = 32'b00000000000000000111011000100001;
assign LUT_2[5282] = 32'b00000000000000010001011001000100;
assign LUT_2[5283] = 32'b00000000000000001110010001011101;
assign LUT_2[5284] = 32'b00000000000000000110111101110000;
assign LUT_2[5285] = 32'b00000000000000000011110110001001;
assign LUT_2[5286] = 32'b00000000000000001101110110101100;
assign LUT_2[5287] = 32'b00000000000000001010101111000101;
assign LUT_2[5288] = 32'b00000000000000000101010001100101;
assign LUT_2[5289] = 32'b00000000000000000010001001111110;
assign LUT_2[5290] = 32'b00000000000000001100001010100001;
assign LUT_2[5291] = 32'b00000000000000001001000010111010;
assign LUT_2[5292] = 32'b00000000000000000001101111001101;
assign LUT_2[5293] = 32'b11111111111111111110100111100110;
assign LUT_2[5294] = 32'b00000000000000001000101000001001;
assign LUT_2[5295] = 32'b00000000000000000101100000100010;
assign LUT_2[5296] = 32'b00000000000000000101000100010010;
assign LUT_2[5297] = 32'b00000000000000000001111100101011;
assign LUT_2[5298] = 32'b00000000000000001011111101001110;
assign LUT_2[5299] = 32'b00000000000000001000110101100111;
assign LUT_2[5300] = 32'b00000000000000000001100001111010;
assign LUT_2[5301] = 32'b11111111111111111110011010010011;
assign LUT_2[5302] = 32'b00000000000000001000011010110110;
assign LUT_2[5303] = 32'b00000000000000000101010011001111;
assign LUT_2[5304] = 32'b11111111111111111111110101101111;
assign LUT_2[5305] = 32'b11111111111111111100101110001000;
assign LUT_2[5306] = 32'b00000000000000000110101110101011;
assign LUT_2[5307] = 32'b00000000000000000011100111000100;
assign LUT_2[5308] = 32'b11111111111111111100010011010111;
assign LUT_2[5309] = 32'b11111111111111111001001011110000;
assign LUT_2[5310] = 32'b00000000000000000011001100010011;
assign LUT_2[5311] = 32'b00000000000000000000000100101100;
assign LUT_2[5312] = 32'b00000000000000000010001101000010;
assign LUT_2[5313] = 32'b11111111111111111111000101011011;
assign LUT_2[5314] = 32'b00000000000000001001000101111110;
assign LUT_2[5315] = 32'b00000000000000000101111110010111;
assign LUT_2[5316] = 32'b11111111111111111110101010101010;
assign LUT_2[5317] = 32'b11111111111111111011100011000011;
assign LUT_2[5318] = 32'b00000000000000000101100011100110;
assign LUT_2[5319] = 32'b00000000000000000010011011111111;
assign LUT_2[5320] = 32'b11111111111111111100111110011111;
assign LUT_2[5321] = 32'b11111111111111111001110110111000;
assign LUT_2[5322] = 32'b00000000000000000011110111011011;
assign LUT_2[5323] = 32'b00000000000000000000101111110100;
assign LUT_2[5324] = 32'b11111111111111111001011100000111;
assign LUT_2[5325] = 32'b11111111111111110110010100100000;
assign LUT_2[5326] = 32'b00000000000000000000010101000011;
assign LUT_2[5327] = 32'b11111111111111111101001101011100;
assign LUT_2[5328] = 32'b11111111111111111100110001001100;
assign LUT_2[5329] = 32'b11111111111111111001101001100101;
assign LUT_2[5330] = 32'b00000000000000000011101010001000;
assign LUT_2[5331] = 32'b00000000000000000000100010100001;
assign LUT_2[5332] = 32'b11111111111111111001001110110100;
assign LUT_2[5333] = 32'b11111111111111110110000111001101;
assign LUT_2[5334] = 32'b00000000000000000000000111110000;
assign LUT_2[5335] = 32'b11111111111111111101000000001001;
assign LUT_2[5336] = 32'b11111111111111110111100010101001;
assign LUT_2[5337] = 32'b11111111111111110100011011000010;
assign LUT_2[5338] = 32'b11111111111111111110011011100101;
assign LUT_2[5339] = 32'b11111111111111111011010011111110;
assign LUT_2[5340] = 32'b11111111111111110100000000010001;
assign LUT_2[5341] = 32'b11111111111111110000111000101010;
assign LUT_2[5342] = 32'b11111111111111111010111001001101;
assign LUT_2[5343] = 32'b11111111111111110111110001100110;
assign LUT_2[5344] = 32'b00000000000000000010101000101011;
assign LUT_2[5345] = 32'b11111111111111111111100001000100;
assign LUT_2[5346] = 32'b00000000000000001001100001100111;
assign LUT_2[5347] = 32'b00000000000000000110011010000000;
assign LUT_2[5348] = 32'b11111111111111111111000110010011;
assign LUT_2[5349] = 32'b11111111111111111011111110101100;
assign LUT_2[5350] = 32'b00000000000000000101111111001111;
assign LUT_2[5351] = 32'b00000000000000000010110111101000;
assign LUT_2[5352] = 32'b11111111111111111101011010001000;
assign LUT_2[5353] = 32'b11111111111111111010010010100001;
assign LUT_2[5354] = 32'b00000000000000000100010011000100;
assign LUT_2[5355] = 32'b00000000000000000001001011011101;
assign LUT_2[5356] = 32'b11111111111111111001110111110000;
assign LUT_2[5357] = 32'b11111111111111110110110000001001;
assign LUT_2[5358] = 32'b00000000000000000000110000101100;
assign LUT_2[5359] = 32'b11111111111111111101101001000101;
assign LUT_2[5360] = 32'b11111111111111111101001100110101;
assign LUT_2[5361] = 32'b11111111111111111010000101001110;
assign LUT_2[5362] = 32'b00000000000000000100000101110001;
assign LUT_2[5363] = 32'b00000000000000000000111110001010;
assign LUT_2[5364] = 32'b11111111111111111001101010011101;
assign LUT_2[5365] = 32'b11111111111111110110100010110110;
assign LUT_2[5366] = 32'b00000000000000000000100011011001;
assign LUT_2[5367] = 32'b11111111111111111101011011110010;
assign LUT_2[5368] = 32'b11111111111111110111111110010010;
assign LUT_2[5369] = 32'b11111111111111110100110110101011;
assign LUT_2[5370] = 32'b11111111111111111110110111001110;
assign LUT_2[5371] = 32'b11111111111111111011101111100111;
assign LUT_2[5372] = 32'b11111111111111110100011011111010;
assign LUT_2[5373] = 32'b11111111111111110001010100010011;
assign LUT_2[5374] = 32'b11111111111111111011010100110110;
assign LUT_2[5375] = 32'b11111111111111111000001101001111;
assign LUT_2[5376] = 32'b00000000000000001001101110110110;
assign LUT_2[5377] = 32'b00000000000000000110100111001111;
assign LUT_2[5378] = 32'b00000000000000010000100111110010;
assign LUT_2[5379] = 32'b00000000000000001101100000001011;
assign LUT_2[5380] = 32'b00000000000000000110001100011110;
assign LUT_2[5381] = 32'b00000000000000000011000100110111;
assign LUT_2[5382] = 32'b00000000000000001101000101011010;
assign LUT_2[5383] = 32'b00000000000000001001111101110011;
assign LUT_2[5384] = 32'b00000000000000000100100000010011;
assign LUT_2[5385] = 32'b00000000000000000001011000101100;
assign LUT_2[5386] = 32'b00000000000000001011011001001111;
assign LUT_2[5387] = 32'b00000000000000001000010001101000;
assign LUT_2[5388] = 32'b00000000000000000000111101111011;
assign LUT_2[5389] = 32'b11111111111111111101110110010100;
assign LUT_2[5390] = 32'b00000000000000000111110110110111;
assign LUT_2[5391] = 32'b00000000000000000100101111010000;
assign LUT_2[5392] = 32'b00000000000000000100010011000000;
assign LUT_2[5393] = 32'b00000000000000000001001011011001;
assign LUT_2[5394] = 32'b00000000000000001011001011111100;
assign LUT_2[5395] = 32'b00000000000000001000000100010101;
assign LUT_2[5396] = 32'b00000000000000000000110000101000;
assign LUT_2[5397] = 32'b11111111111111111101101001000001;
assign LUT_2[5398] = 32'b00000000000000000111101001100100;
assign LUT_2[5399] = 32'b00000000000000000100100001111101;
assign LUT_2[5400] = 32'b11111111111111111111000100011101;
assign LUT_2[5401] = 32'b11111111111111111011111100110110;
assign LUT_2[5402] = 32'b00000000000000000101111101011001;
assign LUT_2[5403] = 32'b00000000000000000010110101110010;
assign LUT_2[5404] = 32'b11111111111111111011100010000101;
assign LUT_2[5405] = 32'b11111111111111111000011010011110;
assign LUT_2[5406] = 32'b00000000000000000010011011000001;
assign LUT_2[5407] = 32'b11111111111111111111010011011010;
assign LUT_2[5408] = 32'b00000000000000001010001010011111;
assign LUT_2[5409] = 32'b00000000000000000111000010111000;
assign LUT_2[5410] = 32'b00000000000000010001000011011011;
assign LUT_2[5411] = 32'b00000000000000001101111011110100;
assign LUT_2[5412] = 32'b00000000000000000110101000000111;
assign LUT_2[5413] = 32'b00000000000000000011100000100000;
assign LUT_2[5414] = 32'b00000000000000001101100001000011;
assign LUT_2[5415] = 32'b00000000000000001010011001011100;
assign LUT_2[5416] = 32'b00000000000000000100111011111100;
assign LUT_2[5417] = 32'b00000000000000000001110100010101;
assign LUT_2[5418] = 32'b00000000000000001011110100111000;
assign LUT_2[5419] = 32'b00000000000000001000101101010001;
assign LUT_2[5420] = 32'b00000000000000000001011001100100;
assign LUT_2[5421] = 32'b11111111111111111110010001111101;
assign LUT_2[5422] = 32'b00000000000000001000010010100000;
assign LUT_2[5423] = 32'b00000000000000000101001010111001;
assign LUT_2[5424] = 32'b00000000000000000100101110101001;
assign LUT_2[5425] = 32'b00000000000000000001100111000010;
assign LUT_2[5426] = 32'b00000000000000001011100111100101;
assign LUT_2[5427] = 32'b00000000000000001000011111111110;
assign LUT_2[5428] = 32'b00000000000000000001001100010001;
assign LUT_2[5429] = 32'b11111111111111111110000100101010;
assign LUT_2[5430] = 32'b00000000000000001000000101001101;
assign LUT_2[5431] = 32'b00000000000000000100111101100110;
assign LUT_2[5432] = 32'b11111111111111111111100000000110;
assign LUT_2[5433] = 32'b11111111111111111100011000011111;
assign LUT_2[5434] = 32'b00000000000000000110011001000010;
assign LUT_2[5435] = 32'b00000000000000000011010001011011;
assign LUT_2[5436] = 32'b11111111111111111011111101101110;
assign LUT_2[5437] = 32'b11111111111111111000110110000111;
assign LUT_2[5438] = 32'b00000000000000000010110110101010;
assign LUT_2[5439] = 32'b11111111111111111111101111000011;
assign LUT_2[5440] = 32'b00000000000000000001110111011001;
assign LUT_2[5441] = 32'b11111111111111111110101111110010;
assign LUT_2[5442] = 32'b00000000000000001000110000010101;
assign LUT_2[5443] = 32'b00000000000000000101101000101110;
assign LUT_2[5444] = 32'b11111111111111111110010101000001;
assign LUT_2[5445] = 32'b11111111111111111011001101011010;
assign LUT_2[5446] = 32'b00000000000000000101001101111101;
assign LUT_2[5447] = 32'b00000000000000000010000110010110;
assign LUT_2[5448] = 32'b11111111111111111100101000110110;
assign LUT_2[5449] = 32'b11111111111111111001100001001111;
assign LUT_2[5450] = 32'b00000000000000000011100001110010;
assign LUT_2[5451] = 32'b00000000000000000000011010001011;
assign LUT_2[5452] = 32'b11111111111111111001000110011110;
assign LUT_2[5453] = 32'b11111111111111110101111110110111;
assign LUT_2[5454] = 32'b11111111111111111111111111011010;
assign LUT_2[5455] = 32'b11111111111111111100110111110011;
assign LUT_2[5456] = 32'b11111111111111111100011011100011;
assign LUT_2[5457] = 32'b11111111111111111001010011111100;
assign LUT_2[5458] = 32'b00000000000000000011010100011111;
assign LUT_2[5459] = 32'b00000000000000000000001100111000;
assign LUT_2[5460] = 32'b11111111111111111000111001001011;
assign LUT_2[5461] = 32'b11111111111111110101110001100100;
assign LUT_2[5462] = 32'b11111111111111111111110010000111;
assign LUT_2[5463] = 32'b11111111111111111100101010100000;
assign LUT_2[5464] = 32'b11111111111111110111001101000000;
assign LUT_2[5465] = 32'b11111111111111110100000101011001;
assign LUT_2[5466] = 32'b11111111111111111110000101111100;
assign LUT_2[5467] = 32'b11111111111111111010111110010101;
assign LUT_2[5468] = 32'b11111111111111110011101010101000;
assign LUT_2[5469] = 32'b11111111111111110000100011000001;
assign LUT_2[5470] = 32'b11111111111111111010100011100100;
assign LUT_2[5471] = 32'b11111111111111110111011011111101;
assign LUT_2[5472] = 32'b00000000000000000010010011000010;
assign LUT_2[5473] = 32'b11111111111111111111001011011011;
assign LUT_2[5474] = 32'b00000000000000001001001011111110;
assign LUT_2[5475] = 32'b00000000000000000110000100010111;
assign LUT_2[5476] = 32'b11111111111111111110110000101010;
assign LUT_2[5477] = 32'b11111111111111111011101001000011;
assign LUT_2[5478] = 32'b00000000000000000101101001100110;
assign LUT_2[5479] = 32'b00000000000000000010100001111111;
assign LUT_2[5480] = 32'b11111111111111111101000100011111;
assign LUT_2[5481] = 32'b11111111111111111001111100111000;
assign LUT_2[5482] = 32'b00000000000000000011111101011011;
assign LUT_2[5483] = 32'b00000000000000000000110101110100;
assign LUT_2[5484] = 32'b11111111111111111001100010000111;
assign LUT_2[5485] = 32'b11111111111111110110011010100000;
assign LUT_2[5486] = 32'b00000000000000000000011011000011;
assign LUT_2[5487] = 32'b11111111111111111101010011011100;
assign LUT_2[5488] = 32'b11111111111111111100110111001100;
assign LUT_2[5489] = 32'b11111111111111111001101111100101;
assign LUT_2[5490] = 32'b00000000000000000011110000001000;
assign LUT_2[5491] = 32'b00000000000000000000101000100001;
assign LUT_2[5492] = 32'b11111111111111111001010100110100;
assign LUT_2[5493] = 32'b11111111111111110110001101001101;
assign LUT_2[5494] = 32'b00000000000000000000001101110000;
assign LUT_2[5495] = 32'b11111111111111111101000110001001;
assign LUT_2[5496] = 32'b11111111111111110111101000101001;
assign LUT_2[5497] = 32'b11111111111111110100100001000010;
assign LUT_2[5498] = 32'b11111111111111111110100001100101;
assign LUT_2[5499] = 32'b11111111111111111011011001111110;
assign LUT_2[5500] = 32'b11111111111111110100000110010001;
assign LUT_2[5501] = 32'b11111111111111110000111110101010;
assign LUT_2[5502] = 32'b11111111111111111010111111001101;
assign LUT_2[5503] = 32'b11111111111111110111110111100110;
assign LUT_2[5504] = 32'b00000000000000001110000011000101;
assign LUT_2[5505] = 32'b00000000000000001010111011011110;
assign LUT_2[5506] = 32'b00000000000000010100111100000001;
assign LUT_2[5507] = 32'b00000000000000010001110100011010;
assign LUT_2[5508] = 32'b00000000000000001010100000101101;
assign LUT_2[5509] = 32'b00000000000000000111011001000110;
assign LUT_2[5510] = 32'b00000000000000010001011001101001;
assign LUT_2[5511] = 32'b00000000000000001110010010000010;
assign LUT_2[5512] = 32'b00000000000000001000110100100010;
assign LUT_2[5513] = 32'b00000000000000000101101100111011;
assign LUT_2[5514] = 32'b00000000000000001111101101011110;
assign LUT_2[5515] = 32'b00000000000000001100100101110111;
assign LUT_2[5516] = 32'b00000000000000000101010010001010;
assign LUT_2[5517] = 32'b00000000000000000010001010100011;
assign LUT_2[5518] = 32'b00000000000000001100001011000110;
assign LUT_2[5519] = 32'b00000000000000001001000011011111;
assign LUT_2[5520] = 32'b00000000000000001000100111001111;
assign LUT_2[5521] = 32'b00000000000000000101011111101000;
assign LUT_2[5522] = 32'b00000000000000001111100000001011;
assign LUT_2[5523] = 32'b00000000000000001100011000100100;
assign LUT_2[5524] = 32'b00000000000000000101000100110111;
assign LUT_2[5525] = 32'b00000000000000000001111101010000;
assign LUT_2[5526] = 32'b00000000000000001011111101110011;
assign LUT_2[5527] = 32'b00000000000000001000110110001100;
assign LUT_2[5528] = 32'b00000000000000000011011000101100;
assign LUT_2[5529] = 32'b00000000000000000000010001000101;
assign LUT_2[5530] = 32'b00000000000000001010010001101000;
assign LUT_2[5531] = 32'b00000000000000000111001010000001;
assign LUT_2[5532] = 32'b11111111111111111111110110010100;
assign LUT_2[5533] = 32'b11111111111111111100101110101101;
assign LUT_2[5534] = 32'b00000000000000000110101111010000;
assign LUT_2[5535] = 32'b00000000000000000011100111101001;
assign LUT_2[5536] = 32'b00000000000000001110011110101110;
assign LUT_2[5537] = 32'b00000000000000001011010111000111;
assign LUT_2[5538] = 32'b00000000000000010101010111101010;
assign LUT_2[5539] = 32'b00000000000000010010010000000011;
assign LUT_2[5540] = 32'b00000000000000001010111100010110;
assign LUT_2[5541] = 32'b00000000000000000111110100101111;
assign LUT_2[5542] = 32'b00000000000000010001110101010010;
assign LUT_2[5543] = 32'b00000000000000001110101101101011;
assign LUT_2[5544] = 32'b00000000000000001001010000001011;
assign LUT_2[5545] = 32'b00000000000000000110001000100100;
assign LUT_2[5546] = 32'b00000000000000010000001001000111;
assign LUT_2[5547] = 32'b00000000000000001101000001100000;
assign LUT_2[5548] = 32'b00000000000000000101101101110011;
assign LUT_2[5549] = 32'b00000000000000000010100110001100;
assign LUT_2[5550] = 32'b00000000000000001100100110101111;
assign LUT_2[5551] = 32'b00000000000000001001011111001000;
assign LUT_2[5552] = 32'b00000000000000001001000010111000;
assign LUT_2[5553] = 32'b00000000000000000101111011010001;
assign LUT_2[5554] = 32'b00000000000000001111111011110100;
assign LUT_2[5555] = 32'b00000000000000001100110100001101;
assign LUT_2[5556] = 32'b00000000000000000101100000100000;
assign LUT_2[5557] = 32'b00000000000000000010011000111001;
assign LUT_2[5558] = 32'b00000000000000001100011001011100;
assign LUT_2[5559] = 32'b00000000000000001001010001110101;
assign LUT_2[5560] = 32'b00000000000000000011110100010101;
assign LUT_2[5561] = 32'b00000000000000000000101100101110;
assign LUT_2[5562] = 32'b00000000000000001010101101010001;
assign LUT_2[5563] = 32'b00000000000000000111100101101010;
assign LUT_2[5564] = 32'b00000000000000000000010001111101;
assign LUT_2[5565] = 32'b11111111111111111101001010010110;
assign LUT_2[5566] = 32'b00000000000000000111001010111001;
assign LUT_2[5567] = 32'b00000000000000000100000011010010;
assign LUT_2[5568] = 32'b00000000000000000110001011101000;
assign LUT_2[5569] = 32'b00000000000000000011000100000001;
assign LUT_2[5570] = 32'b00000000000000001101000100100100;
assign LUT_2[5571] = 32'b00000000000000001001111100111101;
assign LUT_2[5572] = 32'b00000000000000000010101001010000;
assign LUT_2[5573] = 32'b11111111111111111111100001101001;
assign LUT_2[5574] = 32'b00000000000000001001100010001100;
assign LUT_2[5575] = 32'b00000000000000000110011010100101;
assign LUT_2[5576] = 32'b00000000000000000000111101000101;
assign LUT_2[5577] = 32'b11111111111111111101110101011110;
assign LUT_2[5578] = 32'b00000000000000000111110110000001;
assign LUT_2[5579] = 32'b00000000000000000100101110011010;
assign LUT_2[5580] = 32'b11111111111111111101011010101101;
assign LUT_2[5581] = 32'b11111111111111111010010011000110;
assign LUT_2[5582] = 32'b00000000000000000100010011101001;
assign LUT_2[5583] = 32'b00000000000000000001001100000010;
assign LUT_2[5584] = 32'b00000000000000000000101111110010;
assign LUT_2[5585] = 32'b11111111111111111101101000001011;
assign LUT_2[5586] = 32'b00000000000000000111101000101110;
assign LUT_2[5587] = 32'b00000000000000000100100001000111;
assign LUT_2[5588] = 32'b11111111111111111101001101011010;
assign LUT_2[5589] = 32'b11111111111111111010000101110011;
assign LUT_2[5590] = 32'b00000000000000000100000110010110;
assign LUT_2[5591] = 32'b00000000000000000000111110101111;
assign LUT_2[5592] = 32'b11111111111111111011100001001111;
assign LUT_2[5593] = 32'b11111111111111111000011001101000;
assign LUT_2[5594] = 32'b00000000000000000010011010001011;
assign LUT_2[5595] = 32'b11111111111111111111010010100100;
assign LUT_2[5596] = 32'b11111111111111110111111110110111;
assign LUT_2[5597] = 32'b11111111111111110100110111010000;
assign LUT_2[5598] = 32'b11111111111111111110110111110011;
assign LUT_2[5599] = 32'b11111111111111111011110000001100;
assign LUT_2[5600] = 32'b00000000000000000110100111010001;
assign LUT_2[5601] = 32'b00000000000000000011011111101010;
assign LUT_2[5602] = 32'b00000000000000001101100000001101;
assign LUT_2[5603] = 32'b00000000000000001010011000100110;
assign LUT_2[5604] = 32'b00000000000000000011000100111001;
assign LUT_2[5605] = 32'b11111111111111111111111101010010;
assign LUT_2[5606] = 32'b00000000000000001001111101110101;
assign LUT_2[5607] = 32'b00000000000000000110110110001110;
assign LUT_2[5608] = 32'b00000000000000000001011000101110;
assign LUT_2[5609] = 32'b11111111111111111110010001000111;
assign LUT_2[5610] = 32'b00000000000000001000010001101010;
assign LUT_2[5611] = 32'b00000000000000000101001010000011;
assign LUT_2[5612] = 32'b11111111111111111101110110010110;
assign LUT_2[5613] = 32'b11111111111111111010101110101111;
assign LUT_2[5614] = 32'b00000000000000000100101111010010;
assign LUT_2[5615] = 32'b00000000000000000001100111101011;
assign LUT_2[5616] = 32'b00000000000000000001001011011011;
assign LUT_2[5617] = 32'b11111111111111111110000011110100;
assign LUT_2[5618] = 32'b00000000000000001000000100010111;
assign LUT_2[5619] = 32'b00000000000000000100111100110000;
assign LUT_2[5620] = 32'b11111111111111111101101001000011;
assign LUT_2[5621] = 32'b11111111111111111010100001011100;
assign LUT_2[5622] = 32'b00000000000000000100100001111111;
assign LUT_2[5623] = 32'b00000000000000000001011010011000;
assign LUT_2[5624] = 32'b11111111111111111011111100111000;
assign LUT_2[5625] = 32'b11111111111111111000110101010001;
assign LUT_2[5626] = 32'b00000000000000000010110101110100;
assign LUT_2[5627] = 32'b11111111111111111111101110001101;
assign LUT_2[5628] = 32'b11111111111111111000011010100000;
assign LUT_2[5629] = 32'b11111111111111110101010010111001;
assign LUT_2[5630] = 32'b11111111111111111111010011011100;
assign LUT_2[5631] = 32'b11111111111111111100001011110101;
assign LUT_2[5632] = 32'b00000000000000001010100010000010;
assign LUT_2[5633] = 32'b00000000000000000111011010011011;
assign LUT_2[5634] = 32'b00000000000000010001011010111110;
assign LUT_2[5635] = 32'b00000000000000001110010011010111;
assign LUT_2[5636] = 32'b00000000000000000110111111101010;
assign LUT_2[5637] = 32'b00000000000000000011111000000011;
assign LUT_2[5638] = 32'b00000000000000001101111000100110;
assign LUT_2[5639] = 32'b00000000000000001010110000111111;
assign LUT_2[5640] = 32'b00000000000000000101010011011111;
assign LUT_2[5641] = 32'b00000000000000000010001011111000;
assign LUT_2[5642] = 32'b00000000000000001100001100011011;
assign LUT_2[5643] = 32'b00000000000000001001000100110100;
assign LUT_2[5644] = 32'b00000000000000000001110001000111;
assign LUT_2[5645] = 32'b11111111111111111110101001100000;
assign LUT_2[5646] = 32'b00000000000000001000101010000011;
assign LUT_2[5647] = 32'b00000000000000000101100010011100;
assign LUT_2[5648] = 32'b00000000000000000101000110001100;
assign LUT_2[5649] = 32'b00000000000000000001111110100101;
assign LUT_2[5650] = 32'b00000000000000001011111111001000;
assign LUT_2[5651] = 32'b00000000000000001000110111100001;
assign LUT_2[5652] = 32'b00000000000000000001100011110100;
assign LUT_2[5653] = 32'b11111111111111111110011100001101;
assign LUT_2[5654] = 32'b00000000000000001000011100110000;
assign LUT_2[5655] = 32'b00000000000000000101010101001001;
assign LUT_2[5656] = 32'b11111111111111111111110111101001;
assign LUT_2[5657] = 32'b11111111111111111100110000000010;
assign LUT_2[5658] = 32'b00000000000000000110110000100101;
assign LUT_2[5659] = 32'b00000000000000000011101000111110;
assign LUT_2[5660] = 32'b11111111111111111100010101010001;
assign LUT_2[5661] = 32'b11111111111111111001001101101010;
assign LUT_2[5662] = 32'b00000000000000000011001110001101;
assign LUT_2[5663] = 32'b00000000000000000000000110100110;
assign LUT_2[5664] = 32'b00000000000000001010111101101011;
assign LUT_2[5665] = 32'b00000000000000000111110110000100;
assign LUT_2[5666] = 32'b00000000000000010001110110100111;
assign LUT_2[5667] = 32'b00000000000000001110101111000000;
assign LUT_2[5668] = 32'b00000000000000000111011011010011;
assign LUT_2[5669] = 32'b00000000000000000100010011101100;
assign LUT_2[5670] = 32'b00000000000000001110010100001111;
assign LUT_2[5671] = 32'b00000000000000001011001100101000;
assign LUT_2[5672] = 32'b00000000000000000101101111001000;
assign LUT_2[5673] = 32'b00000000000000000010100111100001;
assign LUT_2[5674] = 32'b00000000000000001100101000000100;
assign LUT_2[5675] = 32'b00000000000000001001100000011101;
assign LUT_2[5676] = 32'b00000000000000000010001100110000;
assign LUT_2[5677] = 32'b11111111111111111111000101001001;
assign LUT_2[5678] = 32'b00000000000000001001000101101100;
assign LUT_2[5679] = 32'b00000000000000000101111110000101;
assign LUT_2[5680] = 32'b00000000000000000101100001110101;
assign LUT_2[5681] = 32'b00000000000000000010011010001110;
assign LUT_2[5682] = 32'b00000000000000001100011010110001;
assign LUT_2[5683] = 32'b00000000000000001001010011001010;
assign LUT_2[5684] = 32'b00000000000000000001111111011101;
assign LUT_2[5685] = 32'b11111111111111111110110111110110;
assign LUT_2[5686] = 32'b00000000000000001000111000011001;
assign LUT_2[5687] = 32'b00000000000000000101110000110010;
assign LUT_2[5688] = 32'b00000000000000000000010011010010;
assign LUT_2[5689] = 32'b11111111111111111101001011101011;
assign LUT_2[5690] = 32'b00000000000000000111001100001110;
assign LUT_2[5691] = 32'b00000000000000000100000100100111;
assign LUT_2[5692] = 32'b11111111111111111100110000111010;
assign LUT_2[5693] = 32'b11111111111111111001101001010011;
assign LUT_2[5694] = 32'b00000000000000000011101001110110;
assign LUT_2[5695] = 32'b00000000000000000000100010001111;
assign LUT_2[5696] = 32'b00000000000000000010101010100101;
assign LUT_2[5697] = 32'b11111111111111111111100010111110;
assign LUT_2[5698] = 32'b00000000000000001001100011100001;
assign LUT_2[5699] = 32'b00000000000000000110011011111010;
assign LUT_2[5700] = 32'b11111111111111111111001000001101;
assign LUT_2[5701] = 32'b11111111111111111100000000100110;
assign LUT_2[5702] = 32'b00000000000000000110000001001001;
assign LUT_2[5703] = 32'b00000000000000000010111001100010;
assign LUT_2[5704] = 32'b11111111111111111101011100000010;
assign LUT_2[5705] = 32'b11111111111111111010010100011011;
assign LUT_2[5706] = 32'b00000000000000000100010100111110;
assign LUT_2[5707] = 32'b00000000000000000001001101010111;
assign LUT_2[5708] = 32'b11111111111111111001111001101010;
assign LUT_2[5709] = 32'b11111111111111110110110010000011;
assign LUT_2[5710] = 32'b00000000000000000000110010100110;
assign LUT_2[5711] = 32'b11111111111111111101101010111111;
assign LUT_2[5712] = 32'b11111111111111111101001110101111;
assign LUT_2[5713] = 32'b11111111111111111010000111001000;
assign LUT_2[5714] = 32'b00000000000000000100000111101011;
assign LUT_2[5715] = 32'b00000000000000000001000000000100;
assign LUT_2[5716] = 32'b11111111111111111001101100010111;
assign LUT_2[5717] = 32'b11111111111111110110100100110000;
assign LUT_2[5718] = 32'b00000000000000000000100101010011;
assign LUT_2[5719] = 32'b11111111111111111101011101101100;
assign LUT_2[5720] = 32'b11111111111111111000000000001100;
assign LUT_2[5721] = 32'b11111111111111110100111000100101;
assign LUT_2[5722] = 32'b11111111111111111110111001001000;
assign LUT_2[5723] = 32'b11111111111111111011110001100001;
assign LUT_2[5724] = 32'b11111111111111110100011101110100;
assign LUT_2[5725] = 32'b11111111111111110001010110001101;
assign LUT_2[5726] = 32'b11111111111111111011010110110000;
assign LUT_2[5727] = 32'b11111111111111111000001111001001;
assign LUT_2[5728] = 32'b00000000000000000011000110001110;
assign LUT_2[5729] = 32'b11111111111111111111111110100111;
assign LUT_2[5730] = 32'b00000000000000001001111111001010;
assign LUT_2[5731] = 32'b00000000000000000110110111100011;
assign LUT_2[5732] = 32'b11111111111111111111100011110110;
assign LUT_2[5733] = 32'b11111111111111111100011100001111;
assign LUT_2[5734] = 32'b00000000000000000110011100110010;
assign LUT_2[5735] = 32'b00000000000000000011010101001011;
assign LUT_2[5736] = 32'b11111111111111111101110111101011;
assign LUT_2[5737] = 32'b11111111111111111010110000000100;
assign LUT_2[5738] = 32'b00000000000000000100110000100111;
assign LUT_2[5739] = 32'b00000000000000000001101001000000;
assign LUT_2[5740] = 32'b11111111111111111010010101010011;
assign LUT_2[5741] = 32'b11111111111111110111001101101100;
assign LUT_2[5742] = 32'b00000000000000000001001110001111;
assign LUT_2[5743] = 32'b11111111111111111110000110101000;
assign LUT_2[5744] = 32'b11111111111111111101101010011000;
assign LUT_2[5745] = 32'b11111111111111111010100010110001;
assign LUT_2[5746] = 32'b00000000000000000100100011010100;
assign LUT_2[5747] = 32'b00000000000000000001011011101101;
assign LUT_2[5748] = 32'b11111111111111111010001000000000;
assign LUT_2[5749] = 32'b11111111111111110111000000011001;
assign LUT_2[5750] = 32'b00000000000000000001000000111100;
assign LUT_2[5751] = 32'b11111111111111111101111001010101;
assign LUT_2[5752] = 32'b11111111111111111000011011110101;
assign LUT_2[5753] = 32'b11111111111111110101010100001110;
assign LUT_2[5754] = 32'b11111111111111111111010100110001;
assign LUT_2[5755] = 32'b11111111111111111100001101001010;
assign LUT_2[5756] = 32'b11111111111111110100111001011101;
assign LUT_2[5757] = 32'b11111111111111110001110001110110;
assign LUT_2[5758] = 32'b11111111111111111011110010011001;
assign LUT_2[5759] = 32'b11111111111111111000101010110010;
assign LUT_2[5760] = 32'b00000000000000001110110110010001;
assign LUT_2[5761] = 32'b00000000000000001011101110101010;
assign LUT_2[5762] = 32'b00000000000000010101101111001101;
assign LUT_2[5763] = 32'b00000000000000010010100111100110;
assign LUT_2[5764] = 32'b00000000000000001011010011111001;
assign LUT_2[5765] = 32'b00000000000000001000001100010010;
assign LUT_2[5766] = 32'b00000000000000010010001100110101;
assign LUT_2[5767] = 32'b00000000000000001111000101001110;
assign LUT_2[5768] = 32'b00000000000000001001100111101110;
assign LUT_2[5769] = 32'b00000000000000000110100000000111;
assign LUT_2[5770] = 32'b00000000000000010000100000101010;
assign LUT_2[5771] = 32'b00000000000000001101011001000011;
assign LUT_2[5772] = 32'b00000000000000000110000101010110;
assign LUT_2[5773] = 32'b00000000000000000010111101101111;
assign LUT_2[5774] = 32'b00000000000000001100111110010010;
assign LUT_2[5775] = 32'b00000000000000001001110110101011;
assign LUT_2[5776] = 32'b00000000000000001001011010011011;
assign LUT_2[5777] = 32'b00000000000000000110010010110100;
assign LUT_2[5778] = 32'b00000000000000010000010011010111;
assign LUT_2[5779] = 32'b00000000000000001101001011110000;
assign LUT_2[5780] = 32'b00000000000000000101111000000011;
assign LUT_2[5781] = 32'b00000000000000000010110000011100;
assign LUT_2[5782] = 32'b00000000000000001100110000111111;
assign LUT_2[5783] = 32'b00000000000000001001101001011000;
assign LUT_2[5784] = 32'b00000000000000000100001011111000;
assign LUT_2[5785] = 32'b00000000000000000001000100010001;
assign LUT_2[5786] = 32'b00000000000000001011000100110100;
assign LUT_2[5787] = 32'b00000000000000000111111101001101;
assign LUT_2[5788] = 32'b00000000000000000000101001100000;
assign LUT_2[5789] = 32'b11111111111111111101100001111001;
assign LUT_2[5790] = 32'b00000000000000000111100010011100;
assign LUT_2[5791] = 32'b00000000000000000100011010110101;
assign LUT_2[5792] = 32'b00000000000000001111010001111010;
assign LUT_2[5793] = 32'b00000000000000001100001010010011;
assign LUT_2[5794] = 32'b00000000000000010110001010110110;
assign LUT_2[5795] = 32'b00000000000000010011000011001111;
assign LUT_2[5796] = 32'b00000000000000001011101111100010;
assign LUT_2[5797] = 32'b00000000000000001000100111111011;
assign LUT_2[5798] = 32'b00000000000000010010101000011110;
assign LUT_2[5799] = 32'b00000000000000001111100000110111;
assign LUT_2[5800] = 32'b00000000000000001010000011010111;
assign LUT_2[5801] = 32'b00000000000000000110111011110000;
assign LUT_2[5802] = 32'b00000000000000010000111100010011;
assign LUT_2[5803] = 32'b00000000000000001101110100101100;
assign LUT_2[5804] = 32'b00000000000000000110100000111111;
assign LUT_2[5805] = 32'b00000000000000000011011001011000;
assign LUT_2[5806] = 32'b00000000000000001101011001111011;
assign LUT_2[5807] = 32'b00000000000000001010010010010100;
assign LUT_2[5808] = 32'b00000000000000001001110110000100;
assign LUT_2[5809] = 32'b00000000000000000110101110011101;
assign LUT_2[5810] = 32'b00000000000000010000101111000000;
assign LUT_2[5811] = 32'b00000000000000001101100111011001;
assign LUT_2[5812] = 32'b00000000000000000110010011101100;
assign LUT_2[5813] = 32'b00000000000000000011001100000101;
assign LUT_2[5814] = 32'b00000000000000001101001100101000;
assign LUT_2[5815] = 32'b00000000000000001010000101000001;
assign LUT_2[5816] = 32'b00000000000000000100100111100001;
assign LUT_2[5817] = 32'b00000000000000000001011111111010;
assign LUT_2[5818] = 32'b00000000000000001011100000011101;
assign LUT_2[5819] = 32'b00000000000000001000011000110110;
assign LUT_2[5820] = 32'b00000000000000000001000101001001;
assign LUT_2[5821] = 32'b11111111111111111101111101100010;
assign LUT_2[5822] = 32'b00000000000000000111111110000101;
assign LUT_2[5823] = 32'b00000000000000000100110110011110;
assign LUT_2[5824] = 32'b00000000000000000110111110110100;
assign LUT_2[5825] = 32'b00000000000000000011110111001101;
assign LUT_2[5826] = 32'b00000000000000001101110111110000;
assign LUT_2[5827] = 32'b00000000000000001010110000001001;
assign LUT_2[5828] = 32'b00000000000000000011011100011100;
assign LUT_2[5829] = 32'b00000000000000000000010100110101;
assign LUT_2[5830] = 32'b00000000000000001010010101011000;
assign LUT_2[5831] = 32'b00000000000000000111001101110001;
assign LUT_2[5832] = 32'b00000000000000000001110000010001;
assign LUT_2[5833] = 32'b11111111111111111110101000101010;
assign LUT_2[5834] = 32'b00000000000000001000101001001101;
assign LUT_2[5835] = 32'b00000000000000000101100001100110;
assign LUT_2[5836] = 32'b11111111111111111110001101111001;
assign LUT_2[5837] = 32'b11111111111111111011000110010010;
assign LUT_2[5838] = 32'b00000000000000000101000110110101;
assign LUT_2[5839] = 32'b00000000000000000001111111001110;
assign LUT_2[5840] = 32'b00000000000000000001100010111110;
assign LUT_2[5841] = 32'b11111111111111111110011011010111;
assign LUT_2[5842] = 32'b00000000000000001000011011111010;
assign LUT_2[5843] = 32'b00000000000000000101010100010011;
assign LUT_2[5844] = 32'b11111111111111111110000000100110;
assign LUT_2[5845] = 32'b11111111111111111010111000111111;
assign LUT_2[5846] = 32'b00000000000000000100111001100010;
assign LUT_2[5847] = 32'b00000000000000000001110001111011;
assign LUT_2[5848] = 32'b11111111111111111100010100011011;
assign LUT_2[5849] = 32'b11111111111111111001001100110100;
assign LUT_2[5850] = 32'b00000000000000000011001101010111;
assign LUT_2[5851] = 32'b00000000000000000000000101110000;
assign LUT_2[5852] = 32'b11111111111111111000110010000011;
assign LUT_2[5853] = 32'b11111111111111110101101010011100;
assign LUT_2[5854] = 32'b11111111111111111111101010111111;
assign LUT_2[5855] = 32'b11111111111111111100100011011000;
assign LUT_2[5856] = 32'b00000000000000000111011010011101;
assign LUT_2[5857] = 32'b00000000000000000100010010110110;
assign LUT_2[5858] = 32'b00000000000000001110010011011001;
assign LUT_2[5859] = 32'b00000000000000001011001011110010;
assign LUT_2[5860] = 32'b00000000000000000011111000000101;
assign LUT_2[5861] = 32'b00000000000000000000110000011110;
assign LUT_2[5862] = 32'b00000000000000001010110001000001;
assign LUT_2[5863] = 32'b00000000000000000111101001011010;
assign LUT_2[5864] = 32'b00000000000000000010001011111010;
assign LUT_2[5865] = 32'b11111111111111111111000100010011;
assign LUT_2[5866] = 32'b00000000000000001001000100110110;
assign LUT_2[5867] = 32'b00000000000000000101111101001111;
assign LUT_2[5868] = 32'b11111111111111111110101001100010;
assign LUT_2[5869] = 32'b11111111111111111011100001111011;
assign LUT_2[5870] = 32'b00000000000000000101100010011110;
assign LUT_2[5871] = 32'b00000000000000000010011010110111;
assign LUT_2[5872] = 32'b00000000000000000001111110100111;
assign LUT_2[5873] = 32'b11111111111111111110110111000000;
assign LUT_2[5874] = 32'b00000000000000001000110111100011;
assign LUT_2[5875] = 32'b00000000000000000101101111111100;
assign LUT_2[5876] = 32'b11111111111111111110011100001111;
assign LUT_2[5877] = 32'b11111111111111111011010100101000;
assign LUT_2[5878] = 32'b00000000000000000101010101001011;
assign LUT_2[5879] = 32'b00000000000000000010001101100100;
assign LUT_2[5880] = 32'b11111111111111111100110000000100;
assign LUT_2[5881] = 32'b11111111111111111001101000011101;
assign LUT_2[5882] = 32'b00000000000000000011101001000000;
assign LUT_2[5883] = 32'b00000000000000000000100001011001;
assign LUT_2[5884] = 32'b11111111111111111001001101101100;
assign LUT_2[5885] = 32'b11111111111111110110000110000101;
assign LUT_2[5886] = 32'b00000000000000000000000110101000;
assign LUT_2[5887] = 32'b11111111111111111100111111000001;
assign LUT_2[5888] = 32'b00000000000000001110100000101000;
assign LUT_2[5889] = 32'b00000000000000001011011001000001;
assign LUT_2[5890] = 32'b00000000000000010101011001100100;
assign LUT_2[5891] = 32'b00000000000000010010010001111101;
assign LUT_2[5892] = 32'b00000000000000001010111110010000;
assign LUT_2[5893] = 32'b00000000000000000111110110101001;
assign LUT_2[5894] = 32'b00000000000000010001110111001100;
assign LUT_2[5895] = 32'b00000000000000001110101111100101;
assign LUT_2[5896] = 32'b00000000000000001001010010000101;
assign LUT_2[5897] = 32'b00000000000000000110001010011110;
assign LUT_2[5898] = 32'b00000000000000010000001011000001;
assign LUT_2[5899] = 32'b00000000000000001101000011011010;
assign LUT_2[5900] = 32'b00000000000000000101101111101101;
assign LUT_2[5901] = 32'b00000000000000000010101000000110;
assign LUT_2[5902] = 32'b00000000000000001100101000101001;
assign LUT_2[5903] = 32'b00000000000000001001100001000010;
assign LUT_2[5904] = 32'b00000000000000001001000100110010;
assign LUT_2[5905] = 32'b00000000000000000101111101001011;
assign LUT_2[5906] = 32'b00000000000000001111111101101110;
assign LUT_2[5907] = 32'b00000000000000001100110110000111;
assign LUT_2[5908] = 32'b00000000000000000101100010011010;
assign LUT_2[5909] = 32'b00000000000000000010011010110011;
assign LUT_2[5910] = 32'b00000000000000001100011011010110;
assign LUT_2[5911] = 32'b00000000000000001001010011101111;
assign LUT_2[5912] = 32'b00000000000000000011110110001111;
assign LUT_2[5913] = 32'b00000000000000000000101110101000;
assign LUT_2[5914] = 32'b00000000000000001010101111001011;
assign LUT_2[5915] = 32'b00000000000000000111100111100100;
assign LUT_2[5916] = 32'b00000000000000000000010011110111;
assign LUT_2[5917] = 32'b11111111111111111101001100010000;
assign LUT_2[5918] = 32'b00000000000000000111001100110011;
assign LUT_2[5919] = 32'b00000000000000000100000101001100;
assign LUT_2[5920] = 32'b00000000000000001110111100010001;
assign LUT_2[5921] = 32'b00000000000000001011110100101010;
assign LUT_2[5922] = 32'b00000000000000010101110101001101;
assign LUT_2[5923] = 32'b00000000000000010010101101100110;
assign LUT_2[5924] = 32'b00000000000000001011011001111001;
assign LUT_2[5925] = 32'b00000000000000001000010010010010;
assign LUT_2[5926] = 32'b00000000000000010010010010110101;
assign LUT_2[5927] = 32'b00000000000000001111001011001110;
assign LUT_2[5928] = 32'b00000000000000001001101101101110;
assign LUT_2[5929] = 32'b00000000000000000110100110000111;
assign LUT_2[5930] = 32'b00000000000000010000100110101010;
assign LUT_2[5931] = 32'b00000000000000001101011111000011;
assign LUT_2[5932] = 32'b00000000000000000110001011010110;
assign LUT_2[5933] = 32'b00000000000000000011000011101111;
assign LUT_2[5934] = 32'b00000000000000001101000100010010;
assign LUT_2[5935] = 32'b00000000000000001001111100101011;
assign LUT_2[5936] = 32'b00000000000000001001100000011011;
assign LUT_2[5937] = 32'b00000000000000000110011000110100;
assign LUT_2[5938] = 32'b00000000000000010000011001010111;
assign LUT_2[5939] = 32'b00000000000000001101010001110000;
assign LUT_2[5940] = 32'b00000000000000000101111110000011;
assign LUT_2[5941] = 32'b00000000000000000010110110011100;
assign LUT_2[5942] = 32'b00000000000000001100110110111111;
assign LUT_2[5943] = 32'b00000000000000001001101111011000;
assign LUT_2[5944] = 32'b00000000000000000100010001111000;
assign LUT_2[5945] = 32'b00000000000000000001001010010001;
assign LUT_2[5946] = 32'b00000000000000001011001010110100;
assign LUT_2[5947] = 32'b00000000000000001000000011001101;
assign LUT_2[5948] = 32'b00000000000000000000101111100000;
assign LUT_2[5949] = 32'b11111111111111111101100111111001;
assign LUT_2[5950] = 32'b00000000000000000111101000011100;
assign LUT_2[5951] = 32'b00000000000000000100100000110101;
assign LUT_2[5952] = 32'b00000000000000000110101001001011;
assign LUT_2[5953] = 32'b00000000000000000011100001100100;
assign LUT_2[5954] = 32'b00000000000000001101100010000111;
assign LUT_2[5955] = 32'b00000000000000001010011010100000;
assign LUT_2[5956] = 32'b00000000000000000011000110110011;
assign LUT_2[5957] = 32'b11111111111111111111111111001100;
assign LUT_2[5958] = 32'b00000000000000001001111111101111;
assign LUT_2[5959] = 32'b00000000000000000110111000001000;
assign LUT_2[5960] = 32'b00000000000000000001011010101000;
assign LUT_2[5961] = 32'b11111111111111111110010011000001;
assign LUT_2[5962] = 32'b00000000000000001000010011100100;
assign LUT_2[5963] = 32'b00000000000000000101001011111101;
assign LUT_2[5964] = 32'b11111111111111111101111000010000;
assign LUT_2[5965] = 32'b11111111111111111010110000101001;
assign LUT_2[5966] = 32'b00000000000000000100110001001100;
assign LUT_2[5967] = 32'b00000000000000000001101001100101;
assign LUT_2[5968] = 32'b00000000000000000001001101010101;
assign LUT_2[5969] = 32'b11111111111111111110000101101110;
assign LUT_2[5970] = 32'b00000000000000001000000110010001;
assign LUT_2[5971] = 32'b00000000000000000100111110101010;
assign LUT_2[5972] = 32'b11111111111111111101101010111101;
assign LUT_2[5973] = 32'b11111111111111111010100011010110;
assign LUT_2[5974] = 32'b00000000000000000100100011111001;
assign LUT_2[5975] = 32'b00000000000000000001011100010010;
assign LUT_2[5976] = 32'b11111111111111111011111110110010;
assign LUT_2[5977] = 32'b11111111111111111000110111001011;
assign LUT_2[5978] = 32'b00000000000000000010110111101110;
assign LUT_2[5979] = 32'b11111111111111111111110000000111;
assign LUT_2[5980] = 32'b11111111111111111000011100011010;
assign LUT_2[5981] = 32'b11111111111111110101010100110011;
assign LUT_2[5982] = 32'b11111111111111111111010101010110;
assign LUT_2[5983] = 32'b11111111111111111100001101101111;
assign LUT_2[5984] = 32'b00000000000000000111000100110100;
assign LUT_2[5985] = 32'b00000000000000000011111101001101;
assign LUT_2[5986] = 32'b00000000000000001101111101110000;
assign LUT_2[5987] = 32'b00000000000000001010110110001001;
assign LUT_2[5988] = 32'b00000000000000000011100010011100;
assign LUT_2[5989] = 32'b00000000000000000000011010110101;
assign LUT_2[5990] = 32'b00000000000000001010011011011000;
assign LUT_2[5991] = 32'b00000000000000000111010011110001;
assign LUT_2[5992] = 32'b00000000000000000001110110010001;
assign LUT_2[5993] = 32'b11111111111111111110101110101010;
assign LUT_2[5994] = 32'b00000000000000001000101111001101;
assign LUT_2[5995] = 32'b00000000000000000101100111100110;
assign LUT_2[5996] = 32'b11111111111111111110010011111001;
assign LUT_2[5997] = 32'b11111111111111111011001100010010;
assign LUT_2[5998] = 32'b00000000000000000101001100110101;
assign LUT_2[5999] = 32'b00000000000000000010000101001110;
assign LUT_2[6000] = 32'b00000000000000000001101000111110;
assign LUT_2[6001] = 32'b11111111111111111110100001010111;
assign LUT_2[6002] = 32'b00000000000000001000100001111010;
assign LUT_2[6003] = 32'b00000000000000000101011010010011;
assign LUT_2[6004] = 32'b11111111111111111110000110100110;
assign LUT_2[6005] = 32'b11111111111111111010111110111111;
assign LUT_2[6006] = 32'b00000000000000000100111111100010;
assign LUT_2[6007] = 32'b00000000000000000001110111111011;
assign LUT_2[6008] = 32'b11111111111111111100011010011011;
assign LUT_2[6009] = 32'b11111111111111111001010010110100;
assign LUT_2[6010] = 32'b00000000000000000011010011010111;
assign LUT_2[6011] = 32'b00000000000000000000001011110000;
assign LUT_2[6012] = 32'b11111111111111111000111000000011;
assign LUT_2[6013] = 32'b11111111111111110101110000011100;
assign LUT_2[6014] = 32'b11111111111111111111110000111111;
assign LUT_2[6015] = 32'b11111111111111111100101001011000;
assign LUT_2[6016] = 32'b00000000000000010010110100110111;
assign LUT_2[6017] = 32'b00000000000000001111101101010000;
assign LUT_2[6018] = 32'b00000000000000011001101101110011;
assign LUT_2[6019] = 32'b00000000000000010110100110001100;
assign LUT_2[6020] = 32'b00000000000000001111010010011111;
assign LUT_2[6021] = 32'b00000000000000001100001010111000;
assign LUT_2[6022] = 32'b00000000000000010110001011011011;
assign LUT_2[6023] = 32'b00000000000000010011000011110100;
assign LUT_2[6024] = 32'b00000000000000001101100110010100;
assign LUT_2[6025] = 32'b00000000000000001010011110101101;
assign LUT_2[6026] = 32'b00000000000000010100011111010000;
assign LUT_2[6027] = 32'b00000000000000010001010111101001;
assign LUT_2[6028] = 32'b00000000000000001010000011111100;
assign LUT_2[6029] = 32'b00000000000000000110111100010101;
assign LUT_2[6030] = 32'b00000000000000010000111100111000;
assign LUT_2[6031] = 32'b00000000000000001101110101010001;
assign LUT_2[6032] = 32'b00000000000000001101011001000001;
assign LUT_2[6033] = 32'b00000000000000001010010001011010;
assign LUT_2[6034] = 32'b00000000000000010100010001111101;
assign LUT_2[6035] = 32'b00000000000000010001001010010110;
assign LUT_2[6036] = 32'b00000000000000001001110110101001;
assign LUT_2[6037] = 32'b00000000000000000110101111000010;
assign LUT_2[6038] = 32'b00000000000000010000101111100101;
assign LUT_2[6039] = 32'b00000000000000001101100111111110;
assign LUT_2[6040] = 32'b00000000000000001000001010011110;
assign LUT_2[6041] = 32'b00000000000000000101000010110111;
assign LUT_2[6042] = 32'b00000000000000001111000011011010;
assign LUT_2[6043] = 32'b00000000000000001011111011110011;
assign LUT_2[6044] = 32'b00000000000000000100101000000110;
assign LUT_2[6045] = 32'b00000000000000000001100000011111;
assign LUT_2[6046] = 32'b00000000000000001011100001000010;
assign LUT_2[6047] = 32'b00000000000000001000011001011011;
assign LUT_2[6048] = 32'b00000000000000010011010000100000;
assign LUT_2[6049] = 32'b00000000000000010000001000111001;
assign LUT_2[6050] = 32'b00000000000000011010001001011100;
assign LUT_2[6051] = 32'b00000000000000010111000001110101;
assign LUT_2[6052] = 32'b00000000000000001111101110001000;
assign LUT_2[6053] = 32'b00000000000000001100100110100001;
assign LUT_2[6054] = 32'b00000000000000010110100111000100;
assign LUT_2[6055] = 32'b00000000000000010011011111011101;
assign LUT_2[6056] = 32'b00000000000000001110000001111101;
assign LUT_2[6057] = 32'b00000000000000001010111010010110;
assign LUT_2[6058] = 32'b00000000000000010100111010111001;
assign LUT_2[6059] = 32'b00000000000000010001110011010010;
assign LUT_2[6060] = 32'b00000000000000001010011111100101;
assign LUT_2[6061] = 32'b00000000000000000111010111111110;
assign LUT_2[6062] = 32'b00000000000000010001011000100001;
assign LUT_2[6063] = 32'b00000000000000001110010000111010;
assign LUT_2[6064] = 32'b00000000000000001101110100101010;
assign LUT_2[6065] = 32'b00000000000000001010101101000011;
assign LUT_2[6066] = 32'b00000000000000010100101101100110;
assign LUT_2[6067] = 32'b00000000000000010001100101111111;
assign LUT_2[6068] = 32'b00000000000000001010010010010010;
assign LUT_2[6069] = 32'b00000000000000000111001010101011;
assign LUT_2[6070] = 32'b00000000000000010001001011001110;
assign LUT_2[6071] = 32'b00000000000000001110000011100111;
assign LUT_2[6072] = 32'b00000000000000001000100110000111;
assign LUT_2[6073] = 32'b00000000000000000101011110100000;
assign LUT_2[6074] = 32'b00000000000000001111011111000011;
assign LUT_2[6075] = 32'b00000000000000001100010111011100;
assign LUT_2[6076] = 32'b00000000000000000101000011101111;
assign LUT_2[6077] = 32'b00000000000000000001111100001000;
assign LUT_2[6078] = 32'b00000000000000001011111100101011;
assign LUT_2[6079] = 32'b00000000000000001000110101000100;
assign LUT_2[6080] = 32'b00000000000000001010111101011010;
assign LUT_2[6081] = 32'b00000000000000000111110101110011;
assign LUT_2[6082] = 32'b00000000000000010001110110010110;
assign LUT_2[6083] = 32'b00000000000000001110101110101111;
assign LUT_2[6084] = 32'b00000000000000000111011011000010;
assign LUT_2[6085] = 32'b00000000000000000100010011011011;
assign LUT_2[6086] = 32'b00000000000000001110010011111110;
assign LUT_2[6087] = 32'b00000000000000001011001100010111;
assign LUT_2[6088] = 32'b00000000000000000101101110110111;
assign LUT_2[6089] = 32'b00000000000000000010100111010000;
assign LUT_2[6090] = 32'b00000000000000001100100111110011;
assign LUT_2[6091] = 32'b00000000000000001001100000001100;
assign LUT_2[6092] = 32'b00000000000000000010001100011111;
assign LUT_2[6093] = 32'b11111111111111111111000100111000;
assign LUT_2[6094] = 32'b00000000000000001001000101011011;
assign LUT_2[6095] = 32'b00000000000000000101111101110100;
assign LUT_2[6096] = 32'b00000000000000000101100001100100;
assign LUT_2[6097] = 32'b00000000000000000010011001111101;
assign LUT_2[6098] = 32'b00000000000000001100011010100000;
assign LUT_2[6099] = 32'b00000000000000001001010010111001;
assign LUT_2[6100] = 32'b00000000000000000001111111001100;
assign LUT_2[6101] = 32'b11111111111111111110110111100101;
assign LUT_2[6102] = 32'b00000000000000001000111000001000;
assign LUT_2[6103] = 32'b00000000000000000101110000100001;
assign LUT_2[6104] = 32'b00000000000000000000010011000001;
assign LUT_2[6105] = 32'b11111111111111111101001011011010;
assign LUT_2[6106] = 32'b00000000000000000111001011111101;
assign LUT_2[6107] = 32'b00000000000000000100000100010110;
assign LUT_2[6108] = 32'b11111111111111111100110000101001;
assign LUT_2[6109] = 32'b11111111111111111001101001000010;
assign LUT_2[6110] = 32'b00000000000000000011101001100101;
assign LUT_2[6111] = 32'b00000000000000000000100001111110;
assign LUT_2[6112] = 32'b00000000000000001011011001000011;
assign LUT_2[6113] = 32'b00000000000000001000010001011100;
assign LUT_2[6114] = 32'b00000000000000010010010001111111;
assign LUT_2[6115] = 32'b00000000000000001111001010011000;
assign LUT_2[6116] = 32'b00000000000000000111110110101011;
assign LUT_2[6117] = 32'b00000000000000000100101111000100;
assign LUT_2[6118] = 32'b00000000000000001110101111100111;
assign LUT_2[6119] = 32'b00000000000000001011101000000000;
assign LUT_2[6120] = 32'b00000000000000000110001010100000;
assign LUT_2[6121] = 32'b00000000000000000011000010111001;
assign LUT_2[6122] = 32'b00000000000000001101000011011100;
assign LUT_2[6123] = 32'b00000000000000001001111011110101;
assign LUT_2[6124] = 32'b00000000000000000010101000001000;
assign LUT_2[6125] = 32'b11111111111111111111100000100001;
assign LUT_2[6126] = 32'b00000000000000001001100001000100;
assign LUT_2[6127] = 32'b00000000000000000110011001011101;
assign LUT_2[6128] = 32'b00000000000000000101111101001101;
assign LUT_2[6129] = 32'b00000000000000000010110101100110;
assign LUT_2[6130] = 32'b00000000000000001100110110001001;
assign LUT_2[6131] = 32'b00000000000000001001101110100010;
assign LUT_2[6132] = 32'b00000000000000000010011010110101;
assign LUT_2[6133] = 32'b11111111111111111111010011001110;
assign LUT_2[6134] = 32'b00000000000000001001010011110001;
assign LUT_2[6135] = 32'b00000000000000000110001100001010;
assign LUT_2[6136] = 32'b00000000000000000000101110101010;
assign LUT_2[6137] = 32'b11111111111111111101100111000011;
assign LUT_2[6138] = 32'b00000000000000000111100111100110;
assign LUT_2[6139] = 32'b00000000000000000100011111111111;
assign LUT_2[6140] = 32'b11111111111111111101001100010010;
assign LUT_2[6141] = 32'b11111111111111111010000100101011;
assign LUT_2[6142] = 32'b00000000000000000100000101001110;
assign LUT_2[6143] = 32'b00000000000000000000111101100111;
assign LUT_2[6144] = 32'b11111111111111111010111010000111;
assign LUT_2[6145] = 32'b11111111111111110111110010100000;
assign LUT_2[6146] = 32'b00000000000000000001110011000011;
assign LUT_2[6147] = 32'b11111111111111111110101011011100;
assign LUT_2[6148] = 32'b11111111111111110111010111101111;
assign LUT_2[6149] = 32'b11111111111111110100010000001000;
assign LUT_2[6150] = 32'b11111111111111111110010000101011;
assign LUT_2[6151] = 32'b11111111111111111011001001000100;
assign LUT_2[6152] = 32'b11111111111111110101101011100100;
assign LUT_2[6153] = 32'b11111111111111110010100011111101;
assign LUT_2[6154] = 32'b11111111111111111100100100100000;
assign LUT_2[6155] = 32'b11111111111111111001011100111001;
assign LUT_2[6156] = 32'b11111111111111110010001001001100;
assign LUT_2[6157] = 32'b11111111111111101111000001100101;
assign LUT_2[6158] = 32'b11111111111111111001000010001000;
assign LUT_2[6159] = 32'b11111111111111110101111010100001;
assign LUT_2[6160] = 32'b11111111111111110101011110010001;
assign LUT_2[6161] = 32'b11111111111111110010010110101010;
assign LUT_2[6162] = 32'b11111111111111111100010111001101;
assign LUT_2[6163] = 32'b11111111111111111001001111100110;
assign LUT_2[6164] = 32'b11111111111111110001111011111001;
assign LUT_2[6165] = 32'b11111111111111101110110100010010;
assign LUT_2[6166] = 32'b11111111111111111000110100110101;
assign LUT_2[6167] = 32'b11111111111111110101101101001110;
assign LUT_2[6168] = 32'b11111111111111110000001111101110;
assign LUT_2[6169] = 32'b11111111111111101101001000000111;
assign LUT_2[6170] = 32'b11111111111111110111001000101010;
assign LUT_2[6171] = 32'b11111111111111110100000001000011;
assign LUT_2[6172] = 32'b11111111111111101100101101010110;
assign LUT_2[6173] = 32'b11111111111111101001100101101111;
assign LUT_2[6174] = 32'b11111111111111110011100110010010;
assign LUT_2[6175] = 32'b11111111111111110000011110101011;
assign LUT_2[6176] = 32'b11111111111111111011010101110000;
assign LUT_2[6177] = 32'b11111111111111111000001110001001;
assign LUT_2[6178] = 32'b00000000000000000010001110101100;
assign LUT_2[6179] = 32'b11111111111111111111000111000101;
assign LUT_2[6180] = 32'b11111111111111110111110011011000;
assign LUT_2[6181] = 32'b11111111111111110100101011110001;
assign LUT_2[6182] = 32'b11111111111111111110101100010100;
assign LUT_2[6183] = 32'b11111111111111111011100100101101;
assign LUT_2[6184] = 32'b11111111111111110110000111001101;
assign LUT_2[6185] = 32'b11111111111111110010111111100110;
assign LUT_2[6186] = 32'b11111111111111111101000000001001;
assign LUT_2[6187] = 32'b11111111111111111001111000100010;
assign LUT_2[6188] = 32'b11111111111111110010100100110101;
assign LUT_2[6189] = 32'b11111111111111101111011101001110;
assign LUT_2[6190] = 32'b11111111111111111001011101110001;
assign LUT_2[6191] = 32'b11111111111111110110010110001010;
assign LUT_2[6192] = 32'b11111111111111110101111001111010;
assign LUT_2[6193] = 32'b11111111111111110010110010010011;
assign LUT_2[6194] = 32'b11111111111111111100110010110110;
assign LUT_2[6195] = 32'b11111111111111111001101011001111;
assign LUT_2[6196] = 32'b11111111111111110010010111100010;
assign LUT_2[6197] = 32'b11111111111111101111001111111011;
assign LUT_2[6198] = 32'b11111111111111111001010000011110;
assign LUT_2[6199] = 32'b11111111111111110110001000110111;
assign LUT_2[6200] = 32'b11111111111111110000101011010111;
assign LUT_2[6201] = 32'b11111111111111101101100011110000;
assign LUT_2[6202] = 32'b11111111111111110111100100010011;
assign LUT_2[6203] = 32'b11111111111111110100011100101100;
assign LUT_2[6204] = 32'b11111111111111101101001000111111;
assign LUT_2[6205] = 32'b11111111111111101010000001011000;
assign LUT_2[6206] = 32'b11111111111111110100000001111011;
assign LUT_2[6207] = 32'b11111111111111110000111010010100;
assign LUT_2[6208] = 32'b11111111111111110011000010101010;
assign LUT_2[6209] = 32'b11111111111111101111111011000011;
assign LUT_2[6210] = 32'b11111111111111111001111011100110;
assign LUT_2[6211] = 32'b11111111111111110110110011111111;
assign LUT_2[6212] = 32'b11111111111111101111100000010010;
assign LUT_2[6213] = 32'b11111111111111101100011000101011;
assign LUT_2[6214] = 32'b11111111111111110110011001001110;
assign LUT_2[6215] = 32'b11111111111111110011010001100111;
assign LUT_2[6216] = 32'b11111111111111101101110100000111;
assign LUT_2[6217] = 32'b11111111111111101010101100100000;
assign LUT_2[6218] = 32'b11111111111111110100101101000011;
assign LUT_2[6219] = 32'b11111111111111110001100101011100;
assign LUT_2[6220] = 32'b11111111111111101010010001101111;
assign LUT_2[6221] = 32'b11111111111111100111001010001000;
assign LUT_2[6222] = 32'b11111111111111110001001010101011;
assign LUT_2[6223] = 32'b11111111111111101110000011000100;
assign LUT_2[6224] = 32'b11111111111111101101100110110100;
assign LUT_2[6225] = 32'b11111111111111101010011111001101;
assign LUT_2[6226] = 32'b11111111111111110100011111110000;
assign LUT_2[6227] = 32'b11111111111111110001011000001001;
assign LUT_2[6228] = 32'b11111111111111101010000100011100;
assign LUT_2[6229] = 32'b11111111111111100110111100110101;
assign LUT_2[6230] = 32'b11111111111111110000111101011000;
assign LUT_2[6231] = 32'b11111111111111101101110101110001;
assign LUT_2[6232] = 32'b11111111111111101000011000010001;
assign LUT_2[6233] = 32'b11111111111111100101010000101010;
assign LUT_2[6234] = 32'b11111111111111101111010001001101;
assign LUT_2[6235] = 32'b11111111111111101100001001100110;
assign LUT_2[6236] = 32'b11111111111111100100110101111001;
assign LUT_2[6237] = 32'b11111111111111100001101110010010;
assign LUT_2[6238] = 32'b11111111111111101011101110110101;
assign LUT_2[6239] = 32'b11111111111111101000100111001110;
assign LUT_2[6240] = 32'b11111111111111110011011110010011;
assign LUT_2[6241] = 32'b11111111111111110000010110101100;
assign LUT_2[6242] = 32'b11111111111111111010010111001111;
assign LUT_2[6243] = 32'b11111111111111110111001111101000;
assign LUT_2[6244] = 32'b11111111111111101111111011111011;
assign LUT_2[6245] = 32'b11111111111111101100110100010100;
assign LUT_2[6246] = 32'b11111111111111110110110100110111;
assign LUT_2[6247] = 32'b11111111111111110011101101010000;
assign LUT_2[6248] = 32'b11111111111111101110001111110000;
assign LUT_2[6249] = 32'b11111111111111101011001000001001;
assign LUT_2[6250] = 32'b11111111111111110101001000101100;
assign LUT_2[6251] = 32'b11111111111111110010000001000101;
assign LUT_2[6252] = 32'b11111111111111101010101101011000;
assign LUT_2[6253] = 32'b11111111111111100111100101110001;
assign LUT_2[6254] = 32'b11111111111111110001100110010100;
assign LUT_2[6255] = 32'b11111111111111101110011110101101;
assign LUT_2[6256] = 32'b11111111111111101110000010011101;
assign LUT_2[6257] = 32'b11111111111111101010111010110110;
assign LUT_2[6258] = 32'b11111111111111110100111011011001;
assign LUT_2[6259] = 32'b11111111111111110001110011110010;
assign LUT_2[6260] = 32'b11111111111111101010100000000101;
assign LUT_2[6261] = 32'b11111111111111100111011000011110;
assign LUT_2[6262] = 32'b11111111111111110001011001000001;
assign LUT_2[6263] = 32'b11111111111111101110010001011010;
assign LUT_2[6264] = 32'b11111111111111101000110011111010;
assign LUT_2[6265] = 32'b11111111111111100101101100010011;
assign LUT_2[6266] = 32'b11111111111111101111101100110110;
assign LUT_2[6267] = 32'b11111111111111101100100101001111;
assign LUT_2[6268] = 32'b11111111111111100101010001100010;
assign LUT_2[6269] = 32'b11111111111111100010001001111011;
assign LUT_2[6270] = 32'b11111111111111101100001010011110;
assign LUT_2[6271] = 32'b11111111111111101001000010110111;
assign LUT_2[6272] = 32'b11111111111111111111001110010110;
assign LUT_2[6273] = 32'b11111111111111111100000110101111;
assign LUT_2[6274] = 32'b00000000000000000110000111010010;
assign LUT_2[6275] = 32'b00000000000000000010111111101011;
assign LUT_2[6276] = 32'b11111111111111111011101011111110;
assign LUT_2[6277] = 32'b11111111111111111000100100010111;
assign LUT_2[6278] = 32'b00000000000000000010100100111010;
assign LUT_2[6279] = 32'b11111111111111111111011101010011;
assign LUT_2[6280] = 32'b11111111111111111001111111110011;
assign LUT_2[6281] = 32'b11111111111111110110111000001100;
assign LUT_2[6282] = 32'b00000000000000000000111000101111;
assign LUT_2[6283] = 32'b11111111111111111101110001001000;
assign LUT_2[6284] = 32'b11111111111111110110011101011011;
assign LUT_2[6285] = 32'b11111111111111110011010101110100;
assign LUT_2[6286] = 32'b11111111111111111101010110010111;
assign LUT_2[6287] = 32'b11111111111111111010001110110000;
assign LUT_2[6288] = 32'b11111111111111111001110010100000;
assign LUT_2[6289] = 32'b11111111111111110110101010111001;
assign LUT_2[6290] = 32'b00000000000000000000101011011100;
assign LUT_2[6291] = 32'b11111111111111111101100011110101;
assign LUT_2[6292] = 32'b11111111111111110110010000001000;
assign LUT_2[6293] = 32'b11111111111111110011001000100001;
assign LUT_2[6294] = 32'b11111111111111111101001001000100;
assign LUT_2[6295] = 32'b11111111111111111010000001011101;
assign LUT_2[6296] = 32'b11111111111111110100100011111101;
assign LUT_2[6297] = 32'b11111111111111110001011100010110;
assign LUT_2[6298] = 32'b11111111111111111011011100111001;
assign LUT_2[6299] = 32'b11111111111111111000010101010010;
assign LUT_2[6300] = 32'b11111111111111110001000001100101;
assign LUT_2[6301] = 32'b11111111111111101101111001111110;
assign LUT_2[6302] = 32'b11111111111111110111111010100001;
assign LUT_2[6303] = 32'b11111111111111110100110010111010;
assign LUT_2[6304] = 32'b11111111111111111111101001111111;
assign LUT_2[6305] = 32'b11111111111111111100100010011000;
assign LUT_2[6306] = 32'b00000000000000000110100010111011;
assign LUT_2[6307] = 32'b00000000000000000011011011010100;
assign LUT_2[6308] = 32'b11111111111111111100000111100111;
assign LUT_2[6309] = 32'b11111111111111111001000000000000;
assign LUT_2[6310] = 32'b00000000000000000011000000100011;
assign LUT_2[6311] = 32'b11111111111111111111111000111100;
assign LUT_2[6312] = 32'b11111111111111111010011011011100;
assign LUT_2[6313] = 32'b11111111111111110111010011110101;
assign LUT_2[6314] = 32'b00000000000000000001010100011000;
assign LUT_2[6315] = 32'b11111111111111111110001100110001;
assign LUT_2[6316] = 32'b11111111111111110110111001000100;
assign LUT_2[6317] = 32'b11111111111111110011110001011101;
assign LUT_2[6318] = 32'b11111111111111111101110010000000;
assign LUT_2[6319] = 32'b11111111111111111010101010011001;
assign LUT_2[6320] = 32'b11111111111111111010001110001001;
assign LUT_2[6321] = 32'b11111111111111110111000110100010;
assign LUT_2[6322] = 32'b00000000000000000001000111000101;
assign LUT_2[6323] = 32'b11111111111111111101111111011110;
assign LUT_2[6324] = 32'b11111111111111110110101011110001;
assign LUT_2[6325] = 32'b11111111111111110011100100001010;
assign LUT_2[6326] = 32'b11111111111111111101100100101101;
assign LUT_2[6327] = 32'b11111111111111111010011101000110;
assign LUT_2[6328] = 32'b11111111111111110100111111100110;
assign LUT_2[6329] = 32'b11111111111111110001110111111111;
assign LUT_2[6330] = 32'b11111111111111111011111000100010;
assign LUT_2[6331] = 32'b11111111111111111000110000111011;
assign LUT_2[6332] = 32'b11111111111111110001011101001110;
assign LUT_2[6333] = 32'b11111111111111101110010101100111;
assign LUT_2[6334] = 32'b11111111111111111000010110001010;
assign LUT_2[6335] = 32'b11111111111111110101001110100011;
assign LUT_2[6336] = 32'b11111111111111110111010110111001;
assign LUT_2[6337] = 32'b11111111111111110100001111010010;
assign LUT_2[6338] = 32'b11111111111111111110001111110101;
assign LUT_2[6339] = 32'b11111111111111111011001000001110;
assign LUT_2[6340] = 32'b11111111111111110011110100100001;
assign LUT_2[6341] = 32'b11111111111111110000101100111010;
assign LUT_2[6342] = 32'b11111111111111111010101101011101;
assign LUT_2[6343] = 32'b11111111111111110111100101110110;
assign LUT_2[6344] = 32'b11111111111111110010001000010110;
assign LUT_2[6345] = 32'b11111111111111101111000000101111;
assign LUT_2[6346] = 32'b11111111111111111001000001010010;
assign LUT_2[6347] = 32'b11111111111111110101111001101011;
assign LUT_2[6348] = 32'b11111111111111101110100101111110;
assign LUT_2[6349] = 32'b11111111111111101011011110010111;
assign LUT_2[6350] = 32'b11111111111111110101011110111010;
assign LUT_2[6351] = 32'b11111111111111110010010111010011;
assign LUT_2[6352] = 32'b11111111111111110001111011000011;
assign LUT_2[6353] = 32'b11111111111111101110110011011100;
assign LUT_2[6354] = 32'b11111111111111111000110011111111;
assign LUT_2[6355] = 32'b11111111111111110101101100011000;
assign LUT_2[6356] = 32'b11111111111111101110011000101011;
assign LUT_2[6357] = 32'b11111111111111101011010001000100;
assign LUT_2[6358] = 32'b11111111111111110101010001100111;
assign LUT_2[6359] = 32'b11111111111111110010001010000000;
assign LUT_2[6360] = 32'b11111111111111101100101100100000;
assign LUT_2[6361] = 32'b11111111111111101001100100111001;
assign LUT_2[6362] = 32'b11111111111111110011100101011100;
assign LUT_2[6363] = 32'b11111111111111110000011101110101;
assign LUT_2[6364] = 32'b11111111111111101001001010001000;
assign LUT_2[6365] = 32'b11111111111111100110000010100001;
assign LUT_2[6366] = 32'b11111111111111110000000011000100;
assign LUT_2[6367] = 32'b11111111111111101100111011011101;
assign LUT_2[6368] = 32'b11111111111111110111110010100010;
assign LUT_2[6369] = 32'b11111111111111110100101010111011;
assign LUT_2[6370] = 32'b11111111111111111110101011011110;
assign LUT_2[6371] = 32'b11111111111111111011100011110111;
assign LUT_2[6372] = 32'b11111111111111110100010000001010;
assign LUT_2[6373] = 32'b11111111111111110001001000100011;
assign LUT_2[6374] = 32'b11111111111111111011001001000110;
assign LUT_2[6375] = 32'b11111111111111111000000001011111;
assign LUT_2[6376] = 32'b11111111111111110010100011111111;
assign LUT_2[6377] = 32'b11111111111111101111011100011000;
assign LUT_2[6378] = 32'b11111111111111111001011100111011;
assign LUT_2[6379] = 32'b11111111111111110110010101010100;
assign LUT_2[6380] = 32'b11111111111111101111000001100111;
assign LUT_2[6381] = 32'b11111111111111101011111010000000;
assign LUT_2[6382] = 32'b11111111111111110101111010100011;
assign LUT_2[6383] = 32'b11111111111111110010110010111100;
assign LUT_2[6384] = 32'b11111111111111110010010110101100;
assign LUT_2[6385] = 32'b11111111111111101111001111000101;
assign LUT_2[6386] = 32'b11111111111111111001001111101000;
assign LUT_2[6387] = 32'b11111111111111110110001000000001;
assign LUT_2[6388] = 32'b11111111111111101110110100010100;
assign LUT_2[6389] = 32'b11111111111111101011101100101101;
assign LUT_2[6390] = 32'b11111111111111110101101101010000;
assign LUT_2[6391] = 32'b11111111111111110010100101101001;
assign LUT_2[6392] = 32'b11111111111111101101001000001001;
assign LUT_2[6393] = 32'b11111111111111101010000000100010;
assign LUT_2[6394] = 32'b11111111111111110100000001000101;
assign LUT_2[6395] = 32'b11111111111111110000111001011110;
assign LUT_2[6396] = 32'b11111111111111101001100101110001;
assign LUT_2[6397] = 32'b11111111111111100110011110001010;
assign LUT_2[6398] = 32'b11111111111111110000011110101101;
assign LUT_2[6399] = 32'b11111111111111101101010111000110;
assign LUT_2[6400] = 32'b11111111111111111110111000101101;
assign LUT_2[6401] = 32'b11111111111111111011110001000110;
assign LUT_2[6402] = 32'b00000000000000000101110001101001;
assign LUT_2[6403] = 32'b00000000000000000010101010000010;
assign LUT_2[6404] = 32'b11111111111111111011010110010101;
assign LUT_2[6405] = 32'b11111111111111111000001110101110;
assign LUT_2[6406] = 32'b00000000000000000010001111010001;
assign LUT_2[6407] = 32'b11111111111111111111000111101010;
assign LUT_2[6408] = 32'b11111111111111111001101010001010;
assign LUT_2[6409] = 32'b11111111111111110110100010100011;
assign LUT_2[6410] = 32'b00000000000000000000100011000110;
assign LUT_2[6411] = 32'b11111111111111111101011011011111;
assign LUT_2[6412] = 32'b11111111111111110110000111110010;
assign LUT_2[6413] = 32'b11111111111111110011000000001011;
assign LUT_2[6414] = 32'b11111111111111111101000000101110;
assign LUT_2[6415] = 32'b11111111111111111001111001000111;
assign LUT_2[6416] = 32'b11111111111111111001011100110111;
assign LUT_2[6417] = 32'b11111111111111110110010101010000;
assign LUT_2[6418] = 32'b00000000000000000000010101110011;
assign LUT_2[6419] = 32'b11111111111111111101001110001100;
assign LUT_2[6420] = 32'b11111111111111110101111010011111;
assign LUT_2[6421] = 32'b11111111111111110010110010111000;
assign LUT_2[6422] = 32'b11111111111111111100110011011011;
assign LUT_2[6423] = 32'b11111111111111111001101011110100;
assign LUT_2[6424] = 32'b11111111111111110100001110010100;
assign LUT_2[6425] = 32'b11111111111111110001000110101101;
assign LUT_2[6426] = 32'b11111111111111111011000111010000;
assign LUT_2[6427] = 32'b11111111111111110111111111101001;
assign LUT_2[6428] = 32'b11111111111111110000101011111100;
assign LUT_2[6429] = 32'b11111111111111101101100100010101;
assign LUT_2[6430] = 32'b11111111111111110111100100111000;
assign LUT_2[6431] = 32'b11111111111111110100011101010001;
assign LUT_2[6432] = 32'b11111111111111111111010100010110;
assign LUT_2[6433] = 32'b11111111111111111100001100101111;
assign LUT_2[6434] = 32'b00000000000000000110001101010010;
assign LUT_2[6435] = 32'b00000000000000000011000101101011;
assign LUT_2[6436] = 32'b11111111111111111011110001111110;
assign LUT_2[6437] = 32'b11111111111111111000101010010111;
assign LUT_2[6438] = 32'b00000000000000000010101010111010;
assign LUT_2[6439] = 32'b11111111111111111111100011010011;
assign LUT_2[6440] = 32'b11111111111111111010000101110011;
assign LUT_2[6441] = 32'b11111111111111110110111110001100;
assign LUT_2[6442] = 32'b00000000000000000000111110101111;
assign LUT_2[6443] = 32'b11111111111111111101110111001000;
assign LUT_2[6444] = 32'b11111111111111110110100011011011;
assign LUT_2[6445] = 32'b11111111111111110011011011110100;
assign LUT_2[6446] = 32'b11111111111111111101011100010111;
assign LUT_2[6447] = 32'b11111111111111111010010100110000;
assign LUT_2[6448] = 32'b11111111111111111001111000100000;
assign LUT_2[6449] = 32'b11111111111111110110110000111001;
assign LUT_2[6450] = 32'b00000000000000000000110001011100;
assign LUT_2[6451] = 32'b11111111111111111101101001110101;
assign LUT_2[6452] = 32'b11111111111111110110010110001000;
assign LUT_2[6453] = 32'b11111111111111110011001110100001;
assign LUT_2[6454] = 32'b11111111111111111101001111000100;
assign LUT_2[6455] = 32'b11111111111111111010000111011101;
assign LUT_2[6456] = 32'b11111111111111110100101001111101;
assign LUT_2[6457] = 32'b11111111111111110001100010010110;
assign LUT_2[6458] = 32'b11111111111111111011100010111001;
assign LUT_2[6459] = 32'b11111111111111111000011011010010;
assign LUT_2[6460] = 32'b11111111111111110001000111100101;
assign LUT_2[6461] = 32'b11111111111111101101111111111110;
assign LUT_2[6462] = 32'b11111111111111111000000000100001;
assign LUT_2[6463] = 32'b11111111111111110100111000111010;
assign LUT_2[6464] = 32'b11111111111111110111000001010000;
assign LUT_2[6465] = 32'b11111111111111110011111001101001;
assign LUT_2[6466] = 32'b11111111111111111101111010001100;
assign LUT_2[6467] = 32'b11111111111111111010110010100101;
assign LUT_2[6468] = 32'b11111111111111110011011110111000;
assign LUT_2[6469] = 32'b11111111111111110000010111010001;
assign LUT_2[6470] = 32'b11111111111111111010010111110100;
assign LUT_2[6471] = 32'b11111111111111110111010000001101;
assign LUT_2[6472] = 32'b11111111111111110001110010101101;
assign LUT_2[6473] = 32'b11111111111111101110101011000110;
assign LUT_2[6474] = 32'b11111111111111111000101011101001;
assign LUT_2[6475] = 32'b11111111111111110101100100000010;
assign LUT_2[6476] = 32'b11111111111111101110010000010101;
assign LUT_2[6477] = 32'b11111111111111101011001000101110;
assign LUT_2[6478] = 32'b11111111111111110101001001010001;
assign LUT_2[6479] = 32'b11111111111111110010000001101010;
assign LUT_2[6480] = 32'b11111111111111110001100101011010;
assign LUT_2[6481] = 32'b11111111111111101110011101110011;
assign LUT_2[6482] = 32'b11111111111111111000011110010110;
assign LUT_2[6483] = 32'b11111111111111110101010110101111;
assign LUT_2[6484] = 32'b11111111111111101110000011000010;
assign LUT_2[6485] = 32'b11111111111111101010111011011011;
assign LUT_2[6486] = 32'b11111111111111110100111011111110;
assign LUT_2[6487] = 32'b11111111111111110001110100010111;
assign LUT_2[6488] = 32'b11111111111111101100010110110111;
assign LUT_2[6489] = 32'b11111111111111101001001111010000;
assign LUT_2[6490] = 32'b11111111111111110011001111110011;
assign LUT_2[6491] = 32'b11111111111111110000001000001100;
assign LUT_2[6492] = 32'b11111111111111101000110100011111;
assign LUT_2[6493] = 32'b11111111111111100101101100111000;
assign LUT_2[6494] = 32'b11111111111111101111101101011011;
assign LUT_2[6495] = 32'b11111111111111101100100101110100;
assign LUT_2[6496] = 32'b11111111111111110111011100111001;
assign LUT_2[6497] = 32'b11111111111111110100010101010010;
assign LUT_2[6498] = 32'b11111111111111111110010101110101;
assign LUT_2[6499] = 32'b11111111111111111011001110001110;
assign LUT_2[6500] = 32'b11111111111111110011111010100001;
assign LUT_2[6501] = 32'b11111111111111110000110010111010;
assign LUT_2[6502] = 32'b11111111111111111010110011011101;
assign LUT_2[6503] = 32'b11111111111111110111101011110110;
assign LUT_2[6504] = 32'b11111111111111110010001110010110;
assign LUT_2[6505] = 32'b11111111111111101111000110101111;
assign LUT_2[6506] = 32'b11111111111111111001000111010010;
assign LUT_2[6507] = 32'b11111111111111110101111111101011;
assign LUT_2[6508] = 32'b11111111111111101110101011111110;
assign LUT_2[6509] = 32'b11111111111111101011100100010111;
assign LUT_2[6510] = 32'b11111111111111110101100100111010;
assign LUT_2[6511] = 32'b11111111111111110010011101010011;
assign LUT_2[6512] = 32'b11111111111111110010000001000011;
assign LUT_2[6513] = 32'b11111111111111101110111001011100;
assign LUT_2[6514] = 32'b11111111111111111000111001111111;
assign LUT_2[6515] = 32'b11111111111111110101110010011000;
assign LUT_2[6516] = 32'b11111111111111101110011110101011;
assign LUT_2[6517] = 32'b11111111111111101011010111000100;
assign LUT_2[6518] = 32'b11111111111111110101010111100111;
assign LUT_2[6519] = 32'b11111111111111110010010000000000;
assign LUT_2[6520] = 32'b11111111111111101100110010100000;
assign LUT_2[6521] = 32'b11111111111111101001101010111001;
assign LUT_2[6522] = 32'b11111111111111110011101011011100;
assign LUT_2[6523] = 32'b11111111111111110000100011110101;
assign LUT_2[6524] = 32'b11111111111111101001010000001000;
assign LUT_2[6525] = 32'b11111111111111100110001000100001;
assign LUT_2[6526] = 32'b11111111111111110000001001000100;
assign LUT_2[6527] = 32'b11111111111111101101000001011101;
assign LUT_2[6528] = 32'b00000000000000000011001100111100;
assign LUT_2[6529] = 32'b00000000000000000000000101010101;
assign LUT_2[6530] = 32'b00000000000000001010000101111000;
assign LUT_2[6531] = 32'b00000000000000000110111110010001;
assign LUT_2[6532] = 32'b11111111111111111111101010100100;
assign LUT_2[6533] = 32'b11111111111111111100100010111101;
assign LUT_2[6534] = 32'b00000000000000000110100011100000;
assign LUT_2[6535] = 32'b00000000000000000011011011111001;
assign LUT_2[6536] = 32'b11111111111111111101111110011001;
assign LUT_2[6537] = 32'b11111111111111111010110110110010;
assign LUT_2[6538] = 32'b00000000000000000100110111010101;
assign LUT_2[6539] = 32'b00000000000000000001101111101110;
assign LUT_2[6540] = 32'b11111111111111111010011100000001;
assign LUT_2[6541] = 32'b11111111111111110111010100011010;
assign LUT_2[6542] = 32'b00000000000000000001010100111101;
assign LUT_2[6543] = 32'b11111111111111111110001101010110;
assign LUT_2[6544] = 32'b11111111111111111101110001000110;
assign LUT_2[6545] = 32'b11111111111111111010101001011111;
assign LUT_2[6546] = 32'b00000000000000000100101010000010;
assign LUT_2[6547] = 32'b00000000000000000001100010011011;
assign LUT_2[6548] = 32'b11111111111111111010001110101110;
assign LUT_2[6549] = 32'b11111111111111110111000111000111;
assign LUT_2[6550] = 32'b00000000000000000001000111101010;
assign LUT_2[6551] = 32'b11111111111111111110000000000011;
assign LUT_2[6552] = 32'b11111111111111111000100010100011;
assign LUT_2[6553] = 32'b11111111111111110101011010111100;
assign LUT_2[6554] = 32'b11111111111111111111011011011111;
assign LUT_2[6555] = 32'b11111111111111111100010011111000;
assign LUT_2[6556] = 32'b11111111111111110101000000001011;
assign LUT_2[6557] = 32'b11111111111111110001111000100100;
assign LUT_2[6558] = 32'b11111111111111111011111001000111;
assign LUT_2[6559] = 32'b11111111111111111000110001100000;
assign LUT_2[6560] = 32'b00000000000000000011101000100101;
assign LUT_2[6561] = 32'b00000000000000000000100000111110;
assign LUT_2[6562] = 32'b00000000000000001010100001100001;
assign LUT_2[6563] = 32'b00000000000000000111011001111010;
assign LUT_2[6564] = 32'b00000000000000000000000110001101;
assign LUT_2[6565] = 32'b11111111111111111100111110100110;
assign LUT_2[6566] = 32'b00000000000000000110111111001001;
assign LUT_2[6567] = 32'b00000000000000000011110111100010;
assign LUT_2[6568] = 32'b11111111111111111110011010000010;
assign LUT_2[6569] = 32'b11111111111111111011010010011011;
assign LUT_2[6570] = 32'b00000000000000000101010010111110;
assign LUT_2[6571] = 32'b00000000000000000010001011010111;
assign LUT_2[6572] = 32'b11111111111111111010110111101010;
assign LUT_2[6573] = 32'b11111111111111110111110000000011;
assign LUT_2[6574] = 32'b00000000000000000001110000100110;
assign LUT_2[6575] = 32'b11111111111111111110101000111111;
assign LUT_2[6576] = 32'b11111111111111111110001100101111;
assign LUT_2[6577] = 32'b11111111111111111011000101001000;
assign LUT_2[6578] = 32'b00000000000000000101000101101011;
assign LUT_2[6579] = 32'b00000000000000000001111110000100;
assign LUT_2[6580] = 32'b11111111111111111010101010010111;
assign LUT_2[6581] = 32'b11111111111111110111100010110000;
assign LUT_2[6582] = 32'b00000000000000000001100011010011;
assign LUT_2[6583] = 32'b11111111111111111110011011101100;
assign LUT_2[6584] = 32'b11111111111111111000111110001100;
assign LUT_2[6585] = 32'b11111111111111110101110110100101;
assign LUT_2[6586] = 32'b11111111111111111111110111001000;
assign LUT_2[6587] = 32'b11111111111111111100101111100001;
assign LUT_2[6588] = 32'b11111111111111110101011011110100;
assign LUT_2[6589] = 32'b11111111111111110010010100001101;
assign LUT_2[6590] = 32'b11111111111111111100010100110000;
assign LUT_2[6591] = 32'b11111111111111111001001101001001;
assign LUT_2[6592] = 32'b11111111111111111011010101011111;
assign LUT_2[6593] = 32'b11111111111111111000001101111000;
assign LUT_2[6594] = 32'b00000000000000000010001110011011;
assign LUT_2[6595] = 32'b11111111111111111111000110110100;
assign LUT_2[6596] = 32'b11111111111111110111110011000111;
assign LUT_2[6597] = 32'b11111111111111110100101011100000;
assign LUT_2[6598] = 32'b11111111111111111110101100000011;
assign LUT_2[6599] = 32'b11111111111111111011100100011100;
assign LUT_2[6600] = 32'b11111111111111110110000110111100;
assign LUT_2[6601] = 32'b11111111111111110010111111010101;
assign LUT_2[6602] = 32'b11111111111111111100111111111000;
assign LUT_2[6603] = 32'b11111111111111111001111000010001;
assign LUT_2[6604] = 32'b11111111111111110010100100100100;
assign LUT_2[6605] = 32'b11111111111111101111011100111101;
assign LUT_2[6606] = 32'b11111111111111111001011101100000;
assign LUT_2[6607] = 32'b11111111111111110110010101111001;
assign LUT_2[6608] = 32'b11111111111111110101111001101001;
assign LUT_2[6609] = 32'b11111111111111110010110010000010;
assign LUT_2[6610] = 32'b11111111111111111100110010100101;
assign LUT_2[6611] = 32'b11111111111111111001101010111110;
assign LUT_2[6612] = 32'b11111111111111110010010111010001;
assign LUT_2[6613] = 32'b11111111111111101111001111101010;
assign LUT_2[6614] = 32'b11111111111111111001010000001101;
assign LUT_2[6615] = 32'b11111111111111110110001000100110;
assign LUT_2[6616] = 32'b11111111111111110000101011000110;
assign LUT_2[6617] = 32'b11111111111111101101100011011111;
assign LUT_2[6618] = 32'b11111111111111110111100100000010;
assign LUT_2[6619] = 32'b11111111111111110100011100011011;
assign LUT_2[6620] = 32'b11111111111111101101001000101110;
assign LUT_2[6621] = 32'b11111111111111101010000001000111;
assign LUT_2[6622] = 32'b11111111111111110100000001101010;
assign LUT_2[6623] = 32'b11111111111111110000111010000011;
assign LUT_2[6624] = 32'b11111111111111111011110001001000;
assign LUT_2[6625] = 32'b11111111111111111000101001100001;
assign LUT_2[6626] = 32'b00000000000000000010101010000100;
assign LUT_2[6627] = 32'b11111111111111111111100010011101;
assign LUT_2[6628] = 32'b11111111111111111000001110110000;
assign LUT_2[6629] = 32'b11111111111111110101000111001001;
assign LUT_2[6630] = 32'b11111111111111111111000111101100;
assign LUT_2[6631] = 32'b11111111111111111100000000000101;
assign LUT_2[6632] = 32'b11111111111111110110100010100101;
assign LUT_2[6633] = 32'b11111111111111110011011010111110;
assign LUT_2[6634] = 32'b11111111111111111101011011100001;
assign LUT_2[6635] = 32'b11111111111111111010010011111010;
assign LUT_2[6636] = 32'b11111111111111110011000000001101;
assign LUT_2[6637] = 32'b11111111111111101111111000100110;
assign LUT_2[6638] = 32'b11111111111111111001111001001001;
assign LUT_2[6639] = 32'b11111111111111110110110001100010;
assign LUT_2[6640] = 32'b11111111111111110110010101010010;
assign LUT_2[6641] = 32'b11111111111111110011001101101011;
assign LUT_2[6642] = 32'b11111111111111111101001110001110;
assign LUT_2[6643] = 32'b11111111111111111010000110100111;
assign LUT_2[6644] = 32'b11111111111111110010110010111010;
assign LUT_2[6645] = 32'b11111111111111101111101011010011;
assign LUT_2[6646] = 32'b11111111111111111001101011110110;
assign LUT_2[6647] = 32'b11111111111111110110100100001111;
assign LUT_2[6648] = 32'b11111111111111110001000110101111;
assign LUT_2[6649] = 32'b11111111111111101101111111001000;
assign LUT_2[6650] = 32'b11111111111111110111111111101011;
assign LUT_2[6651] = 32'b11111111111111110100111000000100;
assign LUT_2[6652] = 32'b11111111111111101101100100010111;
assign LUT_2[6653] = 32'b11111111111111101010011100110000;
assign LUT_2[6654] = 32'b11111111111111110100011101010011;
assign LUT_2[6655] = 32'b11111111111111110001010101101100;
assign LUT_2[6656] = 32'b11111111111111111111101011111001;
assign LUT_2[6657] = 32'b11111111111111111100100100010010;
assign LUT_2[6658] = 32'b00000000000000000110100100110101;
assign LUT_2[6659] = 32'b00000000000000000011011101001110;
assign LUT_2[6660] = 32'b11111111111111111100001001100001;
assign LUT_2[6661] = 32'b11111111111111111001000001111010;
assign LUT_2[6662] = 32'b00000000000000000011000010011101;
assign LUT_2[6663] = 32'b11111111111111111111111010110110;
assign LUT_2[6664] = 32'b11111111111111111010011101010110;
assign LUT_2[6665] = 32'b11111111111111110111010101101111;
assign LUT_2[6666] = 32'b00000000000000000001010110010010;
assign LUT_2[6667] = 32'b11111111111111111110001110101011;
assign LUT_2[6668] = 32'b11111111111111110110111010111110;
assign LUT_2[6669] = 32'b11111111111111110011110011010111;
assign LUT_2[6670] = 32'b11111111111111111101110011111010;
assign LUT_2[6671] = 32'b11111111111111111010101100010011;
assign LUT_2[6672] = 32'b11111111111111111010010000000011;
assign LUT_2[6673] = 32'b11111111111111110111001000011100;
assign LUT_2[6674] = 32'b00000000000000000001001000111111;
assign LUT_2[6675] = 32'b11111111111111111110000001011000;
assign LUT_2[6676] = 32'b11111111111111110110101101101011;
assign LUT_2[6677] = 32'b11111111111111110011100110000100;
assign LUT_2[6678] = 32'b11111111111111111101100110100111;
assign LUT_2[6679] = 32'b11111111111111111010011111000000;
assign LUT_2[6680] = 32'b11111111111111110101000001100000;
assign LUT_2[6681] = 32'b11111111111111110001111001111001;
assign LUT_2[6682] = 32'b11111111111111111011111010011100;
assign LUT_2[6683] = 32'b11111111111111111000110010110101;
assign LUT_2[6684] = 32'b11111111111111110001011111001000;
assign LUT_2[6685] = 32'b11111111111111101110010111100001;
assign LUT_2[6686] = 32'b11111111111111111000011000000100;
assign LUT_2[6687] = 32'b11111111111111110101010000011101;
assign LUT_2[6688] = 32'b00000000000000000000000111100010;
assign LUT_2[6689] = 32'b11111111111111111100111111111011;
assign LUT_2[6690] = 32'b00000000000000000111000000011110;
assign LUT_2[6691] = 32'b00000000000000000011111000110111;
assign LUT_2[6692] = 32'b11111111111111111100100101001010;
assign LUT_2[6693] = 32'b11111111111111111001011101100011;
assign LUT_2[6694] = 32'b00000000000000000011011110000110;
assign LUT_2[6695] = 32'b00000000000000000000010110011111;
assign LUT_2[6696] = 32'b11111111111111111010111000111111;
assign LUT_2[6697] = 32'b11111111111111110111110001011000;
assign LUT_2[6698] = 32'b00000000000000000001110001111011;
assign LUT_2[6699] = 32'b11111111111111111110101010010100;
assign LUT_2[6700] = 32'b11111111111111110111010110100111;
assign LUT_2[6701] = 32'b11111111111111110100001111000000;
assign LUT_2[6702] = 32'b11111111111111111110001111100011;
assign LUT_2[6703] = 32'b11111111111111111011000111111100;
assign LUT_2[6704] = 32'b11111111111111111010101011101100;
assign LUT_2[6705] = 32'b11111111111111110111100100000101;
assign LUT_2[6706] = 32'b00000000000000000001100100101000;
assign LUT_2[6707] = 32'b11111111111111111110011101000001;
assign LUT_2[6708] = 32'b11111111111111110111001001010100;
assign LUT_2[6709] = 32'b11111111111111110100000001101101;
assign LUT_2[6710] = 32'b11111111111111111110000010010000;
assign LUT_2[6711] = 32'b11111111111111111010111010101001;
assign LUT_2[6712] = 32'b11111111111111110101011101001001;
assign LUT_2[6713] = 32'b11111111111111110010010101100010;
assign LUT_2[6714] = 32'b11111111111111111100010110000101;
assign LUT_2[6715] = 32'b11111111111111111001001110011110;
assign LUT_2[6716] = 32'b11111111111111110001111010110001;
assign LUT_2[6717] = 32'b11111111111111101110110011001010;
assign LUT_2[6718] = 32'b11111111111111111000110011101101;
assign LUT_2[6719] = 32'b11111111111111110101101100000110;
assign LUT_2[6720] = 32'b11111111111111110111110100011100;
assign LUT_2[6721] = 32'b11111111111111110100101100110101;
assign LUT_2[6722] = 32'b11111111111111111110101101011000;
assign LUT_2[6723] = 32'b11111111111111111011100101110001;
assign LUT_2[6724] = 32'b11111111111111110100010010000100;
assign LUT_2[6725] = 32'b11111111111111110001001010011101;
assign LUT_2[6726] = 32'b11111111111111111011001011000000;
assign LUT_2[6727] = 32'b11111111111111111000000011011001;
assign LUT_2[6728] = 32'b11111111111111110010100101111001;
assign LUT_2[6729] = 32'b11111111111111101111011110010010;
assign LUT_2[6730] = 32'b11111111111111111001011110110101;
assign LUT_2[6731] = 32'b11111111111111110110010111001110;
assign LUT_2[6732] = 32'b11111111111111101111000011100001;
assign LUT_2[6733] = 32'b11111111111111101011111011111010;
assign LUT_2[6734] = 32'b11111111111111110101111100011101;
assign LUT_2[6735] = 32'b11111111111111110010110100110110;
assign LUT_2[6736] = 32'b11111111111111110010011000100110;
assign LUT_2[6737] = 32'b11111111111111101111010000111111;
assign LUT_2[6738] = 32'b11111111111111111001010001100010;
assign LUT_2[6739] = 32'b11111111111111110110001001111011;
assign LUT_2[6740] = 32'b11111111111111101110110110001110;
assign LUT_2[6741] = 32'b11111111111111101011101110100111;
assign LUT_2[6742] = 32'b11111111111111110101101111001010;
assign LUT_2[6743] = 32'b11111111111111110010100111100011;
assign LUT_2[6744] = 32'b11111111111111101101001010000011;
assign LUT_2[6745] = 32'b11111111111111101010000010011100;
assign LUT_2[6746] = 32'b11111111111111110100000010111111;
assign LUT_2[6747] = 32'b11111111111111110000111011011000;
assign LUT_2[6748] = 32'b11111111111111101001100111101011;
assign LUT_2[6749] = 32'b11111111111111100110100000000100;
assign LUT_2[6750] = 32'b11111111111111110000100000100111;
assign LUT_2[6751] = 32'b11111111111111101101011001000000;
assign LUT_2[6752] = 32'b11111111111111111000010000000101;
assign LUT_2[6753] = 32'b11111111111111110101001000011110;
assign LUT_2[6754] = 32'b11111111111111111111001001000001;
assign LUT_2[6755] = 32'b11111111111111111100000001011010;
assign LUT_2[6756] = 32'b11111111111111110100101101101101;
assign LUT_2[6757] = 32'b11111111111111110001100110000110;
assign LUT_2[6758] = 32'b11111111111111111011100110101001;
assign LUT_2[6759] = 32'b11111111111111111000011111000010;
assign LUT_2[6760] = 32'b11111111111111110011000001100010;
assign LUT_2[6761] = 32'b11111111111111101111111001111011;
assign LUT_2[6762] = 32'b11111111111111111001111010011110;
assign LUT_2[6763] = 32'b11111111111111110110110010110111;
assign LUT_2[6764] = 32'b11111111111111101111011111001010;
assign LUT_2[6765] = 32'b11111111111111101100010111100011;
assign LUT_2[6766] = 32'b11111111111111110110011000000110;
assign LUT_2[6767] = 32'b11111111111111110011010000011111;
assign LUT_2[6768] = 32'b11111111111111110010110100001111;
assign LUT_2[6769] = 32'b11111111111111101111101100101000;
assign LUT_2[6770] = 32'b11111111111111111001101101001011;
assign LUT_2[6771] = 32'b11111111111111110110100101100100;
assign LUT_2[6772] = 32'b11111111111111101111010001110111;
assign LUT_2[6773] = 32'b11111111111111101100001010010000;
assign LUT_2[6774] = 32'b11111111111111110110001010110011;
assign LUT_2[6775] = 32'b11111111111111110011000011001100;
assign LUT_2[6776] = 32'b11111111111111101101100101101100;
assign LUT_2[6777] = 32'b11111111111111101010011110000101;
assign LUT_2[6778] = 32'b11111111111111110100011110101000;
assign LUT_2[6779] = 32'b11111111111111110001010111000001;
assign LUT_2[6780] = 32'b11111111111111101010000011010100;
assign LUT_2[6781] = 32'b11111111111111100110111011101101;
assign LUT_2[6782] = 32'b11111111111111110000111100010000;
assign LUT_2[6783] = 32'b11111111111111101101110100101001;
assign LUT_2[6784] = 32'b00000000000000000100000000001000;
assign LUT_2[6785] = 32'b00000000000000000000111000100001;
assign LUT_2[6786] = 32'b00000000000000001010111001000100;
assign LUT_2[6787] = 32'b00000000000000000111110001011101;
assign LUT_2[6788] = 32'b00000000000000000000011101110000;
assign LUT_2[6789] = 32'b11111111111111111101010110001001;
assign LUT_2[6790] = 32'b00000000000000000111010110101100;
assign LUT_2[6791] = 32'b00000000000000000100001111000101;
assign LUT_2[6792] = 32'b11111111111111111110110001100101;
assign LUT_2[6793] = 32'b11111111111111111011101001111110;
assign LUT_2[6794] = 32'b00000000000000000101101010100001;
assign LUT_2[6795] = 32'b00000000000000000010100010111010;
assign LUT_2[6796] = 32'b11111111111111111011001111001101;
assign LUT_2[6797] = 32'b11111111111111111000000111100110;
assign LUT_2[6798] = 32'b00000000000000000010001000001001;
assign LUT_2[6799] = 32'b11111111111111111111000000100010;
assign LUT_2[6800] = 32'b11111111111111111110100100010010;
assign LUT_2[6801] = 32'b11111111111111111011011100101011;
assign LUT_2[6802] = 32'b00000000000000000101011101001110;
assign LUT_2[6803] = 32'b00000000000000000010010101100111;
assign LUT_2[6804] = 32'b11111111111111111011000001111010;
assign LUT_2[6805] = 32'b11111111111111110111111010010011;
assign LUT_2[6806] = 32'b00000000000000000001111010110110;
assign LUT_2[6807] = 32'b11111111111111111110110011001111;
assign LUT_2[6808] = 32'b11111111111111111001010101101111;
assign LUT_2[6809] = 32'b11111111111111110110001110001000;
assign LUT_2[6810] = 32'b00000000000000000000001110101011;
assign LUT_2[6811] = 32'b11111111111111111101000111000100;
assign LUT_2[6812] = 32'b11111111111111110101110011010111;
assign LUT_2[6813] = 32'b11111111111111110010101011110000;
assign LUT_2[6814] = 32'b11111111111111111100101100010011;
assign LUT_2[6815] = 32'b11111111111111111001100100101100;
assign LUT_2[6816] = 32'b00000000000000000100011011110001;
assign LUT_2[6817] = 32'b00000000000000000001010100001010;
assign LUT_2[6818] = 32'b00000000000000001011010100101101;
assign LUT_2[6819] = 32'b00000000000000001000001101000110;
assign LUT_2[6820] = 32'b00000000000000000000111001011001;
assign LUT_2[6821] = 32'b11111111111111111101110001110010;
assign LUT_2[6822] = 32'b00000000000000000111110010010101;
assign LUT_2[6823] = 32'b00000000000000000100101010101110;
assign LUT_2[6824] = 32'b11111111111111111111001101001110;
assign LUT_2[6825] = 32'b11111111111111111100000101100111;
assign LUT_2[6826] = 32'b00000000000000000110000110001010;
assign LUT_2[6827] = 32'b00000000000000000010111110100011;
assign LUT_2[6828] = 32'b11111111111111111011101010110110;
assign LUT_2[6829] = 32'b11111111111111111000100011001111;
assign LUT_2[6830] = 32'b00000000000000000010100011110010;
assign LUT_2[6831] = 32'b11111111111111111111011100001011;
assign LUT_2[6832] = 32'b11111111111111111110111111111011;
assign LUT_2[6833] = 32'b11111111111111111011111000010100;
assign LUT_2[6834] = 32'b00000000000000000101111000110111;
assign LUT_2[6835] = 32'b00000000000000000010110001010000;
assign LUT_2[6836] = 32'b11111111111111111011011101100011;
assign LUT_2[6837] = 32'b11111111111111111000010101111100;
assign LUT_2[6838] = 32'b00000000000000000010010110011111;
assign LUT_2[6839] = 32'b11111111111111111111001110111000;
assign LUT_2[6840] = 32'b11111111111111111001110001011000;
assign LUT_2[6841] = 32'b11111111111111110110101001110001;
assign LUT_2[6842] = 32'b00000000000000000000101010010100;
assign LUT_2[6843] = 32'b11111111111111111101100010101101;
assign LUT_2[6844] = 32'b11111111111111110110001111000000;
assign LUT_2[6845] = 32'b11111111111111110011000111011001;
assign LUT_2[6846] = 32'b11111111111111111101000111111100;
assign LUT_2[6847] = 32'b11111111111111111010000000010101;
assign LUT_2[6848] = 32'b11111111111111111100001000101011;
assign LUT_2[6849] = 32'b11111111111111111001000001000100;
assign LUT_2[6850] = 32'b00000000000000000011000001100111;
assign LUT_2[6851] = 32'b11111111111111111111111010000000;
assign LUT_2[6852] = 32'b11111111111111111000100110010011;
assign LUT_2[6853] = 32'b11111111111111110101011110101100;
assign LUT_2[6854] = 32'b11111111111111111111011111001111;
assign LUT_2[6855] = 32'b11111111111111111100010111101000;
assign LUT_2[6856] = 32'b11111111111111110110111010001000;
assign LUT_2[6857] = 32'b11111111111111110011110010100001;
assign LUT_2[6858] = 32'b11111111111111111101110011000100;
assign LUT_2[6859] = 32'b11111111111111111010101011011101;
assign LUT_2[6860] = 32'b11111111111111110011010111110000;
assign LUT_2[6861] = 32'b11111111111111110000010000001001;
assign LUT_2[6862] = 32'b11111111111111111010010000101100;
assign LUT_2[6863] = 32'b11111111111111110111001001000101;
assign LUT_2[6864] = 32'b11111111111111110110101100110101;
assign LUT_2[6865] = 32'b11111111111111110011100101001110;
assign LUT_2[6866] = 32'b11111111111111111101100101110001;
assign LUT_2[6867] = 32'b11111111111111111010011110001010;
assign LUT_2[6868] = 32'b11111111111111110011001010011101;
assign LUT_2[6869] = 32'b11111111111111110000000010110110;
assign LUT_2[6870] = 32'b11111111111111111010000011011001;
assign LUT_2[6871] = 32'b11111111111111110110111011110010;
assign LUT_2[6872] = 32'b11111111111111110001011110010010;
assign LUT_2[6873] = 32'b11111111111111101110010110101011;
assign LUT_2[6874] = 32'b11111111111111111000010111001110;
assign LUT_2[6875] = 32'b11111111111111110101001111100111;
assign LUT_2[6876] = 32'b11111111111111101101111011111010;
assign LUT_2[6877] = 32'b11111111111111101010110100010011;
assign LUT_2[6878] = 32'b11111111111111110100110100110110;
assign LUT_2[6879] = 32'b11111111111111110001101101001111;
assign LUT_2[6880] = 32'b11111111111111111100100100010100;
assign LUT_2[6881] = 32'b11111111111111111001011100101101;
assign LUT_2[6882] = 32'b00000000000000000011011101010000;
assign LUT_2[6883] = 32'b00000000000000000000010101101001;
assign LUT_2[6884] = 32'b11111111111111111001000001111100;
assign LUT_2[6885] = 32'b11111111111111110101111010010101;
assign LUT_2[6886] = 32'b11111111111111111111111010111000;
assign LUT_2[6887] = 32'b11111111111111111100110011010001;
assign LUT_2[6888] = 32'b11111111111111110111010101110001;
assign LUT_2[6889] = 32'b11111111111111110100001110001010;
assign LUT_2[6890] = 32'b11111111111111111110001110101101;
assign LUT_2[6891] = 32'b11111111111111111011000111000110;
assign LUT_2[6892] = 32'b11111111111111110011110011011001;
assign LUT_2[6893] = 32'b11111111111111110000101011110010;
assign LUT_2[6894] = 32'b11111111111111111010101100010101;
assign LUT_2[6895] = 32'b11111111111111110111100100101110;
assign LUT_2[6896] = 32'b11111111111111110111001000011110;
assign LUT_2[6897] = 32'b11111111111111110100000000110111;
assign LUT_2[6898] = 32'b11111111111111111110000001011010;
assign LUT_2[6899] = 32'b11111111111111111010111001110011;
assign LUT_2[6900] = 32'b11111111111111110011100110000110;
assign LUT_2[6901] = 32'b11111111111111110000011110011111;
assign LUT_2[6902] = 32'b11111111111111111010011111000010;
assign LUT_2[6903] = 32'b11111111111111110111010111011011;
assign LUT_2[6904] = 32'b11111111111111110001111001111011;
assign LUT_2[6905] = 32'b11111111111111101110110010010100;
assign LUT_2[6906] = 32'b11111111111111111000110010110111;
assign LUT_2[6907] = 32'b11111111111111110101101011010000;
assign LUT_2[6908] = 32'b11111111111111101110010111100011;
assign LUT_2[6909] = 32'b11111111111111101011001111111100;
assign LUT_2[6910] = 32'b11111111111111110101010000011111;
assign LUT_2[6911] = 32'b11111111111111110010001000111000;
assign LUT_2[6912] = 32'b00000000000000000011101010011111;
assign LUT_2[6913] = 32'b00000000000000000000100010111000;
assign LUT_2[6914] = 32'b00000000000000001010100011011011;
assign LUT_2[6915] = 32'b00000000000000000111011011110100;
assign LUT_2[6916] = 32'b00000000000000000000001000000111;
assign LUT_2[6917] = 32'b11111111111111111101000000100000;
assign LUT_2[6918] = 32'b00000000000000000111000001000011;
assign LUT_2[6919] = 32'b00000000000000000011111001011100;
assign LUT_2[6920] = 32'b11111111111111111110011011111100;
assign LUT_2[6921] = 32'b11111111111111111011010100010101;
assign LUT_2[6922] = 32'b00000000000000000101010100111000;
assign LUT_2[6923] = 32'b00000000000000000010001101010001;
assign LUT_2[6924] = 32'b11111111111111111010111001100100;
assign LUT_2[6925] = 32'b11111111111111110111110001111101;
assign LUT_2[6926] = 32'b00000000000000000001110010100000;
assign LUT_2[6927] = 32'b11111111111111111110101010111001;
assign LUT_2[6928] = 32'b11111111111111111110001110101001;
assign LUT_2[6929] = 32'b11111111111111111011000111000010;
assign LUT_2[6930] = 32'b00000000000000000101000111100101;
assign LUT_2[6931] = 32'b00000000000000000001111111111110;
assign LUT_2[6932] = 32'b11111111111111111010101100010001;
assign LUT_2[6933] = 32'b11111111111111110111100100101010;
assign LUT_2[6934] = 32'b00000000000000000001100101001101;
assign LUT_2[6935] = 32'b11111111111111111110011101100110;
assign LUT_2[6936] = 32'b11111111111111111001000000000110;
assign LUT_2[6937] = 32'b11111111111111110101111000011111;
assign LUT_2[6938] = 32'b11111111111111111111111001000010;
assign LUT_2[6939] = 32'b11111111111111111100110001011011;
assign LUT_2[6940] = 32'b11111111111111110101011101101110;
assign LUT_2[6941] = 32'b11111111111111110010010110000111;
assign LUT_2[6942] = 32'b11111111111111111100010110101010;
assign LUT_2[6943] = 32'b11111111111111111001001111000011;
assign LUT_2[6944] = 32'b00000000000000000100000110001000;
assign LUT_2[6945] = 32'b00000000000000000000111110100001;
assign LUT_2[6946] = 32'b00000000000000001010111111000100;
assign LUT_2[6947] = 32'b00000000000000000111110111011101;
assign LUT_2[6948] = 32'b00000000000000000000100011110000;
assign LUT_2[6949] = 32'b11111111111111111101011100001001;
assign LUT_2[6950] = 32'b00000000000000000111011100101100;
assign LUT_2[6951] = 32'b00000000000000000100010101000101;
assign LUT_2[6952] = 32'b11111111111111111110110111100101;
assign LUT_2[6953] = 32'b11111111111111111011101111111110;
assign LUT_2[6954] = 32'b00000000000000000101110000100001;
assign LUT_2[6955] = 32'b00000000000000000010101000111010;
assign LUT_2[6956] = 32'b11111111111111111011010101001101;
assign LUT_2[6957] = 32'b11111111111111111000001101100110;
assign LUT_2[6958] = 32'b00000000000000000010001110001001;
assign LUT_2[6959] = 32'b11111111111111111111000110100010;
assign LUT_2[6960] = 32'b11111111111111111110101010010010;
assign LUT_2[6961] = 32'b11111111111111111011100010101011;
assign LUT_2[6962] = 32'b00000000000000000101100011001110;
assign LUT_2[6963] = 32'b00000000000000000010011011100111;
assign LUT_2[6964] = 32'b11111111111111111011000111111010;
assign LUT_2[6965] = 32'b11111111111111111000000000010011;
assign LUT_2[6966] = 32'b00000000000000000010000000110110;
assign LUT_2[6967] = 32'b11111111111111111110111001001111;
assign LUT_2[6968] = 32'b11111111111111111001011011101111;
assign LUT_2[6969] = 32'b11111111111111110110010100001000;
assign LUT_2[6970] = 32'b00000000000000000000010100101011;
assign LUT_2[6971] = 32'b11111111111111111101001101000100;
assign LUT_2[6972] = 32'b11111111111111110101111001010111;
assign LUT_2[6973] = 32'b11111111111111110010110001110000;
assign LUT_2[6974] = 32'b11111111111111111100110010010011;
assign LUT_2[6975] = 32'b11111111111111111001101010101100;
assign LUT_2[6976] = 32'b11111111111111111011110011000010;
assign LUT_2[6977] = 32'b11111111111111111000101011011011;
assign LUT_2[6978] = 32'b00000000000000000010101011111110;
assign LUT_2[6979] = 32'b11111111111111111111100100010111;
assign LUT_2[6980] = 32'b11111111111111111000010000101010;
assign LUT_2[6981] = 32'b11111111111111110101001001000011;
assign LUT_2[6982] = 32'b11111111111111111111001001100110;
assign LUT_2[6983] = 32'b11111111111111111100000001111111;
assign LUT_2[6984] = 32'b11111111111111110110100100011111;
assign LUT_2[6985] = 32'b11111111111111110011011100111000;
assign LUT_2[6986] = 32'b11111111111111111101011101011011;
assign LUT_2[6987] = 32'b11111111111111111010010101110100;
assign LUT_2[6988] = 32'b11111111111111110011000010000111;
assign LUT_2[6989] = 32'b11111111111111101111111010100000;
assign LUT_2[6990] = 32'b11111111111111111001111011000011;
assign LUT_2[6991] = 32'b11111111111111110110110011011100;
assign LUT_2[6992] = 32'b11111111111111110110010111001100;
assign LUT_2[6993] = 32'b11111111111111110011001111100101;
assign LUT_2[6994] = 32'b11111111111111111101010000001000;
assign LUT_2[6995] = 32'b11111111111111111010001000100001;
assign LUT_2[6996] = 32'b11111111111111110010110100110100;
assign LUT_2[6997] = 32'b11111111111111101111101101001101;
assign LUT_2[6998] = 32'b11111111111111111001101101110000;
assign LUT_2[6999] = 32'b11111111111111110110100110001001;
assign LUT_2[7000] = 32'b11111111111111110001001000101001;
assign LUT_2[7001] = 32'b11111111111111101110000001000010;
assign LUT_2[7002] = 32'b11111111111111111000000001100101;
assign LUT_2[7003] = 32'b11111111111111110100111001111110;
assign LUT_2[7004] = 32'b11111111111111101101100110010001;
assign LUT_2[7005] = 32'b11111111111111101010011110101010;
assign LUT_2[7006] = 32'b11111111111111110100011111001101;
assign LUT_2[7007] = 32'b11111111111111110001010111100110;
assign LUT_2[7008] = 32'b11111111111111111100001110101011;
assign LUT_2[7009] = 32'b11111111111111111001000111000100;
assign LUT_2[7010] = 32'b00000000000000000011000111100111;
assign LUT_2[7011] = 32'b00000000000000000000000000000000;
assign LUT_2[7012] = 32'b11111111111111111000101100010011;
assign LUT_2[7013] = 32'b11111111111111110101100100101100;
assign LUT_2[7014] = 32'b11111111111111111111100101001111;
assign LUT_2[7015] = 32'b11111111111111111100011101101000;
assign LUT_2[7016] = 32'b11111111111111110111000000001000;
assign LUT_2[7017] = 32'b11111111111111110011111000100001;
assign LUT_2[7018] = 32'b11111111111111111101111001000100;
assign LUT_2[7019] = 32'b11111111111111111010110001011101;
assign LUT_2[7020] = 32'b11111111111111110011011101110000;
assign LUT_2[7021] = 32'b11111111111111110000010110001001;
assign LUT_2[7022] = 32'b11111111111111111010010110101100;
assign LUT_2[7023] = 32'b11111111111111110111001111000101;
assign LUT_2[7024] = 32'b11111111111111110110110010110101;
assign LUT_2[7025] = 32'b11111111111111110011101011001110;
assign LUT_2[7026] = 32'b11111111111111111101101011110001;
assign LUT_2[7027] = 32'b11111111111111111010100100001010;
assign LUT_2[7028] = 32'b11111111111111110011010000011101;
assign LUT_2[7029] = 32'b11111111111111110000001000110110;
assign LUT_2[7030] = 32'b11111111111111111010001001011001;
assign LUT_2[7031] = 32'b11111111111111110111000001110010;
assign LUT_2[7032] = 32'b11111111111111110001100100010010;
assign LUT_2[7033] = 32'b11111111111111101110011100101011;
assign LUT_2[7034] = 32'b11111111111111111000011101001110;
assign LUT_2[7035] = 32'b11111111111111110101010101100111;
assign LUT_2[7036] = 32'b11111111111111101110000001111010;
assign LUT_2[7037] = 32'b11111111111111101010111010010011;
assign LUT_2[7038] = 32'b11111111111111110100111010110110;
assign LUT_2[7039] = 32'b11111111111111110001110011001111;
assign LUT_2[7040] = 32'b00000000000000000111111110101110;
assign LUT_2[7041] = 32'b00000000000000000100110111000111;
assign LUT_2[7042] = 32'b00000000000000001110110111101010;
assign LUT_2[7043] = 32'b00000000000000001011110000000011;
assign LUT_2[7044] = 32'b00000000000000000100011100010110;
assign LUT_2[7045] = 32'b00000000000000000001010100101111;
assign LUT_2[7046] = 32'b00000000000000001011010101010010;
assign LUT_2[7047] = 32'b00000000000000001000001101101011;
assign LUT_2[7048] = 32'b00000000000000000010110000001011;
assign LUT_2[7049] = 32'b11111111111111111111101000100100;
assign LUT_2[7050] = 32'b00000000000000001001101001000111;
assign LUT_2[7051] = 32'b00000000000000000110100001100000;
assign LUT_2[7052] = 32'b11111111111111111111001101110011;
assign LUT_2[7053] = 32'b11111111111111111100000110001100;
assign LUT_2[7054] = 32'b00000000000000000110000110101111;
assign LUT_2[7055] = 32'b00000000000000000010111111001000;
assign LUT_2[7056] = 32'b00000000000000000010100010111000;
assign LUT_2[7057] = 32'b11111111111111111111011011010001;
assign LUT_2[7058] = 32'b00000000000000001001011011110100;
assign LUT_2[7059] = 32'b00000000000000000110010100001101;
assign LUT_2[7060] = 32'b11111111111111111111000000100000;
assign LUT_2[7061] = 32'b11111111111111111011111000111001;
assign LUT_2[7062] = 32'b00000000000000000101111001011100;
assign LUT_2[7063] = 32'b00000000000000000010110001110101;
assign LUT_2[7064] = 32'b11111111111111111101010100010101;
assign LUT_2[7065] = 32'b11111111111111111010001100101110;
assign LUT_2[7066] = 32'b00000000000000000100001101010001;
assign LUT_2[7067] = 32'b00000000000000000001000101101010;
assign LUT_2[7068] = 32'b11111111111111111001110001111101;
assign LUT_2[7069] = 32'b11111111111111110110101010010110;
assign LUT_2[7070] = 32'b00000000000000000000101010111001;
assign LUT_2[7071] = 32'b11111111111111111101100011010010;
assign LUT_2[7072] = 32'b00000000000000001000011010010111;
assign LUT_2[7073] = 32'b00000000000000000101010010110000;
assign LUT_2[7074] = 32'b00000000000000001111010011010011;
assign LUT_2[7075] = 32'b00000000000000001100001011101100;
assign LUT_2[7076] = 32'b00000000000000000100110111111111;
assign LUT_2[7077] = 32'b00000000000000000001110000011000;
assign LUT_2[7078] = 32'b00000000000000001011110000111011;
assign LUT_2[7079] = 32'b00000000000000001000101001010100;
assign LUT_2[7080] = 32'b00000000000000000011001011110100;
assign LUT_2[7081] = 32'b00000000000000000000000100001101;
assign LUT_2[7082] = 32'b00000000000000001010000100110000;
assign LUT_2[7083] = 32'b00000000000000000110111101001001;
assign LUT_2[7084] = 32'b11111111111111111111101001011100;
assign LUT_2[7085] = 32'b11111111111111111100100001110101;
assign LUT_2[7086] = 32'b00000000000000000110100010011000;
assign LUT_2[7087] = 32'b00000000000000000011011010110001;
assign LUT_2[7088] = 32'b00000000000000000010111110100001;
assign LUT_2[7089] = 32'b11111111111111111111110110111010;
assign LUT_2[7090] = 32'b00000000000000001001110111011101;
assign LUT_2[7091] = 32'b00000000000000000110101111110110;
assign LUT_2[7092] = 32'b11111111111111111111011100001001;
assign LUT_2[7093] = 32'b11111111111111111100010100100010;
assign LUT_2[7094] = 32'b00000000000000000110010101000101;
assign LUT_2[7095] = 32'b00000000000000000011001101011110;
assign LUT_2[7096] = 32'b11111111111111111101101111111110;
assign LUT_2[7097] = 32'b11111111111111111010101000010111;
assign LUT_2[7098] = 32'b00000000000000000100101000111010;
assign LUT_2[7099] = 32'b00000000000000000001100001010011;
assign LUT_2[7100] = 32'b11111111111111111010001101100110;
assign LUT_2[7101] = 32'b11111111111111110111000101111111;
assign LUT_2[7102] = 32'b00000000000000000001000110100010;
assign LUT_2[7103] = 32'b11111111111111111101111110111011;
assign LUT_2[7104] = 32'b00000000000000000000000111010001;
assign LUT_2[7105] = 32'b11111111111111111100111111101010;
assign LUT_2[7106] = 32'b00000000000000000111000000001101;
assign LUT_2[7107] = 32'b00000000000000000011111000100110;
assign LUT_2[7108] = 32'b11111111111111111100100100111001;
assign LUT_2[7109] = 32'b11111111111111111001011101010010;
assign LUT_2[7110] = 32'b00000000000000000011011101110101;
assign LUT_2[7111] = 32'b00000000000000000000010110001110;
assign LUT_2[7112] = 32'b11111111111111111010111000101110;
assign LUT_2[7113] = 32'b11111111111111110111110001000111;
assign LUT_2[7114] = 32'b00000000000000000001110001101010;
assign LUT_2[7115] = 32'b11111111111111111110101010000011;
assign LUT_2[7116] = 32'b11111111111111110111010110010110;
assign LUT_2[7117] = 32'b11111111111111110100001110101111;
assign LUT_2[7118] = 32'b11111111111111111110001111010010;
assign LUT_2[7119] = 32'b11111111111111111011000111101011;
assign LUT_2[7120] = 32'b11111111111111111010101011011011;
assign LUT_2[7121] = 32'b11111111111111110111100011110100;
assign LUT_2[7122] = 32'b00000000000000000001100100010111;
assign LUT_2[7123] = 32'b11111111111111111110011100110000;
assign LUT_2[7124] = 32'b11111111111111110111001001000011;
assign LUT_2[7125] = 32'b11111111111111110100000001011100;
assign LUT_2[7126] = 32'b11111111111111111110000001111111;
assign LUT_2[7127] = 32'b11111111111111111010111010011000;
assign LUT_2[7128] = 32'b11111111111111110101011100111000;
assign LUT_2[7129] = 32'b11111111111111110010010101010001;
assign LUT_2[7130] = 32'b11111111111111111100010101110100;
assign LUT_2[7131] = 32'b11111111111111111001001110001101;
assign LUT_2[7132] = 32'b11111111111111110001111010100000;
assign LUT_2[7133] = 32'b11111111111111101110110010111001;
assign LUT_2[7134] = 32'b11111111111111111000110011011100;
assign LUT_2[7135] = 32'b11111111111111110101101011110101;
assign LUT_2[7136] = 32'b00000000000000000000100010111010;
assign LUT_2[7137] = 32'b11111111111111111101011011010011;
assign LUT_2[7138] = 32'b00000000000000000111011011110110;
assign LUT_2[7139] = 32'b00000000000000000100010100001111;
assign LUT_2[7140] = 32'b11111111111111111101000000100010;
assign LUT_2[7141] = 32'b11111111111111111001111000111011;
assign LUT_2[7142] = 32'b00000000000000000011111001011110;
assign LUT_2[7143] = 32'b00000000000000000000110001110111;
assign LUT_2[7144] = 32'b11111111111111111011010100010111;
assign LUT_2[7145] = 32'b11111111111111111000001100110000;
assign LUT_2[7146] = 32'b00000000000000000010001101010011;
assign LUT_2[7147] = 32'b11111111111111111111000101101100;
assign LUT_2[7148] = 32'b11111111111111110111110001111111;
assign LUT_2[7149] = 32'b11111111111111110100101010011000;
assign LUT_2[7150] = 32'b11111111111111111110101010111011;
assign LUT_2[7151] = 32'b11111111111111111011100011010100;
assign LUT_2[7152] = 32'b11111111111111111011000111000100;
assign LUT_2[7153] = 32'b11111111111111110111111111011101;
assign LUT_2[7154] = 32'b00000000000000000010000000000000;
assign LUT_2[7155] = 32'b11111111111111111110111000011001;
assign LUT_2[7156] = 32'b11111111111111110111100100101100;
assign LUT_2[7157] = 32'b11111111111111110100011101000101;
assign LUT_2[7158] = 32'b11111111111111111110011101101000;
assign LUT_2[7159] = 32'b11111111111111111011010110000001;
assign LUT_2[7160] = 32'b11111111111111110101111000100001;
assign LUT_2[7161] = 32'b11111111111111110010110000111010;
assign LUT_2[7162] = 32'b11111111111111111100110001011101;
assign LUT_2[7163] = 32'b11111111111111111001101001110110;
assign LUT_2[7164] = 32'b11111111111111110010010110001001;
assign LUT_2[7165] = 32'b11111111111111101111001110100010;
assign LUT_2[7166] = 32'b11111111111111111001001111000101;
assign LUT_2[7167] = 32'b11111111111111110110000111011110;
assign LUT_2[7168] = 32'b00000000000000000001100110001100;
assign LUT_2[7169] = 32'b11111111111111111110011110100101;
assign LUT_2[7170] = 32'b00000000000000001000011111001000;
assign LUT_2[7171] = 32'b00000000000000000101010111100001;
assign LUT_2[7172] = 32'b11111111111111111110000011110100;
assign LUT_2[7173] = 32'b11111111111111111010111100001101;
assign LUT_2[7174] = 32'b00000000000000000100111100110000;
assign LUT_2[7175] = 32'b00000000000000000001110101001001;
assign LUT_2[7176] = 32'b11111111111111111100010111101001;
assign LUT_2[7177] = 32'b11111111111111111001010000000010;
assign LUT_2[7178] = 32'b00000000000000000011010000100101;
assign LUT_2[7179] = 32'b00000000000000000000001000111110;
assign LUT_2[7180] = 32'b11111111111111111000110101010001;
assign LUT_2[7181] = 32'b11111111111111110101101101101010;
assign LUT_2[7182] = 32'b11111111111111111111101110001101;
assign LUT_2[7183] = 32'b11111111111111111100100110100110;
assign LUT_2[7184] = 32'b11111111111111111100001010010110;
assign LUT_2[7185] = 32'b11111111111111111001000010101111;
assign LUT_2[7186] = 32'b00000000000000000011000011010010;
assign LUT_2[7187] = 32'b11111111111111111111111011101011;
assign LUT_2[7188] = 32'b11111111111111111000100111111110;
assign LUT_2[7189] = 32'b11111111111111110101100000010111;
assign LUT_2[7190] = 32'b11111111111111111111100000111010;
assign LUT_2[7191] = 32'b11111111111111111100011001010011;
assign LUT_2[7192] = 32'b11111111111111110110111011110011;
assign LUT_2[7193] = 32'b11111111111111110011110100001100;
assign LUT_2[7194] = 32'b11111111111111111101110100101111;
assign LUT_2[7195] = 32'b11111111111111111010101101001000;
assign LUT_2[7196] = 32'b11111111111111110011011001011011;
assign LUT_2[7197] = 32'b11111111111111110000010001110100;
assign LUT_2[7198] = 32'b11111111111111111010010010010111;
assign LUT_2[7199] = 32'b11111111111111110111001010110000;
assign LUT_2[7200] = 32'b00000000000000000010000001110101;
assign LUT_2[7201] = 32'b11111111111111111110111010001110;
assign LUT_2[7202] = 32'b00000000000000001000111010110001;
assign LUT_2[7203] = 32'b00000000000000000101110011001010;
assign LUT_2[7204] = 32'b11111111111111111110011111011101;
assign LUT_2[7205] = 32'b11111111111111111011010111110110;
assign LUT_2[7206] = 32'b00000000000000000101011000011001;
assign LUT_2[7207] = 32'b00000000000000000010010000110010;
assign LUT_2[7208] = 32'b11111111111111111100110011010010;
assign LUT_2[7209] = 32'b11111111111111111001101011101011;
assign LUT_2[7210] = 32'b00000000000000000011101100001110;
assign LUT_2[7211] = 32'b00000000000000000000100100100111;
assign LUT_2[7212] = 32'b11111111111111111001010000111010;
assign LUT_2[7213] = 32'b11111111111111110110001001010011;
assign LUT_2[7214] = 32'b00000000000000000000001001110110;
assign LUT_2[7215] = 32'b11111111111111111101000010001111;
assign LUT_2[7216] = 32'b11111111111111111100100101111111;
assign LUT_2[7217] = 32'b11111111111111111001011110011000;
assign LUT_2[7218] = 32'b00000000000000000011011110111011;
assign LUT_2[7219] = 32'b00000000000000000000010111010100;
assign LUT_2[7220] = 32'b11111111111111111001000011100111;
assign LUT_2[7221] = 32'b11111111111111110101111100000000;
assign LUT_2[7222] = 32'b11111111111111111111111100100011;
assign LUT_2[7223] = 32'b11111111111111111100110100111100;
assign LUT_2[7224] = 32'b11111111111111110111010111011100;
assign LUT_2[7225] = 32'b11111111111111110100001111110101;
assign LUT_2[7226] = 32'b11111111111111111110010000011000;
assign LUT_2[7227] = 32'b11111111111111111011001000110001;
assign LUT_2[7228] = 32'b11111111111111110011110101000100;
assign LUT_2[7229] = 32'b11111111111111110000101101011101;
assign LUT_2[7230] = 32'b11111111111111111010101110000000;
assign LUT_2[7231] = 32'b11111111111111110111100110011001;
assign LUT_2[7232] = 32'b11111111111111111001101110101111;
assign LUT_2[7233] = 32'b11111111111111110110100111001000;
assign LUT_2[7234] = 32'b00000000000000000000100111101011;
assign LUT_2[7235] = 32'b11111111111111111101100000000100;
assign LUT_2[7236] = 32'b11111111111111110110001100010111;
assign LUT_2[7237] = 32'b11111111111111110011000100110000;
assign LUT_2[7238] = 32'b11111111111111111101000101010011;
assign LUT_2[7239] = 32'b11111111111111111001111101101100;
assign LUT_2[7240] = 32'b11111111111111110100100000001100;
assign LUT_2[7241] = 32'b11111111111111110001011000100101;
assign LUT_2[7242] = 32'b11111111111111111011011001001000;
assign LUT_2[7243] = 32'b11111111111111111000010001100001;
assign LUT_2[7244] = 32'b11111111111111110000111101110100;
assign LUT_2[7245] = 32'b11111111111111101101110110001101;
assign LUT_2[7246] = 32'b11111111111111110111110110110000;
assign LUT_2[7247] = 32'b11111111111111110100101111001001;
assign LUT_2[7248] = 32'b11111111111111110100010010111001;
assign LUT_2[7249] = 32'b11111111111111110001001011010010;
assign LUT_2[7250] = 32'b11111111111111111011001011110101;
assign LUT_2[7251] = 32'b11111111111111111000000100001110;
assign LUT_2[7252] = 32'b11111111111111110000110000100001;
assign LUT_2[7253] = 32'b11111111111111101101101000111010;
assign LUT_2[7254] = 32'b11111111111111110111101001011101;
assign LUT_2[7255] = 32'b11111111111111110100100001110110;
assign LUT_2[7256] = 32'b11111111111111101111000100010110;
assign LUT_2[7257] = 32'b11111111111111101011111100101111;
assign LUT_2[7258] = 32'b11111111111111110101111101010010;
assign LUT_2[7259] = 32'b11111111111111110010110101101011;
assign LUT_2[7260] = 32'b11111111111111101011100001111110;
assign LUT_2[7261] = 32'b11111111111111101000011010010111;
assign LUT_2[7262] = 32'b11111111111111110010011010111010;
assign LUT_2[7263] = 32'b11111111111111101111010011010011;
assign LUT_2[7264] = 32'b11111111111111111010001010011000;
assign LUT_2[7265] = 32'b11111111111111110111000010110001;
assign LUT_2[7266] = 32'b00000000000000000001000011010100;
assign LUT_2[7267] = 32'b11111111111111111101111011101101;
assign LUT_2[7268] = 32'b11111111111111110110101000000000;
assign LUT_2[7269] = 32'b11111111111111110011100000011001;
assign LUT_2[7270] = 32'b11111111111111111101100000111100;
assign LUT_2[7271] = 32'b11111111111111111010011001010101;
assign LUT_2[7272] = 32'b11111111111111110100111011110101;
assign LUT_2[7273] = 32'b11111111111111110001110100001110;
assign LUT_2[7274] = 32'b11111111111111111011110100110001;
assign LUT_2[7275] = 32'b11111111111111111000101101001010;
assign LUT_2[7276] = 32'b11111111111111110001011001011101;
assign LUT_2[7277] = 32'b11111111111111101110010001110110;
assign LUT_2[7278] = 32'b11111111111111111000010010011001;
assign LUT_2[7279] = 32'b11111111111111110101001010110010;
assign LUT_2[7280] = 32'b11111111111111110100101110100010;
assign LUT_2[7281] = 32'b11111111111111110001100110111011;
assign LUT_2[7282] = 32'b11111111111111111011100111011110;
assign LUT_2[7283] = 32'b11111111111111111000011111110111;
assign LUT_2[7284] = 32'b11111111111111110001001100001010;
assign LUT_2[7285] = 32'b11111111111111101110000100100011;
assign LUT_2[7286] = 32'b11111111111111111000000101000110;
assign LUT_2[7287] = 32'b11111111111111110100111101011111;
assign LUT_2[7288] = 32'b11111111111111101111011111111111;
assign LUT_2[7289] = 32'b11111111111111101100011000011000;
assign LUT_2[7290] = 32'b11111111111111110110011000111011;
assign LUT_2[7291] = 32'b11111111111111110011010001010100;
assign LUT_2[7292] = 32'b11111111111111101011111101100111;
assign LUT_2[7293] = 32'b11111111111111101000110110000000;
assign LUT_2[7294] = 32'b11111111111111110010110110100011;
assign LUT_2[7295] = 32'b11111111111111101111101110111100;
assign LUT_2[7296] = 32'b00000000000000000101111010011011;
assign LUT_2[7297] = 32'b00000000000000000010110010110100;
assign LUT_2[7298] = 32'b00000000000000001100110011010111;
assign LUT_2[7299] = 32'b00000000000000001001101011110000;
assign LUT_2[7300] = 32'b00000000000000000010011000000011;
assign LUT_2[7301] = 32'b11111111111111111111010000011100;
assign LUT_2[7302] = 32'b00000000000000001001010000111111;
assign LUT_2[7303] = 32'b00000000000000000110001001011000;
assign LUT_2[7304] = 32'b00000000000000000000101011111000;
assign LUT_2[7305] = 32'b11111111111111111101100100010001;
assign LUT_2[7306] = 32'b00000000000000000111100100110100;
assign LUT_2[7307] = 32'b00000000000000000100011101001101;
assign LUT_2[7308] = 32'b11111111111111111101001001100000;
assign LUT_2[7309] = 32'b11111111111111111010000001111001;
assign LUT_2[7310] = 32'b00000000000000000100000010011100;
assign LUT_2[7311] = 32'b00000000000000000000111010110101;
assign LUT_2[7312] = 32'b00000000000000000000011110100101;
assign LUT_2[7313] = 32'b11111111111111111101010110111110;
assign LUT_2[7314] = 32'b00000000000000000111010111100001;
assign LUT_2[7315] = 32'b00000000000000000100001111111010;
assign LUT_2[7316] = 32'b11111111111111111100111100001101;
assign LUT_2[7317] = 32'b11111111111111111001110100100110;
assign LUT_2[7318] = 32'b00000000000000000011110101001001;
assign LUT_2[7319] = 32'b00000000000000000000101101100010;
assign LUT_2[7320] = 32'b11111111111111111011010000000010;
assign LUT_2[7321] = 32'b11111111111111111000001000011011;
assign LUT_2[7322] = 32'b00000000000000000010001000111110;
assign LUT_2[7323] = 32'b11111111111111111111000001010111;
assign LUT_2[7324] = 32'b11111111111111110111101101101010;
assign LUT_2[7325] = 32'b11111111111111110100100110000011;
assign LUT_2[7326] = 32'b11111111111111111110100110100110;
assign LUT_2[7327] = 32'b11111111111111111011011110111111;
assign LUT_2[7328] = 32'b00000000000000000110010110000100;
assign LUT_2[7329] = 32'b00000000000000000011001110011101;
assign LUT_2[7330] = 32'b00000000000000001101001111000000;
assign LUT_2[7331] = 32'b00000000000000001010000111011001;
assign LUT_2[7332] = 32'b00000000000000000010110011101100;
assign LUT_2[7333] = 32'b11111111111111111111101100000101;
assign LUT_2[7334] = 32'b00000000000000001001101100101000;
assign LUT_2[7335] = 32'b00000000000000000110100101000001;
assign LUT_2[7336] = 32'b00000000000000000001000111100001;
assign LUT_2[7337] = 32'b11111111111111111101111111111010;
assign LUT_2[7338] = 32'b00000000000000001000000000011101;
assign LUT_2[7339] = 32'b00000000000000000100111000110110;
assign LUT_2[7340] = 32'b11111111111111111101100101001001;
assign LUT_2[7341] = 32'b11111111111111111010011101100010;
assign LUT_2[7342] = 32'b00000000000000000100011110000101;
assign LUT_2[7343] = 32'b00000000000000000001010110011110;
assign LUT_2[7344] = 32'b00000000000000000000111010001110;
assign LUT_2[7345] = 32'b11111111111111111101110010100111;
assign LUT_2[7346] = 32'b00000000000000000111110011001010;
assign LUT_2[7347] = 32'b00000000000000000100101011100011;
assign LUT_2[7348] = 32'b11111111111111111101010111110110;
assign LUT_2[7349] = 32'b11111111111111111010010000001111;
assign LUT_2[7350] = 32'b00000000000000000100010000110010;
assign LUT_2[7351] = 32'b00000000000000000001001001001011;
assign LUT_2[7352] = 32'b11111111111111111011101011101011;
assign LUT_2[7353] = 32'b11111111111111111000100100000100;
assign LUT_2[7354] = 32'b00000000000000000010100100100111;
assign LUT_2[7355] = 32'b11111111111111111111011101000000;
assign LUT_2[7356] = 32'b11111111111111111000001001010011;
assign LUT_2[7357] = 32'b11111111111111110101000001101100;
assign LUT_2[7358] = 32'b11111111111111111111000010001111;
assign LUT_2[7359] = 32'b11111111111111111011111010101000;
assign LUT_2[7360] = 32'b11111111111111111110000010111110;
assign LUT_2[7361] = 32'b11111111111111111010111011010111;
assign LUT_2[7362] = 32'b00000000000000000100111011111010;
assign LUT_2[7363] = 32'b00000000000000000001110100010011;
assign LUT_2[7364] = 32'b11111111111111111010100000100110;
assign LUT_2[7365] = 32'b11111111111111110111011000111111;
assign LUT_2[7366] = 32'b00000000000000000001011001100010;
assign LUT_2[7367] = 32'b11111111111111111110010001111011;
assign LUT_2[7368] = 32'b11111111111111111000110100011011;
assign LUT_2[7369] = 32'b11111111111111110101101100110100;
assign LUT_2[7370] = 32'b11111111111111111111101101010111;
assign LUT_2[7371] = 32'b11111111111111111100100101110000;
assign LUT_2[7372] = 32'b11111111111111110101010010000011;
assign LUT_2[7373] = 32'b11111111111111110010001010011100;
assign LUT_2[7374] = 32'b11111111111111111100001010111111;
assign LUT_2[7375] = 32'b11111111111111111001000011011000;
assign LUT_2[7376] = 32'b11111111111111111000100111001000;
assign LUT_2[7377] = 32'b11111111111111110101011111100001;
assign LUT_2[7378] = 32'b11111111111111111111100000000100;
assign LUT_2[7379] = 32'b11111111111111111100011000011101;
assign LUT_2[7380] = 32'b11111111111111110101000100110000;
assign LUT_2[7381] = 32'b11111111111111110001111101001001;
assign LUT_2[7382] = 32'b11111111111111111011111101101100;
assign LUT_2[7383] = 32'b11111111111111111000110110000101;
assign LUT_2[7384] = 32'b11111111111111110011011000100101;
assign LUT_2[7385] = 32'b11111111111111110000010000111110;
assign LUT_2[7386] = 32'b11111111111111111010010001100001;
assign LUT_2[7387] = 32'b11111111111111110111001001111010;
assign LUT_2[7388] = 32'b11111111111111101111110110001101;
assign LUT_2[7389] = 32'b11111111111111101100101110100110;
assign LUT_2[7390] = 32'b11111111111111110110101111001001;
assign LUT_2[7391] = 32'b11111111111111110011100111100010;
assign LUT_2[7392] = 32'b11111111111111111110011110100111;
assign LUT_2[7393] = 32'b11111111111111111011010111000000;
assign LUT_2[7394] = 32'b00000000000000000101010111100011;
assign LUT_2[7395] = 32'b00000000000000000010001111111100;
assign LUT_2[7396] = 32'b11111111111111111010111100001111;
assign LUT_2[7397] = 32'b11111111111111110111110100101000;
assign LUT_2[7398] = 32'b00000000000000000001110101001011;
assign LUT_2[7399] = 32'b11111111111111111110101101100100;
assign LUT_2[7400] = 32'b11111111111111111001010000000100;
assign LUT_2[7401] = 32'b11111111111111110110001000011101;
assign LUT_2[7402] = 32'b00000000000000000000001001000000;
assign LUT_2[7403] = 32'b11111111111111111101000001011001;
assign LUT_2[7404] = 32'b11111111111111110101101101101100;
assign LUT_2[7405] = 32'b11111111111111110010100110000101;
assign LUT_2[7406] = 32'b11111111111111111100100110101000;
assign LUT_2[7407] = 32'b11111111111111111001011111000001;
assign LUT_2[7408] = 32'b11111111111111111001000010110001;
assign LUT_2[7409] = 32'b11111111111111110101111011001010;
assign LUT_2[7410] = 32'b11111111111111111111111011101101;
assign LUT_2[7411] = 32'b11111111111111111100110100000110;
assign LUT_2[7412] = 32'b11111111111111110101100000011001;
assign LUT_2[7413] = 32'b11111111111111110010011000110010;
assign LUT_2[7414] = 32'b11111111111111111100011001010101;
assign LUT_2[7415] = 32'b11111111111111111001010001101110;
assign LUT_2[7416] = 32'b11111111111111110011110100001110;
assign LUT_2[7417] = 32'b11111111111111110000101100100111;
assign LUT_2[7418] = 32'b11111111111111111010101101001010;
assign LUT_2[7419] = 32'b11111111111111110111100101100011;
assign LUT_2[7420] = 32'b11111111111111110000010001110110;
assign LUT_2[7421] = 32'b11111111111111101101001010001111;
assign LUT_2[7422] = 32'b11111111111111110111001010110010;
assign LUT_2[7423] = 32'b11111111111111110100000011001011;
assign LUT_2[7424] = 32'b00000000000000000101100100110010;
assign LUT_2[7425] = 32'b00000000000000000010011101001011;
assign LUT_2[7426] = 32'b00000000000000001100011101101110;
assign LUT_2[7427] = 32'b00000000000000001001010110000111;
assign LUT_2[7428] = 32'b00000000000000000010000010011010;
assign LUT_2[7429] = 32'b11111111111111111110111010110011;
assign LUT_2[7430] = 32'b00000000000000001000111011010110;
assign LUT_2[7431] = 32'b00000000000000000101110011101111;
assign LUT_2[7432] = 32'b00000000000000000000010110001111;
assign LUT_2[7433] = 32'b11111111111111111101001110101000;
assign LUT_2[7434] = 32'b00000000000000000111001111001011;
assign LUT_2[7435] = 32'b00000000000000000100000111100100;
assign LUT_2[7436] = 32'b11111111111111111100110011110111;
assign LUT_2[7437] = 32'b11111111111111111001101100010000;
assign LUT_2[7438] = 32'b00000000000000000011101100110011;
assign LUT_2[7439] = 32'b00000000000000000000100101001100;
assign LUT_2[7440] = 32'b00000000000000000000001000111100;
assign LUT_2[7441] = 32'b11111111111111111101000001010101;
assign LUT_2[7442] = 32'b00000000000000000111000001111000;
assign LUT_2[7443] = 32'b00000000000000000011111010010001;
assign LUT_2[7444] = 32'b11111111111111111100100110100100;
assign LUT_2[7445] = 32'b11111111111111111001011110111101;
assign LUT_2[7446] = 32'b00000000000000000011011111100000;
assign LUT_2[7447] = 32'b00000000000000000000010111111001;
assign LUT_2[7448] = 32'b11111111111111111010111010011001;
assign LUT_2[7449] = 32'b11111111111111110111110010110010;
assign LUT_2[7450] = 32'b00000000000000000001110011010101;
assign LUT_2[7451] = 32'b11111111111111111110101011101110;
assign LUT_2[7452] = 32'b11111111111111110111011000000001;
assign LUT_2[7453] = 32'b11111111111111110100010000011010;
assign LUT_2[7454] = 32'b11111111111111111110010000111101;
assign LUT_2[7455] = 32'b11111111111111111011001001010110;
assign LUT_2[7456] = 32'b00000000000000000110000000011011;
assign LUT_2[7457] = 32'b00000000000000000010111000110100;
assign LUT_2[7458] = 32'b00000000000000001100111001010111;
assign LUT_2[7459] = 32'b00000000000000001001110001110000;
assign LUT_2[7460] = 32'b00000000000000000010011110000011;
assign LUT_2[7461] = 32'b11111111111111111111010110011100;
assign LUT_2[7462] = 32'b00000000000000001001010110111111;
assign LUT_2[7463] = 32'b00000000000000000110001111011000;
assign LUT_2[7464] = 32'b00000000000000000000110001111000;
assign LUT_2[7465] = 32'b11111111111111111101101010010001;
assign LUT_2[7466] = 32'b00000000000000000111101010110100;
assign LUT_2[7467] = 32'b00000000000000000100100011001101;
assign LUT_2[7468] = 32'b11111111111111111101001111100000;
assign LUT_2[7469] = 32'b11111111111111111010000111111001;
assign LUT_2[7470] = 32'b00000000000000000100001000011100;
assign LUT_2[7471] = 32'b00000000000000000001000000110101;
assign LUT_2[7472] = 32'b00000000000000000000100100100101;
assign LUT_2[7473] = 32'b11111111111111111101011100111110;
assign LUT_2[7474] = 32'b00000000000000000111011101100001;
assign LUT_2[7475] = 32'b00000000000000000100010101111010;
assign LUT_2[7476] = 32'b11111111111111111101000010001101;
assign LUT_2[7477] = 32'b11111111111111111001111010100110;
assign LUT_2[7478] = 32'b00000000000000000011111011001001;
assign LUT_2[7479] = 32'b00000000000000000000110011100010;
assign LUT_2[7480] = 32'b11111111111111111011010110000010;
assign LUT_2[7481] = 32'b11111111111111111000001110011011;
assign LUT_2[7482] = 32'b00000000000000000010001110111110;
assign LUT_2[7483] = 32'b11111111111111111111000111010111;
assign LUT_2[7484] = 32'b11111111111111110111110011101010;
assign LUT_2[7485] = 32'b11111111111111110100101100000011;
assign LUT_2[7486] = 32'b11111111111111111110101100100110;
assign LUT_2[7487] = 32'b11111111111111111011100100111111;
assign LUT_2[7488] = 32'b11111111111111111101101101010101;
assign LUT_2[7489] = 32'b11111111111111111010100101101110;
assign LUT_2[7490] = 32'b00000000000000000100100110010001;
assign LUT_2[7491] = 32'b00000000000000000001011110101010;
assign LUT_2[7492] = 32'b11111111111111111010001010111101;
assign LUT_2[7493] = 32'b11111111111111110111000011010110;
assign LUT_2[7494] = 32'b00000000000000000001000011111001;
assign LUT_2[7495] = 32'b11111111111111111101111100010010;
assign LUT_2[7496] = 32'b11111111111111111000011110110010;
assign LUT_2[7497] = 32'b11111111111111110101010111001011;
assign LUT_2[7498] = 32'b11111111111111111111010111101110;
assign LUT_2[7499] = 32'b11111111111111111100010000000111;
assign LUT_2[7500] = 32'b11111111111111110100111100011010;
assign LUT_2[7501] = 32'b11111111111111110001110100110011;
assign LUT_2[7502] = 32'b11111111111111111011110101010110;
assign LUT_2[7503] = 32'b11111111111111111000101101101111;
assign LUT_2[7504] = 32'b11111111111111111000010001011111;
assign LUT_2[7505] = 32'b11111111111111110101001001111000;
assign LUT_2[7506] = 32'b11111111111111111111001010011011;
assign LUT_2[7507] = 32'b11111111111111111100000010110100;
assign LUT_2[7508] = 32'b11111111111111110100101111000111;
assign LUT_2[7509] = 32'b11111111111111110001100111100000;
assign LUT_2[7510] = 32'b11111111111111111011101000000011;
assign LUT_2[7511] = 32'b11111111111111111000100000011100;
assign LUT_2[7512] = 32'b11111111111111110011000010111100;
assign LUT_2[7513] = 32'b11111111111111101111111011010101;
assign LUT_2[7514] = 32'b11111111111111111001111011111000;
assign LUT_2[7515] = 32'b11111111111111110110110100010001;
assign LUT_2[7516] = 32'b11111111111111101111100000100100;
assign LUT_2[7517] = 32'b11111111111111101100011000111101;
assign LUT_2[7518] = 32'b11111111111111110110011001100000;
assign LUT_2[7519] = 32'b11111111111111110011010001111001;
assign LUT_2[7520] = 32'b11111111111111111110001000111110;
assign LUT_2[7521] = 32'b11111111111111111011000001010111;
assign LUT_2[7522] = 32'b00000000000000000101000001111010;
assign LUT_2[7523] = 32'b00000000000000000001111010010011;
assign LUT_2[7524] = 32'b11111111111111111010100110100110;
assign LUT_2[7525] = 32'b11111111111111110111011110111111;
assign LUT_2[7526] = 32'b00000000000000000001011111100010;
assign LUT_2[7527] = 32'b11111111111111111110010111111011;
assign LUT_2[7528] = 32'b11111111111111111000111010011011;
assign LUT_2[7529] = 32'b11111111111111110101110010110100;
assign LUT_2[7530] = 32'b11111111111111111111110011010111;
assign LUT_2[7531] = 32'b11111111111111111100101011110000;
assign LUT_2[7532] = 32'b11111111111111110101011000000011;
assign LUT_2[7533] = 32'b11111111111111110010010000011100;
assign LUT_2[7534] = 32'b11111111111111111100010000111111;
assign LUT_2[7535] = 32'b11111111111111111001001001011000;
assign LUT_2[7536] = 32'b11111111111111111000101101001000;
assign LUT_2[7537] = 32'b11111111111111110101100101100001;
assign LUT_2[7538] = 32'b11111111111111111111100110000100;
assign LUT_2[7539] = 32'b11111111111111111100011110011101;
assign LUT_2[7540] = 32'b11111111111111110101001010110000;
assign LUT_2[7541] = 32'b11111111111111110010000011001001;
assign LUT_2[7542] = 32'b11111111111111111100000011101100;
assign LUT_2[7543] = 32'b11111111111111111000111100000101;
assign LUT_2[7544] = 32'b11111111111111110011011110100101;
assign LUT_2[7545] = 32'b11111111111111110000010110111110;
assign LUT_2[7546] = 32'b11111111111111111010010111100001;
assign LUT_2[7547] = 32'b11111111111111110111001111111010;
assign LUT_2[7548] = 32'b11111111111111101111111100001101;
assign LUT_2[7549] = 32'b11111111111111101100110100100110;
assign LUT_2[7550] = 32'b11111111111111110110110101001001;
assign LUT_2[7551] = 32'b11111111111111110011101101100010;
assign LUT_2[7552] = 32'b00000000000000001001111001000001;
assign LUT_2[7553] = 32'b00000000000000000110110001011010;
assign LUT_2[7554] = 32'b00000000000000010000110001111101;
assign LUT_2[7555] = 32'b00000000000000001101101010010110;
assign LUT_2[7556] = 32'b00000000000000000110010110101001;
assign LUT_2[7557] = 32'b00000000000000000011001111000010;
assign LUT_2[7558] = 32'b00000000000000001101001111100101;
assign LUT_2[7559] = 32'b00000000000000001010000111111110;
assign LUT_2[7560] = 32'b00000000000000000100101010011110;
assign LUT_2[7561] = 32'b00000000000000000001100010110111;
assign LUT_2[7562] = 32'b00000000000000001011100011011010;
assign LUT_2[7563] = 32'b00000000000000001000011011110011;
assign LUT_2[7564] = 32'b00000000000000000001001000000110;
assign LUT_2[7565] = 32'b11111111111111111110000000011111;
assign LUT_2[7566] = 32'b00000000000000001000000001000010;
assign LUT_2[7567] = 32'b00000000000000000100111001011011;
assign LUT_2[7568] = 32'b00000000000000000100011101001011;
assign LUT_2[7569] = 32'b00000000000000000001010101100100;
assign LUT_2[7570] = 32'b00000000000000001011010110000111;
assign LUT_2[7571] = 32'b00000000000000001000001110100000;
assign LUT_2[7572] = 32'b00000000000000000000111010110011;
assign LUT_2[7573] = 32'b11111111111111111101110011001100;
assign LUT_2[7574] = 32'b00000000000000000111110011101111;
assign LUT_2[7575] = 32'b00000000000000000100101100001000;
assign LUT_2[7576] = 32'b11111111111111111111001110101000;
assign LUT_2[7577] = 32'b11111111111111111100000111000001;
assign LUT_2[7578] = 32'b00000000000000000110000111100100;
assign LUT_2[7579] = 32'b00000000000000000010111111111101;
assign LUT_2[7580] = 32'b11111111111111111011101100010000;
assign LUT_2[7581] = 32'b11111111111111111000100100101001;
assign LUT_2[7582] = 32'b00000000000000000010100101001100;
assign LUT_2[7583] = 32'b11111111111111111111011101100101;
assign LUT_2[7584] = 32'b00000000000000001010010100101010;
assign LUT_2[7585] = 32'b00000000000000000111001101000011;
assign LUT_2[7586] = 32'b00000000000000010001001101100110;
assign LUT_2[7587] = 32'b00000000000000001110000101111111;
assign LUT_2[7588] = 32'b00000000000000000110110010010010;
assign LUT_2[7589] = 32'b00000000000000000011101010101011;
assign LUT_2[7590] = 32'b00000000000000001101101011001110;
assign LUT_2[7591] = 32'b00000000000000001010100011100111;
assign LUT_2[7592] = 32'b00000000000000000101000110000111;
assign LUT_2[7593] = 32'b00000000000000000001111110100000;
assign LUT_2[7594] = 32'b00000000000000001011111111000011;
assign LUT_2[7595] = 32'b00000000000000001000110111011100;
assign LUT_2[7596] = 32'b00000000000000000001100011101111;
assign LUT_2[7597] = 32'b11111111111111111110011100001000;
assign LUT_2[7598] = 32'b00000000000000001000011100101011;
assign LUT_2[7599] = 32'b00000000000000000101010101000100;
assign LUT_2[7600] = 32'b00000000000000000100111000110100;
assign LUT_2[7601] = 32'b00000000000000000001110001001101;
assign LUT_2[7602] = 32'b00000000000000001011110001110000;
assign LUT_2[7603] = 32'b00000000000000001000101010001001;
assign LUT_2[7604] = 32'b00000000000000000001010110011100;
assign LUT_2[7605] = 32'b11111111111111111110001110110101;
assign LUT_2[7606] = 32'b00000000000000001000001111011000;
assign LUT_2[7607] = 32'b00000000000000000101000111110001;
assign LUT_2[7608] = 32'b11111111111111111111101010010001;
assign LUT_2[7609] = 32'b11111111111111111100100010101010;
assign LUT_2[7610] = 32'b00000000000000000110100011001101;
assign LUT_2[7611] = 32'b00000000000000000011011011100110;
assign LUT_2[7612] = 32'b11111111111111111100000111111001;
assign LUT_2[7613] = 32'b11111111111111111001000000010010;
assign LUT_2[7614] = 32'b00000000000000000011000000110101;
assign LUT_2[7615] = 32'b11111111111111111111111001001110;
assign LUT_2[7616] = 32'b00000000000000000010000001100100;
assign LUT_2[7617] = 32'b11111111111111111110111001111101;
assign LUT_2[7618] = 32'b00000000000000001000111010100000;
assign LUT_2[7619] = 32'b00000000000000000101110010111001;
assign LUT_2[7620] = 32'b11111111111111111110011111001100;
assign LUT_2[7621] = 32'b11111111111111111011010111100101;
assign LUT_2[7622] = 32'b00000000000000000101011000001000;
assign LUT_2[7623] = 32'b00000000000000000010010000100001;
assign LUT_2[7624] = 32'b11111111111111111100110011000001;
assign LUT_2[7625] = 32'b11111111111111111001101011011010;
assign LUT_2[7626] = 32'b00000000000000000011101011111101;
assign LUT_2[7627] = 32'b00000000000000000000100100010110;
assign LUT_2[7628] = 32'b11111111111111111001010000101001;
assign LUT_2[7629] = 32'b11111111111111110110001001000010;
assign LUT_2[7630] = 32'b00000000000000000000001001100101;
assign LUT_2[7631] = 32'b11111111111111111101000001111110;
assign LUT_2[7632] = 32'b11111111111111111100100101101110;
assign LUT_2[7633] = 32'b11111111111111111001011110000111;
assign LUT_2[7634] = 32'b00000000000000000011011110101010;
assign LUT_2[7635] = 32'b00000000000000000000010111000011;
assign LUT_2[7636] = 32'b11111111111111111001000011010110;
assign LUT_2[7637] = 32'b11111111111111110101111011101111;
assign LUT_2[7638] = 32'b11111111111111111111111100010010;
assign LUT_2[7639] = 32'b11111111111111111100110100101011;
assign LUT_2[7640] = 32'b11111111111111110111010111001011;
assign LUT_2[7641] = 32'b11111111111111110100001111100100;
assign LUT_2[7642] = 32'b11111111111111111110010000000111;
assign LUT_2[7643] = 32'b11111111111111111011001000100000;
assign LUT_2[7644] = 32'b11111111111111110011110100110011;
assign LUT_2[7645] = 32'b11111111111111110000101101001100;
assign LUT_2[7646] = 32'b11111111111111111010101101101111;
assign LUT_2[7647] = 32'b11111111111111110111100110001000;
assign LUT_2[7648] = 32'b00000000000000000010011101001101;
assign LUT_2[7649] = 32'b11111111111111111111010101100110;
assign LUT_2[7650] = 32'b00000000000000001001010110001001;
assign LUT_2[7651] = 32'b00000000000000000110001110100010;
assign LUT_2[7652] = 32'b11111111111111111110111010110101;
assign LUT_2[7653] = 32'b11111111111111111011110011001110;
assign LUT_2[7654] = 32'b00000000000000000101110011110001;
assign LUT_2[7655] = 32'b00000000000000000010101100001010;
assign LUT_2[7656] = 32'b11111111111111111101001110101010;
assign LUT_2[7657] = 32'b11111111111111111010000111000011;
assign LUT_2[7658] = 32'b00000000000000000100000111100110;
assign LUT_2[7659] = 32'b00000000000000000000111111111111;
assign LUT_2[7660] = 32'b11111111111111111001101100010010;
assign LUT_2[7661] = 32'b11111111111111110110100100101011;
assign LUT_2[7662] = 32'b00000000000000000000100101001110;
assign LUT_2[7663] = 32'b11111111111111111101011101100111;
assign LUT_2[7664] = 32'b11111111111111111101000001010111;
assign LUT_2[7665] = 32'b11111111111111111001111001110000;
assign LUT_2[7666] = 32'b00000000000000000011111010010011;
assign LUT_2[7667] = 32'b00000000000000000000110010101100;
assign LUT_2[7668] = 32'b11111111111111111001011110111111;
assign LUT_2[7669] = 32'b11111111111111110110010111011000;
assign LUT_2[7670] = 32'b00000000000000000000010111111011;
assign LUT_2[7671] = 32'b11111111111111111101010000010100;
assign LUT_2[7672] = 32'b11111111111111110111110010110100;
assign LUT_2[7673] = 32'b11111111111111110100101011001101;
assign LUT_2[7674] = 32'b11111111111111111110101011110000;
assign LUT_2[7675] = 32'b11111111111111111011100100001001;
assign LUT_2[7676] = 32'b11111111111111110100010000011100;
assign LUT_2[7677] = 32'b11111111111111110001001000110101;
assign LUT_2[7678] = 32'b11111111111111111011001001011000;
assign LUT_2[7679] = 32'b11111111111111111000000001110001;
assign LUT_2[7680] = 32'b00000000000000000110010111111110;
assign LUT_2[7681] = 32'b00000000000000000011010000010111;
assign LUT_2[7682] = 32'b00000000000000001101010000111010;
assign LUT_2[7683] = 32'b00000000000000001010001001010011;
assign LUT_2[7684] = 32'b00000000000000000010110101100110;
assign LUT_2[7685] = 32'b11111111111111111111101101111111;
assign LUT_2[7686] = 32'b00000000000000001001101110100010;
assign LUT_2[7687] = 32'b00000000000000000110100110111011;
assign LUT_2[7688] = 32'b00000000000000000001001001011011;
assign LUT_2[7689] = 32'b11111111111111111110000001110100;
assign LUT_2[7690] = 32'b00000000000000001000000010010111;
assign LUT_2[7691] = 32'b00000000000000000100111010110000;
assign LUT_2[7692] = 32'b11111111111111111101100111000011;
assign LUT_2[7693] = 32'b11111111111111111010011111011100;
assign LUT_2[7694] = 32'b00000000000000000100011111111111;
assign LUT_2[7695] = 32'b00000000000000000001011000011000;
assign LUT_2[7696] = 32'b00000000000000000000111100001000;
assign LUT_2[7697] = 32'b11111111111111111101110100100001;
assign LUT_2[7698] = 32'b00000000000000000111110101000100;
assign LUT_2[7699] = 32'b00000000000000000100101101011101;
assign LUT_2[7700] = 32'b11111111111111111101011001110000;
assign LUT_2[7701] = 32'b11111111111111111010010010001001;
assign LUT_2[7702] = 32'b00000000000000000100010010101100;
assign LUT_2[7703] = 32'b00000000000000000001001011000101;
assign LUT_2[7704] = 32'b11111111111111111011101101100101;
assign LUT_2[7705] = 32'b11111111111111111000100101111110;
assign LUT_2[7706] = 32'b00000000000000000010100110100001;
assign LUT_2[7707] = 32'b11111111111111111111011110111010;
assign LUT_2[7708] = 32'b11111111111111111000001011001101;
assign LUT_2[7709] = 32'b11111111111111110101000011100110;
assign LUT_2[7710] = 32'b11111111111111111111000100001001;
assign LUT_2[7711] = 32'b11111111111111111011111100100010;
assign LUT_2[7712] = 32'b00000000000000000110110011100111;
assign LUT_2[7713] = 32'b00000000000000000011101100000000;
assign LUT_2[7714] = 32'b00000000000000001101101100100011;
assign LUT_2[7715] = 32'b00000000000000001010100100111100;
assign LUT_2[7716] = 32'b00000000000000000011010001001111;
assign LUT_2[7717] = 32'b00000000000000000000001001101000;
assign LUT_2[7718] = 32'b00000000000000001010001010001011;
assign LUT_2[7719] = 32'b00000000000000000111000010100100;
assign LUT_2[7720] = 32'b00000000000000000001100101000100;
assign LUT_2[7721] = 32'b11111111111111111110011101011101;
assign LUT_2[7722] = 32'b00000000000000001000011110000000;
assign LUT_2[7723] = 32'b00000000000000000101010110011001;
assign LUT_2[7724] = 32'b11111111111111111110000010101100;
assign LUT_2[7725] = 32'b11111111111111111010111011000101;
assign LUT_2[7726] = 32'b00000000000000000100111011101000;
assign LUT_2[7727] = 32'b00000000000000000001110100000001;
assign LUT_2[7728] = 32'b00000000000000000001010111110001;
assign LUT_2[7729] = 32'b11111111111111111110010000001010;
assign LUT_2[7730] = 32'b00000000000000001000010000101101;
assign LUT_2[7731] = 32'b00000000000000000101001001000110;
assign LUT_2[7732] = 32'b11111111111111111101110101011001;
assign LUT_2[7733] = 32'b11111111111111111010101101110010;
assign LUT_2[7734] = 32'b00000000000000000100101110010101;
assign LUT_2[7735] = 32'b00000000000000000001100110101110;
assign LUT_2[7736] = 32'b11111111111111111100001001001110;
assign LUT_2[7737] = 32'b11111111111111111001000001100111;
assign LUT_2[7738] = 32'b00000000000000000011000010001010;
assign LUT_2[7739] = 32'b11111111111111111111111010100011;
assign LUT_2[7740] = 32'b11111111111111111000100110110110;
assign LUT_2[7741] = 32'b11111111111111110101011111001111;
assign LUT_2[7742] = 32'b11111111111111111111011111110010;
assign LUT_2[7743] = 32'b11111111111111111100011000001011;
assign LUT_2[7744] = 32'b11111111111111111110100000100001;
assign LUT_2[7745] = 32'b11111111111111111011011000111010;
assign LUT_2[7746] = 32'b00000000000000000101011001011101;
assign LUT_2[7747] = 32'b00000000000000000010010001110110;
assign LUT_2[7748] = 32'b11111111111111111010111110001001;
assign LUT_2[7749] = 32'b11111111111111110111110110100010;
assign LUT_2[7750] = 32'b00000000000000000001110111000101;
assign LUT_2[7751] = 32'b11111111111111111110101111011110;
assign LUT_2[7752] = 32'b11111111111111111001010001111110;
assign LUT_2[7753] = 32'b11111111111111110110001010010111;
assign LUT_2[7754] = 32'b00000000000000000000001010111010;
assign LUT_2[7755] = 32'b11111111111111111101000011010011;
assign LUT_2[7756] = 32'b11111111111111110101101111100110;
assign LUT_2[7757] = 32'b11111111111111110010100111111111;
assign LUT_2[7758] = 32'b11111111111111111100101000100010;
assign LUT_2[7759] = 32'b11111111111111111001100000111011;
assign LUT_2[7760] = 32'b11111111111111111001000100101011;
assign LUT_2[7761] = 32'b11111111111111110101111101000100;
assign LUT_2[7762] = 32'b11111111111111111111111101100111;
assign LUT_2[7763] = 32'b11111111111111111100110110000000;
assign LUT_2[7764] = 32'b11111111111111110101100010010011;
assign LUT_2[7765] = 32'b11111111111111110010011010101100;
assign LUT_2[7766] = 32'b11111111111111111100011011001111;
assign LUT_2[7767] = 32'b11111111111111111001010011101000;
assign LUT_2[7768] = 32'b11111111111111110011110110001000;
assign LUT_2[7769] = 32'b11111111111111110000101110100001;
assign LUT_2[7770] = 32'b11111111111111111010101111000100;
assign LUT_2[7771] = 32'b11111111111111110111100111011101;
assign LUT_2[7772] = 32'b11111111111111110000010011110000;
assign LUT_2[7773] = 32'b11111111111111101101001100001001;
assign LUT_2[7774] = 32'b11111111111111110111001100101100;
assign LUT_2[7775] = 32'b11111111111111110100000101000101;
assign LUT_2[7776] = 32'b11111111111111111110111100001010;
assign LUT_2[7777] = 32'b11111111111111111011110100100011;
assign LUT_2[7778] = 32'b00000000000000000101110101000110;
assign LUT_2[7779] = 32'b00000000000000000010101101011111;
assign LUT_2[7780] = 32'b11111111111111111011011001110010;
assign LUT_2[7781] = 32'b11111111111111111000010010001011;
assign LUT_2[7782] = 32'b00000000000000000010010010101110;
assign LUT_2[7783] = 32'b11111111111111111111001011000111;
assign LUT_2[7784] = 32'b11111111111111111001101101100111;
assign LUT_2[7785] = 32'b11111111111111110110100110000000;
assign LUT_2[7786] = 32'b00000000000000000000100110100011;
assign LUT_2[7787] = 32'b11111111111111111101011110111100;
assign LUT_2[7788] = 32'b11111111111111110110001011001111;
assign LUT_2[7789] = 32'b11111111111111110011000011101000;
assign LUT_2[7790] = 32'b11111111111111111101000100001011;
assign LUT_2[7791] = 32'b11111111111111111001111100100100;
assign LUT_2[7792] = 32'b11111111111111111001100000010100;
assign LUT_2[7793] = 32'b11111111111111110110011000101101;
assign LUT_2[7794] = 32'b00000000000000000000011001010000;
assign LUT_2[7795] = 32'b11111111111111111101010001101001;
assign LUT_2[7796] = 32'b11111111111111110101111101111100;
assign LUT_2[7797] = 32'b11111111111111110010110110010101;
assign LUT_2[7798] = 32'b11111111111111111100110110111000;
assign LUT_2[7799] = 32'b11111111111111111001101111010001;
assign LUT_2[7800] = 32'b11111111111111110100010001110001;
assign LUT_2[7801] = 32'b11111111111111110001001010001010;
assign LUT_2[7802] = 32'b11111111111111111011001010101101;
assign LUT_2[7803] = 32'b11111111111111111000000011000110;
assign LUT_2[7804] = 32'b11111111111111110000101111011001;
assign LUT_2[7805] = 32'b11111111111111101101100111110010;
assign LUT_2[7806] = 32'b11111111111111110111101000010101;
assign LUT_2[7807] = 32'b11111111111111110100100000101110;
assign LUT_2[7808] = 32'b00000000000000001010101100001101;
assign LUT_2[7809] = 32'b00000000000000000111100100100110;
assign LUT_2[7810] = 32'b00000000000000010001100101001001;
assign LUT_2[7811] = 32'b00000000000000001110011101100010;
assign LUT_2[7812] = 32'b00000000000000000111001001110101;
assign LUT_2[7813] = 32'b00000000000000000100000010001110;
assign LUT_2[7814] = 32'b00000000000000001110000010110001;
assign LUT_2[7815] = 32'b00000000000000001010111011001010;
assign LUT_2[7816] = 32'b00000000000000000101011101101010;
assign LUT_2[7817] = 32'b00000000000000000010010110000011;
assign LUT_2[7818] = 32'b00000000000000001100010110100110;
assign LUT_2[7819] = 32'b00000000000000001001001110111111;
assign LUT_2[7820] = 32'b00000000000000000001111011010010;
assign LUT_2[7821] = 32'b11111111111111111110110011101011;
assign LUT_2[7822] = 32'b00000000000000001000110100001110;
assign LUT_2[7823] = 32'b00000000000000000101101100100111;
assign LUT_2[7824] = 32'b00000000000000000101010000010111;
assign LUT_2[7825] = 32'b00000000000000000010001000110000;
assign LUT_2[7826] = 32'b00000000000000001100001001010011;
assign LUT_2[7827] = 32'b00000000000000001001000001101100;
assign LUT_2[7828] = 32'b00000000000000000001101101111111;
assign LUT_2[7829] = 32'b11111111111111111110100110011000;
assign LUT_2[7830] = 32'b00000000000000001000100110111011;
assign LUT_2[7831] = 32'b00000000000000000101011111010100;
assign LUT_2[7832] = 32'b00000000000000000000000001110100;
assign LUT_2[7833] = 32'b11111111111111111100111010001101;
assign LUT_2[7834] = 32'b00000000000000000110111010110000;
assign LUT_2[7835] = 32'b00000000000000000011110011001001;
assign LUT_2[7836] = 32'b11111111111111111100011111011100;
assign LUT_2[7837] = 32'b11111111111111111001010111110101;
assign LUT_2[7838] = 32'b00000000000000000011011000011000;
assign LUT_2[7839] = 32'b00000000000000000000010000110001;
assign LUT_2[7840] = 32'b00000000000000001011000111110110;
assign LUT_2[7841] = 32'b00000000000000001000000000001111;
assign LUT_2[7842] = 32'b00000000000000010010000000110010;
assign LUT_2[7843] = 32'b00000000000000001110111001001011;
assign LUT_2[7844] = 32'b00000000000000000111100101011110;
assign LUT_2[7845] = 32'b00000000000000000100011101110111;
assign LUT_2[7846] = 32'b00000000000000001110011110011010;
assign LUT_2[7847] = 32'b00000000000000001011010110110011;
assign LUT_2[7848] = 32'b00000000000000000101111001010011;
assign LUT_2[7849] = 32'b00000000000000000010110001101100;
assign LUT_2[7850] = 32'b00000000000000001100110010001111;
assign LUT_2[7851] = 32'b00000000000000001001101010101000;
assign LUT_2[7852] = 32'b00000000000000000010010110111011;
assign LUT_2[7853] = 32'b11111111111111111111001111010100;
assign LUT_2[7854] = 32'b00000000000000001001001111110111;
assign LUT_2[7855] = 32'b00000000000000000110001000010000;
assign LUT_2[7856] = 32'b00000000000000000101101100000000;
assign LUT_2[7857] = 32'b00000000000000000010100100011001;
assign LUT_2[7858] = 32'b00000000000000001100100100111100;
assign LUT_2[7859] = 32'b00000000000000001001011101010101;
assign LUT_2[7860] = 32'b00000000000000000010001001101000;
assign LUT_2[7861] = 32'b11111111111111111111000010000001;
assign LUT_2[7862] = 32'b00000000000000001001000010100100;
assign LUT_2[7863] = 32'b00000000000000000101111010111101;
assign LUT_2[7864] = 32'b00000000000000000000011101011101;
assign LUT_2[7865] = 32'b11111111111111111101010101110110;
assign LUT_2[7866] = 32'b00000000000000000111010110011001;
assign LUT_2[7867] = 32'b00000000000000000100001110110010;
assign LUT_2[7868] = 32'b11111111111111111100111011000101;
assign LUT_2[7869] = 32'b11111111111111111001110011011110;
assign LUT_2[7870] = 32'b00000000000000000011110100000001;
assign LUT_2[7871] = 32'b00000000000000000000101100011010;
assign LUT_2[7872] = 32'b00000000000000000010110100110000;
assign LUT_2[7873] = 32'b11111111111111111111101101001001;
assign LUT_2[7874] = 32'b00000000000000001001101101101100;
assign LUT_2[7875] = 32'b00000000000000000110100110000101;
assign LUT_2[7876] = 32'b11111111111111111111010010011000;
assign LUT_2[7877] = 32'b11111111111111111100001010110001;
assign LUT_2[7878] = 32'b00000000000000000110001011010100;
assign LUT_2[7879] = 32'b00000000000000000011000011101101;
assign LUT_2[7880] = 32'b11111111111111111101100110001101;
assign LUT_2[7881] = 32'b11111111111111111010011110100110;
assign LUT_2[7882] = 32'b00000000000000000100011111001001;
assign LUT_2[7883] = 32'b00000000000000000001010111100010;
assign LUT_2[7884] = 32'b11111111111111111010000011110101;
assign LUT_2[7885] = 32'b11111111111111110110111100001110;
assign LUT_2[7886] = 32'b00000000000000000000111100110001;
assign LUT_2[7887] = 32'b11111111111111111101110101001010;
assign LUT_2[7888] = 32'b11111111111111111101011000111010;
assign LUT_2[7889] = 32'b11111111111111111010010001010011;
assign LUT_2[7890] = 32'b00000000000000000100010001110110;
assign LUT_2[7891] = 32'b00000000000000000001001010001111;
assign LUT_2[7892] = 32'b11111111111111111001110110100010;
assign LUT_2[7893] = 32'b11111111111111110110101110111011;
assign LUT_2[7894] = 32'b00000000000000000000101111011110;
assign LUT_2[7895] = 32'b11111111111111111101100111110111;
assign LUT_2[7896] = 32'b11111111111111111000001010010111;
assign LUT_2[7897] = 32'b11111111111111110101000010110000;
assign LUT_2[7898] = 32'b11111111111111111111000011010011;
assign LUT_2[7899] = 32'b11111111111111111011111011101100;
assign LUT_2[7900] = 32'b11111111111111110100100111111111;
assign LUT_2[7901] = 32'b11111111111111110001100000011000;
assign LUT_2[7902] = 32'b11111111111111111011100000111011;
assign LUT_2[7903] = 32'b11111111111111111000011001010100;
assign LUT_2[7904] = 32'b00000000000000000011010000011001;
assign LUT_2[7905] = 32'b00000000000000000000001000110010;
assign LUT_2[7906] = 32'b00000000000000001010001001010101;
assign LUT_2[7907] = 32'b00000000000000000111000001101110;
assign LUT_2[7908] = 32'b11111111111111111111101110000001;
assign LUT_2[7909] = 32'b11111111111111111100100110011010;
assign LUT_2[7910] = 32'b00000000000000000110100110111101;
assign LUT_2[7911] = 32'b00000000000000000011011111010110;
assign LUT_2[7912] = 32'b11111111111111111110000001110110;
assign LUT_2[7913] = 32'b11111111111111111010111010001111;
assign LUT_2[7914] = 32'b00000000000000000100111010110010;
assign LUT_2[7915] = 32'b00000000000000000001110011001011;
assign LUT_2[7916] = 32'b11111111111111111010011111011110;
assign LUT_2[7917] = 32'b11111111111111110111010111110111;
assign LUT_2[7918] = 32'b00000000000000000001011000011010;
assign LUT_2[7919] = 32'b11111111111111111110010000110011;
assign LUT_2[7920] = 32'b11111111111111111101110100100011;
assign LUT_2[7921] = 32'b11111111111111111010101100111100;
assign LUT_2[7922] = 32'b00000000000000000100101101011111;
assign LUT_2[7923] = 32'b00000000000000000001100101111000;
assign LUT_2[7924] = 32'b11111111111111111010010010001011;
assign LUT_2[7925] = 32'b11111111111111110111001010100100;
assign LUT_2[7926] = 32'b00000000000000000001001011000111;
assign LUT_2[7927] = 32'b11111111111111111110000011100000;
assign LUT_2[7928] = 32'b11111111111111111000100110000000;
assign LUT_2[7929] = 32'b11111111111111110101011110011001;
assign LUT_2[7930] = 32'b11111111111111111111011110111100;
assign LUT_2[7931] = 32'b11111111111111111100010111010101;
assign LUT_2[7932] = 32'b11111111111111110101000011101000;
assign LUT_2[7933] = 32'b11111111111111110001111100000001;
assign LUT_2[7934] = 32'b11111111111111111011111100100100;
assign LUT_2[7935] = 32'b11111111111111111000110100111101;
assign LUT_2[7936] = 32'b00000000000000001010010110100100;
assign LUT_2[7937] = 32'b00000000000000000111001110111101;
assign LUT_2[7938] = 32'b00000000000000010001001111100000;
assign LUT_2[7939] = 32'b00000000000000001110000111111001;
assign LUT_2[7940] = 32'b00000000000000000110110100001100;
assign LUT_2[7941] = 32'b00000000000000000011101100100101;
assign LUT_2[7942] = 32'b00000000000000001101101101001000;
assign LUT_2[7943] = 32'b00000000000000001010100101100001;
assign LUT_2[7944] = 32'b00000000000000000101001000000001;
assign LUT_2[7945] = 32'b00000000000000000010000000011010;
assign LUT_2[7946] = 32'b00000000000000001100000000111101;
assign LUT_2[7947] = 32'b00000000000000001000111001010110;
assign LUT_2[7948] = 32'b00000000000000000001100101101001;
assign LUT_2[7949] = 32'b11111111111111111110011110000010;
assign LUT_2[7950] = 32'b00000000000000001000011110100101;
assign LUT_2[7951] = 32'b00000000000000000101010110111110;
assign LUT_2[7952] = 32'b00000000000000000100111010101110;
assign LUT_2[7953] = 32'b00000000000000000001110011000111;
assign LUT_2[7954] = 32'b00000000000000001011110011101010;
assign LUT_2[7955] = 32'b00000000000000001000101100000011;
assign LUT_2[7956] = 32'b00000000000000000001011000010110;
assign LUT_2[7957] = 32'b11111111111111111110010000101111;
assign LUT_2[7958] = 32'b00000000000000001000010001010010;
assign LUT_2[7959] = 32'b00000000000000000101001001101011;
assign LUT_2[7960] = 32'b11111111111111111111101100001011;
assign LUT_2[7961] = 32'b11111111111111111100100100100100;
assign LUT_2[7962] = 32'b00000000000000000110100101000111;
assign LUT_2[7963] = 32'b00000000000000000011011101100000;
assign LUT_2[7964] = 32'b11111111111111111100001001110011;
assign LUT_2[7965] = 32'b11111111111111111001000010001100;
assign LUT_2[7966] = 32'b00000000000000000011000010101111;
assign LUT_2[7967] = 32'b11111111111111111111111011001000;
assign LUT_2[7968] = 32'b00000000000000001010110010001101;
assign LUT_2[7969] = 32'b00000000000000000111101010100110;
assign LUT_2[7970] = 32'b00000000000000010001101011001001;
assign LUT_2[7971] = 32'b00000000000000001110100011100010;
assign LUT_2[7972] = 32'b00000000000000000111001111110101;
assign LUT_2[7973] = 32'b00000000000000000100001000001110;
assign LUT_2[7974] = 32'b00000000000000001110001000110001;
assign LUT_2[7975] = 32'b00000000000000001011000001001010;
assign LUT_2[7976] = 32'b00000000000000000101100011101010;
assign LUT_2[7977] = 32'b00000000000000000010011100000011;
assign LUT_2[7978] = 32'b00000000000000001100011100100110;
assign LUT_2[7979] = 32'b00000000000000001001010100111111;
assign LUT_2[7980] = 32'b00000000000000000010000001010010;
assign LUT_2[7981] = 32'b11111111111111111110111001101011;
assign LUT_2[7982] = 32'b00000000000000001000111010001110;
assign LUT_2[7983] = 32'b00000000000000000101110010100111;
assign LUT_2[7984] = 32'b00000000000000000101010110010111;
assign LUT_2[7985] = 32'b00000000000000000010001110110000;
assign LUT_2[7986] = 32'b00000000000000001100001111010011;
assign LUT_2[7987] = 32'b00000000000000001001000111101100;
assign LUT_2[7988] = 32'b00000000000000000001110011111111;
assign LUT_2[7989] = 32'b11111111111111111110101100011000;
assign LUT_2[7990] = 32'b00000000000000001000101100111011;
assign LUT_2[7991] = 32'b00000000000000000101100101010100;
assign LUT_2[7992] = 32'b00000000000000000000000111110100;
assign LUT_2[7993] = 32'b11111111111111111101000000001101;
assign LUT_2[7994] = 32'b00000000000000000111000000110000;
assign LUT_2[7995] = 32'b00000000000000000011111001001001;
assign LUT_2[7996] = 32'b11111111111111111100100101011100;
assign LUT_2[7997] = 32'b11111111111111111001011101110101;
assign LUT_2[7998] = 32'b00000000000000000011011110011000;
assign LUT_2[7999] = 32'b00000000000000000000010110110001;
assign LUT_2[8000] = 32'b00000000000000000010011111000111;
assign LUT_2[8001] = 32'b11111111111111111111010111100000;
assign LUT_2[8002] = 32'b00000000000000001001011000000011;
assign LUT_2[8003] = 32'b00000000000000000110010000011100;
assign LUT_2[8004] = 32'b11111111111111111110111100101111;
assign LUT_2[8005] = 32'b11111111111111111011110101001000;
assign LUT_2[8006] = 32'b00000000000000000101110101101011;
assign LUT_2[8007] = 32'b00000000000000000010101110000100;
assign LUT_2[8008] = 32'b11111111111111111101010000100100;
assign LUT_2[8009] = 32'b11111111111111111010001000111101;
assign LUT_2[8010] = 32'b00000000000000000100001001100000;
assign LUT_2[8011] = 32'b00000000000000000001000001111001;
assign LUT_2[8012] = 32'b11111111111111111001101110001100;
assign LUT_2[8013] = 32'b11111111111111110110100110100101;
assign LUT_2[8014] = 32'b00000000000000000000100111001000;
assign LUT_2[8015] = 32'b11111111111111111101011111100001;
assign LUT_2[8016] = 32'b11111111111111111101000011010001;
assign LUT_2[8017] = 32'b11111111111111111001111011101010;
assign LUT_2[8018] = 32'b00000000000000000011111100001101;
assign LUT_2[8019] = 32'b00000000000000000000110100100110;
assign LUT_2[8020] = 32'b11111111111111111001100000111001;
assign LUT_2[8021] = 32'b11111111111111110110011001010010;
assign LUT_2[8022] = 32'b00000000000000000000011001110101;
assign LUT_2[8023] = 32'b11111111111111111101010010001110;
assign LUT_2[8024] = 32'b11111111111111110111110100101110;
assign LUT_2[8025] = 32'b11111111111111110100101101000111;
assign LUT_2[8026] = 32'b11111111111111111110101101101010;
assign LUT_2[8027] = 32'b11111111111111111011100110000011;
assign LUT_2[8028] = 32'b11111111111111110100010010010110;
assign LUT_2[8029] = 32'b11111111111111110001001010101111;
assign LUT_2[8030] = 32'b11111111111111111011001011010010;
assign LUT_2[8031] = 32'b11111111111111111000000011101011;
assign LUT_2[8032] = 32'b00000000000000000010111010110000;
assign LUT_2[8033] = 32'b11111111111111111111110011001001;
assign LUT_2[8034] = 32'b00000000000000001001110011101100;
assign LUT_2[8035] = 32'b00000000000000000110101100000101;
assign LUT_2[8036] = 32'b11111111111111111111011000011000;
assign LUT_2[8037] = 32'b11111111111111111100010000110001;
assign LUT_2[8038] = 32'b00000000000000000110010001010100;
assign LUT_2[8039] = 32'b00000000000000000011001001101101;
assign LUT_2[8040] = 32'b11111111111111111101101100001101;
assign LUT_2[8041] = 32'b11111111111111111010100100100110;
assign LUT_2[8042] = 32'b00000000000000000100100101001001;
assign LUT_2[8043] = 32'b00000000000000000001011101100010;
assign LUT_2[8044] = 32'b11111111111111111010001001110101;
assign LUT_2[8045] = 32'b11111111111111110111000010001110;
assign LUT_2[8046] = 32'b00000000000000000001000010110001;
assign LUT_2[8047] = 32'b11111111111111111101111011001010;
assign LUT_2[8048] = 32'b11111111111111111101011110111010;
assign LUT_2[8049] = 32'b11111111111111111010010111010011;
assign LUT_2[8050] = 32'b00000000000000000100010111110110;
assign LUT_2[8051] = 32'b00000000000000000001010000001111;
assign LUT_2[8052] = 32'b11111111111111111001111100100010;
assign LUT_2[8053] = 32'b11111111111111110110110100111011;
assign LUT_2[8054] = 32'b00000000000000000000110101011110;
assign LUT_2[8055] = 32'b11111111111111111101101101110111;
assign LUT_2[8056] = 32'b11111111111111111000010000010111;
assign LUT_2[8057] = 32'b11111111111111110101001000110000;
assign LUT_2[8058] = 32'b11111111111111111111001001010011;
assign LUT_2[8059] = 32'b11111111111111111100000001101100;
assign LUT_2[8060] = 32'b11111111111111110100101101111111;
assign LUT_2[8061] = 32'b11111111111111110001100110011000;
assign LUT_2[8062] = 32'b11111111111111111011100110111011;
assign LUT_2[8063] = 32'b11111111111111111000011111010100;
assign LUT_2[8064] = 32'b00000000000000001110101010110011;
assign LUT_2[8065] = 32'b00000000000000001011100011001100;
assign LUT_2[8066] = 32'b00000000000000010101100011101111;
assign LUT_2[8067] = 32'b00000000000000010010011100001000;
assign LUT_2[8068] = 32'b00000000000000001011001000011011;
assign LUT_2[8069] = 32'b00000000000000001000000000110100;
assign LUT_2[8070] = 32'b00000000000000010010000001010111;
assign LUT_2[8071] = 32'b00000000000000001110111001110000;
assign LUT_2[8072] = 32'b00000000000000001001011100010000;
assign LUT_2[8073] = 32'b00000000000000000110010100101001;
assign LUT_2[8074] = 32'b00000000000000010000010101001100;
assign LUT_2[8075] = 32'b00000000000000001101001101100101;
assign LUT_2[8076] = 32'b00000000000000000101111001111000;
assign LUT_2[8077] = 32'b00000000000000000010110010010001;
assign LUT_2[8078] = 32'b00000000000000001100110010110100;
assign LUT_2[8079] = 32'b00000000000000001001101011001101;
assign LUT_2[8080] = 32'b00000000000000001001001110111101;
assign LUT_2[8081] = 32'b00000000000000000110000111010110;
assign LUT_2[8082] = 32'b00000000000000010000000111111001;
assign LUT_2[8083] = 32'b00000000000000001101000000010010;
assign LUT_2[8084] = 32'b00000000000000000101101100100101;
assign LUT_2[8085] = 32'b00000000000000000010100100111110;
assign LUT_2[8086] = 32'b00000000000000001100100101100001;
assign LUT_2[8087] = 32'b00000000000000001001011101111010;
assign LUT_2[8088] = 32'b00000000000000000100000000011010;
assign LUT_2[8089] = 32'b00000000000000000000111000110011;
assign LUT_2[8090] = 32'b00000000000000001010111001010110;
assign LUT_2[8091] = 32'b00000000000000000111110001101111;
assign LUT_2[8092] = 32'b00000000000000000000011110000010;
assign LUT_2[8093] = 32'b11111111111111111101010110011011;
assign LUT_2[8094] = 32'b00000000000000000111010110111110;
assign LUT_2[8095] = 32'b00000000000000000100001111010111;
assign LUT_2[8096] = 32'b00000000000000001111000110011100;
assign LUT_2[8097] = 32'b00000000000000001011111110110101;
assign LUT_2[8098] = 32'b00000000000000010101111111011000;
assign LUT_2[8099] = 32'b00000000000000010010110111110001;
assign LUT_2[8100] = 32'b00000000000000001011100100000100;
assign LUT_2[8101] = 32'b00000000000000001000011100011101;
assign LUT_2[8102] = 32'b00000000000000010010011101000000;
assign LUT_2[8103] = 32'b00000000000000001111010101011001;
assign LUT_2[8104] = 32'b00000000000000001001110111111001;
assign LUT_2[8105] = 32'b00000000000000000110110000010010;
assign LUT_2[8106] = 32'b00000000000000010000110000110101;
assign LUT_2[8107] = 32'b00000000000000001101101001001110;
assign LUT_2[8108] = 32'b00000000000000000110010101100001;
assign LUT_2[8109] = 32'b00000000000000000011001101111010;
assign LUT_2[8110] = 32'b00000000000000001101001110011101;
assign LUT_2[8111] = 32'b00000000000000001010000110110110;
assign LUT_2[8112] = 32'b00000000000000001001101010100110;
assign LUT_2[8113] = 32'b00000000000000000110100010111111;
assign LUT_2[8114] = 32'b00000000000000010000100011100010;
assign LUT_2[8115] = 32'b00000000000000001101011011111011;
assign LUT_2[8116] = 32'b00000000000000000110001000001110;
assign LUT_2[8117] = 32'b00000000000000000011000000100111;
assign LUT_2[8118] = 32'b00000000000000001101000001001010;
assign LUT_2[8119] = 32'b00000000000000001001111001100011;
assign LUT_2[8120] = 32'b00000000000000000100011100000011;
assign LUT_2[8121] = 32'b00000000000000000001010100011100;
assign LUT_2[8122] = 32'b00000000000000001011010100111111;
assign LUT_2[8123] = 32'b00000000000000001000001101011000;
assign LUT_2[8124] = 32'b00000000000000000000111001101011;
assign LUT_2[8125] = 32'b11111111111111111101110010000100;
assign LUT_2[8126] = 32'b00000000000000000111110010100111;
assign LUT_2[8127] = 32'b00000000000000000100101011000000;
assign LUT_2[8128] = 32'b00000000000000000110110011010110;
assign LUT_2[8129] = 32'b00000000000000000011101011101111;
assign LUT_2[8130] = 32'b00000000000000001101101100010010;
assign LUT_2[8131] = 32'b00000000000000001010100100101011;
assign LUT_2[8132] = 32'b00000000000000000011010000111110;
assign LUT_2[8133] = 32'b00000000000000000000001001010111;
assign LUT_2[8134] = 32'b00000000000000001010001001111010;
assign LUT_2[8135] = 32'b00000000000000000111000010010011;
assign LUT_2[8136] = 32'b00000000000000000001100100110011;
assign LUT_2[8137] = 32'b11111111111111111110011101001100;
assign LUT_2[8138] = 32'b00000000000000001000011101101111;
assign LUT_2[8139] = 32'b00000000000000000101010110001000;
assign LUT_2[8140] = 32'b11111111111111111110000010011011;
assign LUT_2[8141] = 32'b11111111111111111010111010110100;
assign LUT_2[8142] = 32'b00000000000000000100111011010111;
assign LUT_2[8143] = 32'b00000000000000000001110011110000;
assign LUT_2[8144] = 32'b00000000000000000001010111100000;
assign LUT_2[8145] = 32'b11111111111111111110001111111001;
assign LUT_2[8146] = 32'b00000000000000001000010000011100;
assign LUT_2[8147] = 32'b00000000000000000101001000110101;
assign LUT_2[8148] = 32'b11111111111111111101110101001000;
assign LUT_2[8149] = 32'b11111111111111111010101101100001;
assign LUT_2[8150] = 32'b00000000000000000100101110000100;
assign LUT_2[8151] = 32'b00000000000000000001100110011101;
assign LUT_2[8152] = 32'b11111111111111111100001000111101;
assign LUT_2[8153] = 32'b11111111111111111001000001010110;
assign LUT_2[8154] = 32'b00000000000000000011000001111001;
assign LUT_2[8155] = 32'b11111111111111111111111010010010;
assign LUT_2[8156] = 32'b11111111111111111000100110100101;
assign LUT_2[8157] = 32'b11111111111111110101011110111110;
assign LUT_2[8158] = 32'b11111111111111111111011111100001;
assign LUT_2[8159] = 32'b11111111111111111100010111111010;
assign LUT_2[8160] = 32'b00000000000000000111001110111111;
assign LUT_2[8161] = 32'b00000000000000000100000111011000;
assign LUT_2[8162] = 32'b00000000000000001110000111111011;
assign LUT_2[8163] = 32'b00000000000000001011000000010100;
assign LUT_2[8164] = 32'b00000000000000000011101100100111;
assign LUT_2[8165] = 32'b00000000000000000000100101000000;
assign LUT_2[8166] = 32'b00000000000000001010100101100011;
assign LUT_2[8167] = 32'b00000000000000000111011101111100;
assign LUT_2[8168] = 32'b00000000000000000010000000011100;
assign LUT_2[8169] = 32'b11111111111111111110111000110101;
assign LUT_2[8170] = 32'b00000000000000001000111001011000;
assign LUT_2[8171] = 32'b00000000000000000101110001110001;
assign LUT_2[8172] = 32'b11111111111111111110011110000100;
assign LUT_2[8173] = 32'b11111111111111111011010110011101;
assign LUT_2[8174] = 32'b00000000000000000101010111000000;
assign LUT_2[8175] = 32'b00000000000000000010001111011001;
assign LUT_2[8176] = 32'b00000000000000000001110011001001;
assign LUT_2[8177] = 32'b11111111111111111110101011100010;
assign LUT_2[8178] = 32'b00000000000000001000101100000101;
assign LUT_2[8179] = 32'b00000000000000000101100100011110;
assign LUT_2[8180] = 32'b11111111111111111110010000110001;
assign LUT_2[8181] = 32'b11111111111111111011001001001010;
assign LUT_2[8182] = 32'b00000000000000000101001001101101;
assign LUT_2[8183] = 32'b00000000000000000010000010000110;
assign LUT_2[8184] = 32'b11111111111111111100100100100110;
assign LUT_2[8185] = 32'b11111111111111111001011100111111;
assign LUT_2[8186] = 32'b00000000000000000011011101100010;
assign LUT_2[8187] = 32'b00000000000000000000010101111011;
assign LUT_2[8188] = 32'b11111111111111111001000010001110;
assign LUT_2[8189] = 32'b11111111111111110101111010100111;
assign LUT_2[8190] = 32'b11111111111111111111111011001010;
assign LUT_2[8191] = 32'b11111111111111111100110011100011;
assign LUT_2[8192] = 32'b11111111111111111001010101111110;
assign LUT_2[8193] = 32'b11111111111111110110001110010111;
assign LUT_2[8194] = 32'b00000000000000000000001110111010;
assign LUT_2[8195] = 32'b11111111111111111101000111010011;
assign LUT_2[8196] = 32'b11111111111111110101110011100110;
assign LUT_2[8197] = 32'b11111111111111110010101011111111;
assign LUT_2[8198] = 32'b11111111111111111100101100100010;
assign LUT_2[8199] = 32'b11111111111111111001100100111011;
assign LUT_2[8200] = 32'b11111111111111110100000111011011;
assign LUT_2[8201] = 32'b11111111111111110000111111110100;
assign LUT_2[8202] = 32'b11111111111111111011000000010111;
assign LUT_2[8203] = 32'b11111111111111110111111000110000;
assign LUT_2[8204] = 32'b11111111111111110000100101000011;
assign LUT_2[8205] = 32'b11111111111111101101011101011100;
assign LUT_2[8206] = 32'b11111111111111110111011101111111;
assign LUT_2[8207] = 32'b11111111111111110100010110011000;
assign LUT_2[8208] = 32'b11111111111111110011111010001000;
assign LUT_2[8209] = 32'b11111111111111110000110010100001;
assign LUT_2[8210] = 32'b11111111111111111010110011000100;
assign LUT_2[8211] = 32'b11111111111111110111101011011101;
assign LUT_2[8212] = 32'b11111111111111110000010111110000;
assign LUT_2[8213] = 32'b11111111111111101101010000001001;
assign LUT_2[8214] = 32'b11111111111111110111010000101100;
assign LUT_2[8215] = 32'b11111111111111110100001001000101;
assign LUT_2[8216] = 32'b11111111111111101110101011100101;
assign LUT_2[8217] = 32'b11111111111111101011100011111110;
assign LUT_2[8218] = 32'b11111111111111110101100100100001;
assign LUT_2[8219] = 32'b11111111111111110010011100111010;
assign LUT_2[8220] = 32'b11111111111111101011001001001101;
assign LUT_2[8221] = 32'b11111111111111101000000001100110;
assign LUT_2[8222] = 32'b11111111111111110010000010001001;
assign LUT_2[8223] = 32'b11111111111111101110111010100010;
assign LUT_2[8224] = 32'b11111111111111111001110001100111;
assign LUT_2[8225] = 32'b11111111111111110110101010000000;
assign LUT_2[8226] = 32'b00000000000000000000101010100011;
assign LUT_2[8227] = 32'b11111111111111111101100010111100;
assign LUT_2[8228] = 32'b11111111111111110110001111001111;
assign LUT_2[8229] = 32'b11111111111111110011000111101000;
assign LUT_2[8230] = 32'b11111111111111111101001000001011;
assign LUT_2[8231] = 32'b11111111111111111010000000100100;
assign LUT_2[8232] = 32'b11111111111111110100100011000100;
assign LUT_2[8233] = 32'b11111111111111110001011011011101;
assign LUT_2[8234] = 32'b11111111111111111011011100000000;
assign LUT_2[8235] = 32'b11111111111111111000010100011001;
assign LUT_2[8236] = 32'b11111111111111110001000000101100;
assign LUT_2[8237] = 32'b11111111111111101101111001000101;
assign LUT_2[8238] = 32'b11111111111111110111111001101000;
assign LUT_2[8239] = 32'b11111111111111110100110010000001;
assign LUT_2[8240] = 32'b11111111111111110100010101110001;
assign LUT_2[8241] = 32'b11111111111111110001001110001010;
assign LUT_2[8242] = 32'b11111111111111111011001110101101;
assign LUT_2[8243] = 32'b11111111111111111000000111000110;
assign LUT_2[8244] = 32'b11111111111111110000110011011001;
assign LUT_2[8245] = 32'b11111111111111101101101011110010;
assign LUT_2[8246] = 32'b11111111111111110111101100010101;
assign LUT_2[8247] = 32'b11111111111111110100100100101110;
assign LUT_2[8248] = 32'b11111111111111101111000111001110;
assign LUT_2[8249] = 32'b11111111111111101011111111100111;
assign LUT_2[8250] = 32'b11111111111111110110000000001010;
assign LUT_2[8251] = 32'b11111111111111110010111000100011;
assign LUT_2[8252] = 32'b11111111111111101011100100110110;
assign LUT_2[8253] = 32'b11111111111111101000011101001111;
assign LUT_2[8254] = 32'b11111111111111110010011101110010;
assign LUT_2[8255] = 32'b11111111111111101111010110001011;
assign LUT_2[8256] = 32'b11111111111111110001011110100001;
assign LUT_2[8257] = 32'b11111111111111101110010110111010;
assign LUT_2[8258] = 32'b11111111111111111000010111011101;
assign LUT_2[8259] = 32'b11111111111111110101001111110110;
assign LUT_2[8260] = 32'b11111111111111101101111100001001;
assign LUT_2[8261] = 32'b11111111111111101010110100100010;
assign LUT_2[8262] = 32'b11111111111111110100110101000101;
assign LUT_2[8263] = 32'b11111111111111110001101101011110;
assign LUT_2[8264] = 32'b11111111111111101100001111111110;
assign LUT_2[8265] = 32'b11111111111111101001001000010111;
assign LUT_2[8266] = 32'b11111111111111110011001000111010;
assign LUT_2[8267] = 32'b11111111111111110000000001010011;
assign LUT_2[8268] = 32'b11111111111111101000101101100110;
assign LUT_2[8269] = 32'b11111111111111100101100101111111;
assign LUT_2[8270] = 32'b11111111111111101111100110100010;
assign LUT_2[8271] = 32'b11111111111111101100011110111011;
assign LUT_2[8272] = 32'b11111111111111101100000010101011;
assign LUT_2[8273] = 32'b11111111111111101000111011000100;
assign LUT_2[8274] = 32'b11111111111111110010111011100111;
assign LUT_2[8275] = 32'b11111111111111101111110100000000;
assign LUT_2[8276] = 32'b11111111111111101000100000010011;
assign LUT_2[8277] = 32'b11111111111111100101011000101100;
assign LUT_2[8278] = 32'b11111111111111101111011001001111;
assign LUT_2[8279] = 32'b11111111111111101100010001101000;
assign LUT_2[8280] = 32'b11111111111111100110110100001000;
assign LUT_2[8281] = 32'b11111111111111100011101100100001;
assign LUT_2[8282] = 32'b11111111111111101101101101000100;
assign LUT_2[8283] = 32'b11111111111111101010100101011101;
assign LUT_2[8284] = 32'b11111111111111100011010001110000;
assign LUT_2[8285] = 32'b11111111111111100000001010001001;
assign LUT_2[8286] = 32'b11111111111111101010001010101100;
assign LUT_2[8287] = 32'b11111111111111100111000011000101;
assign LUT_2[8288] = 32'b11111111111111110001111010001010;
assign LUT_2[8289] = 32'b11111111111111101110110010100011;
assign LUT_2[8290] = 32'b11111111111111111000110011000110;
assign LUT_2[8291] = 32'b11111111111111110101101011011111;
assign LUT_2[8292] = 32'b11111111111111101110010111110010;
assign LUT_2[8293] = 32'b11111111111111101011010000001011;
assign LUT_2[8294] = 32'b11111111111111110101010000101110;
assign LUT_2[8295] = 32'b11111111111111110010001001000111;
assign LUT_2[8296] = 32'b11111111111111101100101011100111;
assign LUT_2[8297] = 32'b11111111111111101001100100000000;
assign LUT_2[8298] = 32'b11111111111111110011100100100011;
assign LUT_2[8299] = 32'b11111111111111110000011100111100;
assign LUT_2[8300] = 32'b11111111111111101001001001001111;
assign LUT_2[8301] = 32'b11111111111111100110000001101000;
assign LUT_2[8302] = 32'b11111111111111110000000010001011;
assign LUT_2[8303] = 32'b11111111111111101100111010100100;
assign LUT_2[8304] = 32'b11111111111111101100011110010100;
assign LUT_2[8305] = 32'b11111111111111101001010110101101;
assign LUT_2[8306] = 32'b11111111111111110011010111010000;
assign LUT_2[8307] = 32'b11111111111111110000001111101001;
assign LUT_2[8308] = 32'b11111111111111101000111011111100;
assign LUT_2[8309] = 32'b11111111111111100101110100010101;
assign LUT_2[8310] = 32'b11111111111111101111110100111000;
assign LUT_2[8311] = 32'b11111111111111101100101101010001;
assign LUT_2[8312] = 32'b11111111111111100111001111110001;
assign LUT_2[8313] = 32'b11111111111111100100001000001010;
assign LUT_2[8314] = 32'b11111111111111101110001000101101;
assign LUT_2[8315] = 32'b11111111111111101011000001000110;
assign LUT_2[8316] = 32'b11111111111111100011101101011001;
assign LUT_2[8317] = 32'b11111111111111100000100101110010;
assign LUT_2[8318] = 32'b11111111111111101010100110010101;
assign LUT_2[8319] = 32'b11111111111111100111011110101110;
assign LUT_2[8320] = 32'b11111111111111111101101010001101;
assign LUT_2[8321] = 32'b11111111111111111010100010100110;
assign LUT_2[8322] = 32'b00000000000000000100100011001001;
assign LUT_2[8323] = 32'b00000000000000000001011011100010;
assign LUT_2[8324] = 32'b11111111111111111010000111110101;
assign LUT_2[8325] = 32'b11111111111111110111000000001110;
assign LUT_2[8326] = 32'b00000000000000000001000000110001;
assign LUT_2[8327] = 32'b11111111111111111101111001001010;
assign LUT_2[8328] = 32'b11111111111111111000011011101010;
assign LUT_2[8329] = 32'b11111111111111110101010100000011;
assign LUT_2[8330] = 32'b11111111111111111111010100100110;
assign LUT_2[8331] = 32'b11111111111111111100001100111111;
assign LUT_2[8332] = 32'b11111111111111110100111001010010;
assign LUT_2[8333] = 32'b11111111111111110001110001101011;
assign LUT_2[8334] = 32'b11111111111111111011110010001110;
assign LUT_2[8335] = 32'b11111111111111111000101010100111;
assign LUT_2[8336] = 32'b11111111111111111000001110010111;
assign LUT_2[8337] = 32'b11111111111111110101000110110000;
assign LUT_2[8338] = 32'b11111111111111111111000111010011;
assign LUT_2[8339] = 32'b11111111111111111011111111101100;
assign LUT_2[8340] = 32'b11111111111111110100101011111111;
assign LUT_2[8341] = 32'b11111111111111110001100100011000;
assign LUT_2[8342] = 32'b11111111111111111011100100111011;
assign LUT_2[8343] = 32'b11111111111111111000011101010100;
assign LUT_2[8344] = 32'b11111111111111110010111111110100;
assign LUT_2[8345] = 32'b11111111111111101111111000001101;
assign LUT_2[8346] = 32'b11111111111111111001111000110000;
assign LUT_2[8347] = 32'b11111111111111110110110001001001;
assign LUT_2[8348] = 32'b11111111111111101111011101011100;
assign LUT_2[8349] = 32'b11111111111111101100010101110101;
assign LUT_2[8350] = 32'b11111111111111110110010110011000;
assign LUT_2[8351] = 32'b11111111111111110011001110110001;
assign LUT_2[8352] = 32'b11111111111111111110000101110110;
assign LUT_2[8353] = 32'b11111111111111111010111110001111;
assign LUT_2[8354] = 32'b00000000000000000100111110110010;
assign LUT_2[8355] = 32'b00000000000000000001110111001011;
assign LUT_2[8356] = 32'b11111111111111111010100011011110;
assign LUT_2[8357] = 32'b11111111111111110111011011110111;
assign LUT_2[8358] = 32'b00000000000000000001011100011010;
assign LUT_2[8359] = 32'b11111111111111111110010100110011;
assign LUT_2[8360] = 32'b11111111111111111000110111010011;
assign LUT_2[8361] = 32'b11111111111111110101101111101100;
assign LUT_2[8362] = 32'b11111111111111111111110000001111;
assign LUT_2[8363] = 32'b11111111111111111100101000101000;
assign LUT_2[8364] = 32'b11111111111111110101010100111011;
assign LUT_2[8365] = 32'b11111111111111110010001101010100;
assign LUT_2[8366] = 32'b11111111111111111100001101110111;
assign LUT_2[8367] = 32'b11111111111111111001000110010000;
assign LUT_2[8368] = 32'b11111111111111111000101010000000;
assign LUT_2[8369] = 32'b11111111111111110101100010011001;
assign LUT_2[8370] = 32'b11111111111111111111100010111100;
assign LUT_2[8371] = 32'b11111111111111111100011011010101;
assign LUT_2[8372] = 32'b11111111111111110101000111101000;
assign LUT_2[8373] = 32'b11111111111111110010000000000001;
assign LUT_2[8374] = 32'b11111111111111111100000000100100;
assign LUT_2[8375] = 32'b11111111111111111000111000111101;
assign LUT_2[8376] = 32'b11111111111111110011011011011101;
assign LUT_2[8377] = 32'b11111111111111110000010011110110;
assign LUT_2[8378] = 32'b11111111111111111010010100011001;
assign LUT_2[8379] = 32'b11111111111111110111001100110010;
assign LUT_2[8380] = 32'b11111111111111101111111001000101;
assign LUT_2[8381] = 32'b11111111111111101100110001011110;
assign LUT_2[8382] = 32'b11111111111111110110110010000001;
assign LUT_2[8383] = 32'b11111111111111110011101010011010;
assign LUT_2[8384] = 32'b11111111111111110101110010110000;
assign LUT_2[8385] = 32'b11111111111111110010101011001001;
assign LUT_2[8386] = 32'b11111111111111111100101011101100;
assign LUT_2[8387] = 32'b11111111111111111001100100000101;
assign LUT_2[8388] = 32'b11111111111111110010010000011000;
assign LUT_2[8389] = 32'b11111111111111101111001000110001;
assign LUT_2[8390] = 32'b11111111111111111001001001010100;
assign LUT_2[8391] = 32'b11111111111111110110000001101101;
assign LUT_2[8392] = 32'b11111111111111110000100100001101;
assign LUT_2[8393] = 32'b11111111111111101101011100100110;
assign LUT_2[8394] = 32'b11111111111111110111011101001001;
assign LUT_2[8395] = 32'b11111111111111110100010101100010;
assign LUT_2[8396] = 32'b11111111111111101101000001110101;
assign LUT_2[8397] = 32'b11111111111111101001111010001110;
assign LUT_2[8398] = 32'b11111111111111110011111010110001;
assign LUT_2[8399] = 32'b11111111111111110000110011001010;
assign LUT_2[8400] = 32'b11111111111111110000010110111010;
assign LUT_2[8401] = 32'b11111111111111101101001111010011;
assign LUT_2[8402] = 32'b11111111111111110111001111110110;
assign LUT_2[8403] = 32'b11111111111111110100001000001111;
assign LUT_2[8404] = 32'b11111111111111101100110100100010;
assign LUT_2[8405] = 32'b11111111111111101001101100111011;
assign LUT_2[8406] = 32'b11111111111111110011101101011110;
assign LUT_2[8407] = 32'b11111111111111110000100101110111;
assign LUT_2[8408] = 32'b11111111111111101011001000010111;
assign LUT_2[8409] = 32'b11111111111111101000000000110000;
assign LUT_2[8410] = 32'b11111111111111110010000001010011;
assign LUT_2[8411] = 32'b11111111111111101110111001101100;
assign LUT_2[8412] = 32'b11111111111111100111100101111111;
assign LUT_2[8413] = 32'b11111111111111100100011110011000;
assign LUT_2[8414] = 32'b11111111111111101110011110111011;
assign LUT_2[8415] = 32'b11111111111111101011010111010100;
assign LUT_2[8416] = 32'b11111111111111110110001110011001;
assign LUT_2[8417] = 32'b11111111111111110011000110110010;
assign LUT_2[8418] = 32'b11111111111111111101000111010101;
assign LUT_2[8419] = 32'b11111111111111111001111111101110;
assign LUT_2[8420] = 32'b11111111111111110010101100000001;
assign LUT_2[8421] = 32'b11111111111111101111100100011010;
assign LUT_2[8422] = 32'b11111111111111111001100100111101;
assign LUT_2[8423] = 32'b11111111111111110110011101010110;
assign LUT_2[8424] = 32'b11111111111111110000111111110110;
assign LUT_2[8425] = 32'b11111111111111101101111000001111;
assign LUT_2[8426] = 32'b11111111111111110111111000110010;
assign LUT_2[8427] = 32'b11111111111111110100110001001011;
assign LUT_2[8428] = 32'b11111111111111101101011101011110;
assign LUT_2[8429] = 32'b11111111111111101010010101110111;
assign LUT_2[8430] = 32'b11111111111111110100010110011010;
assign LUT_2[8431] = 32'b11111111111111110001001110110011;
assign LUT_2[8432] = 32'b11111111111111110000110010100011;
assign LUT_2[8433] = 32'b11111111111111101101101010111100;
assign LUT_2[8434] = 32'b11111111111111110111101011011111;
assign LUT_2[8435] = 32'b11111111111111110100100011111000;
assign LUT_2[8436] = 32'b11111111111111101101010000001011;
assign LUT_2[8437] = 32'b11111111111111101010001000100100;
assign LUT_2[8438] = 32'b11111111111111110100001001000111;
assign LUT_2[8439] = 32'b11111111111111110001000001100000;
assign LUT_2[8440] = 32'b11111111111111101011100100000000;
assign LUT_2[8441] = 32'b11111111111111101000011100011001;
assign LUT_2[8442] = 32'b11111111111111110010011100111100;
assign LUT_2[8443] = 32'b11111111111111101111010101010101;
assign LUT_2[8444] = 32'b11111111111111101000000001101000;
assign LUT_2[8445] = 32'b11111111111111100100111010000001;
assign LUT_2[8446] = 32'b11111111111111101110111010100100;
assign LUT_2[8447] = 32'b11111111111111101011110010111101;
assign LUT_2[8448] = 32'b11111111111111111101010100100100;
assign LUT_2[8449] = 32'b11111111111111111010001100111101;
assign LUT_2[8450] = 32'b00000000000000000100001101100000;
assign LUT_2[8451] = 32'b00000000000000000001000101111001;
assign LUT_2[8452] = 32'b11111111111111111001110010001100;
assign LUT_2[8453] = 32'b11111111111111110110101010100101;
assign LUT_2[8454] = 32'b00000000000000000000101011001000;
assign LUT_2[8455] = 32'b11111111111111111101100011100001;
assign LUT_2[8456] = 32'b11111111111111111000000110000001;
assign LUT_2[8457] = 32'b11111111111111110100111110011010;
assign LUT_2[8458] = 32'b11111111111111111110111110111101;
assign LUT_2[8459] = 32'b11111111111111111011110111010110;
assign LUT_2[8460] = 32'b11111111111111110100100011101001;
assign LUT_2[8461] = 32'b11111111111111110001011100000010;
assign LUT_2[8462] = 32'b11111111111111111011011100100101;
assign LUT_2[8463] = 32'b11111111111111111000010100111110;
assign LUT_2[8464] = 32'b11111111111111110111111000101110;
assign LUT_2[8465] = 32'b11111111111111110100110001000111;
assign LUT_2[8466] = 32'b11111111111111111110110001101010;
assign LUT_2[8467] = 32'b11111111111111111011101010000011;
assign LUT_2[8468] = 32'b11111111111111110100010110010110;
assign LUT_2[8469] = 32'b11111111111111110001001110101111;
assign LUT_2[8470] = 32'b11111111111111111011001111010010;
assign LUT_2[8471] = 32'b11111111111111111000000111101011;
assign LUT_2[8472] = 32'b11111111111111110010101010001011;
assign LUT_2[8473] = 32'b11111111111111101111100010100100;
assign LUT_2[8474] = 32'b11111111111111111001100011000111;
assign LUT_2[8475] = 32'b11111111111111110110011011100000;
assign LUT_2[8476] = 32'b11111111111111101111000111110011;
assign LUT_2[8477] = 32'b11111111111111101100000000001100;
assign LUT_2[8478] = 32'b11111111111111110110000000101111;
assign LUT_2[8479] = 32'b11111111111111110010111001001000;
assign LUT_2[8480] = 32'b11111111111111111101110000001101;
assign LUT_2[8481] = 32'b11111111111111111010101000100110;
assign LUT_2[8482] = 32'b00000000000000000100101001001001;
assign LUT_2[8483] = 32'b00000000000000000001100001100010;
assign LUT_2[8484] = 32'b11111111111111111010001101110101;
assign LUT_2[8485] = 32'b11111111111111110111000110001110;
assign LUT_2[8486] = 32'b00000000000000000001000110110001;
assign LUT_2[8487] = 32'b11111111111111111101111111001010;
assign LUT_2[8488] = 32'b11111111111111111000100001101010;
assign LUT_2[8489] = 32'b11111111111111110101011010000011;
assign LUT_2[8490] = 32'b11111111111111111111011010100110;
assign LUT_2[8491] = 32'b11111111111111111100010010111111;
assign LUT_2[8492] = 32'b11111111111111110100111111010010;
assign LUT_2[8493] = 32'b11111111111111110001110111101011;
assign LUT_2[8494] = 32'b11111111111111111011111000001110;
assign LUT_2[8495] = 32'b11111111111111111000110000100111;
assign LUT_2[8496] = 32'b11111111111111111000010100010111;
assign LUT_2[8497] = 32'b11111111111111110101001100110000;
assign LUT_2[8498] = 32'b11111111111111111111001101010011;
assign LUT_2[8499] = 32'b11111111111111111100000101101100;
assign LUT_2[8500] = 32'b11111111111111110100110001111111;
assign LUT_2[8501] = 32'b11111111111111110001101010011000;
assign LUT_2[8502] = 32'b11111111111111111011101010111011;
assign LUT_2[8503] = 32'b11111111111111111000100011010100;
assign LUT_2[8504] = 32'b11111111111111110011000101110100;
assign LUT_2[8505] = 32'b11111111111111101111111110001101;
assign LUT_2[8506] = 32'b11111111111111111001111110110000;
assign LUT_2[8507] = 32'b11111111111111110110110111001001;
assign LUT_2[8508] = 32'b11111111111111101111100011011100;
assign LUT_2[8509] = 32'b11111111111111101100011011110101;
assign LUT_2[8510] = 32'b11111111111111110110011100011000;
assign LUT_2[8511] = 32'b11111111111111110011010100110001;
assign LUT_2[8512] = 32'b11111111111111110101011101000111;
assign LUT_2[8513] = 32'b11111111111111110010010101100000;
assign LUT_2[8514] = 32'b11111111111111111100010110000011;
assign LUT_2[8515] = 32'b11111111111111111001001110011100;
assign LUT_2[8516] = 32'b11111111111111110001111010101111;
assign LUT_2[8517] = 32'b11111111111111101110110011001000;
assign LUT_2[8518] = 32'b11111111111111111000110011101011;
assign LUT_2[8519] = 32'b11111111111111110101101100000100;
assign LUT_2[8520] = 32'b11111111111111110000001110100100;
assign LUT_2[8521] = 32'b11111111111111101101000110111101;
assign LUT_2[8522] = 32'b11111111111111110111000111100000;
assign LUT_2[8523] = 32'b11111111111111110011111111111001;
assign LUT_2[8524] = 32'b11111111111111101100101100001100;
assign LUT_2[8525] = 32'b11111111111111101001100100100101;
assign LUT_2[8526] = 32'b11111111111111110011100101001000;
assign LUT_2[8527] = 32'b11111111111111110000011101100001;
assign LUT_2[8528] = 32'b11111111111111110000000001010001;
assign LUT_2[8529] = 32'b11111111111111101100111001101010;
assign LUT_2[8530] = 32'b11111111111111110110111010001101;
assign LUT_2[8531] = 32'b11111111111111110011110010100110;
assign LUT_2[8532] = 32'b11111111111111101100011110111001;
assign LUT_2[8533] = 32'b11111111111111101001010111010010;
assign LUT_2[8534] = 32'b11111111111111110011010111110101;
assign LUT_2[8535] = 32'b11111111111111110000010000001110;
assign LUT_2[8536] = 32'b11111111111111101010110010101110;
assign LUT_2[8537] = 32'b11111111111111100111101011000111;
assign LUT_2[8538] = 32'b11111111111111110001101011101010;
assign LUT_2[8539] = 32'b11111111111111101110100100000011;
assign LUT_2[8540] = 32'b11111111111111100111010000010110;
assign LUT_2[8541] = 32'b11111111111111100100001000101111;
assign LUT_2[8542] = 32'b11111111111111101110001001010010;
assign LUT_2[8543] = 32'b11111111111111101011000001101011;
assign LUT_2[8544] = 32'b11111111111111110101111000110000;
assign LUT_2[8545] = 32'b11111111111111110010110001001001;
assign LUT_2[8546] = 32'b11111111111111111100110001101100;
assign LUT_2[8547] = 32'b11111111111111111001101010000101;
assign LUT_2[8548] = 32'b11111111111111110010010110011000;
assign LUT_2[8549] = 32'b11111111111111101111001110110001;
assign LUT_2[8550] = 32'b11111111111111111001001111010100;
assign LUT_2[8551] = 32'b11111111111111110110000111101101;
assign LUT_2[8552] = 32'b11111111111111110000101010001101;
assign LUT_2[8553] = 32'b11111111111111101101100010100110;
assign LUT_2[8554] = 32'b11111111111111110111100011001001;
assign LUT_2[8555] = 32'b11111111111111110100011011100010;
assign LUT_2[8556] = 32'b11111111111111101101000111110101;
assign LUT_2[8557] = 32'b11111111111111101010000000001110;
assign LUT_2[8558] = 32'b11111111111111110100000000110001;
assign LUT_2[8559] = 32'b11111111111111110000111001001010;
assign LUT_2[8560] = 32'b11111111111111110000011100111010;
assign LUT_2[8561] = 32'b11111111111111101101010101010011;
assign LUT_2[8562] = 32'b11111111111111110111010101110110;
assign LUT_2[8563] = 32'b11111111111111110100001110001111;
assign LUT_2[8564] = 32'b11111111111111101100111010100010;
assign LUT_2[8565] = 32'b11111111111111101001110010111011;
assign LUT_2[8566] = 32'b11111111111111110011110011011110;
assign LUT_2[8567] = 32'b11111111111111110000101011110111;
assign LUT_2[8568] = 32'b11111111111111101011001110010111;
assign LUT_2[8569] = 32'b11111111111111101000000110110000;
assign LUT_2[8570] = 32'b11111111111111110010000111010011;
assign LUT_2[8571] = 32'b11111111111111101110111111101100;
assign LUT_2[8572] = 32'b11111111111111100111101011111111;
assign LUT_2[8573] = 32'b11111111111111100100100100011000;
assign LUT_2[8574] = 32'b11111111111111101110100100111011;
assign LUT_2[8575] = 32'b11111111111111101011011101010100;
assign LUT_2[8576] = 32'b00000000000000000001101000110011;
assign LUT_2[8577] = 32'b11111111111111111110100001001100;
assign LUT_2[8578] = 32'b00000000000000001000100001101111;
assign LUT_2[8579] = 32'b00000000000000000101011010001000;
assign LUT_2[8580] = 32'b11111111111111111110000110011011;
assign LUT_2[8581] = 32'b11111111111111111010111110110100;
assign LUT_2[8582] = 32'b00000000000000000100111111010111;
assign LUT_2[8583] = 32'b00000000000000000001110111110000;
assign LUT_2[8584] = 32'b11111111111111111100011010010000;
assign LUT_2[8585] = 32'b11111111111111111001010010101001;
assign LUT_2[8586] = 32'b00000000000000000011010011001100;
assign LUT_2[8587] = 32'b00000000000000000000001011100101;
assign LUT_2[8588] = 32'b11111111111111111000110111111000;
assign LUT_2[8589] = 32'b11111111111111110101110000010001;
assign LUT_2[8590] = 32'b11111111111111111111110000110100;
assign LUT_2[8591] = 32'b11111111111111111100101001001101;
assign LUT_2[8592] = 32'b11111111111111111100001100111101;
assign LUT_2[8593] = 32'b11111111111111111001000101010110;
assign LUT_2[8594] = 32'b00000000000000000011000101111001;
assign LUT_2[8595] = 32'b11111111111111111111111110010010;
assign LUT_2[8596] = 32'b11111111111111111000101010100101;
assign LUT_2[8597] = 32'b11111111111111110101100010111110;
assign LUT_2[8598] = 32'b11111111111111111111100011100001;
assign LUT_2[8599] = 32'b11111111111111111100011011111010;
assign LUT_2[8600] = 32'b11111111111111110110111110011010;
assign LUT_2[8601] = 32'b11111111111111110011110110110011;
assign LUT_2[8602] = 32'b11111111111111111101110111010110;
assign LUT_2[8603] = 32'b11111111111111111010101111101111;
assign LUT_2[8604] = 32'b11111111111111110011011100000010;
assign LUT_2[8605] = 32'b11111111111111110000010100011011;
assign LUT_2[8606] = 32'b11111111111111111010010100111110;
assign LUT_2[8607] = 32'b11111111111111110111001101010111;
assign LUT_2[8608] = 32'b00000000000000000010000100011100;
assign LUT_2[8609] = 32'b11111111111111111110111100110101;
assign LUT_2[8610] = 32'b00000000000000001000111101011000;
assign LUT_2[8611] = 32'b00000000000000000101110101110001;
assign LUT_2[8612] = 32'b11111111111111111110100010000100;
assign LUT_2[8613] = 32'b11111111111111111011011010011101;
assign LUT_2[8614] = 32'b00000000000000000101011011000000;
assign LUT_2[8615] = 32'b00000000000000000010010011011001;
assign LUT_2[8616] = 32'b11111111111111111100110101111001;
assign LUT_2[8617] = 32'b11111111111111111001101110010010;
assign LUT_2[8618] = 32'b00000000000000000011101110110101;
assign LUT_2[8619] = 32'b00000000000000000000100111001110;
assign LUT_2[8620] = 32'b11111111111111111001010011100001;
assign LUT_2[8621] = 32'b11111111111111110110001011111010;
assign LUT_2[8622] = 32'b00000000000000000000001100011101;
assign LUT_2[8623] = 32'b11111111111111111101000100110110;
assign LUT_2[8624] = 32'b11111111111111111100101000100110;
assign LUT_2[8625] = 32'b11111111111111111001100000111111;
assign LUT_2[8626] = 32'b00000000000000000011100001100010;
assign LUT_2[8627] = 32'b00000000000000000000011001111011;
assign LUT_2[8628] = 32'b11111111111111111001000110001110;
assign LUT_2[8629] = 32'b11111111111111110101111110100111;
assign LUT_2[8630] = 32'b11111111111111111111111111001010;
assign LUT_2[8631] = 32'b11111111111111111100110111100011;
assign LUT_2[8632] = 32'b11111111111111110111011010000011;
assign LUT_2[8633] = 32'b11111111111111110100010010011100;
assign LUT_2[8634] = 32'b11111111111111111110010010111111;
assign LUT_2[8635] = 32'b11111111111111111011001011011000;
assign LUT_2[8636] = 32'b11111111111111110011110111101011;
assign LUT_2[8637] = 32'b11111111111111110000110000000100;
assign LUT_2[8638] = 32'b11111111111111111010110000100111;
assign LUT_2[8639] = 32'b11111111111111110111101001000000;
assign LUT_2[8640] = 32'b11111111111111111001110001010110;
assign LUT_2[8641] = 32'b11111111111111110110101001101111;
assign LUT_2[8642] = 32'b00000000000000000000101010010010;
assign LUT_2[8643] = 32'b11111111111111111101100010101011;
assign LUT_2[8644] = 32'b11111111111111110110001110111110;
assign LUT_2[8645] = 32'b11111111111111110011000111010111;
assign LUT_2[8646] = 32'b11111111111111111101000111111010;
assign LUT_2[8647] = 32'b11111111111111111010000000010011;
assign LUT_2[8648] = 32'b11111111111111110100100010110011;
assign LUT_2[8649] = 32'b11111111111111110001011011001100;
assign LUT_2[8650] = 32'b11111111111111111011011011101111;
assign LUT_2[8651] = 32'b11111111111111111000010100001000;
assign LUT_2[8652] = 32'b11111111111111110001000000011011;
assign LUT_2[8653] = 32'b11111111111111101101111000110100;
assign LUT_2[8654] = 32'b11111111111111110111111001010111;
assign LUT_2[8655] = 32'b11111111111111110100110001110000;
assign LUT_2[8656] = 32'b11111111111111110100010101100000;
assign LUT_2[8657] = 32'b11111111111111110001001101111001;
assign LUT_2[8658] = 32'b11111111111111111011001110011100;
assign LUT_2[8659] = 32'b11111111111111111000000110110101;
assign LUT_2[8660] = 32'b11111111111111110000110011001000;
assign LUT_2[8661] = 32'b11111111111111101101101011100001;
assign LUT_2[8662] = 32'b11111111111111110111101100000100;
assign LUT_2[8663] = 32'b11111111111111110100100100011101;
assign LUT_2[8664] = 32'b11111111111111101111000110111101;
assign LUT_2[8665] = 32'b11111111111111101011111111010110;
assign LUT_2[8666] = 32'b11111111111111110101111111111001;
assign LUT_2[8667] = 32'b11111111111111110010111000010010;
assign LUT_2[8668] = 32'b11111111111111101011100100100101;
assign LUT_2[8669] = 32'b11111111111111101000011100111110;
assign LUT_2[8670] = 32'b11111111111111110010011101100001;
assign LUT_2[8671] = 32'b11111111111111101111010101111010;
assign LUT_2[8672] = 32'b11111111111111111010001100111111;
assign LUT_2[8673] = 32'b11111111111111110111000101011000;
assign LUT_2[8674] = 32'b00000000000000000001000101111011;
assign LUT_2[8675] = 32'b11111111111111111101111110010100;
assign LUT_2[8676] = 32'b11111111111111110110101010100111;
assign LUT_2[8677] = 32'b11111111111111110011100011000000;
assign LUT_2[8678] = 32'b11111111111111111101100011100011;
assign LUT_2[8679] = 32'b11111111111111111010011011111100;
assign LUT_2[8680] = 32'b11111111111111110100111110011100;
assign LUT_2[8681] = 32'b11111111111111110001110110110101;
assign LUT_2[8682] = 32'b11111111111111111011110111011000;
assign LUT_2[8683] = 32'b11111111111111111000101111110001;
assign LUT_2[8684] = 32'b11111111111111110001011100000100;
assign LUT_2[8685] = 32'b11111111111111101110010100011101;
assign LUT_2[8686] = 32'b11111111111111111000010101000000;
assign LUT_2[8687] = 32'b11111111111111110101001101011001;
assign LUT_2[8688] = 32'b11111111111111110100110001001001;
assign LUT_2[8689] = 32'b11111111111111110001101001100010;
assign LUT_2[8690] = 32'b11111111111111111011101010000101;
assign LUT_2[8691] = 32'b11111111111111111000100010011110;
assign LUT_2[8692] = 32'b11111111111111110001001110110001;
assign LUT_2[8693] = 32'b11111111111111101110000111001010;
assign LUT_2[8694] = 32'b11111111111111111000000111101101;
assign LUT_2[8695] = 32'b11111111111111110101000000000110;
assign LUT_2[8696] = 32'b11111111111111101111100010100110;
assign LUT_2[8697] = 32'b11111111111111101100011010111111;
assign LUT_2[8698] = 32'b11111111111111110110011011100010;
assign LUT_2[8699] = 32'b11111111111111110011010011111011;
assign LUT_2[8700] = 32'b11111111111111101100000000001110;
assign LUT_2[8701] = 32'b11111111111111101000111000100111;
assign LUT_2[8702] = 32'b11111111111111110010111001001010;
assign LUT_2[8703] = 32'b11111111111111101111110001100011;
assign LUT_2[8704] = 32'b11111111111111111110000111110000;
assign LUT_2[8705] = 32'b11111111111111111011000000001001;
assign LUT_2[8706] = 32'b00000000000000000101000000101100;
assign LUT_2[8707] = 32'b00000000000000000001111001000101;
assign LUT_2[8708] = 32'b11111111111111111010100101011000;
assign LUT_2[8709] = 32'b11111111111111110111011101110001;
assign LUT_2[8710] = 32'b00000000000000000001011110010100;
assign LUT_2[8711] = 32'b11111111111111111110010110101101;
assign LUT_2[8712] = 32'b11111111111111111000111001001101;
assign LUT_2[8713] = 32'b11111111111111110101110001100110;
assign LUT_2[8714] = 32'b11111111111111111111110010001001;
assign LUT_2[8715] = 32'b11111111111111111100101010100010;
assign LUT_2[8716] = 32'b11111111111111110101010110110101;
assign LUT_2[8717] = 32'b11111111111111110010001111001110;
assign LUT_2[8718] = 32'b11111111111111111100001111110001;
assign LUT_2[8719] = 32'b11111111111111111001001000001010;
assign LUT_2[8720] = 32'b11111111111111111000101011111010;
assign LUT_2[8721] = 32'b11111111111111110101100100010011;
assign LUT_2[8722] = 32'b11111111111111111111100100110110;
assign LUT_2[8723] = 32'b11111111111111111100011101001111;
assign LUT_2[8724] = 32'b11111111111111110101001001100010;
assign LUT_2[8725] = 32'b11111111111111110010000001111011;
assign LUT_2[8726] = 32'b11111111111111111100000010011110;
assign LUT_2[8727] = 32'b11111111111111111000111010110111;
assign LUT_2[8728] = 32'b11111111111111110011011101010111;
assign LUT_2[8729] = 32'b11111111111111110000010101110000;
assign LUT_2[8730] = 32'b11111111111111111010010110010011;
assign LUT_2[8731] = 32'b11111111111111110111001110101100;
assign LUT_2[8732] = 32'b11111111111111101111111010111111;
assign LUT_2[8733] = 32'b11111111111111101100110011011000;
assign LUT_2[8734] = 32'b11111111111111110110110011111011;
assign LUT_2[8735] = 32'b11111111111111110011101100010100;
assign LUT_2[8736] = 32'b11111111111111111110100011011001;
assign LUT_2[8737] = 32'b11111111111111111011011011110010;
assign LUT_2[8738] = 32'b00000000000000000101011100010101;
assign LUT_2[8739] = 32'b00000000000000000010010100101110;
assign LUT_2[8740] = 32'b11111111111111111011000001000001;
assign LUT_2[8741] = 32'b11111111111111110111111001011010;
assign LUT_2[8742] = 32'b00000000000000000001111001111101;
assign LUT_2[8743] = 32'b11111111111111111110110010010110;
assign LUT_2[8744] = 32'b11111111111111111001010100110110;
assign LUT_2[8745] = 32'b11111111111111110110001101001111;
assign LUT_2[8746] = 32'b00000000000000000000001101110010;
assign LUT_2[8747] = 32'b11111111111111111101000110001011;
assign LUT_2[8748] = 32'b11111111111111110101110010011110;
assign LUT_2[8749] = 32'b11111111111111110010101010110111;
assign LUT_2[8750] = 32'b11111111111111111100101011011010;
assign LUT_2[8751] = 32'b11111111111111111001100011110011;
assign LUT_2[8752] = 32'b11111111111111111001000111100011;
assign LUT_2[8753] = 32'b11111111111111110101111111111100;
assign LUT_2[8754] = 32'b00000000000000000000000000011111;
assign LUT_2[8755] = 32'b11111111111111111100111000111000;
assign LUT_2[8756] = 32'b11111111111111110101100101001011;
assign LUT_2[8757] = 32'b11111111111111110010011101100100;
assign LUT_2[8758] = 32'b11111111111111111100011110000111;
assign LUT_2[8759] = 32'b11111111111111111001010110100000;
assign LUT_2[8760] = 32'b11111111111111110011111001000000;
assign LUT_2[8761] = 32'b11111111111111110000110001011001;
assign LUT_2[8762] = 32'b11111111111111111010110001111100;
assign LUT_2[8763] = 32'b11111111111111110111101010010101;
assign LUT_2[8764] = 32'b11111111111111110000010110101000;
assign LUT_2[8765] = 32'b11111111111111101101001111000001;
assign LUT_2[8766] = 32'b11111111111111110111001111100100;
assign LUT_2[8767] = 32'b11111111111111110100000111111101;
assign LUT_2[8768] = 32'b11111111111111110110010000010011;
assign LUT_2[8769] = 32'b11111111111111110011001000101100;
assign LUT_2[8770] = 32'b11111111111111111101001001001111;
assign LUT_2[8771] = 32'b11111111111111111010000001101000;
assign LUT_2[8772] = 32'b11111111111111110010101101111011;
assign LUT_2[8773] = 32'b11111111111111101111100110010100;
assign LUT_2[8774] = 32'b11111111111111111001100110110111;
assign LUT_2[8775] = 32'b11111111111111110110011111010000;
assign LUT_2[8776] = 32'b11111111111111110001000001110000;
assign LUT_2[8777] = 32'b11111111111111101101111010001001;
assign LUT_2[8778] = 32'b11111111111111110111111010101100;
assign LUT_2[8779] = 32'b11111111111111110100110011000101;
assign LUT_2[8780] = 32'b11111111111111101101011111011000;
assign LUT_2[8781] = 32'b11111111111111101010010111110001;
assign LUT_2[8782] = 32'b11111111111111110100011000010100;
assign LUT_2[8783] = 32'b11111111111111110001010000101101;
assign LUT_2[8784] = 32'b11111111111111110000110100011101;
assign LUT_2[8785] = 32'b11111111111111101101101100110110;
assign LUT_2[8786] = 32'b11111111111111110111101101011001;
assign LUT_2[8787] = 32'b11111111111111110100100101110010;
assign LUT_2[8788] = 32'b11111111111111101101010010000101;
assign LUT_2[8789] = 32'b11111111111111101010001010011110;
assign LUT_2[8790] = 32'b11111111111111110100001011000001;
assign LUT_2[8791] = 32'b11111111111111110001000011011010;
assign LUT_2[8792] = 32'b11111111111111101011100101111010;
assign LUT_2[8793] = 32'b11111111111111101000011110010011;
assign LUT_2[8794] = 32'b11111111111111110010011110110110;
assign LUT_2[8795] = 32'b11111111111111101111010111001111;
assign LUT_2[8796] = 32'b11111111111111101000000011100010;
assign LUT_2[8797] = 32'b11111111111111100100111011111011;
assign LUT_2[8798] = 32'b11111111111111101110111100011110;
assign LUT_2[8799] = 32'b11111111111111101011110100110111;
assign LUT_2[8800] = 32'b11111111111111110110101011111100;
assign LUT_2[8801] = 32'b11111111111111110011100100010101;
assign LUT_2[8802] = 32'b11111111111111111101100100111000;
assign LUT_2[8803] = 32'b11111111111111111010011101010001;
assign LUT_2[8804] = 32'b11111111111111110011001001100100;
assign LUT_2[8805] = 32'b11111111111111110000000001111101;
assign LUT_2[8806] = 32'b11111111111111111010000010100000;
assign LUT_2[8807] = 32'b11111111111111110110111010111001;
assign LUT_2[8808] = 32'b11111111111111110001011101011001;
assign LUT_2[8809] = 32'b11111111111111101110010101110010;
assign LUT_2[8810] = 32'b11111111111111111000010110010101;
assign LUT_2[8811] = 32'b11111111111111110101001110101110;
assign LUT_2[8812] = 32'b11111111111111101101111011000001;
assign LUT_2[8813] = 32'b11111111111111101010110011011010;
assign LUT_2[8814] = 32'b11111111111111110100110011111101;
assign LUT_2[8815] = 32'b11111111111111110001101100010110;
assign LUT_2[8816] = 32'b11111111111111110001010000000110;
assign LUT_2[8817] = 32'b11111111111111101110001000011111;
assign LUT_2[8818] = 32'b11111111111111111000001001000010;
assign LUT_2[8819] = 32'b11111111111111110101000001011011;
assign LUT_2[8820] = 32'b11111111111111101101101101101110;
assign LUT_2[8821] = 32'b11111111111111101010100110000111;
assign LUT_2[8822] = 32'b11111111111111110100100110101010;
assign LUT_2[8823] = 32'b11111111111111110001011111000011;
assign LUT_2[8824] = 32'b11111111111111101100000001100011;
assign LUT_2[8825] = 32'b11111111111111101000111001111100;
assign LUT_2[8826] = 32'b11111111111111110010111010011111;
assign LUT_2[8827] = 32'b11111111111111101111110010111000;
assign LUT_2[8828] = 32'b11111111111111101000011111001011;
assign LUT_2[8829] = 32'b11111111111111100101010111100100;
assign LUT_2[8830] = 32'b11111111111111101111011000000111;
assign LUT_2[8831] = 32'b11111111111111101100010000100000;
assign LUT_2[8832] = 32'b00000000000000000010011011111111;
assign LUT_2[8833] = 32'b11111111111111111111010100011000;
assign LUT_2[8834] = 32'b00000000000000001001010100111011;
assign LUT_2[8835] = 32'b00000000000000000110001101010100;
assign LUT_2[8836] = 32'b11111111111111111110111001100111;
assign LUT_2[8837] = 32'b11111111111111111011110010000000;
assign LUT_2[8838] = 32'b00000000000000000101110010100011;
assign LUT_2[8839] = 32'b00000000000000000010101010111100;
assign LUT_2[8840] = 32'b11111111111111111101001101011100;
assign LUT_2[8841] = 32'b11111111111111111010000101110101;
assign LUT_2[8842] = 32'b00000000000000000100000110011000;
assign LUT_2[8843] = 32'b00000000000000000000111110110001;
assign LUT_2[8844] = 32'b11111111111111111001101011000100;
assign LUT_2[8845] = 32'b11111111111111110110100011011101;
assign LUT_2[8846] = 32'b00000000000000000000100100000000;
assign LUT_2[8847] = 32'b11111111111111111101011100011001;
assign LUT_2[8848] = 32'b11111111111111111101000000001001;
assign LUT_2[8849] = 32'b11111111111111111001111000100010;
assign LUT_2[8850] = 32'b00000000000000000011111001000101;
assign LUT_2[8851] = 32'b00000000000000000000110001011110;
assign LUT_2[8852] = 32'b11111111111111111001011101110001;
assign LUT_2[8853] = 32'b11111111111111110110010110001010;
assign LUT_2[8854] = 32'b00000000000000000000010110101101;
assign LUT_2[8855] = 32'b11111111111111111101001111000110;
assign LUT_2[8856] = 32'b11111111111111110111110001100110;
assign LUT_2[8857] = 32'b11111111111111110100101001111111;
assign LUT_2[8858] = 32'b11111111111111111110101010100010;
assign LUT_2[8859] = 32'b11111111111111111011100010111011;
assign LUT_2[8860] = 32'b11111111111111110100001111001110;
assign LUT_2[8861] = 32'b11111111111111110001000111100111;
assign LUT_2[8862] = 32'b11111111111111111011001000001010;
assign LUT_2[8863] = 32'b11111111111111111000000000100011;
assign LUT_2[8864] = 32'b00000000000000000010110111101000;
assign LUT_2[8865] = 32'b11111111111111111111110000000001;
assign LUT_2[8866] = 32'b00000000000000001001110000100100;
assign LUT_2[8867] = 32'b00000000000000000110101000111101;
assign LUT_2[8868] = 32'b11111111111111111111010101010000;
assign LUT_2[8869] = 32'b11111111111111111100001101101001;
assign LUT_2[8870] = 32'b00000000000000000110001110001100;
assign LUT_2[8871] = 32'b00000000000000000011000110100101;
assign LUT_2[8872] = 32'b11111111111111111101101001000101;
assign LUT_2[8873] = 32'b11111111111111111010100001011110;
assign LUT_2[8874] = 32'b00000000000000000100100010000001;
assign LUT_2[8875] = 32'b00000000000000000001011010011010;
assign LUT_2[8876] = 32'b11111111111111111010000110101101;
assign LUT_2[8877] = 32'b11111111111111110110111111000110;
assign LUT_2[8878] = 32'b00000000000000000000111111101001;
assign LUT_2[8879] = 32'b11111111111111111101111000000010;
assign LUT_2[8880] = 32'b11111111111111111101011011110010;
assign LUT_2[8881] = 32'b11111111111111111010010100001011;
assign LUT_2[8882] = 32'b00000000000000000100010100101110;
assign LUT_2[8883] = 32'b00000000000000000001001101000111;
assign LUT_2[8884] = 32'b11111111111111111001111001011010;
assign LUT_2[8885] = 32'b11111111111111110110110001110011;
assign LUT_2[8886] = 32'b00000000000000000000110010010110;
assign LUT_2[8887] = 32'b11111111111111111101101010101111;
assign LUT_2[8888] = 32'b11111111111111111000001101001111;
assign LUT_2[8889] = 32'b11111111111111110101000101101000;
assign LUT_2[8890] = 32'b11111111111111111111000110001011;
assign LUT_2[8891] = 32'b11111111111111111011111110100100;
assign LUT_2[8892] = 32'b11111111111111110100101010110111;
assign LUT_2[8893] = 32'b11111111111111110001100011010000;
assign LUT_2[8894] = 32'b11111111111111111011100011110011;
assign LUT_2[8895] = 32'b11111111111111111000011100001100;
assign LUT_2[8896] = 32'b11111111111111111010100100100010;
assign LUT_2[8897] = 32'b11111111111111110111011100111011;
assign LUT_2[8898] = 32'b00000000000000000001011101011110;
assign LUT_2[8899] = 32'b11111111111111111110010101110111;
assign LUT_2[8900] = 32'b11111111111111110111000010001010;
assign LUT_2[8901] = 32'b11111111111111110011111010100011;
assign LUT_2[8902] = 32'b11111111111111111101111011000110;
assign LUT_2[8903] = 32'b11111111111111111010110011011111;
assign LUT_2[8904] = 32'b11111111111111110101010101111111;
assign LUT_2[8905] = 32'b11111111111111110010001110011000;
assign LUT_2[8906] = 32'b11111111111111111100001110111011;
assign LUT_2[8907] = 32'b11111111111111111001000111010100;
assign LUT_2[8908] = 32'b11111111111111110001110011100111;
assign LUT_2[8909] = 32'b11111111111111101110101100000000;
assign LUT_2[8910] = 32'b11111111111111111000101100100011;
assign LUT_2[8911] = 32'b11111111111111110101100100111100;
assign LUT_2[8912] = 32'b11111111111111110101001000101100;
assign LUT_2[8913] = 32'b11111111111111110010000001000101;
assign LUT_2[8914] = 32'b11111111111111111100000001101000;
assign LUT_2[8915] = 32'b11111111111111111000111010000001;
assign LUT_2[8916] = 32'b11111111111111110001100110010100;
assign LUT_2[8917] = 32'b11111111111111101110011110101101;
assign LUT_2[8918] = 32'b11111111111111111000011111010000;
assign LUT_2[8919] = 32'b11111111111111110101010111101001;
assign LUT_2[8920] = 32'b11111111111111101111111010001001;
assign LUT_2[8921] = 32'b11111111111111101100110010100010;
assign LUT_2[8922] = 32'b11111111111111110110110011000101;
assign LUT_2[8923] = 32'b11111111111111110011101011011110;
assign LUT_2[8924] = 32'b11111111111111101100010111110001;
assign LUT_2[8925] = 32'b11111111111111101001010000001010;
assign LUT_2[8926] = 32'b11111111111111110011010000101101;
assign LUT_2[8927] = 32'b11111111111111110000001001000110;
assign LUT_2[8928] = 32'b11111111111111111011000000001011;
assign LUT_2[8929] = 32'b11111111111111110111111000100100;
assign LUT_2[8930] = 32'b00000000000000000001111001000111;
assign LUT_2[8931] = 32'b11111111111111111110110001100000;
assign LUT_2[8932] = 32'b11111111111111110111011101110011;
assign LUT_2[8933] = 32'b11111111111111110100010110001100;
assign LUT_2[8934] = 32'b11111111111111111110010110101111;
assign LUT_2[8935] = 32'b11111111111111111011001111001000;
assign LUT_2[8936] = 32'b11111111111111110101110001101000;
assign LUT_2[8937] = 32'b11111111111111110010101010000001;
assign LUT_2[8938] = 32'b11111111111111111100101010100100;
assign LUT_2[8939] = 32'b11111111111111111001100010111101;
assign LUT_2[8940] = 32'b11111111111111110010001111010000;
assign LUT_2[8941] = 32'b11111111111111101111000111101001;
assign LUT_2[8942] = 32'b11111111111111111001001000001100;
assign LUT_2[8943] = 32'b11111111111111110110000000100101;
assign LUT_2[8944] = 32'b11111111111111110101100100010101;
assign LUT_2[8945] = 32'b11111111111111110010011100101110;
assign LUT_2[8946] = 32'b11111111111111111100011101010001;
assign LUT_2[8947] = 32'b11111111111111111001010101101010;
assign LUT_2[8948] = 32'b11111111111111110010000001111101;
assign LUT_2[8949] = 32'b11111111111111101110111010010110;
assign LUT_2[8950] = 32'b11111111111111111000111010111001;
assign LUT_2[8951] = 32'b11111111111111110101110011010010;
assign LUT_2[8952] = 32'b11111111111111110000010101110010;
assign LUT_2[8953] = 32'b11111111111111101101001110001011;
assign LUT_2[8954] = 32'b11111111111111110111001110101110;
assign LUT_2[8955] = 32'b11111111111111110100000111000111;
assign LUT_2[8956] = 32'b11111111111111101100110011011010;
assign LUT_2[8957] = 32'b11111111111111101001101011110011;
assign LUT_2[8958] = 32'b11111111111111110011101100010110;
assign LUT_2[8959] = 32'b11111111111111110000100100101111;
assign LUT_2[8960] = 32'b00000000000000000010000110010110;
assign LUT_2[8961] = 32'b11111111111111111110111110101111;
assign LUT_2[8962] = 32'b00000000000000001000111111010010;
assign LUT_2[8963] = 32'b00000000000000000101110111101011;
assign LUT_2[8964] = 32'b11111111111111111110100011111110;
assign LUT_2[8965] = 32'b11111111111111111011011100010111;
assign LUT_2[8966] = 32'b00000000000000000101011100111010;
assign LUT_2[8967] = 32'b00000000000000000010010101010011;
assign LUT_2[8968] = 32'b11111111111111111100110111110011;
assign LUT_2[8969] = 32'b11111111111111111001110000001100;
assign LUT_2[8970] = 32'b00000000000000000011110000101111;
assign LUT_2[8971] = 32'b00000000000000000000101001001000;
assign LUT_2[8972] = 32'b11111111111111111001010101011011;
assign LUT_2[8973] = 32'b11111111111111110110001101110100;
assign LUT_2[8974] = 32'b00000000000000000000001110010111;
assign LUT_2[8975] = 32'b11111111111111111101000110110000;
assign LUT_2[8976] = 32'b11111111111111111100101010100000;
assign LUT_2[8977] = 32'b11111111111111111001100010111001;
assign LUT_2[8978] = 32'b00000000000000000011100011011100;
assign LUT_2[8979] = 32'b00000000000000000000011011110101;
assign LUT_2[8980] = 32'b11111111111111111001001000001000;
assign LUT_2[8981] = 32'b11111111111111110110000000100001;
assign LUT_2[8982] = 32'b00000000000000000000000001000100;
assign LUT_2[8983] = 32'b11111111111111111100111001011101;
assign LUT_2[8984] = 32'b11111111111111110111011011111101;
assign LUT_2[8985] = 32'b11111111111111110100010100010110;
assign LUT_2[8986] = 32'b11111111111111111110010100111001;
assign LUT_2[8987] = 32'b11111111111111111011001101010010;
assign LUT_2[8988] = 32'b11111111111111110011111001100101;
assign LUT_2[8989] = 32'b11111111111111110000110001111110;
assign LUT_2[8990] = 32'b11111111111111111010110010100001;
assign LUT_2[8991] = 32'b11111111111111110111101010111010;
assign LUT_2[8992] = 32'b00000000000000000010100001111111;
assign LUT_2[8993] = 32'b11111111111111111111011010011000;
assign LUT_2[8994] = 32'b00000000000000001001011010111011;
assign LUT_2[8995] = 32'b00000000000000000110010011010100;
assign LUT_2[8996] = 32'b11111111111111111110111111100111;
assign LUT_2[8997] = 32'b11111111111111111011111000000000;
assign LUT_2[8998] = 32'b00000000000000000101111000100011;
assign LUT_2[8999] = 32'b00000000000000000010110000111100;
assign LUT_2[9000] = 32'b11111111111111111101010011011100;
assign LUT_2[9001] = 32'b11111111111111111010001011110101;
assign LUT_2[9002] = 32'b00000000000000000100001100011000;
assign LUT_2[9003] = 32'b00000000000000000001000100110001;
assign LUT_2[9004] = 32'b11111111111111111001110001000100;
assign LUT_2[9005] = 32'b11111111111111110110101001011101;
assign LUT_2[9006] = 32'b00000000000000000000101010000000;
assign LUT_2[9007] = 32'b11111111111111111101100010011001;
assign LUT_2[9008] = 32'b11111111111111111101000110001001;
assign LUT_2[9009] = 32'b11111111111111111001111110100010;
assign LUT_2[9010] = 32'b00000000000000000011111111000101;
assign LUT_2[9011] = 32'b00000000000000000000110111011110;
assign LUT_2[9012] = 32'b11111111111111111001100011110001;
assign LUT_2[9013] = 32'b11111111111111110110011100001010;
assign LUT_2[9014] = 32'b00000000000000000000011100101101;
assign LUT_2[9015] = 32'b11111111111111111101010101000110;
assign LUT_2[9016] = 32'b11111111111111110111110111100110;
assign LUT_2[9017] = 32'b11111111111111110100101111111111;
assign LUT_2[9018] = 32'b11111111111111111110110000100010;
assign LUT_2[9019] = 32'b11111111111111111011101000111011;
assign LUT_2[9020] = 32'b11111111111111110100010101001110;
assign LUT_2[9021] = 32'b11111111111111110001001101100111;
assign LUT_2[9022] = 32'b11111111111111111011001110001010;
assign LUT_2[9023] = 32'b11111111111111111000000110100011;
assign LUT_2[9024] = 32'b11111111111111111010001110111001;
assign LUT_2[9025] = 32'b11111111111111110111000111010010;
assign LUT_2[9026] = 32'b00000000000000000001000111110101;
assign LUT_2[9027] = 32'b11111111111111111110000000001110;
assign LUT_2[9028] = 32'b11111111111111110110101100100001;
assign LUT_2[9029] = 32'b11111111111111110011100100111010;
assign LUT_2[9030] = 32'b11111111111111111101100101011101;
assign LUT_2[9031] = 32'b11111111111111111010011101110110;
assign LUT_2[9032] = 32'b11111111111111110101000000010110;
assign LUT_2[9033] = 32'b11111111111111110001111000101111;
assign LUT_2[9034] = 32'b11111111111111111011111001010010;
assign LUT_2[9035] = 32'b11111111111111111000110001101011;
assign LUT_2[9036] = 32'b11111111111111110001011101111110;
assign LUT_2[9037] = 32'b11111111111111101110010110010111;
assign LUT_2[9038] = 32'b11111111111111111000010110111010;
assign LUT_2[9039] = 32'b11111111111111110101001111010011;
assign LUT_2[9040] = 32'b11111111111111110100110011000011;
assign LUT_2[9041] = 32'b11111111111111110001101011011100;
assign LUT_2[9042] = 32'b11111111111111111011101011111111;
assign LUT_2[9043] = 32'b11111111111111111000100100011000;
assign LUT_2[9044] = 32'b11111111111111110001010000101011;
assign LUT_2[9045] = 32'b11111111111111101110001001000100;
assign LUT_2[9046] = 32'b11111111111111111000001001100111;
assign LUT_2[9047] = 32'b11111111111111110101000010000000;
assign LUT_2[9048] = 32'b11111111111111101111100100100000;
assign LUT_2[9049] = 32'b11111111111111101100011100111001;
assign LUT_2[9050] = 32'b11111111111111110110011101011100;
assign LUT_2[9051] = 32'b11111111111111110011010101110101;
assign LUT_2[9052] = 32'b11111111111111101100000010001000;
assign LUT_2[9053] = 32'b11111111111111101000111010100001;
assign LUT_2[9054] = 32'b11111111111111110010111011000100;
assign LUT_2[9055] = 32'b11111111111111101111110011011101;
assign LUT_2[9056] = 32'b11111111111111111010101010100010;
assign LUT_2[9057] = 32'b11111111111111110111100010111011;
assign LUT_2[9058] = 32'b00000000000000000001100011011110;
assign LUT_2[9059] = 32'b11111111111111111110011011110111;
assign LUT_2[9060] = 32'b11111111111111110111001000001010;
assign LUT_2[9061] = 32'b11111111111111110100000000100011;
assign LUT_2[9062] = 32'b11111111111111111110000001000110;
assign LUT_2[9063] = 32'b11111111111111111010111001011111;
assign LUT_2[9064] = 32'b11111111111111110101011011111111;
assign LUT_2[9065] = 32'b11111111111111110010010100011000;
assign LUT_2[9066] = 32'b11111111111111111100010100111011;
assign LUT_2[9067] = 32'b11111111111111111001001101010100;
assign LUT_2[9068] = 32'b11111111111111110001111001100111;
assign LUT_2[9069] = 32'b11111111111111101110110010000000;
assign LUT_2[9070] = 32'b11111111111111111000110010100011;
assign LUT_2[9071] = 32'b11111111111111110101101010111100;
assign LUT_2[9072] = 32'b11111111111111110101001110101100;
assign LUT_2[9073] = 32'b11111111111111110010000111000101;
assign LUT_2[9074] = 32'b11111111111111111100000111101000;
assign LUT_2[9075] = 32'b11111111111111111001000000000001;
assign LUT_2[9076] = 32'b11111111111111110001101100010100;
assign LUT_2[9077] = 32'b11111111111111101110100100101101;
assign LUT_2[9078] = 32'b11111111111111111000100101010000;
assign LUT_2[9079] = 32'b11111111111111110101011101101001;
assign LUT_2[9080] = 32'b11111111111111110000000000001001;
assign LUT_2[9081] = 32'b11111111111111101100111000100010;
assign LUT_2[9082] = 32'b11111111111111110110111001000101;
assign LUT_2[9083] = 32'b11111111111111110011110001011110;
assign LUT_2[9084] = 32'b11111111111111101100011101110001;
assign LUT_2[9085] = 32'b11111111111111101001010110001010;
assign LUT_2[9086] = 32'b11111111111111110011010110101101;
assign LUT_2[9087] = 32'b11111111111111110000001111000110;
assign LUT_2[9088] = 32'b00000000000000000110011010100101;
assign LUT_2[9089] = 32'b00000000000000000011010010111110;
assign LUT_2[9090] = 32'b00000000000000001101010011100001;
assign LUT_2[9091] = 32'b00000000000000001010001011111010;
assign LUT_2[9092] = 32'b00000000000000000010111000001101;
assign LUT_2[9093] = 32'b11111111111111111111110000100110;
assign LUT_2[9094] = 32'b00000000000000001001110001001001;
assign LUT_2[9095] = 32'b00000000000000000110101001100010;
assign LUT_2[9096] = 32'b00000000000000000001001100000010;
assign LUT_2[9097] = 32'b11111111111111111110000100011011;
assign LUT_2[9098] = 32'b00000000000000001000000100111110;
assign LUT_2[9099] = 32'b00000000000000000100111101010111;
assign LUT_2[9100] = 32'b11111111111111111101101001101010;
assign LUT_2[9101] = 32'b11111111111111111010100010000011;
assign LUT_2[9102] = 32'b00000000000000000100100010100110;
assign LUT_2[9103] = 32'b00000000000000000001011010111111;
assign LUT_2[9104] = 32'b00000000000000000000111110101111;
assign LUT_2[9105] = 32'b11111111111111111101110111001000;
assign LUT_2[9106] = 32'b00000000000000000111110111101011;
assign LUT_2[9107] = 32'b00000000000000000100110000000100;
assign LUT_2[9108] = 32'b11111111111111111101011100010111;
assign LUT_2[9109] = 32'b11111111111111111010010100110000;
assign LUT_2[9110] = 32'b00000000000000000100010101010011;
assign LUT_2[9111] = 32'b00000000000000000001001101101100;
assign LUT_2[9112] = 32'b11111111111111111011110000001100;
assign LUT_2[9113] = 32'b11111111111111111000101000100101;
assign LUT_2[9114] = 32'b00000000000000000010101001001000;
assign LUT_2[9115] = 32'b11111111111111111111100001100001;
assign LUT_2[9116] = 32'b11111111111111111000001101110100;
assign LUT_2[9117] = 32'b11111111111111110101000110001101;
assign LUT_2[9118] = 32'b11111111111111111111000110110000;
assign LUT_2[9119] = 32'b11111111111111111011111111001001;
assign LUT_2[9120] = 32'b00000000000000000110110110001110;
assign LUT_2[9121] = 32'b00000000000000000011101110100111;
assign LUT_2[9122] = 32'b00000000000000001101101111001010;
assign LUT_2[9123] = 32'b00000000000000001010100111100011;
assign LUT_2[9124] = 32'b00000000000000000011010011110110;
assign LUT_2[9125] = 32'b00000000000000000000001100001111;
assign LUT_2[9126] = 32'b00000000000000001010001100110010;
assign LUT_2[9127] = 32'b00000000000000000111000101001011;
assign LUT_2[9128] = 32'b00000000000000000001100111101011;
assign LUT_2[9129] = 32'b11111111111111111110100000000100;
assign LUT_2[9130] = 32'b00000000000000001000100000100111;
assign LUT_2[9131] = 32'b00000000000000000101011001000000;
assign LUT_2[9132] = 32'b11111111111111111110000101010011;
assign LUT_2[9133] = 32'b11111111111111111010111101101100;
assign LUT_2[9134] = 32'b00000000000000000100111110001111;
assign LUT_2[9135] = 32'b00000000000000000001110110101000;
assign LUT_2[9136] = 32'b00000000000000000001011010011000;
assign LUT_2[9137] = 32'b11111111111111111110010010110001;
assign LUT_2[9138] = 32'b00000000000000001000010011010100;
assign LUT_2[9139] = 32'b00000000000000000101001011101101;
assign LUT_2[9140] = 32'b11111111111111111101111000000000;
assign LUT_2[9141] = 32'b11111111111111111010110000011001;
assign LUT_2[9142] = 32'b00000000000000000100110000111100;
assign LUT_2[9143] = 32'b00000000000000000001101001010101;
assign LUT_2[9144] = 32'b11111111111111111100001011110101;
assign LUT_2[9145] = 32'b11111111111111111001000100001110;
assign LUT_2[9146] = 32'b00000000000000000011000100110001;
assign LUT_2[9147] = 32'b11111111111111111111111101001010;
assign LUT_2[9148] = 32'b11111111111111111000101001011101;
assign LUT_2[9149] = 32'b11111111111111110101100001110110;
assign LUT_2[9150] = 32'b11111111111111111111100010011001;
assign LUT_2[9151] = 32'b11111111111111111100011010110010;
assign LUT_2[9152] = 32'b11111111111111111110100011001000;
assign LUT_2[9153] = 32'b11111111111111111011011011100001;
assign LUT_2[9154] = 32'b00000000000000000101011100000100;
assign LUT_2[9155] = 32'b00000000000000000010010100011101;
assign LUT_2[9156] = 32'b11111111111111111011000000110000;
assign LUT_2[9157] = 32'b11111111111111110111111001001001;
assign LUT_2[9158] = 32'b00000000000000000001111001101100;
assign LUT_2[9159] = 32'b11111111111111111110110010000101;
assign LUT_2[9160] = 32'b11111111111111111001010100100101;
assign LUT_2[9161] = 32'b11111111111111110110001100111110;
assign LUT_2[9162] = 32'b00000000000000000000001101100001;
assign LUT_2[9163] = 32'b11111111111111111101000101111010;
assign LUT_2[9164] = 32'b11111111111111110101110010001101;
assign LUT_2[9165] = 32'b11111111111111110010101010100110;
assign LUT_2[9166] = 32'b11111111111111111100101011001001;
assign LUT_2[9167] = 32'b11111111111111111001100011100010;
assign LUT_2[9168] = 32'b11111111111111111001000111010010;
assign LUT_2[9169] = 32'b11111111111111110101111111101011;
assign LUT_2[9170] = 32'b00000000000000000000000000001110;
assign LUT_2[9171] = 32'b11111111111111111100111000100111;
assign LUT_2[9172] = 32'b11111111111111110101100100111010;
assign LUT_2[9173] = 32'b11111111111111110010011101010011;
assign LUT_2[9174] = 32'b11111111111111111100011101110110;
assign LUT_2[9175] = 32'b11111111111111111001010110001111;
assign LUT_2[9176] = 32'b11111111111111110011111000101111;
assign LUT_2[9177] = 32'b11111111111111110000110001001000;
assign LUT_2[9178] = 32'b11111111111111111010110001101011;
assign LUT_2[9179] = 32'b11111111111111110111101010000100;
assign LUT_2[9180] = 32'b11111111111111110000010110010111;
assign LUT_2[9181] = 32'b11111111111111101101001110110000;
assign LUT_2[9182] = 32'b11111111111111110111001111010011;
assign LUT_2[9183] = 32'b11111111111111110100000111101100;
assign LUT_2[9184] = 32'b11111111111111111110111110110001;
assign LUT_2[9185] = 32'b11111111111111111011110111001010;
assign LUT_2[9186] = 32'b00000000000000000101110111101101;
assign LUT_2[9187] = 32'b00000000000000000010110000000110;
assign LUT_2[9188] = 32'b11111111111111111011011100011001;
assign LUT_2[9189] = 32'b11111111111111111000010100110010;
assign LUT_2[9190] = 32'b00000000000000000010010101010101;
assign LUT_2[9191] = 32'b11111111111111111111001101101110;
assign LUT_2[9192] = 32'b11111111111111111001110000001110;
assign LUT_2[9193] = 32'b11111111111111110110101000100111;
assign LUT_2[9194] = 32'b00000000000000000000101001001010;
assign LUT_2[9195] = 32'b11111111111111111101100001100011;
assign LUT_2[9196] = 32'b11111111111111110110001101110110;
assign LUT_2[9197] = 32'b11111111111111110011000110001111;
assign LUT_2[9198] = 32'b11111111111111111101000110110010;
assign LUT_2[9199] = 32'b11111111111111111001111111001011;
assign LUT_2[9200] = 32'b11111111111111111001100010111011;
assign LUT_2[9201] = 32'b11111111111111110110011011010100;
assign LUT_2[9202] = 32'b00000000000000000000011011110111;
assign LUT_2[9203] = 32'b11111111111111111101010100010000;
assign LUT_2[9204] = 32'b11111111111111110110000000100011;
assign LUT_2[9205] = 32'b11111111111111110010111000111100;
assign LUT_2[9206] = 32'b11111111111111111100111001011111;
assign LUT_2[9207] = 32'b11111111111111111001110001111000;
assign LUT_2[9208] = 32'b11111111111111110100010100011000;
assign LUT_2[9209] = 32'b11111111111111110001001100110001;
assign LUT_2[9210] = 32'b11111111111111111011001101010100;
assign LUT_2[9211] = 32'b11111111111111111000000101101101;
assign LUT_2[9212] = 32'b11111111111111110000110010000000;
assign LUT_2[9213] = 32'b11111111111111101101101010011001;
assign LUT_2[9214] = 32'b11111111111111110111101010111100;
assign LUT_2[9215] = 32'b11111111111111110100100011010101;
assign LUT_2[9216] = 32'b00000000000000000000000010000011;
assign LUT_2[9217] = 32'b11111111111111111100111010011100;
assign LUT_2[9218] = 32'b00000000000000000110111010111111;
assign LUT_2[9219] = 32'b00000000000000000011110011011000;
assign LUT_2[9220] = 32'b11111111111111111100011111101011;
assign LUT_2[9221] = 32'b11111111111111111001011000000100;
assign LUT_2[9222] = 32'b00000000000000000011011000100111;
assign LUT_2[9223] = 32'b00000000000000000000010001000000;
assign LUT_2[9224] = 32'b11111111111111111010110011100000;
assign LUT_2[9225] = 32'b11111111111111110111101011111001;
assign LUT_2[9226] = 32'b00000000000000000001101100011100;
assign LUT_2[9227] = 32'b11111111111111111110100100110101;
assign LUT_2[9228] = 32'b11111111111111110111010001001000;
assign LUT_2[9229] = 32'b11111111111111110100001001100001;
assign LUT_2[9230] = 32'b11111111111111111110001010000100;
assign LUT_2[9231] = 32'b11111111111111111011000010011101;
assign LUT_2[9232] = 32'b11111111111111111010100110001101;
assign LUT_2[9233] = 32'b11111111111111110111011110100110;
assign LUT_2[9234] = 32'b00000000000000000001011111001001;
assign LUT_2[9235] = 32'b11111111111111111110010111100010;
assign LUT_2[9236] = 32'b11111111111111110111000011110101;
assign LUT_2[9237] = 32'b11111111111111110011111100001110;
assign LUT_2[9238] = 32'b11111111111111111101111100110001;
assign LUT_2[9239] = 32'b11111111111111111010110101001010;
assign LUT_2[9240] = 32'b11111111111111110101010111101010;
assign LUT_2[9241] = 32'b11111111111111110010010000000011;
assign LUT_2[9242] = 32'b11111111111111111100010000100110;
assign LUT_2[9243] = 32'b11111111111111111001001000111111;
assign LUT_2[9244] = 32'b11111111111111110001110101010010;
assign LUT_2[9245] = 32'b11111111111111101110101101101011;
assign LUT_2[9246] = 32'b11111111111111111000101110001110;
assign LUT_2[9247] = 32'b11111111111111110101100110100111;
assign LUT_2[9248] = 32'b00000000000000000000011101101100;
assign LUT_2[9249] = 32'b11111111111111111101010110000101;
assign LUT_2[9250] = 32'b00000000000000000111010110101000;
assign LUT_2[9251] = 32'b00000000000000000100001111000001;
assign LUT_2[9252] = 32'b11111111111111111100111011010100;
assign LUT_2[9253] = 32'b11111111111111111001110011101101;
assign LUT_2[9254] = 32'b00000000000000000011110100010000;
assign LUT_2[9255] = 32'b00000000000000000000101100101001;
assign LUT_2[9256] = 32'b11111111111111111011001111001001;
assign LUT_2[9257] = 32'b11111111111111111000000111100010;
assign LUT_2[9258] = 32'b00000000000000000010001000000101;
assign LUT_2[9259] = 32'b11111111111111111111000000011110;
assign LUT_2[9260] = 32'b11111111111111110111101100110001;
assign LUT_2[9261] = 32'b11111111111111110100100101001010;
assign LUT_2[9262] = 32'b11111111111111111110100101101101;
assign LUT_2[9263] = 32'b11111111111111111011011110000110;
assign LUT_2[9264] = 32'b11111111111111111011000001110110;
assign LUT_2[9265] = 32'b11111111111111110111111010001111;
assign LUT_2[9266] = 32'b00000000000000000001111010110010;
assign LUT_2[9267] = 32'b11111111111111111110110011001011;
assign LUT_2[9268] = 32'b11111111111111110111011111011110;
assign LUT_2[9269] = 32'b11111111111111110100010111110111;
assign LUT_2[9270] = 32'b11111111111111111110011000011010;
assign LUT_2[9271] = 32'b11111111111111111011010000110011;
assign LUT_2[9272] = 32'b11111111111111110101110011010011;
assign LUT_2[9273] = 32'b11111111111111110010101011101100;
assign LUT_2[9274] = 32'b11111111111111111100101100001111;
assign LUT_2[9275] = 32'b11111111111111111001100100101000;
assign LUT_2[9276] = 32'b11111111111111110010010000111011;
assign LUT_2[9277] = 32'b11111111111111101111001001010100;
assign LUT_2[9278] = 32'b11111111111111111001001001110111;
assign LUT_2[9279] = 32'b11111111111111110110000010010000;
assign LUT_2[9280] = 32'b11111111111111111000001010100110;
assign LUT_2[9281] = 32'b11111111111111110101000010111111;
assign LUT_2[9282] = 32'b11111111111111111111000011100010;
assign LUT_2[9283] = 32'b11111111111111111011111011111011;
assign LUT_2[9284] = 32'b11111111111111110100101000001110;
assign LUT_2[9285] = 32'b11111111111111110001100000100111;
assign LUT_2[9286] = 32'b11111111111111111011100001001010;
assign LUT_2[9287] = 32'b11111111111111111000011001100011;
assign LUT_2[9288] = 32'b11111111111111110010111100000011;
assign LUT_2[9289] = 32'b11111111111111101111110100011100;
assign LUT_2[9290] = 32'b11111111111111111001110100111111;
assign LUT_2[9291] = 32'b11111111111111110110101101011000;
assign LUT_2[9292] = 32'b11111111111111101111011001101011;
assign LUT_2[9293] = 32'b11111111111111101100010010000100;
assign LUT_2[9294] = 32'b11111111111111110110010010100111;
assign LUT_2[9295] = 32'b11111111111111110011001011000000;
assign LUT_2[9296] = 32'b11111111111111110010101110110000;
assign LUT_2[9297] = 32'b11111111111111101111100111001001;
assign LUT_2[9298] = 32'b11111111111111111001100111101100;
assign LUT_2[9299] = 32'b11111111111111110110100000000101;
assign LUT_2[9300] = 32'b11111111111111101111001100011000;
assign LUT_2[9301] = 32'b11111111111111101100000100110001;
assign LUT_2[9302] = 32'b11111111111111110110000101010100;
assign LUT_2[9303] = 32'b11111111111111110010111101101101;
assign LUT_2[9304] = 32'b11111111111111101101100000001101;
assign LUT_2[9305] = 32'b11111111111111101010011000100110;
assign LUT_2[9306] = 32'b11111111111111110100011001001001;
assign LUT_2[9307] = 32'b11111111111111110001010001100010;
assign LUT_2[9308] = 32'b11111111111111101001111101110101;
assign LUT_2[9309] = 32'b11111111111111100110110110001110;
assign LUT_2[9310] = 32'b11111111111111110000110110110001;
assign LUT_2[9311] = 32'b11111111111111101101101111001010;
assign LUT_2[9312] = 32'b11111111111111111000100110001111;
assign LUT_2[9313] = 32'b11111111111111110101011110101000;
assign LUT_2[9314] = 32'b11111111111111111111011111001011;
assign LUT_2[9315] = 32'b11111111111111111100010111100100;
assign LUT_2[9316] = 32'b11111111111111110101000011110111;
assign LUT_2[9317] = 32'b11111111111111110001111100010000;
assign LUT_2[9318] = 32'b11111111111111111011111100110011;
assign LUT_2[9319] = 32'b11111111111111111000110101001100;
assign LUT_2[9320] = 32'b11111111111111110011010111101100;
assign LUT_2[9321] = 32'b11111111111111110000010000000101;
assign LUT_2[9322] = 32'b11111111111111111010010000101000;
assign LUT_2[9323] = 32'b11111111111111110111001001000001;
assign LUT_2[9324] = 32'b11111111111111101111110101010100;
assign LUT_2[9325] = 32'b11111111111111101100101101101101;
assign LUT_2[9326] = 32'b11111111111111110110101110010000;
assign LUT_2[9327] = 32'b11111111111111110011100110101001;
assign LUT_2[9328] = 32'b11111111111111110011001010011001;
assign LUT_2[9329] = 32'b11111111111111110000000010110010;
assign LUT_2[9330] = 32'b11111111111111111010000011010101;
assign LUT_2[9331] = 32'b11111111111111110110111011101110;
assign LUT_2[9332] = 32'b11111111111111101111101000000001;
assign LUT_2[9333] = 32'b11111111111111101100100000011010;
assign LUT_2[9334] = 32'b11111111111111110110100000111101;
assign LUT_2[9335] = 32'b11111111111111110011011001010110;
assign LUT_2[9336] = 32'b11111111111111101101111011110110;
assign LUT_2[9337] = 32'b11111111111111101010110100001111;
assign LUT_2[9338] = 32'b11111111111111110100110100110010;
assign LUT_2[9339] = 32'b11111111111111110001101101001011;
assign LUT_2[9340] = 32'b11111111111111101010011001011110;
assign LUT_2[9341] = 32'b11111111111111100111010001110111;
assign LUT_2[9342] = 32'b11111111111111110001010010011010;
assign LUT_2[9343] = 32'b11111111111111101110001010110011;
assign LUT_2[9344] = 32'b00000000000000000100010110010010;
assign LUT_2[9345] = 32'b00000000000000000001001110101011;
assign LUT_2[9346] = 32'b00000000000000001011001111001110;
assign LUT_2[9347] = 32'b00000000000000001000000111100111;
assign LUT_2[9348] = 32'b00000000000000000000110011111010;
assign LUT_2[9349] = 32'b11111111111111111101101100010011;
assign LUT_2[9350] = 32'b00000000000000000111101100110110;
assign LUT_2[9351] = 32'b00000000000000000100100101001111;
assign LUT_2[9352] = 32'b11111111111111111111000111101111;
assign LUT_2[9353] = 32'b11111111111111111100000000001000;
assign LUT_2[9354] = 32'b00000000000000000110000000101011;
assign LUT_2[9355] = 32'b00000000000000000010111001000100;
assign LUT_2[9356] = 32'b11111111111111111011100101010111;
assign LUT_2[9357] = 32'b11111111111111111000011101110000;
assign LUT_2[9358] = 32'b00000000000000000010011110010011;
assign LUT_2[9359] = 32'b11111111111111111111010110101100;
assign LUT_2[9360] = 32'b11111111111111111110111010011100;
assign LUT_2[9361] = 32'b11111111111111111011110010110101;
assign LUT_2[9362] = 32'b00000000000000000101110011011000;
assign LUT_2[9363] = 32'b00000000000000000010101011110001;
assign LUT_2[9364] = 32'b11111111111111111011011000000100;
assign LUT_2[9365] = 32'b11111111111111111000010000011101;
assign LUT_2[9366] = 32'b00000000000000000010010001000000;
assign LUT_2[9367] = 32'b11111111111111111111001001011001;
assign LUT_2[9368] = 32'b11111111111111111001101011111001;
assign LUT_2[9369] = 32'b11111111111111110110100100010010;
assign LUT_2[9370] = 32'b00000000000000000000100100110101;
assign LUT_2[9371] = 32'b11111111111111111101011101001110;
assign LUT_2[9372] = 32'b11111111111111110110001001100001;
assign LUT_2[9373] = 32'b11111111111111110011000001111010;
assign LUT_2[9374] = 32'b11111111111111111101000010011101;
assign LUT_2[9375] = 32'b11111111111111111001111010110110;
assign LUT_2[9376] = 32'b00000000000000000100110001111011;
assign LUT_2[9377] = 32'b00000000000000000001101010010100;
assign LUT_2[9378] = 32'b00000000000000001011101010110111;
assign LUT_2[9379] = 32'b00000000000000001000100011010000;
assign LUT_2[9380] = 32'b00000000000000000001001111100011;
assign LUT_2[9381] = 32'b11111111111111111110000111111100;
assign LUT_2[9382] = 32'b00000000000000001000001000011111;
assign LUT_2[9383] = 32'b00000000000000000101000000111000;
assign LUT_2[9384] = 32'b11111111111111111111100011011000;
assign LUT_2[9385] = 32'b11111111111111111100011011110001;
assign LUT_2[9386] = 32'b00000000000000000110011100010100;
assign LUT_2[9387] = 32'b00000000000000000011010100101101;
assign LUT_2[9388] = 32'b11111111111111111100000001000000;
assign LUT_2[9389] = 32'b11111111111111111000111001011001;
assign LUT_2[9390] = 32'b00000000000000000010111001111100;
assign LUT_2[9391] = 32'b11111111111111111111110010010101;
assign LUT_2[9392] = 32'b11111111111111111111010110000101;
assign LUT_2[9393] = 32'b11111111111111111100001110011110;
assign LUT_2[9394] = 32'b00000000000000000110001111000001;
assign LUT_2[9395] = 32'b00000000000000000011000111011010;
assign LUT_2[9396] = 32'b11111111111111111011110011101101;
assign LUT_2[9397] = 32'b11111111111111111000101100000110;
assign LUT_2[9398] = 32'b00000000000000000010101100101001;
assign LUT_2[9399] = 32'b11111111111111111111100101000010;
assign LUT_2[9400] = 32'b11111111111111111010000111100010;
assign LUT_2[9401] = 32'b11111111111111110110111111111011;
assign LUT_2[9402] = 32'b00000000000000000001000000011110;
assign LUT_2[9403] = 32'b11111111111111111101111000110111;
assign LUT_2[9404] = 32'b11111111111111110110100101001010;
assign LUT_2[9405] = 32'b11111111111111110011011101100011;
assign LUT_2[9406] = 32'b11111111111111111101011110000110;
assign LUT_2[9407] = 32'b11111111111111111010010110011111;
assign LUT_2[9408] = 32'b11111111111111111100011110110101;
assign LUT_2[9409] = 32'b11111111111111111001010111001110;
assign LUT_2[9410] = 32'b00000000000000000011010111110001;
assign LUT_2[9411] = 32'b00000000000000000000010000001010;
assign LUT_2[9412] = 32'b11111111111111111000111100011101;
assign LUT_2[9413] = 32'b11111111111111110101110100110110;
assign LUT_2[9414] = 32'b11111111111111111111110101011001;
assign LUT_2[9415] = 32'b11111111111111111100101101110010;
assign LUT_2[9416] = 32'b11111111111111110111010000010010;
assign LUT_2[9417] = 32'b11111111111111110100001000101011;
assign LUT_2[9418] = 32'b11111111111111111110001001001110;
assign LUT_2[9419] = 32'b11111111111111111011000001100111;
assign LUT_2[9420] = 32'b11111111111111110011101101111010;
assign LUT_2[9421] = 32'b11111111111111110000100110010011;
assign LUT_2[9422] = 32'b11111111111111111010100110110110;
assign LUT_2[9423] = 32'b11111111111111110111011111001111;
assign LUT_2[9424] = 32'b11111111111111110111000010111111;
assign LUT_2[9425] = 32'b11111111111111110011111011011000;
assign LUT_2[9426] = 32'b11111111111111111101111011111011;
assign LUT_2[9427] = 32'b11111111111111111010110100010100;
assign LUT_2[9428] = 32'b11111111111111110011100000100111;
assign LUT_2[9429] = 32'b11111111111111110000011001000000;
assign LUT_2[9430] = 32'b11111111111111111010011001100011;
assign LUT_2[9431] = 32'b11111111111111110111010001111100;
assign LUT_2[9432] = 32'b11111111111111110001110100011100;
assign LUT_2[9433] = 32'b11111111111111101110101100110101;
assign LUT_2[9434] = 32'b11111111111111111000101101011000;
assign LUT_2[9435] = 32'b11111111111111110101100101110001;
assign LUT_2[9436] = 32'b11111111111111101110010010000100;
assign LUT_2[9437] = 32'b11111111111111101011001010011101;
assign LUT_2[9438] = 32'b11111111111111110101001011000000;
assign LUT_2[9439] = 32'b11111111111111110010000011011001;
assign LUT_2[9440] = 32'b11111111111111111100111010011110;
assign LUT_2[9441] = 32'b11111111111111111001110010110111;
assign LUT_2[9442] = 32'b00000000000000000011110011011010;
assign LUT_2[9443] = 32'b00000000000000000000101011110011;
assign LUT_2[9444] = 32'b11111111111111111001011000000110;
assign LUT_2[9445] = 32'b11111111111111110110010000011111;
assign LUT_2[9446] = 32'b00000000000000000000010001000010;
assign LUT_2[9447] = 32'b11111111111111111101001001011011;
assign LUT_2[9448] = 32'b11111111111111110111101011111011;
assign LUT_2[9449] = 32'b11111111111111110100100100010100;
assign LUT_2[9450] = 32'b11111111111111111110100100110111;
assign LUT_2[9451] = 32'b11111111111111111011011101010000;
assign LUT_2[9452] = 32'b11111111111111110100001001100011;
assign LUT_2[9453] = 32'b11111111111111110001000001111100;
assign LUT_2[9454] = 32'b11111111111111111011000010011111;
assign LUT_2[9455] = 32'b11111111111111110111111010111000;
assign LUT_2[9456] = 32'b11111111111111110111011110101000;
assign LUT_2[9457] = 32'b11111111111111110100010111000001;
assign LUT_2[9458] = 32'b11111111111111111110010111100100;
assign LUT_2[9459] = 32'b11111111111111111011001111111101;
assign LUT_2[9460] = 32'b11111111111111110011111100010000;
assign LUT_2[9461] = 32'b11111111111111110000110100101001;
assign LUT_2[9462] = 32'b11111111111111111010110101001100;
assign LUT_2[9463] = 32'b11111111111111110111101101100101;
assign LUT_2[9464] = 32'b11111111111111110010010000000101;
assign LUT_2[9465] = 32'b11111111111111101111001000011110;
assign LUT_2[9466] = 32'b11111111111111111001001001000001;
assign LUT_2[9467] = 32'b11111111111111110110000001011010;
assign LUT_2[9468] = 32'b11111111111111101110101101101101;
assign LUT_2[9469] = 32'b11111111111111101011100110000110;
assign LUT_2[9470] = 32'b11111111111111110101100110101001;
assign LUT_2[9471] = 32'b11111111111111110010011111000010;
assign LUT_2[9472] = 32'b00000000000000000100000000101001;
assign LUT_2[9473] = 32'b00000000000000000000111001000010;
assign LUT_2[9474] = 32'b00000000000000001010111001100101;
assign LUT_2[9475] = 32'b00000000000000000111110001111110;
assign LUT_2[9476] = 32'b00000000000000000000011110010001;
assign LUT_2[9477] = 32'b11111111111111111101010110101010;
assign LUT_2[9478] = 32'b00000000000000000111010111001101;
assign LUT_2[9479] = 32'b00000000000000000100001111100110;
assign LUT_2[9480] = 32'b11111111111111111110110010000110;
assign LUT_2[9481] = 32'b11111111111111111011101010011111;
assign LUT_2[9482] = 32'b00000000000000000101101011000010;
assign LUT_2[9483] = 32'b00000000000000000010100011011011;
assign LUT_2[9484] = 32'b11111111111111111011001111101110;
assign LUT_2[9485] = 32'b11111111111111111000001000000111;
assign LUT_2[9486] = 32'b00000000000000000010001000101010;
assign LUT_2[9487] = 32'b11111111111111111111000001000011;
assign LUT_2[9488] = 32'b11111111111111111110100100110011;
assign LUT_2[9489] = 32'b11111111111111111011011101001100;
assign LUT_2[9490] = 32'b00000000000000000101011101101111;
assign LUT_2[9491] = 32'b00000000000000000010010110001000;
assign LUT_2[9492] = 32'b11111111111111111011000010011011;
assign LUT_2[9493] = 32'b11111111111111110111111010110100;
assign LUT_2[9494] = 32'b00000000000000000001111011010111;
assign LUT_2[9495] = 32'b11111111111111111110110011110000;
assign LUT_2[9496] = 32'b11111111111111111001010110010000;
assign LUT_2[9497] = 32'b11111111111111110110001110101001;
assign LUT_2[9498] = 32'b00000000000000000000001111001100;
assign LUT_2[9499] = 32'b11111111111111111101000111100101;
assign LUT_2[9500] = 32'b11111111111111110101110011111000;
assign LUT_2[9501] = 32'b11111111111111110010101100010001;
assign LUT_2[9502] = 32'b11111111111111111100101100110100;
assign LUT_2[9503] = 32'b11111111111111111001100101001101;
assign LUT_2[9504] = 32'b00000000000000000100011100010010;
assign LUT_2[9505] = 32'b00000000000000000001010100101011;
assign LUT_2[9506] = 32'b00000000000000001011010101001110;
assign LUT_2[9507] = 32'b00000000000000001000001101100111;
assign LUT_2[9508] = 32'b00000000000000000000111001111010;
assign LUT_2[9509] = 32'b11111111111111111101110010010011;
assign LUT_2[9510] = 32'b00000000000000000111110010110110;
assign LUT_2[9511] = 32'b00000000000000000100101011001111;
assign LUT_2[9512] = 32'b11111111111111111111001101101111;
assign LUT_2[9513] = 32'b11111111111111111100000110001000;
assign LUT_2[9514] = 32'b00000000000000000110000110101011;
assign LUT_2[9515] = 32'b00000000000000000010111111000100;
assign LUT_2[9516] = 32'b11111111111111111011101011010111;
assign LUT_2[9517] = 32'b11111111111111111000100011110000;
assign LUT_2[9518] = 32'b00000000000000000010100100010011;
assign LUT_2[9519] = 32'b11111111111111111111011100101100;
assign LUT_2[9520] = 32'b11111111111111111111000000011100;
assign LUT_2[9521] = 32'b11111111111111111011111000110101;
assign LUT_2[9522] = 32'b00000000000000000101111001011000;
assign LUT_2[9523] = 32'b00000000000000000010110001110001;
assign LUT_2[9524] = 32'b11111111111111111011011110000100;
assign LUT_2[9525] = 32'b11111111111111111000010110011101;
assign LUT_2[9526] = 32'b00000000000000000010010111000000;
assign LUT_2[9527] = 32'b11111111111111111111001111011001;
assign LUT_2[9528] = 32'b11111111111111111001110001111001;
assign LUT_2[9529] = 32'b11111111111111110110101010010010;
assign LUT_2[9530] = 32'b00000000000000000000101010110101;
assign LUT_2[9531] = 32'b11111111111111111101100011001110;
assign LUT_2[9532] = 32'b11111111111111110110001111100001;
assign LUT_2[9533] = 32'b11111111111111110011000111111010;
assign LUT_2[9534] = 32'b11111111111111111101001000011101;
assign LUT_2[9535] = 32'b11111111111111111010000000110110;
assign LUT_2[9536] = 32'b11111111111111111100001001001100;
assign LUT_2[9537] = 32'b11111111111111111001000001100101;
assign LUT_2[9538] = 32'b00000000000000000011000010001000;
assign LUT_2[9539] = 32'b11111111111111111111111010100001;
assign LUT_2[9540] = 32'b11111111111111111000100110110100;
assign LUT_2[9541] = 32'b11111111111111110101011111001101;
assign LUT_2[9542] = 32'b11111111111111111111011111110000;
assign LUT_2[9543] = 32'b11111111111111111100011000001001;
assign LUT_2[9544] = 32'b11111111111111110110111010101001;
assign LUT_2[9545] = 32'b11111111111111110011110011000010;
assign LUT_2[9546] = 32'b11111111111111111101110011100101;
assign LUT_2[9547] = 32'b11111111111111111010101011111110;
assign LUT_2[9548] = 32'b11111111111111110011011000010001;
assign LUT_2[9549] = 32'b11111111111111110000010000101010;
assign LUT_2[9550] = 32'b11111111111111111010010001001101;
assign LUT_2[9551] = 32'b11111111111111110111001001100110;
assign LUT_2[9552] = 32'b11111111111111110110101101010110;
assign LUT_2[9553] = 32'b11111111111111110011100101101111;
assign LUT_2[9554] = 32'b11111111111111111101100110010010;
assign LUT_2[9555] = 32'b11111111111111111010011110101011;
assign LUT_2[9556] = 32'b11111111111111110011001010111110;
assign LUT_2[9557] = 32'b11111111111111110000000011010111;
assign LUT_2[9558] = 32'b11111111111111111010000011111010;
assign LUT_2[9559] = 32'b11111111111111110110111100010011;
assign LUT_2[9560] = 32'b11111111111111110001011110110011;
assign LUT_2[9561] = 32'b11111111111111101110010111001100;
assign LUT_2[9562] = 32'b11111111111111111000010111101111;
assign LUT_2[9563] = 32'b11111111111111110101010000001000;
assign LUT_2[9564] = 32'b11111111111111101101111100011011;
assign LUT_2[9565] = 32'b11111111111111101010110100110100;
assign LUT_2[9566] = 32'b11111111111111110100110101010111;
assign LUT_2[9567] = 32'b11111111111111110001101101110000;
assign LUT_2[9568] = 32'b11111111111111111100100100110101;
assign LUT_2[9569] = 32'b11111111111111111001011101001110;
assign LUT_2[9570] = 32'b00000000000000000011011101110001;
assign LUT_2[9571] = 32'b00000000000000000000010110001010;
assign LUT_2[9572] = 32'b11111111111111111001000010011101;
assign LUT_2[9573] = 32'b11111111111111110101111010110110;
assign LUT_2[9574] = 32'b11111111111111111111111011011001;
assign LUT_2[9575] = 32'b11111111111111111100110011110010;
assign LUT_2[9576] = 32'b11111111111111110111010110010010;
assign LUT_2[9577] = 32'b11111111111111110100001110101011;
assign LUT_2[9578] = 32'b11111111111111111110001111001110;
assign LUT_2[9579] = 32'b11111111111111111011000111100111;
assign LUT_2[9580] = 32'b11111111111111110011110011111010;
assign LUT_2[9581] = 32'b11111111111111110000101100010011;
assign LUT_2[9582] = 32'b11111111111111111010101100110110;
assign LUT_2[9583] = 32'b11111111111111110111100101001111;
assign LUT_2[9584] = 32'b11111111111111110111001000111111;
assign LUT_2[9585] = 32'b11111111111111110100000001011000;
assign LUT_2[9586] = 32'b11111111111111111110000001111011;
assign LUT_2[9587] = 32'b11111111111111111010111010010100;
assign LUT_2[9588] = 32'b11111111111111110011100110100111;
assign LUT_2[9589] = 32'b11111111111111110000011111000000;
assign LUT_2[9590] = 32'b11111111111111111010011111100011;
assign LUT_2[9591] = 32'b11111111111111110111010111111100;
assign LUT_2[9592] = 32'b11111111111111110001111010011100;
assign LUT_2[9593] = 32'b11111111111111101110110010110101;
assign LUT_2[9594] = 32'b11111111111111111000110011011000;
assign LUT_2[9595] = 32'b11111111111111110101101011110001;
assign LUT_2[9596] = 32'b11111111111111101110011000000100;
assign LUT_2[9597] = 32'b11111111111111101011010000011101;
assign LUT_2[9598] = 32'b11111111111111110101010001000000;
assign LUT_2[9599] = 32'b11111111111111110010001001011001;
assign LUT_2[9600] = 32'b00000000000000001000010100111000;
assign LUT_2[9601] = 32'b00000000000000000101001101010001;
assign LUT_2[9602] = 32'b00000000000000001111001101110100;
assign LUT_2[9603] = 32'b00000000000000001100000110001101;
assign LUT_2[9604] = 32'b00000000000000000100110010100000;
assign LUT_2[9605] = 32'b00000000000000000001101010111001;
assign LUT_2[9606] = 32'b00000000000000001011101011011100;
assign LUT_2[9607] = 32'b00000000000000001000100011110101;
assign LUT_2[9608] = 32'b00000000000000000011000110010101;
assign LUT_2[9609] = 32'b11111111111111111111111110101110;
assign LUT_2[9610] = 32'b00000000000000001001111111010001;
assign LUT_2[9611] = 32'b00000000000000000110110111101010;
assign LUT_2[9612] = 32'b11111111111111111111100011111101;
assign LUT_2[9613] = 32'b11111111111111111100011100010110;
assign LUT_2[9614] = 32'b00000000000000000110011100111001;
assign LUT_2[9615] = 32'b00000000000000000011010101010010;
assign LUT_2[9616] = 32'b00000000000000000010111001000010;
assign LUT_2[9617] = 32'b11111111111111111111110001011011;
assign LUT_2[9618] = 32'b00000000000000001001110001111110;
assign LUT_2[9619] = 32'b00000000000000000110101010010111;
assign LUT_2[9620] = 32'b11111111111111111111010110101010;
assign LUT_2[9621] = 32'b11111111111111111100001111000011;
assign LUT_2[9622] = 32'b00000000000000000110001111100110;
assign LUT_2[9623] = 32'b00000000000000000011000111111111;
assign LUT_2[9624] = 32'b11111111111111111101101010011111;
assign LUT_2[9625] = 32'b11111111111111111010100010111000;
assign LUT_2[9626] = 32'b00000000000000000100100011011011;
assign LUT_2[9627] = 32'b00000000000000000001011011110100;
assign LUT_2[9628] = 32'b11111111111111111010001000000111;
assign LUT_2[9629] = 32'b11111111111111110111000000100000;
assign LUT_2[9630] = 32'b00000000000000000001000001000011;
assign LUT_2[9631] = 32'b11111111111111111101111001011100;
assign LUT_2[9632] = 32'b00000000000000001000110000100001;
assign LUT_2[9633] = 32'b00000000000000000101101000111010;
assign LUT_2[9634] = 32'b00000000000000001111101001011101;
assign LUT_2[9635] = 32'b00000000000000001100100001110110;
assign LUT_2[9636] = 32'b00000000000000000101001110001001;
assign LUT_2[9637] = 32'b00000000000000000010000110100010;
assign LUT_2[9638] = 32'b00000000000000001100000111000101;
assign LUT_2[9639] = 32'b00000000000000001000111111011110;
assign LUT_2[9640] = 32'b00000000000000000011100001111110;
assign LUT_2[9641] = 32'b00000000000000000000011010010111;
assign LUT_2[9642] = 32'b00000000000000001010011010111010;
assign LUT_2[9643] = 32'b00000000000000000111010011010011;
assign LUT_2[9644] = 32'b11111111111111111111111111100110;
assign LUT_2[9645] = 32'b11111111111111111100110111111111;
assign LUT_2[9646] = 32'b00000000000000000110111000100010;
assign LUT_2[9647] = 32'b00000000000000000011110000111011;
assign LUT_2[9648] = 32'b00000000000000000011010100101011;
assign LUT_2[9649] = 32'b00000000000000000000001101000100;
assign LUT_2[9650] = 32'b00000000000000001010001101100111;
assign LUT_2[9651] = 32'b00000000000000000111000110000000;
assign LUT_2[9652] = 32'b11111111111111111111110010010011;
assign LUT_2[9653] = 32'b11111111111111111100101010101100;
assign LUT_2[9654] = 32'b00000000000000000110101011001111;
assign LUT_2[9655] = 32'b00000000000000000011100011101000;
assign LUT_2[9656] = 32'b11111111111111111110000110001000;
assign LUT_2[9657] = 32'b11111111111111111010111110100001;
assign LUT_2[9658] = 32'b00000000000000000100111111000100;
assign LUT_2[9659] = 32'b00000000000000000001110111011101;
assign LUT_2[9660] = 32'b11111111111111111010100011110000;
assign LUT_2[9661] = 32'b11111111111111110111011100001001;
assign LUT_2[9662] = 32'b00000000000000000001011100101100;
assign LUT_2[9663] = 32'b11111111111111111110010101000101;
assign LUT_2[9664] = 32'b00000000000000000000011101011011;
assign LUT_2[9665] = 32'b11111111111111111101010101110100;
assign LUT_2[9666] = 32'b00000000000000000111010110010111;
assign LUT_2[9667] = 32'b00000000000000000100001110110000;
assign LUT_2[9668] = 32'b11111111111111111100111011000011;
assign LUT_2[9669] = 32'b11111111111111111001110011011100;
assign LUT_2[9670] = 32'b00000000000000000011110011111111;
assign LUT_2[9671] = 32'b00000000000000000000101100011000;
assign LUT_2[9672] = 32'b11111111111111111011001110111000;
assign LUT_2[9673] = 32'b11111111111111111000000111010001;
assign LUT_2[9674] = 32'b00000000000000000010000111110100;
assign LUT_2[9675] = 32'b11111111111111111111000000001101;
assign LUT_2[9676] = 32'b11111111111111110111101100100000;
assign LUT_2[9677] = 32'b11111111111111110100100100111001;
assign LUT_2[9678] = 32'b11111111111111111110100101011100;
assign LUT_2[9679] = 32'b11111111111111111011011101110101;
assign LUT_2[9680] = 32'b11111111111111111011000001100101;
assign LUT_2[9681] = 32'b11111111111111110111111001111110;
assign LUT_2[9682] = 32'b00000000000000000001111010100001;
assign LUT_2[9683] = 32'b11111111111111111110110010111010;
assign LUT_2[9684] = 32'b11111111111111110111011111001101;
assign LUT_2[9685] = 32'b11111111111111110100010111100110;
assign LUT_2[9686] = 32'b11111111111111111110011000001001;
assign LUT_2[9687] = 32'b11111111111111111011010000100010;
assign LUT_2[9688] = 32'b11111111111111110101110011000010;
assign LUT_2[9689] = 32'b11111111111111110010101011011011;
assign LUT_2[9690] = 32'b11111111111111111100101011111110;
assign LUT_2[9691] = 32'b11111111111111111001100100010111;
assign LUT_2[9692] = 32'b11111111111111110010010000101010;
assign LUT_2[9693] = 32'b11111111111111101111001001000011;
assign LUT_2[9694] = 32'b11111111111111111001001001100110;
assign LUT_2[9695] = 32'b11111111111111110110000001111111;
assign LUT_2[9696] = 32'b00000000000000000000111001000100;
assign LUT_2[9697] = 32'b11111111111111111101110001011101;
assign LUT_2[9698] = 32'b00000000000000000111110010000000;
assign LUT_2[9699] = 32'b00000000000000000100101010011001;
assign LUT_2[9700] = 32'b11111111111111111101010110101100;
assign LUT_2[9701] = 32'b11111111111111111010001111000101;
assign LUT_2[9702] = 32'b00000000000000000100001111101000;
assign LUT_2[9703] = 32'b00000000000000000001001000000001;
assign LUT_2[9704] = 32'b11111111111111111011101010100001;
assign LUT_2[9705] = 32'b11111111111111111000100010111010;
assign LUT_2[9706] = 32'b00000000000000000010100011011101;
assign LUT_2[9707] = 32'b11111111111111111111011011110110;
assign LUT_2[9708] = 32'b11111111111111111000001000001001;
assign LUT_2[9709] = 32'b11111111111111110101000000100010;
assign LUT_2[9710] = 32'b11111111111111111111000001000101;
assign LUT_2[9711] = 32'b11111111111111111011111001011110;
assign LUT_2[9712] = 32'b11111111111111111011011101001110;
assign LUT_2[9713] = 32'b11111111111111111000010101100111;
assign LUT_2[9714] = 32'b00000000000000000010010110001010;
assign LUT_2[9715] = 32'b11111111111111111111001110100011;
assign LUT_2[9716] = 32'b11111111111111110111111010110110;
assign LUT_2[9717] = 32'b11111111111111110100110011001111;
assign LUT_2[9718] = 32'b11111111111111111110110011110010;
assign LUT_2[9719] = 32'b11111111111111111011101100001011;
assign LUT_2[9720] = 32'b11111111111111110110001110101011;
assign LUT_2[9721] = 32'b11111111111111110011000111000100;
assign LUT_2[9722] = 32'b11111111111111111101000111100111;
assign LUT_2[9723] = 32'b11111111111111111010000000000000;
assign LUT_2[9724] = 32'b11111111111111110010101100010011;
assign LUT_2[9725] = 32'b11111111111111101111100100101100;
assign LUT_2[9726] = 32'b11111111111111111001100101001111;
assign LUT_2[9727] = 32'b11111111111111110110011101101000;
assign LUT_2[9728] = 32'b00000000000000000100110011110101;
assign LUT_2[9729] = 32'b00000000000000000001101100001110;
assign LUT_2[9730] = 32'b00000000000000001011101100110001;
assign LUT_2[9731] = 32'b00000000000000001000100101001010;
assign LUT_2[9732] = 32'b00000000000000000001010001011101;
assign LUT_2[9733] = 32'b11111111111111111110001001110110;
assign LUT_2[9734] = 32'b00000000000000001000001010011001;
assign LUT_2[9735] = 32'b00000000000000000101000010110010;
assign LUT_2[9736] = 32'b11111111111111111111100101010010;
assign LUT_2[9737] = 32'b11111111111111111100011101101011;
assign LUT_2[9738] = 32'b00000000000000000110011110001110;
assign LUT_2[9739] = 32'b00000000000000000011010110100111;
assign LUT_2[9740] = 32'b11111111111111111100000010111010;
assign LUT_2[9741] = 32'b11111111111111111000111011010011;
assign LUT_2[9742] = 32'b00000000000000000010111011110110;
assign LUT_2[9743] = 32'b11111111111111111111110100001111;
assign LUT_2[9744] = 32'b11111111111111111111010111111111;
assign LUT_2[9745] = 32'b11111111111111111100010000011000;
assign LUT_2[9746] = 32'b00000000000000000110010000111011;
assign LUT_2[9747] = 32'b00000000000000000011001001010100;
assign LUT_2[9748] = 32'b11111111111111111011110101100111;
assign LUT_2[9749] = 32'b11111111111111111000101110000000;
assign LUT_2[9750] = 32'b00000000000000000010101110100011;
assign LUT_2[9751] = 32'b11111111111111111111100110111100;
assign LUT_2[9752] = 32'b11111111111111111010001001011100;
assign LUT_2[9753] = 32'b11111111111111110111000001110101;
assign LUT_2[9754] = 32'b00000000000000000001000010011000;
assign LUT_2[9755] = 32'b11111111111111111101111010110001;
assign LUT_2[9756] = 32'b11111111111111110110100111000100;
assign LUT_2[9757] = 32'b11111111111111110011011111011101;
assign LUT_2[9758] = 32'b11111111111111111101100000000000;
assign LUT_2[9759] = 32'b11111111111111111010011000011001;
assign LUT_2[9760] = 32'b00000000000000000101001111011110;
assign LUT_2[9761] = 32'b00000000000000000010000111110111;
assign LUT_2[9762] = 32'b00000000000000001100001000011010;
assign LUT_2[9763] = 32'b00000000000000001001000000110011;
assign LUT_2[9764] = 32'b00000000000000000001101101000110;
assign LUT_2[9765] = 32'b11111111111111111110100101011111;
assign LUT_2[9766] = 32'b00000000000000001000100110000010;
assign LUT_2[9767] = 32'b00000000000000000101011110011011;
assign LUT_2[9768] = 32'b00000000000000000000000000111011;
assign LUT_2[9769] = 32'b11111111111111111100111001010100;
assign LUT_2[9770] = 32'b00000000000000000110111001110111;
assign LUT_2[9771] = 32'b00000000000000000011110010010000;
assign LUT_2[9772] = 32'b11111111111111111100011110100011;
assign LUT_2[9773] = 32'b11111111111111111001010110111100;
assign LUT_2[9774] = 32'b00000000000000000011010111011111;
assign LUT_2[9775] = 32'b00000000000000000000001111111000;
assign LUT_2[9776] = 32'b11111111111111111111110011101000;
assign LUT_2[9777] = 32'b11111111111111111100101100000001;
assign LUT_2[9778] = 32'b00000000000000000110101100100100;
assign LUT_2[9779] = 32'b00000000000000000011100100111101;
assign LUT_2[9780] = 32'b11111111111111111100010001010000;
assign LUT_2[9781] = 32'b11111111111111111001001001101001;
assign LUT_2[9782] = 32'b00000000000000000011001010001100;
assign LUT_2[9783] = 32'b00000000000000000000000010100101;
assign LUT_2[9784] = 32'b11111111111111111010100101000101;
assign LUT_2[9785] = 32'b11111111111111110111011101011110;
assign LUT_2[9786] = 32'b00000000000000000001011110000001;
assign LUT_2[9787] = 32'b11111111111111111110010110011010;
assign LUT_2[9788] = 32'b11111111111111110111000010101101;
assign LUT_2[9789] = 32'b11111111111111110011111011000110;
assign LUT_2[9790] = 32'b11111111111111111101111011101001;
assign LUT_2[9791] = 32'b11111111111111111010110100000010;
assign LUT_2[9792] = 32'b11111111111111111100111100011000;
assign LUT_2[9793] = 32'b11111111111111111001110100110001;
assign LUT_2[9794] = 32'b00000000000000000011110101010100;
assign LUT_2[9795] = 32'b00000000000000000000101101101101;
assign LUT_2[9796] = 32'b11111111111111111001011010000000;
assign LUT_2[9797] = 32'b11111111111111110110010010011001;
assign LUT_2[9798] = 32'b00000000000000000000010010111100;
assign LUT_2[9799] = 32'b11111111111111111101001011010101;
assign LUT_2[9800] = 32'b11111111111111110111101101110101;
assign LUT_2[9801] = 32'b11111111111111110100100110001110;
assign LUT_2[9802] = 32'b11111111111111111110100110110001;
assign LUT_2[9803] = 32'b11111111111111111011011111001010;
assign LUT_2[9804] = 32'b11111111111111110100001011011101;
assign LUT_2[9805] = 32'b11111111111111110001000011110110;
assign LUT_2[9806] = 32'b11111111111111111011000100011001;
assign LUT_2[9807] = 32'b11111111111111110111111100110010;
assign LUT_2[9808] = 32'b11111111111111110111100000100010;
assign LUT_2[9809] = 32'b11111111111111110100011000111011;
assign LUT_2[9810] = 32'b11111111111111111110011001011110;
assign LUT_2[9811] = 32'b11111111111111111011010001110111;
assign LUT_2[9812] = 32'b11111111111111110011111110001010;
assign LUT_2[9813] = 32'b11111111111111110000110110100011;
assign LUT_2[9814] = 32'b11111111111111111010110111000110;
assign LUT_2[9815] = 32'b11111111111111110111101111011111;
assign LUT_2[9816] = 32'b11111111111111110010010001111111;
assign LUT_2[9817] = 32'b11111111111111101111001010011000;
assign LUT_2[9818] = 32'b11111111111111111001001010111011;
assign LUT_2[9819] = 32'b11111111111111110110000011010100;
assign LUT_2[9820] = 32'b11111111111111101110101111100111;
assign LUT_2[9821] = 32'b11111111111111101011101000000000;
assign LUT_2[9822] = 32'b11111111111111110101101000100011;
assign LUT_2[9823] = 32'b11111111111111110010100000111100;
assign LUT_2[9824] = 32'b11111111111111111101011000000001;
assign LUT_2[9825] = 32'b11111111111111111010010000011010;
assign LUT_2[9826] = 32'b00000000000000000100010000111101;
assign LUT_2[9827] = 32'b00000000000000000001001001010110;
assign LUT_2[9828] = 32'b11111111111111111001110101101001;
assign LUT_2[9829] = 32'b11111111111111110110101110000010;
assign LUT_2[9830] = 32'b00000000000000000000101110100101;
assign LUT_2[9831] = 32'b11111111111111111101100110111110;
assign LUT_2[9832] = 32'b11111111111111111000001001011110;
assign LUT_2[9833] = 32'b11111111111111110101000001110111;
assign LUT_2[9834] = 32'b11111111111111111111000010011010;
assign LUT_2[9835] = 32'b11111111111111111011111010110011;
assign LUT_2[9836] = 32'b11111111111111110100100111000110;
assign LUT_2[9837] = 32'b11111111111111110001011111011111;
assign LUT_2[9838] = 32'b11111111111111111011100000000010;
assign LUT_2[9839] = 32'b11111111111111111000011000011011;
assign LUT_2[9840] = 32'b11111111111111110111111100001011;
assign LUT_2[9841] = 32'b11111111111111110100110100100100;
assign LUT_2[9842] = 32'b11111111111111111110110101000111;
assign LUT_2[9843] = 32'b11111111111111111011101101100000;
assign LUT_2[9844] = 32'b11111111111111110100011001110011;
assign LUT_2[9845] = 32'b11111111111111110001010010001100;
assign LUT_2[9846] = 32'b11111111111111111011010010101111;
assign LUT_2[9847] = 32'b11111111111111111000001011001000;
assign LUT_2[9848] = 32'b11111111111111110010101101101000;
assign LUT_2[9849] = 32'b11111111111111101111100110000001;
assign LUT_2[9850] = 32'b11111111111111111001100110100100;
assign LUT_2[9851] = 32'b11111111111111110110011110111101;
assign LUT_2[9852] = 32'b11111111111111101111001011010000;
assign LUT_2[9853] = 32'b11111111111111101100000011101001;
assign LUT_2[9854] = 32'b11111111111111110110000100001100;
assign LUT_2[9855] = 32'b11111111111111110010111100100101;
assign LUT_2[9856] = 32'b00000000000000001001001000000100;
assign LUT_2[9857] = 32'b00000000000000000110000000011101;
assign LUT_2[9858] = 32'b00000000000000010000000001000000;
assign LUT_2[9859] = 32'b00000000000000001100111001011001;
assign LUT_2[9860] = 32'b00000000000000000101100101101100;
assign LUT_2[9861] = 32'b00000000000000000010011110000101;
assign LUT_2[9862] = 32'b00000000000000001100011110101000;
assign LUT_2[9863] = 32'b00000000000000001001010111000001;
assign LUT_2[9864] = 32'b00000000000000000011111001100001;
assign LUT_2[9865] = 32'b00000000000000000000110001111010;
assign LUT_2[9866] = 32'b00000000000000001010110010011101;
assign LUT_2[9867] = 32'b00000000000000000111101010110110;
assign LUT_2[9868] = 32'b00000000000000000000010111001001;
assign LUT_2[9869] = 32'b11111111111111111101001111100010;
assign LUT_2[9870] = 32'b00000000000000000111010000000101;
assign LUT_2[9871] = 32'b00000000000000000100001000011110;
assign LUT_2[9872] = 32'b00000000000000000011101100001110;
assign LUT_2[9873] = 32'b00000000000000000000100100100111;
assign LUT_2[9874] = 32'b00000000000000001010100101001010;
assign LUT_2[9875] = 32'b00000000000000000111011101100011;
assign LUT_2[9876] = 32'b00000000000000000000001001110110;
assign LUT_2[9877] = 32'b11111111111111111101000010001111;
assign LUT_2[9878] = 32'b00000000000000000111000010110010;
assign LUT_2[9879] = 32'b00000000000000000011111011001011;
assign LUT_2[9880] = 32'b11111111111111111110011101101011;
assign LUT_2[9881] = 32'b11111111111111111011010110000100;
assign LUT_2[9882] = 32'b00000000000000000101010110100111;
assign LUT_2[9883] = 32'b00000000000000000010001111000000;
assign LUT_2[9884] = 32'b11111111111111111010111011010011;
assign LUT_2[9885] = 32'b11111111111111110111110011101100;
assign LUT_2[9886] = 32'b00000000000000000001110100001111;
assign LUT_2[9887] = 32'b11111111111111111110101100101000;
assign LUT_2[9888] = 32'b00000000000000001001100011101101;
assign LUT_2[9889] = 32'b00000000000000000110011100000110;
assign LUT_2[9890] = 32'b00000000000000010000011100101001;
assign LUT_2[9891] = 32'b00000000000000001101010101000010;
assign LUT_2[9892] = 32'b00000000000000000110000001010101;
assign LUT_2[9893] = 32'b00000000000000000010111001101110;
assign LUT_2[9894] = 32'b00000000000000001100111010010001;
assign LUT_2[9895] = 32'b00000000000000001001110010101010;
assign LUT_2[9896] = 32'b00000000000000000100010101001010;
assign LUT_2[9897] = 32'b00000000000000000001001101100011;
assign LUT_2[9898] = 32'b00000000000000001011001110000110;
assign LUT_2[9899] = 32'b00000000000000001000000110011111;
assign LUT_2[9900] = 32'b00000000000000000000110010110010;
assign LUT_2[9901] = 32'b11111111111111111101101011001011;
assign LUT_2[9902] = 32'b00000000000000000111101011101110;
assign LUT_2[9903] = 32'b00000000000000000100100100000111;
assign LUT_2[9904] = 32'b00000000000000000100000111110111;
assign LUT_2[9905] = 32'b00000000000000000001000000010000;
assign LUT_2[9906] = 32'b00000000000000001011000000110011;
assign LUT_2[9907] = 32'b00000000000000000111111001001100;
assign LUT_2[9908] = 32'b00000000000000000000100101011111;
assign LUT_2[9909] = 32'b11111111111111111101011101111000;
assign LUT_2[9910] = 32'b00000000000000000111011110011011;
assign LUT_2[9911] = 32'b00000000000000000100010110110100;
assign LUT_2[9912] = 32'b11111111111111111110111001010100;
assign LUT_2[9913] = 32'b11111111111111111011110001101101;
assign LUT_2[9914] = 32'b00000000000000000101110010010000;
assign LUT_2[9915] = 32'b00000000000000000010101010101001;
assign LUT_2[9916] = 32'b11111111111111111011010110111100;
assign LUT_2[9917] = 32'b11111111111111111000001111010101;
assign LUT_2[9918] = 32'b00000000000000000010001111111000;
assign LUT_2[9919] = 32'b11111111111111111111001000010001;
assign LUT_2[9920] = 32'b00000000000000000001010000100111;
assign LUT_2[9921] = 32'b11111111111111111110001001000000;
assign LUT_2[9922] = 32'b00000000000000001000001001100011;
assign LUT_2[9923] = 32'b00000000000000000101000001111100;
assign LUT_2[9924] = 32'b11111111111111111101101110001111;
assign LUT_2[9925] = 32'b11111111111111111010100110101000;
assign LUT_2[9926] = 32'b00000000000000000100100111001011;
assign LUT_2[9927] = 32'b00000000000000000001011111100100;
assign LUT_2[9928] = 32'b11111111111111111100000010000100;
assign LUT_2[9929] = 32'b11111111111111111000111010011101;
assign LUT_2[9930] = 32'b00000000000000000010111011000000;
assign LUT_2[9931] = 32'b11111111111111111111110011011001;
assign LUT_2[9932] = 32'b11111111111111111000011111101100;
assign LUT_2[9933] = 32'b11111111111111110101011000000101;
assign LUT_2[9934] = 32'b11111111111111111111011000101000;
assign LUT_2[9935] = 32'b11111111111111111100010001000001;
assign LUT_2[9936] = 32'b11111111111111111011110100110001;
assign LUT_2[9937] = 32'b11111111111111111000101101001010;
assign LUT_2[9938] = 32'b00000000000000000010101101101101;
assign LUT_2[9939] = 32'b11111111111111111111100110000110;
assign LUT_2[9940] = 32'b11111111111111111000010010011001;
assign LUT_2[9941] = 32'b11111111111111110101001010110010;
assign LUT_2[9942] = 32'b11111111111111111111001011010101;
assign LUT_2[9943] = 32'b11111111111111111100000011101110;
assign LUT_2[9944] = 32'b11111111111111110110100110001110;
assign LUT_2[9945] = 32'b11111111111111110011011110100111;
assign LUT_2[9946] = 32'b11111111111111111101011111001010;
assign LUT_2[9947] = 32'b11111111111111111010010111100011;
assign LUT_2[9948] = 32'b11111111111111110011000011110110;
assign LUT_2[9949] = 32'b11111111111111101111111100001111;
assign LUT_2[9950] = 32'b11111111111111111001111100110010;
assign LUT_2[9951] = 32'b11111111111111110110110101001011;
assign LUT_2[9952] = 32'b00000000000000000001101100010000;
assign LUT_2[9953] = 32'b11111111111111111110100100101001;
assign LUT_2[9954] = 32'b00000000000000001000100101001100;
assign LUT_2[9955] = 32'b00000000000000000101011101100101;
assign LUT_2[9956] = 32'b11111111111111111110001001111000;
assign LUT_2[9957] = 32'b11111111111111111011000010010001;
assign LUT_2[9958] = 32'b00000000000000000101000010110100;
assign LUT_2[9959] = 32'b00000000000000000001111011001101;
assign LUT_2[9960] = 32'b11111111111111111100011101101101;
assign LUT_2[9961] = 32'b11111111111111111001010110000110;
assign LUT_2[9962] = 32'b00000000000000000011010110101001;
assign LUT_2[9963] = 32'b00000000000000000000001111000010;
assign LUT_2[9964] = 32'b11111111111111111000111011010101;
assign LUT_2[9965] = 32'b11111111111111110101110011101110;
assign LUT_2[9966] = 32'b11111111111111111111110100010001;
assign LUT_2[9967] = 32'b11111111111111111100101100101010;
assign LUT_2[9968] = 32'b11111111111111111100010000011010;
assign LUT_2[9969] = 32'b11111111111111111001001000110011;
assign LUT_2[9970] = 32'b00000000000000000011001001010110;
assign LUT_2[9971] = 32'b00000000000000000000000001101111;
assign LUT_2[9972] = 32'b11111111111111111000101110000010;
assign LUT_2[9973] = 32'b11111111111111110101100110011011;
assign LUT_2[9974] = 32'b11111111111111111111100110111110;
assign LUT_2[9975] = 32'b11111111111111111100011111010111;
assign LUT_2[9976] = 32'b11111111111111110111000001110111;
assign LUT_2[9977] = 32'b11111111111111110011111010010000;
assign LUT_2[9978] = 32'b11111111111111111101111010110011;
assign LUT_2[9979] = 32'b11111111111111111010110011001100;
assign LUT_2[9980] = 32'b11111111111111110011011111011111;
assign LUT_2[9981] = 32'b11111111111111110000010111111000;
assign LUT_2[9982] = 32'b11111111111111111010011000011011;
assign LUT_2[9983] = 32'b11111111111111110111010000110100;
assign LUT_2[9984] = 32'b00000000000000001000110010011011;
assign LUT_2[9985] = 32'b00000000000000000101101010110100;
assign LUT_2[9986] = 32'b00000000000000001111101011010111;
assign LUT_2[9987] = 32'b00000000000000001100100011110000;
assign LUT_2[9988] = 32'b00000000000000000101010000000011;
assign LUT_2[9989] = 32'b00000000000000000010001000011100;
assign LUT_2[9990] = 32'b00000000000000001100001000111111;
assign LUT_2[9991] = 32'b00000000000000001001000001011000;
assign LUT_2[9992] = 32'b00000000000000000011100011111000;
assign LUT_2[9993] = 32'b00000000000000000000011100010001;
assign LUT_2[9994] = 32'b00000000000000001010011100110100;
assign LUT_2[9995] = 32'b00000000000000000111010101001101;
assign LUT_2[9996] = 32'b00000000000000000000000001100000;
assign LUT_2[9997] = 32'b11111111111111111100111001111001;
assign LUT_2[9998] = 32'b00000000000000000110111010011100;
assign LUT_2[9999] = 32'b00000000000000000011110010110101;
assign LUT_2[10000] = 32'b00000000000000000011010110100101;
assign LUT_2[10001] = 32'b00000000000000000000001110111110;
assign LUT_2[10002] = 32'b00000000000000001010001111100001;
assign LUT_2[10003] = 32'b00000000000000000111000111111010;
assign LUT_2[10004] = 32'b11111111111111111111110100001101;
assign LUT_2[10005] = 32'b11111111111111111100101100100110;
assign LUT_2[10006] = 32'b00000000000000000110101101001001;
assign LUT_2[10007] = 32'b00000000000000000011100101100010;
assign LUT_2[10008] = 32'b11111111111111111110001000000010;
assign LUT_2[10009] = 32'b11111111111111111011000000011011;
assign LUT_2[10010] = 32'b00000000000000000101000000111110;
assign LUT_2[10011] = 32'b00000000000000000001111001010111;
assign LUT_2[10012] = 32'b11111111111111111010100101101010;
assign LUT_2[10013] = 32'b11111111111111110111011110000011;
assign LUT_2[10014] = 32'b00000000000000000001011110100110;
assign LUT_2[10015] = 32'b11111111111111111110010110111111;
assign LUT_2[10016] = 32'b00000000000000001001001110000100;
assign LUT_2[10017] = 32'b00000000000000000110000110011101;
assign LUT_2[10018] = 32'b00000000000000010000000111000000;
assign LUT_2[10019] = 32'b00000000000000001100111111011001;
assign LUT_2[10020] = 32'b00000000000000000101101011101100;
assign LUT_2[10021] = 32'b00000000000000000010100100000101;
assign LUT_2[10022] = 32'b00000000000000001100100100101000;
assign LUT_2[10023] = 32'b00000000000000001001011101000001;
assign LUT_2[10024] = 32'b00000000000000000011111111100001;
assign LUT_2[10025] = 32'b00000000000000000000110111111010;
assign LUT_2[10026] = 32'b00000000000000001010111000011101;
assign LUT_2[10027] = 32'b00000000000000000111110000110110;
assign LUT_2[10028] = 32'b00000000000000000000011101001001;
assign LUT_2[10029] = 32'b11111111111111111101010101100010;
assign LUT_2[10030] = 32'b00000000000000000111010110000101;
assign LUT_2[10031] = 32'b00000000000000000100001110011110;
assign LUT_2[10032] = 32'b00000000000000000011110010001110;
assign LUT_2[10033] = 32'b00000000000000000000101010100111;
assign LUT_2[10034] = 32'b00000000000000001010101011001010;
assign LUT_2[10035] = 32'b00000000000000000111100011100011;
assign LUT_2[10036] = 32'b00000000000000000000001111110110;
assign LUT_2[10037] = 32'b11111111111111111101001000001111;
assign LUT_2[10038] = 32'b00000000000000000111001000110010;
assign LUT_2[10039] = 32'b00000000000000000100000001001011;
assign LUT_2[10040] = 32'b11111111111111111110100011101011;
assign LUT_2[10041] = 32'b11111111111111111011011100000100;
assign LUT_2[10042] = 32'b00000000000000000101011100100111;
assign LUT_2[10043] = 32'b00000000000000000010010101000000;
assign LUT_2[10044] = 32'b11111111111111111011000001010011;
assign LUT_2[10045] = 32'b11111111111111110111111001101100;
assign LUT_2[10046] = 32'b00000000000000000001111010001111;
assign LUT_2[10047] = 32'b11111111111111111110110010101000;
assign LUT_2[10048] = 32'b00000000000000000000111010111110;
assign LUT_2[10049] = 32'b11111111111111111101110011010111;
assign LUT_2[10050] = 32'b00000000000000000111110011111010;
assign LUT_2[10051] = 32'b00000000000000000100101100010011;
assign LUT_2[10052] = 32'b11111111111111111101011000100110;
assign LUT_2[10053] = 32'b11111111111111111010010000111111;
assign LUT_2[10054] = 32'b00000000000000000100010001100010;
assign LUT_2[10055] = 32'b00000000000000000001001001111011;
assign LUT_2[10056] = 32'b11111111111111111011101100011011;
assign LUT_2[10057] = 32'b11111111111111111000100100110100;
assign LUT_2[10058] = 32'b00000000000000000010100101010111;
assign LUT_2[10059] = 32'b11111111111111111111011101110000;
assign LUT_2[10060] = 32'b11111111111111111000001010000011;
assign LUT_2[10061] = 32'b11111111111111110101000010011100;
assign LUT_2[10062] = 32'b11111111111111111111000010111111;
assign LUT_2[10063] = 32'b11111111111111111011111011011000;
assign LUT_2[10064] = 32'b11111111111111111011011111001000;
assign LUT_2[10065] = 32'b11111111111111111000010111100001;
assign LUT_2[10066] = 32'b00000000000000000010011000000100;
assign LUT_2[10067] = 32'b11111111111111111111010000011101;
assign LUT_2[10068] = 32'b11111111111111110111111100110000;
assign LUT_2[10069] = 32'b11111111111111110100110101001001;
assign LUT_2[10070] = 32'b11111111111111111110110101101100;
assign LUT_2[10071] = 32'b11111111111111111011101110000101;
assign LUT_2[10072] = 32'b11111111111111110110010000100101;
assign LUT_2[10073] = 32'b11111111111111110011001000111110;
assign LUT_2[10074] = 32'b11111111111111111101001001100001;
assign LUT_2[10075] = 32'b11111111111111111010000001111010;
assign LUT_2[10076] = 32'b11111111111111110010101110001101;
assign LUT_2[10077] = 32'b11111111111111101111100110100110;
assign LUT_2[10078] = 32'b11111111111111111001100111001001;
assign LUT_2[10079] = 32'b11111111111111110110011111100010;
assign LUT_2[10080] = 32'b00000000000000000001010110100111;
assign LUT_2[10081] = 32'b11111111111111111110001111000000;
assign LUT_2[10082] = 32'b00000000000000001000001111100011;
assign LUT_2[10083] = 32'b00000000000000000101000111111100;
assign LUT_2[10084] = 32'b11111111111111111101110100001111;
assign LUT_2[10085] = 32'b11111111111111111010101100101000;
assign LUT_2[10086] = 32'b00000000000000000100101101001011;
assign LUT_2[10087] = 32'b00000000000000000001100101100100;
assign LUT_2[10088] = 32'b11111111111111111100001000000100;
assign LUT_2[10089] = 32'b11111111111111111001000000011101;
assign LUT_2[10090] = 32'b00000000000000000011000001000000;
assign LUT_2[10091] = 32'b11111111111111111111111001011001;
assign LUT_2[10092] = 32'b11111111111111111000100101101100;
assign LUT_2[10093] = 32'b11111111111111110101011110000101;
assign LUT_2[10094] = 32'b11111111111111111111011110101000;
assign LUT_2[10095] = 32'b11111111111111111100010111000001;
assign LUT_2[10096] = 32'b11111111111111111011111010110001;
assign LUT_2[10097] = 32'b11111111111111111000110011001010;
assign LUT_2[10098] = 32'b00000000000000000010110011101101;
assign LUT_2[10099] = 32'b11111111111111111111101100000110;
assign LUT_2[10100] = 32'b11111111111111111000011000011001;
assign LUT_2[10101] = 32'b11111111111111110101010000110010;
assign LUT_2[10102] = 32'b11111111111111111111010001010101;
assign LUT_2[10103] = 32'b11111111111111111100001001101110;
assign LUT_2[10104] = 32'b11111111111111110110101100001110;
assign LUT_2[10105] = 32'b11111111111111110011100100100111;
assign LUT_2[10106] = 32'b11111111111111111101100101001010;
assign LUT_2[10107] = 32'b11111111111111111010011101100011;
assign LUT_2[10108] = 32'b11111111111111110011001001110110;
assign LUT_2[10109] = 32'b11111111111111110000000010001111;
assign LUT_2[10110] = 32'b11111111111111111010000010110010;
assign LUT_2[10111] = 32'b11111111111111110110111011001011;
assign LUT_2[10112] = 32'b00000000000000001101000110101010;
assign LUT_2[10113] = 32'b00000000000000001001111111000011;
assign LUT_2[10114] = 32'b00000000000000010011111111100110;
assign LUT_2[10115] = 32'b00000000000000010000110111111111;
assign LUT_2[10116] = 32'b00000000000000001001100100010010;
assign LUT_2[10117] = 32'b00000000000000000110011100101011;
assign LUT_2[10118] = 32'b00000000000000010000011101001110;
assign LUT_2[10119] = 32'b00000000000000001101010101100111;
assign LUT_2[10120] = 32'b00000000000000000111111000000111;
assign LUT_2[10121] = 32'b00000000000000000100110000100000;
assign LUT_2[10122] = 32'b00000000000000001110110001000011;
assign LUT_2[10123] = 32'b00000000000000001011101001011100;
assign LUT_2[10124] = 32'b00000000000000000100010101101111;
assign LUT_2[10125] = 32'b00000000000000000001001110001000;
assign LUT_2[10126] = 32'b00000000000000001011001110101011;
assign LUT_2[10127] = 32'b00000000000000001000000111000100;
assign LUT_2[10128] = 32'b00000000000000000111101010110100;
assign LUT_2[10129] = 32'b00000000000000000100100011001101;
assign LUT_2[10130] = 32'b00000000000000001110100011110000;
assign LUT_2[10131] = 32'b00000000000000001011011100001001;
assign LUT_2[10132] = 32'b00000000000000000100001000011100;
assign LUT_2[10133] = 32'b00000000000000000001000000110101;
assign LUT_2[10134] = 32'b00000000000000001011000001011000;
assign LUT_2[10135] = 32'b00000000000000000111111001110001;
assign LUT_2[10136] = 32'b00000000000000000010011100010001;
assign LUT_2[10137] = 32'b11111111111111111111010100101010;
assign LUT_2[10138] = 32'b00000000000000001001010101001101;
assign LUT_2[10139] = 32'b00000000000000000110001101100110;
assign LUT_2[10140] = 32'b11111111111111111110111001111001;
assign LUT_2[10141] = 32'b11111111111111111011110010010010;
assign LUT_2[10142] = 32'b00000000000000000101110010110101;
assign LUT_2[10143] = 32'b00000000000000000010101011001110;
assign LUT_2[10144] = 32'b00000000000000001101100010010011;
assign LUT_2[10145] = 32'b00000000000000001010011010101100;
assign LUT_2[10146] = 32'b00000000000000010100011011001111;
assign LUT_2[10147] = 32'b00000000000000010001010011101000;
assign LUT_2[10148] = 32'b00000000000000001001111111111011;
assign LUT_2[10149] = 32'b00000000000000000110111000010100;
assign LUT_2[10150] = 32'b00000000000000010000111000110111;
assign LUT_2[10151] = 32'b00000000000000001101110001010000;
assign LUT_2[10152] = 32'b00000000000000001000010011110000;
assign LUT_2[10153] = 32'b00000000000000000101001100001001;
assign LUT_2[10154] = 32'b00000000000000001111001100101100;
assign LUT_2[10155] = 32'b00000000000000001100000101000101;
assign LUT_2[10156] = 32'b00000000000000000100110001011000;
assign LUT_2[10157] = 32'b00000000000000000001101001110001;
assign LUT_2[10158] = 32'b00000000000000001011101010010100;
assign LUT_2[10159] = 32'b00000000000000001000100010101101;
assign LUT_2[10160] = 32'b00000000000000001000000110011101;
assign LUT_2[10161] = 32'b00000000000000000100111110110110;
assign LUT_2[10162] = 32'b00000000000000001110111111011001;
assign LUT_2[10163] = 32'b00000000000000001011110111110010;
assign LUT_2[10164] = 32'b00000000000000000100100100000101;
assign LUT_2[10165] = 32'b00000000000000000001011100011110;
assign LUT_2[10166] = 32'b00000000000000001011011101000001;
assign LUT_2[10167] = 32'b00000000000000001000010101011010;
assign LUT_2[10168] = 32'b00000000000000000010110111111010;
assign LUT_2[10169] = 32'b11111111111111111111110000010011;
assign LUT_2[10170] = 32'b00000000000000001001110000110110;
assign LUT_2[10171] = 32'b00000000000000000110101001001111;
assign LUT_2[10172] = 32'b11111111111111111111010101100010;
assign LUT_2[10173] = 32'b11111111111111111100001101111011;
assign LUT_2[10174] = 32'b00000000000000000110001110011110;
assign LUT_2[10175] = 32'b00000000000000000011000110110111;
assign LUT_2[10176] = 32'b00000000000000000101001111001101;
assign LUT_2[10177] = 32'b00000000000000000010000111100110;
assign LUT_2[10178] = 32'b00000000000000001100001000001001;
assign LUT_2[10179] = 32'b00000000000000001001000000100010;
assign LUT_2[10180] = 32'b00000000000000000001101100110101;
assign LUT_2[10181] = 32'b11111111111111111110100101001110;
assign LUT_2[10182] = 32'b00000000000000001000100101110001;
assign LUT_2[10183] = 32'b00000000000000000101011110001010;
assign LUT_2[10184] = 32'b00000000000000000000000000101010;
assign LUT_2[10185] = 32'b11111111111111111100111001000011;
assign LUT_2[10186] = 32'b00000000000000000110111001100110;
assign LUT_2[10187] = 32'b00000000000000000011110001111111;
assign LUT_2[10188] = 32'b11111111111111111100011110010010;
assign LUT_2[10189] = 32'b11111111111111111001010110101011;
assign LUT_2[10190] = 32'b00000000000000000011010111001110;
assign LUT_2[10191] = 32'b00000000000000000000001111100111;
assign LUT_2[10192] = 32'b11111111111111111111110011010111;
assign LUT_2[10193] = 32'b11111111111111111100101011110000;
assign LUT_2[10194] = 32'b00000000000000000110101100010011;
assign LUT_2[10195] = 32'b00000000000000000011100100101100;
assign LUT_2[10196] = 32'b11111111111111111100010000111111;
assign LUT_2[10197] = 32'b11111111111111111001001001011000;
assign LUT_2[10198] = 32'b00000000000000000011001001111011;
assign LUT_2[10199] = 32'b00000000000000000000000010010100;
assign LUT_2[10200] = 32'b11111111111111111010100100110100;
assign LUT_2[10201] = 32'b11111111111111110111011101001101;
assign LUT_2[10202] = 32'b00000000000000000001011101110000;
assign LUT_2[10203] = 32'b11111111111111111110010110001001;
assign LUT_2[10204] = 32'b11111111111111110111000010011100;
assign LUT_2[10205] = 32'b11111111111111110011111010110101;
assign LUT_2[10206] = 32'b11111111111111111101111011011000;
assign LUT_2[10207] = 32'b11111111111111111010110011110001;
assign LUT_2[10208] = 32'b00000000000000000101101010110110;
assign LUT_2[10209] = 32'b00000000000000000010100011001111;
assign LUT_2[10210] = 32'b00000000000000001100100011110010;
assign LUT_2[10211] = 32'b00000000000000001001011100001011;
assign LUT_2[10212] = 32'b00000000000000000010001000011110;
assign LUT_2[10213] = 32'b11111111111111111111000000110111;
assign LUT_2[10214] = 32'b00000000000000001001000001011010;
assign LUT_2[10215] = 32'b00000000000000000101111001110011;
assign LUT_2[10216] = 32'b00000000000000000000011100010011;
assign LUT_2[10217] = 32'b11111111111111111101010100101100;
assign LUT_2[10218] = 32'b00000000000000000111010101001111;
assign LUT_2[10219] = 32'b00000000000000000100001101101000;
assign LUT_2[10220] = 32'b11111111111111111100111001111011;
assign LUT_2[10221] = 32'b11111111111111111001110010010100;
assign LUT_2[10222] = 32'b00000000000000000011110010110111;
assign LUT_2[10223] = 32'b00000000000000000000101011010000;
assign LUT_2[10224] = 32'b00000000000000000000001111000000;
assign LUT_2[10225] = 32'b11111111111111111101000111011001;
assign LUT_2[10226] = 32'b00000000000000000111000111111100;
assign LUT_2[10227] = 32'b00000000000000000100000000010101;
assign LUT_2[10228] = 32'b11111111111111111100101100101000;
assign LUT_2[10229] = 32'b11111111111111111001100101000001;
assign LUT_2[10230] = 32'b00000000000000000011100101100100;
assign LUT_2[10231] = 32'b00000000000000000000011101111101;
assign LUT_2[10232] = 32'b11111111111111111011000000011101;
assign LUT_2[10233] = 32'b11111111111111110111111000110110;
assign LUT_2[10234] = 32'b00000000000000000001111001011001;
assign LUT_2[10235] = 32'b11111111111111111110110001110010;
assign LUT_2[10236] = 32'b11111111111111110111011110000101;
assign LUT_2[10237] = 32'b11111111111111110100010110011110;
assign LUT_2[10238] = 32'b11111111111111111110010111000001;
assign LUT_2[10239] = 32'b11111111111111111011001111011010;
assign LUT_2[10240] = 32'b11111111111111110101001011111010;
assign LUT_2[10241] = 32'b11111111111111110010000100010011;
assign LUT_2[10242] = 32'b11111111111111111100000100110110;
assign LUT_2[10243] = 32'b11111111111111111000111101001111;
assign LUT_2[10244] = 32'b11111111111111110001101001100010;
assign LUT_2[10245] = 32'b11111111111111101110100001111011;
assign LUT_2[10246] = 32'b11111111111111111000100010011110;
assign LUT_2[10247] = 32'b11111111111111110101011010110111;
assign LUT_2[10248] = 32'b11111111111111101111111101010111;
assign LUT_2[10249] = 32'b11111111111111101100110101110000;
assign LUT_2[10250] = 32'b11111111111111110110110110010011;
assign LUT_2[10251] = 32'b11111111111111110011101110101100;
assign LUT_2[10252] = 32'b11111111111111101100011010111111;
assign LUT_2[10253] = 32'b11111111111111101001010011011000;
assign LUT_2[10254] = 32'b11111111111111110011010011111011;
assign LUT_2[10255] = 32'b11111111111111110000001100010100;
assign LUT_2[10256] = 32'b11111111111111101111110000000100;
assign LUT_2[10257] = 32'b11111111111111101100101000011101;
assign LUT_2[10258] = 32'b11111111111111110110101001000000;
assign LUT_2[10259] = 32'b11111111111111110011100001011001;
assign LUT_2[10260] = 32'b11111111111111101100001101101100;
assign LUT_2[10261] = 32'b11111111111111101001000110000101;
assign LUT_2[10262] = 32'b11111111111111110011000110101000;
assign LUT_2[10263] = 32'b11111111111111101111111111000001;
assign LUT_2[10264] = 32'b11111111111111101010100001100001;
assign LUT_2[10265] = 32'b11111111111111100111011001111010;
assign LUT_2[10266] = 32'b11111111111111110001011010011101;
assign LUT_2[10267] = 32'b11111111111111101110010010110110;
assign LUT_2[10268] = 32'b11111111111111100110111111001001;
assign LUT_2[10269] = 32'b11111111111111100011110111100010;
assign LUT_2[10270] = 32'b11111111111111101101111000000101;
assign LUT_2[10271] = 32'b11111111111111101010110000011110;
assign LUT_2[10272] = 32'b11111111111111110101100111100011;
assign LUT_2[10273] = 32'b11111111111111110010011111111100;
assign LUT_2[10274] = 32'b11111111111111111100100000011111;
assign LUT_2[10275] = 32'b11111111111111111001011000111000;
assign LUT_2[10276] = 32'b11111111111111110010000101001011;
assign LUT_2[10277] = 32'b11111111111111101110111101100100;
assign LUT_2[10278] = 32'b11111111111111111000111110000111;
assign LUT_2[10279] = 32'b11111111111111110101110110100000;
assign LUT_2[10280] = 32'b11111111111111110000011001000000;
assign LUT_2[10281] = 32'b11111111111111101101010001011001;
assign LUT_2[10282] = 32'b11111111111111110111010001111100;
assign LUT_2[10283] = 32'b11111111111111110100001010010101;
assign LUT_2[10284] = 32'b11111111111111101100110110101000;
assign LUT_2[10285] = 32'b11111111111111101001101111000001;
assign LUT_2[10286] = 32'b11111111111111110011101111100100;
assign LUT_2[10287] = 32'b11111111111111110000100111111101;
assign LUT_2[10288] = 32'b11111111111111110000001011101101;
assign LUT_2[10289] = 32'b11111111111111101101000100000110;
assign LUT_2[10290] = 32'b11111111111111110111000100101001;
assign LUT_2[10291] = 32'b11111111111111110011111101000010;
assign LUT_2[10292] = 32'b11111111111111101100101001010101;
assign LUT_2[10293] = 32'b11111111111111101001100001101110;
assign LUT_2[10294] = 32'b11111111111111110011100010010001;
assign LUT_2[10295] = 32'b11111111111111110000011010101010;
assign LUT_2[10296] = 32'b11111111111111101010111101001010;
assign LUT_2[10297] = 32'b11111111111111100111110101100011;
assign LUT_2[10298] = 32'b11111111111111110001110110000110;
assign LUT_2[10299] = 32'b11111111111111101110101110011111;
assign LUT_2[10300] = 32'b11111111111111100111011010110010;
assign LUT_2[10301] = 32'b11111111111111100100010011001011;
assign LUT_2[10302] = 32'b11111111111111101110010011101110;
assign LUT_2[10303] = 32'b11111111111111101011001100000111;
assign LUT_2[10304] = 32'b11111111111111101101010100011101;
assign LUT_2[10305] = 32'b11111111111111101010001100110110;
assign LUT_2[10306] = 32'b11111111111111110100001101011001;
assign LUT_2[10307] = 32'b11111111111111110001000101110010;
assign LUT_2[10308] = 32'b11111111111111101001110010000101;
assign LUT_2[10309] = 32'b11111111111111100110101010011110;
assign LUT_2[10310] = 32'b11111111111111110000101011000001;
assign LUT_2[10311] = 32'b11111111111111101101100011011010;
assign LUT_2[10312] = 32'b11111111111111101000000101111010;
assign LUT_2[10313] = 32'b11111111111111100100111110010011;
assign LUT_2[10314] = 32'b11111111111111101110111110110110;
assign LUT_2[10315] = 32'b11111111111111101011110111001111;
assign LUT_2[10316] = 32'b11111111111111100100100011100010;
assign LUT_2[10317] = 32'b11111111111111100001011011111011;
assign LUT_2[10318] = 32'b11111111111111101011011100011110;
assign LUT_2[10319] = 32'b11111111111111101000010100110111;
assign LUT_2[10320] = 32'b11111111111111100111111000100111;
assign LUT_2[10321] = 32'b11111111111111100100110001000000;
assign LUT_2[10322] = 32'b11111111111111101110110001100011;
assign LUT_2[10323] = 32'b11111111111111101011101001111100;
assign LUT_2[10324] = 32'b11111111111111100100010110001111;
assign LUT_2[10325] = 32'b11111111111111100001001110101000;
assign LUT_2[10326] = 32'b11111111111111101011001111001011;
assign LUT_2[10327] = 32'b11111111111111101000000111100100;
assign LUT_2[10328] = 32'b11111111111111100010101010000100;
assign LUT_2[10329] = 32'b11111111111111011111100010011101;
assign LUT_2[10330] = 32'b11111111111111101001100011000000;
assign LUT_2[10331] = 32'b11111111111111100110011011011001;
assign LUT_2[10332] = 32'b11111111111111011111000111101100;
assign LUT_2[10333] = 32'b11111111111111011100000000000101;
assign LUT_2[10334] = 32'b11111111111111100110000000101000;
assign LUT_2[10335] = 32'b11111111111111100010111001000001;
assign LUT_2[10336] = 32'b11111111111111101101110000000110;
assign LUT_2[10337] = 32'b11111111111111101010101000011111;
assign LUT_2[10338] = 32'b11111111111111110100101001000010;
assign LUT_2[10339] = 32'b11111111111111110001100001011011;
assign LUT_2[10340] = 32'b11111111111111101010001101101110;
assign LUT_2[10341] = 32'b11111111111111100111000110000111;
assign LUT_2[10342] = 32'b11111111111111110001000110101010;
assign LUT_2[10343] = 32'b11111111111111101101111111000011;
assign LUT_2[10344] = 32'b11111111111111101000100001100011;
assign LUT_2[10345] = 32'b11111111111111100101011001111100;
assign LUT_2[10346] = 32'b11111111111111101111011010011111;
assign LUT_2[10347] = 32'b11111111111111101100010010111000;
assign LUT_2[10348] = 32'b11111111111111100100111111001011;
assign LUT_2[10349] = 32'b11111111111111100001110111100100;
assign LUT_2[10350] = 32'b11111111111111101011111000000111;
assign LUT_2[10351] = 32'b11111111111111101000110000100000;
assign LUT_2[10352] = 32'b11111111111111101000010100010000;
assign LUT_2[10353] = 32'b11111111111111100101001100101001;
assign LUT_2[10354] = 32'b11111111111111101111001101001100;
assign LUT_2[10355] = 32'b11111111111111101100000101100101;
assign LUT_2[10356] = 32'b11111111111111100100110001111000;
assign LUT_2[10357] = 32'b11111111111111100001101010010001;
assign LUT_2[10358] = 32'b11111111111111101011101010110100;
assign LUT_2[10359] = 32'b11111111111111101000100011001101;
assign LUT_2[10360] = 32'b11111111111111100011000101101101;
assign LUT_2[10361] = 32'b11111111111111011111111110000110;
assign LUT_2[10362] = 32'b11111111111111101001111110101001;
assign LUT_2[10363] = 32'b11111111111111100110110111000010;
assign LUT_2[10364] = 32'b11111111111111011111100011010101;
assign LUT_2[10365] = 32'b11111111111111011100011011101110;
assign LUT_2[10366] = 32'b11111111111111100110011100010001;
assign LUT_2[10367] = 32'b11111111111111100011010100101010;
assign LUT_2[10368] = 32'b11111111111111111001100000001001;
assign LUT_2[10369] = 32'b11111111111111110110011000100010;
assign LUT_2[10370] = 32'b00000000000000000000011001000101;
assign LUT_2[10371] = 32'b11111111111111111101010001011110;
assign LUT_2[10372] = 32'b11111111111111110101111101110001;
assign LUT_2[10373] = 32'b11111111111111110010110110001010;
assign LUT_2[10374] = 32'b11111111111111111100110110101101;
assign LUT_2[10375] = 32'b11111111111111111001101111000110;
assign LUT_2[10376] = 32'b11111111111111110100010001100110;
assign LUT_2[10377] = 32'b11111111111111110001001001111111;
assign LUT_2[10378] = 32'b11111111111111111011001010100010;
assign LUT_2[10379] = 32'b11111111111111111000000010111011;
assign LUT_2[10380] = 32'b11111111111111110000101111001110;
assign LUT_2[10381] = 32'b11111111111111101101100111100111;
assign LUT_2[10382] = 32'b11111111111111110111101000001010;
assign LUT_2[10383] = 32'b11111111111111110100100000100011;
assign LUT_2[10384] = 32'b11111111111111110100000100010011;
assign LUT_2[10385] = 32'b11111111111111110000111100101100;
assign LUT_2[10386] = 32'b11111111111111111010111101001111;
assign LUT_2[10387] = 32'b11111111111111110111110101101000;
assign LUT_2[10388] = 32'b11111111111111110000100001111011;
assign LUT_2[10389] = 32'b11111111111111101101011010010100;
assign LUT_2[10390] = 32'b11111111111111110111011010110111;
assign LUT_2[10391] = 32'b11111111111111110100010011010000;
assign LUT_2[10392] = 32'b11111111111111101110110101110000;
assign LUT_2[10393] = 32'b11111111111111101011101110001001;
assign LUT_2[10394] = 32'b11111111111111110101101110101100;
assign LUT_2[10395] = 32'b11111111111111110010100111000101;
assign LUT_2[10396] = 32'b11111111111111101011010011011000;
assign LUT_2[10397] = 32'b11111111111111101000001011110001;
assign LUT_2[10398] = 32'b11111111111111110010001100010100;
assign LUT_2[10399] = 32'b11111111111111101111000100101101;
assign LUT_2[10400] = 32'b11111111111111111001111011110010;
assign LUT_2[10401] = 32'b11111111111111110110110100001011;
assign LUT_2[10402] = 32'b00000000000000000000110100101110;
assign LUT_2[10403] = 32'b11111111111111111101101101000111;
assign LUT_2[10404] = 32'b11111111111111110110011001011010;
assign LUT_2[10405] = 32'b11111111111111110011010001110011;
assign LUT_2[10406] = 32'b11111111111111111101010010010110;
assign LUT_2[10407] = 32'b11111111111111111010001010101111;
assign LUT_2[10408] = 32'b11111111111111110100101101001111;
assign LUT_2[10409] = 32'b11111111111111110001100101101000;
assign LUT_2[10410] = 32'b11111111111111111011100110001011;
assign LUT_2[10411] = 32'b11111111111111111000011110100100;
assign LUT_2[10412] = 32'b11111111111111110001001010110111;
assign LUT_2[10413] = 32'b11111111111111101110000011010000;
assign LUT_2[10414] = 32'b11111111111111111000000011110011;
assign LUT_2[10415] = 32'b11111111111111110100111100001100;
assign LUT_2[10416] = 32'b11111111111111110100011111111100;
assign LUT_2[10417] = 32'b11111111111111110001011000010101;
assign LUT_2[10418] = 32'b11111111111111111011011000111000;
assign LUT_2[10419] = 32'b11111111111111111000010001010001;
assign LUT_2[10420] = 32'b11111111111111110000111101100100;
assign LUT_2[10421] = 32'b11111111111111101101110101111101;
assign LUT_2[10422] = 32'b11111111111111110111110110100000;
assign LUT_2[10423] = 32'b11111111111111110100101110111001;
assign LUT_2[10424] = 32'b11111111111111101111010001011001;
assign LUT_2[10425] = 32'b11111111111111101100001001110010;
assign LUT_2[10426] = 32'b11111111111111110110001010010101;
assign LUT_2[10427] = 32'b11111111111111110011000010101110;
assign LUT_2[10428] = 32'b11111111111111101011101111000001;
assign LUT_2[10429] = 32'b11111111111111101000100111011010;
assign LUT_2[10430] = 32'b11111111111111110010100111111101;
assign LUT_2[10431] = 32'b11111111111111101111100000010110;
assign LUT_2[10432] = 32'b11111111111111110001101000101100;
assign LUT_2[10433] = 32'b11111111111111101110100001000101;
assign LUT_2[10434] = 32'b11111111111111111000100001101000;
assign LUT_2[10435] = 32'b11111111111111110101011010000001;
assign LUT_2[10436] = 32'b11111111111111101110000110010100;
assign LUT_2[10437] = 32'b11111111111111101010111110101101;
assign LUT_2[10438] = 32'b11111111111111110100111111010000;
assign LUT_2[10439] = 32'b11111111111111110001110111101001;
assign LUT_2[10440] = 32'b11111111111111101100011010001001;
assign LUT_2[10441] = 32'b11111111111111101001010010100010;
assign LUT_2[10442] = 32'b11111111111111110011010011000101;
assign LUT_2[10443] = 32'b11111111111111110000001011011110;
assign LUT_2[10444] = 32'b11111111111111101000110111110001;
assign LUT_2[10445] = 32'b11111111111111100101110000001010;
assign LUT_2[10446] = 32'b11111111111111101111110000101101;
assign LUT_2[10447] = 32'b11111111111111101100101001000110;
assign LUT_2[10448] = 32'b11111111111111101100001100110110;
assign LUT_2[10449] = 32'b11111111111111101001000101001111;
assign LUT_2[10450] = 32'b11111111111111110011000101110010;
assign LUT_2[10451] = 32'b11111111111111101111111110001011;
assign LUT_2[10452] = 32'b11111111111111101000101010011110;
assign LUT_2[10453] = 32'b11111111111111100101100010110111;
assign LUT_2[10454] = 32'b11111111111111101111100011011010;
assign LUT_2[10455] = 32'b11111111111111101100011011110011;
assign LUT_2[10456] = 32'b11111111111111100110111110010011;
assign LUT_2[10457] = 32'b11111111111111100011110110101100;
assign LUT_2[10458] = 32'b11111111111111101101110111001111;
assign LUT_2[10459] = 32'b11111111111111101010101111101000;
assign LUT_2[10460] = 32'b11111111111111100011011011111011;
assign LUT_2[10461] = 32'b11111111111111100000010100010100;
assign LUT_2[10462] = 32'b11111111111111101010010100110111;
assign LUT_2[10463] = 32'b11111111111111100111001101010000;
assign LUT_2[10464] = 32'b11111111111111110010000100010101;
assign LUT_2[10465] = 32'b11111111111111101110111100101110;
assign LUT_2[10466] = 32'b11111111111111111000111101010001;
assign LUT_2[10467] = 32'b11111111111111110101110101101010;
assign LUT_2[10468] = 32'b11111111111111101110100001111101;
assign LUT_2[10469] = 32'b11111111111111101011011010010110;
assign LUT_2[10470] = 32'b11111111111111110101011010111001;
assign LUT_2[10471] = 32'b11111111111111110010010011010010;
assign LUT_2[10472] = 32'b11111111111111101100110101110010;
assign LUT_2[10473] = 32'b11111111111111101001101110001011;
assign LUT_2[10474] = 32'b11111111111111110011101110101110;
assign LUT_2[10475] = 32'b11111111111111110000100111000111;
assign LUT_2[10476] = 32'b11111111111111101001010011011010;
assign LUT_2[10477] = 32'b11111111111111100110001011110011;
assign LUT_2[10478] = 32'b11111111111111110000001100010110;
assign LUT_2[10479] = 32'b11111111111111101101000100101111;
assign LUT_2[10480] = 32'b11111111111111101100101000011111;
assign LUT_2[10481] = 32'b11111111111111101001100000111000;
assign LUT_2[10482] = 32'b11111111111111110011100001011011;
assign LUT_2[10483] = 32'b11111111111111110000011001110100;
assign LUT_2[10484] = 32'b11111111111111101001000110000111;
assign LUT_2[10485] = 32'b11111111111111100101111110100000;
assign LUT_2[10486] = 32'b11111111111111101111111111000011;
assign LUT_2[10487] = 32'b11111111111111101100110111011100;
assign LUT_2[10488] = 32'b11111111111111100111011001111100;
assign LUT_2[10489] = 32'b11111111111111100100010010010101;
assign LUT_2[10490] = 32'b11111111111111101110010010111000;
assign LUT_2[10491] = 32'b11111111111111101011001011010001;
assign LUT_2[10492] = 32'b11111111111111100011110111100100;
assign LUT_2[10493] = 32'b11111111111111100000101111111101;
assign LUT_2[10494] = 32'b11111111111111101010110000100000;
assign LUT_2[10495] = 32'b11111111111111100111101000111001;
assign LUT_2[10496] = 32'b11111111111111111001001010100000;
assign LUT_2[10497] = 32'b11111111111111110110000010111001;
assign LUT_2[10498] = 32'b00000000000000000000000011011100;
assign LUT_2[10499] = 32'b11111111111111111100111011110101;
assign LUT_2[10500] = 32'b11111111111111110101101000001000;
assign LUT_2[10501] = 32'b11111111111111110010100000100001;
assign LUT_2[10502] = 32'b11111111111111111100100001000100;
assign LUT_2[10503] = 32'b11111111111111111001011001011101;
assign LUT_2[10504] = 32'b11111111111111110011111011111101;
assign LUT_2[10505] = 32'b11111111111111110000110100010110;
assign LUT_2[10506] = 32'b11111111111111111010110100111001;
assign LUT_2[10507] = 32'b11111111111111110111101101010010;
assign LUT_2[10508] = 32'b11111111111111110000011001100101;
assign LUT_2[10509] = 32'b11111111111111101101010001111110;
assign LUT_2[10510] = 32'b11111111111111110111010010100001;
assign LUT_2[10511] = 32'b11111111111111110100001010111010;
assign LUT_2[10512] = 32'b11111111111111110011101110101010;
assign LUT_2[10513] = 32'b11111111111111110000100111000011;
assign LUT_2[10514] = 32'b11111111111111111010100111100110;
assign LUT_2[10515] = 32'b11111111111111110111011111111111;
assign LUT_2[10516] = 32'b11111111111111110000001100010010;
assign LUT_2[10517] = 32'b11111111111111101101000100101011;
assign LUT_2[10518] = 32'b11111111111111110111000101001110;
assign LUT_2[10519] = 32'b11111111111111110011111101100111;
assign LUT_2[10520] = 32'b11111111111111101110100000000111;
assign LUT_2[10521] = 32'b11111111111111101011011000100000;
assign LUT_2[10522] = 32'b11111111111111110101011001000011;
assign LUT_2[10523] = 32'b11111111111111110010010001011100;
assign LUT_2[10524] = 32'b11111111111111101010111101101111;
assign LUT_2[10525] = 32'b11111111111111100111110110001000;
assign LUT_2[10526] = 32'b11111111111111110001110110101011;
assign LUT_2[10527] = 32'b11111111111111101110101111000100;
assign LUT_2[10528] = 32'b11111111111111111001100110001001;
assign LUT_2[10529] = 32'b11111111111111110110011110100010;
assign LUT_2[10530] = 32'b00000000000000000000011111000101;
assign LUT_2[10531] = 32'b11111111111111111101010111011110;
assign LUT_2[10532] = 32'b11111111111111110110000011110001;
assign LUT_2[10533] = 32'b11111111111111110010111100001010;
assign LUT_2[10534] = 32'b11111111111111111100111100101101;
assign LUT_2[10535] = 32'b11111111111111111001110101000110;
assign LUT_2[10536] = 32'b11111111111111110100010111100110;
assign LUT_2[10537] = 32'b11111111111111110001001111111111;
assign LUT_2[10538] = 32'b11111111111111111011010000100010;
assign LUT_2[10539] = 32'b11111111111111111000001000111011;
assign LUT_2[10540] = 32'b11111111111111110000110101001110;
assign LUT_2[10541] = 32'b11111111111111101101101101100111;
assign LUT_2[10542] = 32'b11111111111111110111101110001010;
assign LUT_2[10543] = 32'b11111111111111110100100110100011;
assign LUT_2[10544] = 32'b11111111111111110100001010010011;
assign LUT_2[10545] = 32'b11111111111111110001000010101100;
assign LUT_2[10546] = 32'b11111111111111111011000011001111;
assign LUT_2[10547] = 32'b11111111111111110111111011101000;
assign LUT_2[10548] = 32'b11111111111111110000100111111011;
assign LUT_2[10549] = 32'b11111111111111101101100000010100;
assign LUT_2[10550] = 32'b11111111111111110111100000110111;
assign LUT_2[10551] = 32'b11111111111111110100011001010000;
assign LUT_2[10552] = 32'b11111111111111101110111011110000;
assign LUT_2[10553] = 32'b11111111111111101011110100001001;
assign LUT_2[10554] = 32'b11111111111111110101110100101100;
assign LUT_2[10555] = 32'b11111111111111110010101101000101;
assign LUT_2[10556] = 32'b11111111111111101011011001011000;
assign LUT_2[10557] = 32'b11111111111111101000010001110001;
assign LUT_2[10558] = 32'b11111111111111110010010010010100;
assign LUT_2[10559] = 32'b11111111111111101111001010101101;
assign LUT_2[10560] = 32'b11111111111111110001010011000011;
assign LUT_2[10561] = 32'b11111111111111101110001011011100;
assign LUT_2[10562] = 32'b11111111111111111000001011111111;
assign LUT_2[10563] = 32'b11111111111111110101000100011000;
assign LUT_2[10564] = 32'b11111111111111101101110000101011;
assign LUT_2[10565] = 32'b11111111111111101010101001000100;
assign LUT_2[10566] = 32'b11111111111111110100101001100111;
assign LUT_2[10567] = 32'b11111111111111110001100010000000;
assign LUT_2[10568] = 32'b11111111111111101100000100100000;
assign LUT_2[10569] = 32'b11111111111111101000111100111001;
assign LUT_2[10570] = 32'b11111111111111110010111101011100;
assign LUT_2[10571] = 32'b11111111111111101111110101110101;
assign LUT_2[10572] = 32'b11111111111111101000100010001000;
assign LUT_2[10573] = 32'b11111111111111100101011010100001;
assign LUT_2[10574] = 32'b11111111111111101111011011000100;
assign LUT_2[10575] = 32'b11111111111111101100010011011101;
assign LUT_2[10576] = 32'b11111111111111101011110111001101;
assign LUT_2[10577] = 32'b11111111111111101000101111100110;
assign LUT_2[10578] = 32'b11111111111111110010110000001001;
assign LUT_2[10579] = 32'b11111111111111101111101000100010;
assign LUT_2[10580] = 32'b11111111111111101000010100110101;
assign LUT_2[10581] = 32'b11111111111111100101001101001110;
assign LUT_2[10582] = 32'b11111111111111101111001101110001;
assign LUT_2[10583] = 32'b11111111111111101100000110001010;
assign LUT_2[10584] = 32'b11111111111111100110101000101010;
assign LUT_2[10585] = 32'b11111111111111100011100001000011;
assign LUT_2[10586] = 32'b11111111111111101101100001100110;
assign LUT_2[10587] = 32'b11111111111111101010011001111111;
assign LUT_2[10588] = 32'b11111111111111100011000110010010;
assign LUT_2[10589] = 32'b11111111111111011111111110101011;
assign LUT_2[10590] = 32'b11111111111111101001111111001110;
assign LUT_2[10591] = 32'b11111111111111100110110111100111;
assign LUT_2[10592] = 32'b11111111111111110001101110101100;
assign LUT_2[10593] = 32'b11111111111111101110100111000101;
assign LUT_2[10594] = 32'b11111111111111111000100111101000;
assign LUT_2[10595] = 32'b11111111111111110101100000000001;
assign LUT_2[10596] = 32'b11111111111111101110001100010100;
assign LUT_2[10597] = 32'b11111111111111101011000100101101;
assign LUT_2[10598] = 32'b11111111111111110101000101010000;
assign LUT_2[10599] = 32'b11111111111111110001111101101001;
assign LUT_2[10600] = 32'b11111111111111101100100000001001;
assign LUT_2[10601] = 32'b11111111111111101001011000100010;
assign LUT_2[10602] = 32'b11111111111111110011011001000101;
assign LUT_2[10603] = 32'b11111111111111110000010001011110;
assign LUT_2[10604] = 32'b11111111111111101000111101110001;
assign LUT_2[10605] = 32'b11111111111111100101110110001010;
assign LUT_2[10606] = 32'b11111111111111101111110110101101;
assign LUT_2[10607] = 32'b11111111111111101100101111000110;
assign LUT_2[10608] = 32'b11111111111111101100010010110110;
assign LUT_2[10609] = 32'b11111111111111101001001011001111;
assign LUT_2[10610] = 32'b11111111111111110011001011110010;
assign LUT_2[10611] = 32'b11111111111111110000000100001011;
assign LUT_2[10612] = 32'b11111111111111101000110000011110;
assign LUT_2[10613] = 32'b11111111111111100101101000110111;
assign LUT_2[10614] = 32'b11111111111111101111101001011010;
assign LUT_2[10615] = 32'b11111111111111101100100001110011;
assign LUT_2[10616] = 32'b11111111111111100111000100010011;
assign LUT_2[10617] = 32'b11111111111111100011111100101100;
assign LUT_2[10618] = 32'b11111111111111101101111101001111;
assign LUT_2[10619] = 32'b11111111111111101010110101101000;
assign LUT_2[10620] = 32'b11111111111111100011100001111011;
assign LUT_2[10621] = 32'b11111111111111100000011010010100;
assign LUT_2[10622] = 32'b11111111111111101010011010110111;
assign LUT_2[10623] = 32'b11111111111111100111010011010000;
assign LUT_2[10624] = 32'b11111111111111111101011110101111;
assign LUT_2[10625] = 32'b11111111111111111010010111001000;
assign LUT_2[10626] = 32'b00000000000000000100010111101011;
assign LUT_2[10627] = 32'b00000000000000000001010000000100;
assign LUT_2[10628] = 32'b11111111111111111001111100010111;
assign LUT_2[10629] = 32'b11111111111111110110110100110000;
assign LUT_2[10630] = 32'b00000000000000000000110101010011;
assign LUT_2[10631] = 32'b11111111111111111101101101101100;
assign LUT_2[10632] = 32'b11111111111111111000010000001100;
assign LUT_2[10633] = 32'b11111111111111110101001000100101;
assign LUT_2[10634] = 32'b11111111111111111111001001001000;
assign LUT_2[10635] = 32'b11111111111111111100000001100001;
assign LUT_2[10636] = 32'b11111111111111110100101101110100;
assign LUT_2[10637] = 32'b11111111111111110001100110001101;
assign LUT_2[10638] = 32'b11111111111111111011100110110000;
assign LUT_2[10639] = 32'b11111111111111111000011111001001;
assign LUT_2[10640] = 32'b11111111111111111000000010111001;
assign LUT_2[10641] = 32'b11111111111111110100111011010010;
assign LUT_2[10642] = 32'b11111111111111111110111011110101;
assign LUT_2[10643] = 32'b11111111111111111011110100001110;
assign LUT_2[10644] = 32'b11111111111111110100100000100001;
assign LUT_2[10645] = 32'b11111111111111110001011000111010;
assign LUT_2[10646] = 32'b11111111111111111011011001011101;
assign LUT_2[10647] = 32'b11111111111111111000010001110110;
assign LUT_2[10648] = 32'b11111111111111110010110100010110;
assign LUT_2[10649] = 32'b11111111111111101111101100101111;
assign LUT_2[10650] = 32'b11111111111111111001101101010010;
assign LUT_2[10651] = 32'b11111111111111110110100101101011;
assign LUT_2[10652] = 32'b11111111111111101111010001111110;
assign LUT_2[10653] = 32'b11111111111111101100001010010111;
assign LUT_2[10654] = 32'b11111111111111110110001010111010;
assign LUT_2[10655] = 32'b11111111111111110011000011010011;
assign LUT_2[10656] = 32'b11111111111111111101111010011000;
assign LUT_2[10657] = 32'b11111111111111111010110010110001;
assign LUT_2[10658] = 32'b00000000000000000100110011010100;
assign LUT_2[10659] = 32'b00000000000000000001101011101101;
assign LUT_2[10660] = 32'b11111111111111111010011000000000;
assign LUT_2[10661] = 32'b11111111111111110111010000011001;
assign LUT_2[10662] = 32'b00000000000000000001010000111100;
assign LUT_2[10663] = 32'b11111111111111111110001001010101;
assign LUT_2[10664] = 32'b11111111111111111000101011110101;
assign LUT_2[10665] = 32'b11111111111111110101100100001110;
assign LUT_2[10666] = 32'b11111111111111111111100100110001;
assign LUT_2[10667] = 32'b11111111111111111100011101001010;
assign LUT_2[10668] = 32'b11111111111111110101001001011101;
assign LUT_2[10669] = 32'b11111111111111110010000001110110;
assign LUT_2[10670] = 32'b11111111111111111100000010011001;
assign LUT_2[10671] = 32'b11111111111111111000111010110010;
assign LUT_2[10672] = 32'b11111111111111111000011110100010;
assign LUT_2[10673] = 32'b11111111111111110101010110111011;
assign LUT_2[10674] = 32'b11111111111111111111010111011110;
assign LUT_2[10675] = 32'b11111111111111111100001111110111;
assign LUT_2[10676] = 32'b11111111111111110100111100001010;
assign LUT_2[10677] = 32'b11111111111111110001110100100011;
assign LUT_2[10678] = 32'b11111111111111111011110101000110;
assign LUT_2[10679] = 32'b11111111111111111000101101011111;
assign LUT_2[10680] = 32'b11111111111111110011001111111111;
assign LUT_2[10681] = 32'b11111111111111110000001000011000;
assign LUT_2[10682] = 32'b11111111111111111010001000111011;
assign LUT_2[10683] = 32'b11111111111111110111000001010100;
assign LUT_2[10684] = 32'b11111111111111101111101101100111;
assign LUT_2[10685] = 32'b11111111111111101100100110000000;
assign LUT_2[10686] = 32'b11111111111111110110100110100011;
assign LUT_2[10687] = 32'b11111111111111110011011110111100;
assign LUT_2[10688] = 32'b11111111111111110101100111010010;
assign LUT_2[10689] = 32'b11111111111111110010011111101011;
assign LUT_2[10690] = 32'b11111111111111111100100000001110;
assign LUT_2[10691] = 32'b11111111111111111001011000100111;
assign LUT_2[10692] = 32'b11111111111111110010000100111010;
assign LUT_2[10693] = 32'b11111111111111101110111101010011;
assign LUT_2[10694] = 32'b11111111111111111000111101110110;
assign LUT_2[10695] = 32'b11111111111111110101110110001111;
assign LUT_2[10696] = 32'b11111111111111110000011000101111;
assign LUT_2[10697] = 32'b11111111111111101101010001001000;
assign LUT_2[10698] = 32'b11111111111111110111010001101011;
assign LUT_2[10699] = 32'b11111111111111110100001010000100;
assign LUT_2[10700] = 32'b11111111111111101100110110010111;
assign LUT_2[10701] = 32'b11111111111111101001101110110000;
assign LUT_2[10702] = 32'b11111111111111110011101111010011;
assign LUT_2[10703] = 32'b11111111111111110000100111101100;
assign LUT_2[10704] = 32'b11111111111111110000001011011100;
assign LUT_2[10705] = 32'b11111111111111101101000011110101;
assign LUT_2[10706] = 32'b11111111111111110111000100011000;
assign LUT_2[10707] = 32'b11111111111111110011111100110001;
assign LUT_2[10708] = 32'b11111111111111101100101001000100;
assign LUT_2[10709] = 32'b11111111111111101001100001011101;
assign LUT_2[10710] = 32'b11111111111111110011100010000000;
assign LUT_2[10711] = 32'b11111111111111110000011010011001;
assign LUT_2[10712] = 32'b11111111111111101010111100111001;
assign LUT_2[10713] = 32'b11111111111111100111110101010010;
assign LUT_2[10714] = 32'b11111111111111110001110101110101;
assign LUT_2[10715] = 32'b11111111111111101110101110001110;
assign LUT_2[10716] = 32'b11111111111111100111011010100001;
assign LUT_2[10717] = 32'b11111111111111100100010010111010;
assign LUT_2[10718] = 32'b11111111111111101110010011011101;
assign LUT_2[10719] = 32'b11111111111111101011001011110110;
assign LUT_2[10720] = 32'b11111111111111110110000010111011;
assign LUT_2[10721] = 32'b11111111111111110010111011010100;
assign LUT_2[10722] = 32'b11111111111111111100111011110111;
assign LUT_2[10723] = 32'b11111111111111111001110100010000;
assign LUT_2[10724] = 32'b11111111111111110010100000100011;
assign LUT_2[10725] = 32'b11111111111111101111011000111100;
assign LUT_2[10726] = 32'b11111111111111111001011001011111;
assign LUT_2[10727] = 32'b11111111111111110110010001111000;
assign LUT_2[10728] = 32'b11111111111111110000110100011000;
assign LUT_2[10729] = 32'b11111111111111101101101100110001;
assign LUT_2[10730] = 32'b11111111111111110111101101010100;
assign LUT_2[10731] = 32'b11111111111111110100100101101101;
assign LUT_2[10732] = 32'b11111111111111101101010010000000;
assign LUT_2[10733] = 32'b11111111111111101010001010011001;
assign LUT_2[10734] = 32'b11111111111111110100001010111100;
assign LUT_2[10735] = 32'b11111111111111110001000011010101;
assign LUT_2[10736] = 32'b11111111111111110000100111000101;
assign LUT_2[10737] = 32'b11111111111111101101011111011110;
assign LUT_2[10738] = 32'b11111111111111110111100000000001;
assign LUT_2[10739] = 32'b11111111111111110100011000011010;
assign LUT_2[10740] = 32'b11111111111111101101000100101101;
assign LUT_2[10741] = 32'b11111111111111101001111101000110;
assign LUT_2[10742] = 32'b11111111111111110011111101101001;
assign LUT_2[10743] = 32'b11111111111111110000110110000010;
assign LUT_2[10744] = 32'b11111111111111101011011000100010;
assign LUT_2[10745] = 32'b11111111111111101000010000111011;
assign LUT_2[10746] = 32'b11111111111111110010010001011110;
assign LUT_2[10747] = 32'b11111111111111101111001001110111;
assign LUT_2[10748] = 32'b11111111111111100111110110001010;
assign LUT_2[10749] = 32'b11111111111111100100101110100011;
assign LUT_2[10750] = 32'b11111111111111101110101111000110;
assign LUT_2[10751] = 32'b11111111111111101011100111011111;
assign LUT_2[10752] = 32'b11111111111111111001111101101100;
assign LUT_2[10753] = 32'b11111111111111110110110110000101;
assign LUT_2[10754] = 32'b00000000000000000000110110101000;
assign LUT_2[10755] = 32'b11111111111111111101101111000001;
assign LUT_2[10756] = 32'b11111111111111110110011011010100;
assign LUT_2[10757] = 32'b11111111111111110011010011101101;
assign LUT_2[10758] = 32'b11111111111111111101010100010000;
assign LUT_2[10759] = 32'b11111111111111111010001100101001;
assign LUT_2[10760] = 32'b11111111111111110100101111001001;
assign LUT_2[10761] = 32'b11111111111111110001100111100010;
assign LUT_2[10762] = 32'b11111111111111111011101000000101;
assign LUT_2[10763] = 32'b11111111111111111000100000011110;
assign LUT_2[10764] = 32'b11111111111111110001001100110001;
assign LUT_2[10765] = 32'b11111111111111101110000101001010;
assign LUT_2[10766] = 32'b11111111111111111000000101101101;
assign LUT_2[10767] = 32'b11111111111111110100111110000110;
assign LUT_2[10768] = 32'b11111111111111110100100001110110;
assign LUT_2[10769] = 32'b11111111111111110001011010001111;
assign LUT_2[10770] = 32'b11111111111111111011011010110010;
assign LUT_2[10771] = 32'b11111111111111111000010011001011;
assign LUT_2[10772] = 32'b11111111111111110000111111011110;
assign LUT_2[10773] = 32'b11111111111111101101110111110111;
assign LUT_2[10774] = 32'b11111111111111110111111000011010;
assign LUT_2[10775] = 32'b11111111111111110100110000110011;
assign LUT_2[10776] = 32'b11111111111111101111010011010011;
assign LUT_2[10777] = 32'b11111111111111101100001011101100;
assign LUT_2[10778] = 32'b11111111111111110110001100001111;
assign LUT_2[10779] = 32'b11111111111111110011000100101000;
assign LUT_2[10780] = 32'b11111111111111101011110000111011;
assign LUT_2[10781] = 32'b11111111111111101000101001010100;
assign LUT_2[10782] = 32'b11111111111111110010101001110111;
assign LUT_2[10783] = 32'b11111111111111101111100010010000;
assign LUT_2[10784] = 32'b11111111111111111010011001010101;
assign LUT_2[10785] = 32'b11111111111111110111010001101110;
assign LUT_2[10786] = 32'b00000000000000000001010010010001;
assign LUT_2[10787] = 32'b11111111111111111110001010101010;
assign LUT_2[10788] = 32'b11111111111111110110110110111101;
assign LUT_2[10789] = 32'b11111111111111110011101111010110;
assign LUT_2[10790] = 32'b11111111111111111101101111111001;
assign LUT_2[10791] = 32'b11111111111111111010101000010010;
assign LUT_2[10792] = 32'b11111111111111110101001010110010;
assign LUT_2[10793] = 32'b11111111111111110010000011001011;
assign LUT_2[10794] = 32'b11111111111111111100000011101110;
assign LUT_2[10795] = 32'b11111111111111111000111100000111;
assign LUT_2[10796] = 32'b11111111111111110001101000011010;
assign LUT_2[10797] = 32'b11111111111111101110100000110011;
assign LUT_2[10798] = 32'b11111111111111111000100001010110;
assign LUT_2[10799] = 32'b11111111111111110101011001101111;
assign LUT_2[10800] = 32'b11111111111111110100111101011111;
assign LUT_2[10801] = 32'b11111111111111110001110101111000;
assign LUT_2[10802] = 32'b11111111111111111011110110011011;
assign LUT_2[10803] = 32'b11111111111111111000101110110100;
assign LUT_2[10804] = 32'b11111111111111110001011011000111;
assign LUT_2[10805] = 32'b11111111111111101110010011100000;
assign LUT_2[10806] = 32'b11111111111111111000010100000011;
assign LUT_2[10807] = 32'b11111111111111110101001100011100;
assign LUT_2[10808] = 32'b11111111111111101111101110111100;
assign LUT_2[10809] = 32'b11111111111111101100100111010101;
assign LUT_2[10810] = 32'b11111111111111110110100111111000;
assign LUT_2[10811] = 32'b11111111111111110011100000010001;
assign LUT_2[10812] = 32'b11111111111111101100001100100100;
assign LUT_2[10813] = 32'b11111111111111101001000100111101;
assign LUT_2[10814] = 32'b11111111111111110011000101100000;
assign LUT_2[10815] = 32'b11111111111111101111111101111001;
assign LUT_2[10816] = 32'b11111111111111110010000110001111;
assign LUT_2[10817] = 32'b11111111111111101110111110101000;
assign LUT_2[10818] = 32'b11111111111111111000111111001011;
assign LUT_2[10819] = 32'b11111111111111110101110111100100;
assign LUT_2[10820] = 32'b11111111111111101110100011110111;
assign LUT_2[10821] = 32'b11111111111111101011011100010000;
assign LUT_2[10822] = 32'b11111111111111110101011100110011;
assign LUT_2[10823] = 32'b11111111111111110010010101001100;
assign LUT_2[10824] = 32'b11111111111111101100110111101100;
assign LUT_2[10825] = 32'b11111111111111101001110000000101;
assign LUT_2[10826] = 32'b11111111111111110011110000101000;
assign LUT_2[10827] = 32'b11111111111111110000101001000001;
assign LUT_2[10828] = 32'b11111111111111101001010101010100;
assign LUT_2[10829] = 32'b11111111111111100110001101101101;
assign LUT_2[10830] = 32'b11111111111111110000001110010000;
assign LUT_2[10831] = 32'b11111111111111101101000110101001;
assign LUT_2[10832] = 32'b11111111111111101100101010011001;
assign LUT_2[10833] = 32'b11111111111111101001100010110010;
assign LUT_2[10834] = 32'b11111111111111110011100011010101;
assign LUT_2[10835] = 32'b11111111111111110000011011101110;
assign LUT_2[10836] = 32'b11111111111111101001001000000001;
assign LUT_2[10837] = 32'b11111111111111100110000000011010;
assign LUT_2[10838] = 32'b11111111111111110000000000111101;
assign LUT_2[10839] = 32'b11111111111111101100111001010110;
assign LUT_2[10840] = 32'b11111111111111100111011011110110;
assign LUT_2[10841] = 32'b11111111111111100100010100001111;
assign LUT_2[10842] = 32'b11111111111111101110010100110010;
assign LUT_2[10843] = 32'b11111111111111101011001101001011;
assign LUT_2[10844] = 32'b11111111111111100011111001011110;
assign LUT_2[10845] = 32'b11111111111111100000110001110111;
assign LUT_2[10846] = 32'b11111111111111101010110010011010;
assign LUT_2[10847] = 32'b11111111111111100111101010110011;
assign LUT_2[10848] = 32'b11111111111111110010100001111000;
assign LUT_2[10849] = 32'b11111111111111101111011010010001;
assign LUT_2[10850] = 32'b11111111111111111001011010110100;
assign LUT_2[10851] = 32'b11111111111111110110010011001101;
assign LUT_2[10852] = 32'b11111111111111101110111111100000;
assign LUT_2[10853] = 32'b11111111111111101011110111111001;
assign LUT_2[10854] = 32'b11111111111111110101111000011100;
assign LUT_2[10855] = 32'b11111111111111110010110000110101;
assign LUT_2[10856] = 32'b11111111111111101101010011010101;
assign LUT_2[10857] = 32'b11111111111111101010001011101110;
assign LUT_2[10858] = 32'b11111111111111110100001100010001;
assign LUT_2[10859] = 32'b11111111111111110001000100101010;
assign LUT_2[10860] = 32'b11111111111111101001110000111101;
assign LUT_2[10861] = 32'b11111111111111100110101001010110;
assign LUT_2[10862] = 32'b11111111111111110000101001111001;
assign LUT_2[10863] = 32'b11111111111111101101100010010010;
assign LUT_2[10864] = 32'b11111111111111101101000110000010;
assign LUT_2[10865] = 32'b11111111111111101001111110011011;
assign LUT_2[10866] = 32'b11111111111111110011111110111110;
assign LUT_2[10867] = 32'b11111111111111110000110111010111;
assign LUT_2[10868] = 32'b11111111111111101001100011101010;
assign LUT_2[10869] = 32'b11111111111111100110011100000011;
assign LUT_2[10870] = 32'b11111111111111110000011100100110;
assign LUT_2[10871] = 32'b11111111111111101101010100111111;
assign LUT_2[10872] = 32'b11111111111111100111110111011111;
assign LUT_2[10873] = 32'b11111111111111100100101111111000;
assign LUT_2[10874] = 32'b11111111111111101110110000011011;
assign LUT_2[10875] = 32'b11111111111111101011101000110100;
assign LUT_2[10876] = 32'b11111111111111100100010101000111;
assign LUT_2[10877] = 32'b11111111111111100001001101100000;
assign LUT_2[10878] = 32'b11111111111111101011001110000011;
assign LUT_2[10879] = 32'b11111111111111101000000110011100;
assign LUT_2[10880] = 32'b11111111111111111110010001111011;
assign LUT_2[10881] = 32'b11111111111111111011001010010100;
assign LUT_2[10882] = 32'b00000000000000000101001010110111;
assign LUT_2[10883] = 32'b00000000000000000010000011010000;
assign LUT_2[10884] = 32'b11111111111111111010101111100011;
assign LUT_2[10885] = 32'b11111111111111110111100111111100;
assign LUT_2[10886] = 32'b00000000000000000001101000011111;
assign LUT_2[10887] = 32'b11111111111111111110100000111000;
assign LUT_2[10888] = 32'b11111111111111111001000011011000;
assign LUT_2[10889] = 32'b11111111111111110101111011110001;
assign LUT_2[10890] = 32'b11111111111111111111111100010100;
assign LUT_2[10891] = 32'b11111111111111111100110100101101;
assign LUT_2[10892] = 32'b11111111111111110101100001000000;
assign LUT_2[10893] = 32'b11111111111111110010011001011001;
assign LUT_2[10894] = 32'b11111111111111111100011001111100;
assign LUT_2[10895] = 32'b11111111111111111001010010010101;
assign LUT_2[10896] = 32'b11111111111111111000110110000101;
assign LUT_2[10897] = 32'b11111111111111110101101110011110;
assign LUT_2[10898] = 32'b11111111111111111111101111000001;
assign LUT_2[10899] = 32'b11111111111111111100100111011010;
assign LUT_2[10900] = 32'b11111111111111110101010011101101;
assign LUT_2[10901] = 32'b11111111111111110010001100000110;
assign LUT_2[10902] = 32'b11111111111111111100001100101001;
assign LUT_2[10903] = 32'b11111111111111111001000101000010;
assign LUT_2[10904] = 32'b11111111111111110011100111100010;
assign LUT_2[10905] = 32'b11111111111111110000011111111011;
assign LUT_2[10906] = 32'b11111111111111111010100000011110;
assign LUT_2[10907] = 32'b11111111111111110111011000110111;
assign LUT_2[10908] = 32'b11111111111111110000000101001010;
assign LUT_2[10909] = 32'b11111111111111101100111101100011;
assign LUT_2[10910] = 32'b11111111111111110110111110000110;
assign LUT_2[10911] = 32'b11111111111111110011110110011111;
assign LUT_2[10912] = 32'b11111111111111111110101101100100;
assign LUT_2[10913] = 32'b11111111111111111011100101111101;
assign LUT_2[10914] = 32'b00000000000000000101100110100000;
assign LUT_2[10915] = 32'b00000000000000000010011110111001;
assign LUT_2[10916] = 32'b11111111111111111011001011001100;
assign LUT_2[10917] = 32'b11111111111111111000000011100101;
assign LUT_2[10918] = 32'b00000000000000000010000100001000;
assign LUT_2[10919] = 32'b11111111111111111110111100100001;
assign LUT_2[10920] = 32'b11111111111111111001011111000001;
assign LUT_2[10921] = 32'b11111111111111110110010111011010;
assign LUT_2[10922] = 32'b00000000000000000000010111111101;
assign LUT_2[10923] = 32'b11111111111111111101010000010110;
assign LUT_2[10924] = 32'b11111111111111110101111100101001;
assign LUT_2[10925] = 32'b11111111111111110010110101000010;
assign LUT_2[10926] = 32'b11111111111111111100110101100101;
assign LUT_2[10927] = 32'b11111111111111111001101101111110;
assign LUT_2[10928] = 32'b11111111111111111001010001101110;
assign LUT_2[10929] = 32'b11111111111111110110001010000111;
assign LUT_2[10930] = 32'b00000000000000000000001010101010;
assign LUT_2[10931] = 32'b11111111111111111101000011000011;
assign LUT_2[10932] = 32'b11111111111111110101101111010110;
assign LUT_2[10933] = 32'b11111111111111110010100111101111;
assign LUT_2[10934] = 32'b11111111111111111100101000010010;
assign LUT_2[10935] = 32'b11111111111111111001100000101011;
assign LUT_2[10936] = 32'b11111111111111110100000011001011;
assign LUT_2[10937] = 32'b11111111111111110000111011100100;
assign LUT_2[10938] = 32'b11111111111111111010111100000111;
assign LUT_2[10939] = 32'b11111111111111110111110100100000;
assign LUT_2[10940] = 32'b11111111111111110000100000110011;
assign LUT_2[10941] = 32'b11111111111111101101011001001100;
assign LUT_2[10942] = 32'b11111111111111110111011001101111;
assign LUT_2[10943] = 32'b11111111111111110100010010001000;
assign LUT_2[10944] = 32'b11111111111111110110011010011110;
assign LUT_2[10945] = 32'b11111111111111110011010010110111;
assign LUT_2[10946] = 32'b11111111111111111101010011011010;
assign LUT_2[10947] = 32'b11111111111111111010001011110011;
assign LUT_2[10948] = 32'b11111111111111110010111000000110;
assign LUT_2[10949] = 32'b11111111111111101111110000011111;
assign LUT_2[10950] = 32'b11111111111111111001110001000010;
assign LUT_2[10951] = 32'b11111111111111110110101001011011;
assign LUT_2[10952] = 32'b11111111111111110001001011111011;
assign LUT_2[10953] = 32'b11111111111111101110000100010100;
assign LUT_2[10954] = 32'b11111111111111111000000100110111;
assign LUT_2[10955] = 32'b11111111111111110100111101010000;
assign LUT_2[10956] = 32'b11111111111111101101101001100011;
assign LUT_2[10957] = 32'b11111111111111101010100001111100;
assign LUT_2[10958] = 32'b11111111111111110100100010011111;
assign LUT_2[10959] = 32'b11111111111111110001011010111000;
assign LUT_2[10960] = 32'b11111111111111110000111110101000;
assign LUT_2[10961] = 32'b11111111111111101101110111000001;
assign LUT_2[10962] = 32'b11111111111111110111110111100100;
assign LUT_2[10963] = 32'b11111111111111110100101111111101;
assign LUT_2[10964] = 32'b11111111111111101101011100010000;
assign LUT_2[10965] = 32'b11111111111111101010010100101001;
assign LUT_2[10966] = 32'b11111111111111110100010101001100;
assign LUT_2[10967] = 32'b11111111111111110001001101100101;
assign LUT_2[10968] = 32'b11111111111111101011110000000101;
assign LUT_2[10969] = 32'b11111111111111101000101000011110;
assign LUT_2[10970] = 32'b11111111111111110010101001000001;
assign LUT_2[10971] = 32'b11111111111111101111100001011010;
assign LUT_2[10972] = 32'b11111111111111101000001101101101;
assign LUT_2[10973] = 32'b11111111111111100101000110000110;
assign LUT_2[10974] = 32'b11111111111111101111000110101001;
assign LUT_2[10975] = 32'b11111111111111101011111111000010;
assign LUT_2[10976] = 32'b11111111111111110110110110000111;
assign LUT_2[10977] = 32'b11111111111111110011101110100000;
assign LUT_2[10978] = 32'b11111111111111111101101111000011;
assign LUT_2[10979] = 32'b11111111111111111010100111011100;
assign LUT_2[10980] = 32'b11111111111111110011010011101111;
assign LUT_2[10981] = 32'b11111111111111110000001100001000;
assign LUT_2[10982] = 32'b11111111111111111010001100101011;
assign LUT_2[10983] = 32'b11111111111111110111000101000100;
assign LUT_2[10984] = 32'b11111111111111110001100111100100;
assign LUT_2[10985] = 32'b11111111111111101110011111111101;
assign LUT_2[10986] = 32'b11111111111111111000100000100000;
assign LUT_2[10987] = 32'b11111111111111110101011000111001;
assign LUT_2[10988] = 32'b11111111111111101110000101001100;
assign LUT_2[10989] = 32'b11111111111111101010111101100101;
assign LUT_2[10990] = 32'b11111111111111110100111110001000;
assign LUT_2[10991] = 32'b11111111111111110001110110100001;
assign LUT_2[10992] = 32'b11111111111111110001011010010001;
assign LUT_2[10993] = 32'b11111111111111101110010010101010;
assign LUT_2[10994] = 32'b11111111111111111000010011001101;
assign LUT_2[10995] = 32'b11111111111111110101001011100110;
assign LUT_2[10996] = 32'b11111111111111101101110111111001;
assign LUT_2[10997] = 32'b11111111111111101010110000010010;
assign LUT_2[10998] = 32'b11111111111111110100110000110101;
assign LUT_2[10999] = 32'b11111111111111110001101001001110;
assign LUT_2[11000] = 32'b11111111111111101100001011101110;
assign LUT_2[11001] = 32'b11111111111111101001000100000111;
assign LUT_2[11002] = 32'b11111111111111110011000100101010;
assign LUT_2[11003] = 32'b11111111111111101111111101000011;
assign LUT_2[11004] = 32'b11111111111111101000101001010110;
assign LUT_2[11005] = 32'b11111111111111100101100001101111;
assign LUT_2[11006] = 32'b11111111111111101111100010010010;
assign LUT_2[11007] = 32'b11111111111111101100011010101011;
assign LUT_2[11008] = 32'b11111111111111111101111100010010;
assign LUT_2[11009] = 32'b11111111111111111010110100101011;
assign LUT_2[11010] = 32'b00000000000000000100110101001110;
assign LUT_2[11011] = 32'b00000000000000000001101101100111;
assign LUT_2[11012] = 32'b11111111111111111010011001111010;
assign LUT_2[11013] = 32'b11111111111111110111010010010011;
assign LUT_2[11014] = 32'b00000000000000000001010010110110;
assign LUT_2[11015] = 32'b11111111111111111110001011001111;
assign LUT_2[11016] = 32'b11111111111111111000101101101111;
assign LUT_2[11017] = 32'b11111111111111110101100110001000;
assign LUT_2[11018] = 32'b11111111111111111111100110101011;
assign LUT_2[11019] = 32'b11111111111111111100011111000100;
assign LUT_2[11020] = 32'b11111111111111110101001011010111;
assign LUT_2[11021] = 32'b11111111111111110010000011110000;
assign LUT_2[11022] = 32'b11111111111111111100000100010011;
assign LUT_2[11023] = 32'b11111111111111111000111100101100;
assign LUT_2[11024] = 32'b11111111111111111000100000011100;
assign LUT_2[11025] = 32'b11111111111111110101011000110101;
assign LUT_2[11026] = 32'b11111111111111111111011001011000;
assign LUT_2[11027] = 32'b11111111111111111100010001110001;
assign LUT_2[11028] = 32'b11111111111111110100111110000100;
assign LUT_2[11029] = 32'b11111111111111110001110110011101;
assign LUT_2[11030] = 32'b11111111111111111011110111000000;
assign LUT_2[11031] = 32'b11111111111111111000101111011001;
assign LUT_2[11032] = 32'b11111111111111110011010001111001;
assign LUT_2[11033] = 32'b11111111111111110000001010010010;
assign LUT_2[11034] = 32'b11111111111111111010001010110101;
assign LUT_2[11035] = 32'b11111111111111110111000011001110;
assign LUT_2[11036] = 32'b11111111111111101111101111100001;
assign LUT_2[11037] = 32'b11111111111111101100100111111010;
assign LUT_2[11038] = 32'b11111111111111110110101000011101;
assign LUT_2[11039] = 32'b11111111111111110011100000110110;
assign LUT_2[11040] = 32'b11111111111111111110010111111011;
assign LUT_2[11041] = 32'b11111111111111111011010000010100;
assign LUT_2[11042] = 32'b00000000000000000101010000110111;
assign LUT_2[11043] = 32'b00000000000000000010001001010000;
assign LUT_2[11044] = 32'b11111111111111111010110101100011;
assign LUT_2[11045] = 32'b11111111111111110111101101111100;
assign LUT_2[11046] = 32'b00000000000000000001101110011111;
assign LUT_2[11047] = 32'b11111111111111111110100110111000;
assign LUT_2[11048] = 32'b11111111111111111001001001011000;
assign LUT_2[11049] = 32'b11111111111111110110000001110001;
assign LUT_2[11050] = 32'b00000000000000000000000010010100;
assign LUT_2[11051] = 32'b11111111111111111100111010101101;
assign LUT_2[11052] = 32'b11111111111111110101100111000000;
assign LUT_2[11053] = 32'b11111111111111110010011111011001;
assign LUT_2[11054] = 32'b11111111111111111100011111111100;
assign LUT_2[11055] = 32'b11111111111111111001011000010101;
assign LUT_2[11056] = 32'b11111111111111111000111100000101;
assign LUT_2[11057] = 32'b11111111111111110101110100011110;
assign LUT_2[11058] = 32'b11111111111111111111110101000001;
assign LUT_2[11059] = 32'b11111111111111111100101101011010;
assign LUT_2[11060] = 32'b11111111111111110101011001101101;
assign LUT_2[11061] = 32'b11111111111111110010010010000110;
assign LUT_2[11062] = 32'b11111111111111111100010010101001;
assign LUT_2[11063] = 32'b11111111111111111001001011000010;
assign LUT_2[11064] = 32'b11111111111111110011101101100010;
assign LUT_2[11065] = 32'b11111111111111110000100101111011;
assign LUT_2[11066] = 32'b11111111111111111010100110011110;
assign LUT_2[11067] = 32'b11111111111111110111011110110111;
assign LUT_2[11068] = 32'b11111111111111110000001011001010;
assign LUT_2[11069] = 32'b11111111111111101101000011100011;
assign LUT_2[11070] = 32'b11111111111111110111000100000110;
assign LUT_2[11071] = 32'b11111111111111110011111100011111;
assign LUT_2[11072] = 32'b11111111111111110110000100110101;
assign LUT_2[11073] = 32'b11111111111111110010111101001110;
assign LUT_2[11074] = 32'b11111111111111111100111101110001;
assign LUT_2[11075] = 32'b11111111111111111001110110001010;
assign LUT_2[11076] = 32'b11111111111111110010100010011101;
assign LUT_2[11077] = 32'b11111111111111101111011010110110;
assign LUT_2[11078] = 32'b11111111111111111001011011011001;
assign LUT_2[11079] = 32'b11111111111111110110010011110010;
assign LUT_2[11080] = 32'b11111111111111110000110110010010;
assign LUT_2[11081] = 32'b11111111111111101101101110101011;
assign LUT_2[11082] = 32'b11111111111111110111101111001110;
assign LUT_2[11083] = 32'b11111111111111110100100111100111;
assign LUT_2[11084] = 32'b11111111111111101101010011111010;
assign LUT_2[11085] = 32'b11111111111111101010001100010011;
assign LUT_2[11086] = 32'b11111111111111110100001100110110;
assign LUT_2[11087] = 32'b11111111111111110001000101001111;
assign LUT_2[11088] = 32'b11111111111111110000101000111111;
assign LUT_2[11089] = 32'b11111111111111101101100001011000;
assign LUT_2[11090] = 32'b11111111111111110111100001111011;
assign LUT_2[11091] = 32'b11111111111111110100011010010100;
assign LUT_2[11092] = 32'b11111111111111101101000110100111;
assign LUT_2[11093] = 32'b11111111111111101001111111000000;
assign LUT_2[11094] = 32'b11111111111111110011111111100011;
assign LUT_2[11095] = 32'b11111111111111110000110111111100;
assign LUT_2[11096] = 32'b11111111111111101011011010011100;
assign LUT_2[11097] = 32'b11111111111111101000010010110101;
assign LUT_2[11098] = 32'b11111111111111110010010011011000;
assign LUT_2[11099] = 32'b11111111111111101111001011110001;
assign LUT_2[11100] = 32'b11111111111111100111111000000100;
assign LUT_2[11101] = 32'b11111111111111100100110000011101;
assign LUT_2[11102] = 32'b11111111111111101110110001000000;
assign LUT_2[11103] = 32'b11111111111111101011101001011001;
assign LUT_2[11104] = 32'b11111111111111110110100000011110;
assign LUT_2[11105] = 32'b11111111111111110011011000110111;
assign LUT_2[11106] = 32'b11111111111111111101011001011010;
assign LUT_2[11107] = 32'b11111111111111111010010001110011;
assign LUT_2[11108] = 32'b11111111111111110010111110000110;
assign LUT_2[11109] = 32'b11111111111111101111110110011111;
assign LUT_2[11110] = 32'b11111111111111111001110111000010;
assign LUT_2[11111] = 32'b11111111111111110110101111011011;
assign LUT_2[11112] = 32'b11111111111111110001010001111011;
assign LUT_2[11113] = 32'b11111111111111101110001010010100;
assign LUT_2[11114] = 32'b11111111111111111000001010110111;
assign LUT_2[11115] = 32'b11111111111111110101000011010000;
assign LUT_2[11116] = 32'b11111111111111101101101111100011;
assign LUT_2[11117] = 32'b11111111111111101010100111111100;
assign LUT_2[11118] = 32'b11111111111111110100101000011111;
assign LUT_2[11119] = 32'b11111111111111110001100000111000;
assign LUT_2[11120] = 32'b11111111111111110001000100101000;
assign LUT_2[11121] = 32'b11111111111111101101111101000001;
assign LUT_2[11122] = 32'b11111111111111110111111101100100;
assign LUT_2[11123] = 32'b11111111111111110100110101111101;
assign LUT_2[11124] = 32'b11111111111111101101100010010000;
assign LUT_2[11125] = 32'b11111111111111101010011010101001;
assign LUT_2[11126] = 32'b11111111111111110100011011001100;
assign LUT_2[11127] = 32'b11111111111111110001010011100101;
assign LUT_2[11128] = 32'b11111111111111101011110110000101;
assign LUT_2[11129] = 32'b11111111111111101000101110011110;
assign LUT_2[11130] = 32'b11111111111111110010101111000001;
assign LUT_2[11131] = 32'b11111111111111101111100111011010;
assign LUT_2[11132] = 32'b11111111111111101000010011101101;
assign LUT_2[11133] = 32'b11111111111111100101001100000110;
assign LUT_2[11134] = 32'b11111111111111101111001100101001;
assign LUT_2[11135] = 32'b11111111111111101100000101000010;
assign LUT_2[11136] = 32'b00000000000000000010010000100001;
assign LUT_2[11137] = 32'b11111111111111111111001000111010;
assign LUT_2[11138] = 32'b00000000000000001001001001011101;
assign LUT_2[11139] = 32'b00000000000000000110000001110110;
assign LUT_2[11140] = 32'b11111111111111111110101110001001;
assign LUT_2[11141] = 32'b11111111111111111011100110100010;
assign LUT_2[11142] = 32'b00000000000000000101100111000101;
assign LUT_2[11143] = 32'b00000000000000000010011111011110;
assign LUT_2[11144] = 32'b11111111111111111101000001111110;
assign LUT_2[11145] = 32'b11111111111111111001111010010111;
assign LUT_2[11146] = 32'b00000000000000000011111010111010;
assign LUT_2[11147] = 32'b00000000000000000000110011010011;
assign LUT_2[11148] = 32'b11111111111111111001011111100110;
assign LUT_2[11149] = 32'b11111111111111110110010111111111;
assign LUT_2[11150] = 32'b00000000000000000000011000100010;
assign LUT_2[11151] = 32'b11111111111111111101010000111011;
assign LUT_2[11152] = 32'b11111111111111111100110100101011;
assign LUT_2[11153] = 32'b11111111111111111001101101000100;
assign LUT_2[11154] = 32'b00000000000000000011101101100111;
assign LUT_2[11155] = 32'b00000000000000000000100110000000;
assign LUT_2[11156] = 32'b11111111111111111001010010010011;
assign LUT_2[11157] = 32'b11111111111111110110001010101100;
assign LUT_2[11158] = 32'b00000000000000000000001011001111;
assign LUT_2[11159] = 32'b11111111111111111101000011101000;
assign LUT_2[11160] = 32'b11111111111111110111100110001000;
assign LUT_2[11161] = 32'b11111111111111110100011110100001;
assign LUT_2[11162] = 32'b11111111111111111110011111000100;
assign LUT_2[11163] = 32'b11111111111111111011010111011101;
assign LUT_2[11164] = 32'b11111111111111110100000011110000;
assign LUT_2[11165] = 32'b11111111111111110000111100001001;
assign LUT_2[11166] = 32'b11111111111111111010111100101100;
assign LUT_2[11167] = 32'b11111111111111110111110101000101;
assign LUT_2[11168] = 32'b00000000000000000010101100001010;
assign LUT_2[11169] = 32'b11111111111111111111100100100011;
assign LUT_2[11170] = 32'b00000000000000001001100101000110;
assign LUT_2[11171] = 32'b00000000000000000110011101011111;
assign LUT_2[11172] = 32'b11111111111111111111001001110010;
assign LUT_2[11173] = 32'b11111111111111111100000010001011;
assign LUT_2[11174] = 32'b00000000000000000110000010101110;
assign LUT_2[11175] = 32'b00000000000000000010111011000111;
assign LUT_2[11176] = 32'b11111111111111111101011101100111;
assign LUT_2[11177] = 32'b11111111111111111010010110000000;
assign LUT_2[11178] = 32'b00000000000000000100010110100011;
assign LUT_2[11179] = 32'b00000000000000000001001110111100;
assign LUT_2[11180] = 32'b11111111111111111001111011001111;
assign LUT_2[11181] = 32'b11111111111111110110110011101000;
assign LUT_2[11182] = 32'b00000000000000000000110100001011;
assign LUT_2[11183] = 32'b11111111111111111101101100100100;
assign LUT_2[11184] = 32'b11111111111111111101010000010100;
assign LUT_2[11185] = 32'b11111111111111111010001000101101;
assign LUT_2[11186] = 32'b00000000000000000100001001010000;
assign LUT_2[11187] = 32'b00000000000000000001000001101001;
assign LUT_2[11188] = 32'b11111111111111111001101101111100;
assign LUT_2[11189] = 32'b11111111111111110110100110010101;
assign LUT_2[11190] = 32'b00000000000000000000100110111000;
assign LUT_2[11191] = 32'b11111111111111111101011111010001;
assign LUT_2[11192] = 32'b11111111111111111000000001110001;
assign LUT_2[11193] = 32'b11111111111111110100111010001010;
assign LUT_2[11194] = 32'b11111111111111111110111010101101;
assign LUT_2[11195] = 32'b11111111111111111011110011000110;
assign LUT_2[11196] = 32'b11111111111111110100011111011001;
assign LUT_2[11197] = 32'b11111111111111110001010111110010;
assign LUT_2[11198] = 32'b11111111111111111011011000010101;
assign LUT_2[11199] = 32'b11111111111111111000010000101110;
assign LUT_2[11200] = 32'b11111111111111111010011001000100;
assign LUT_2[11201] = 32'b11111111111111110111010001011101;
assign LUT_2[11202] = 32'b00000000000000000001010010000000;
assign LUT_2[11203] = 32'b11111111111111111110001010011001;
assign LUT_2[11204] = 32'b11111111111111110110110110101100;
assign LUT_2[11205] = 32'b11111111111111110011101111000101;
assign LUT_2[11206] = 32'b11111111111111111101101111101000;
assign LUT_2[11207] = 32'b11111111111111111010101000000001;
assign LUT_2[11208] = 32'b11111111111111110101001010100001;
assign LUT_2[11209] = 32'b11111111111111110010000010111010;
assign LUT_2[11210] = 32'b11111111111111111100000011011101;
assign LUT_2[11211] = 32'b11111111111111111000111011110110;
assign LUT_2[11212] = 32'b11111111111111110001101000001001;
assign LUT_2[11213] = 32'b11111111111111101110100000100010;
assign LUT_2[11214] = 32'b11111111111111111000100001000101;
assign LUT_2[11215] = 32'b11111111111111110101011001011110;
assign LUT_2[11216] = 32'b11111111111111110100111101001110;
assign LUT_2[11217] = 32'b11111111111111110001110101100111;
assign LUT_2[11218] = 32'b11111111111111111011110110001010;
assign LUT_2[11219] = 32'b11111111111111111000101110100011;
assign LUT_2[11220] = 32'b11111111111111110001011010110110;
assign LUT_2[11221] = 32'b11111111111111101110010011001111;
assign LUT_2[11222] = 32'b11111111111111111000010011110010;
assign LUT_2[11223] = 32'b11111111111111110101001100001011;
assign LUT_2[11224] = 32'b11111111111111101111101110101011;
assign LUT_2[11225] = 32'b11111111111111101100100111000100;
assign LUT_2[11226] = 32'b11111111111111110110100111100111;
assign LUT_2[11227] = 32'b11111111111111110011100000000000;
assign LUT_2[11228] = 32'b11111111111111101100001100010011;
assign LUT_2[11229] = 32'b11111111111111101001000100101100;
assign LUT_2[11230] = 32'b11111111111111110011000101001111;
assign LUT_2[11231] = 32'b11111111111111101111111101101000;
assign LUT_2[11232] = 32'b11111111111111111010110100101101;
assign LUT_2[11233] = 32'b11111111111111110111101101000110;
assign LUT_2[11234] = 32'b00000000000000000001101101101001;
assign LUT_2[11235] = 32'b11111111111111111110100110000010;
assign LUT_2[11236] = 32'b11111111111111110111010010010101;
assign LUT_2[11237] = 32'b11111111111111110100001010101110;
assign LUT_2[11238] = 32'b11111111111111111110001011010001;
assign LUT_2[11239] = 32'b11111111111111111011000011101010;
assign LUT_2[11240] = 32'b11111111111111110101100110001010;
assign LUT_2[11241] = 32'b11111111111111110010011110100011;
assign LUT_2[11242] = 32'b11111111111111111100011111000110;
assign LUT_2[11243] = 32'b11111111111111111001010111011111;
assign LUT_2[11244] = 32'b11111111111111110010000011110010;
assign LUT_2[11245] = 32'b11111111111111101110111100001011;
assign LUT_2[11246] = 32'b11111111111111111000111100101110;
assign LUT_2[11247] = 32'b11111111111111110101110101000111;
assign LUT_2[11248] = 32'b11111111111111110101011000110111;
assign LUT_2[11249] = 32'b11111111111111110010010001010000;
assign LUT_2[11250] = 32'b11111111111111111100010001110011;
assign LUT_2[11251] = 32'b11111111111111111001001010001100;
assign LUT_2[11252] = 32'b11111111111111110001110110011111;
assign LUT_2[11253] = 32'b11111111111111101110101110111000;
assign LUT_2[11254] = 32'b11111111111111111000101111011011;
assign LUT_2[11255] = 32'b11111111111111110101100111110100;
assign LUT_2[11256] = 32'b11111111111111110000001010010100;
assign LUT_2[11257] = 32'b11111111111111101101000010101101;
assign LUT_2[11258] = 32'b11111111111111110111000011010000;
assign LUT_2[11259] = 32'b11111111111111110011111011101001;
assign LUT_2[11260] = 32'b11111111111111101100100111111100;
assign LUT_2[11261] = 32'b11111111111111101001100000010101;
assign LUT_2[11262] = 32'b11111111111111110011100000111000;
assign LUT_2[11263] = 32'b11111111111111110000011001010001;
assign LUT_2[11264] = 32'b11111111111111111011110111111111;
assign LUT_2[11265] = 32'b11111111111111111000110000011000;
assign LUT_2[11266] = 32'b00000000000000000010110000111011;
assign LUT_2[11267] = 32'b11111111111111111111101001010100;
assign LUT_2[11268] = 32'b11111111111111111000010101100111;
assign LUT_2[11269] = 32'b11111111111111110101001110000000;
assign LUT_2[11270] = 32'b11111111111111111111001110100011;
assign LUT_2[11271] = 32'b11111111111111111100000110111100;
assign LUT_2[11272] = 32'b11111111111111110110101001011100;
assign LUT_2[11273] = 32'b11111111111111110011100001110101;
assign LUT_2[11274] = 32'b11111111111111111101100010011000;
assign LUT_2[11275] = 32'b11111111111111111010011010110001;
assign LUT_2[11276] = 32'b11111111111111110011000111000100;
assign LUT_2[11277] = 32'b11111111111111101111111111011101;
assign LUT_2[11278] = 32'b11111111111111111010000000000000;
assign LUT_2[11279] = 32'b11111111111111110110111000011001;
assign LUT_2[11280] = 32'b11111111111111110110011100001001;
assign LUT_2[11281] = 32'b11111111111111110011010100100010;
assign LUT_2[11282] = 32'b11111111111111111101010101000101;
assign LUT_2[11283] = 32'b11111111111111111010001101011110;
assign LUT_2[11284] = 32'b11111111111111110010111001110001;
assign LUT_2[11285] = 32'b11111111111111101111110010001010;
assign LUT_2[11286] = 32'b11111111111111111001110010101101;
assign LUT_2[11287] = 32'b11111111111111110110101011000110;
assign LUT_2[11288] = 32'b11111111111111110001001101100110;
assign LUT_2[11289] = 32'b11111111111111101110000101111111;
assign LUT_2[11290] = 32'b11111111111111111000000110100010;
assign LUT_2[11291] = 32'b11111111111111110100111110111011;
assign LUT_2[11292] = 32'b11111111111111101101101011001110;
assign LUT_2[11293] = 32'b11111111111111101010100011100111;
assign LUT_2[11294] = 32'b11111111111111110100100100001010;
assign LUT_2[11295] = 32'b11111111111111110001011100100011;
assign LUT_2[11296] = 32'b11111111111111111100010011101000;
assign LUT_2[11297] = 32'b11111111111111111001001100000001;
assign LUT_2[11298] = 32'b00000000000000000011001100100100;
assign LUT_2[11299] = 32'b00000000000000000000000100111101;
assign LUT_2[11300] = 32'b11111111111111111000110001010000;
assign LUT_2[11301] = 32'b11111111111111110101101001101001;
assign LUT_2[11302] = 32'b11111111111111111111101010001100;
assign LUT_2[11303] = 32'b11111111111111111100100010100101;
assign LUT_2[11304] = 32'b11111111111111110111000101000101;
assign LUT_2[11305] = 32'b11111111111111110011111101011110;
assign LUT_2[11306] = 32'b11111111111111111101111110000001;
assign LUT_2[11307] = 32'b11111111111111111010110110011010;
assign LUT_2[11308] = 32'b11111111111111110011100010101101;
assign LUT_2[11309] = 32'b11111111111111110000011011000110;
assign LUT_2[11310] = 32'b11111111111111111010011011101001;
assign LUT_2[11311] = 32'b11111111111111110111010100000010;
assign LUT_2[11312] = 32'b11111111111111110110110111110010;
assign LUT_2[11313] = 32'b11111111111111110011110000001011;
assign LUT_2[11314] = 32'b11111111111111111101110000101110;
assign LUT_2[11315] = 32'b11111111111111111010101001000111;
assign LUT_2[11316] = 32'b11111111111111110011010101011010;
assign LUT_2[11317] = 32'b11111111111111110000001101110011;
assign LUT_2[11318] = 32'b11111111111111111010001110010110;
assign LUT_2[11319] = 32'b11111111111111110111000110101111;
assign LUT_2[11320] = 32'b11111111111111110001101001001111;
assign LUT_2[11321] = 32'b11111111111111101110100001101000;
assign LUT_2[11322] = 32'b11111111111111111000100010001011;
assign LUT_2[11323] = 32'b11111111111111110101011010100100;
assign LUT_2[11324] = 32'b11111111111111101110000110110111;
assign LUT_2[11325] = 32'b11111111111111101010111111010000;
assign LUT_2[11326] = 32'b11111111111111110100111111110011;
assign LUT_2[11327] = 32'b11111111111111110001111000001100;
assign LUT_2[11328] = 32'b11111111111111110100000000100010;
assign LUT_2[11329] = 32'b11111111111111110000111000111011;
assign LUT_2[11330] = 32'b11111111111111111010111001011110;
assign LUT_2[11331] = 32'b11111111111111110111110001110111;
assign LUT_2[11332] = 32'b11111111111111110000011110001010;
assign LUT_2[11333] = 32'b11111111111111101101010110100011;
assign LUT_2[11334] = 32'b11111111111111110111010111000110;
assign LUT_2[11335] = 32'b11111111111111110100001111011111;
assign LUT_2[11336] = 32'b11111111111111101110110001111111;
assign LUT_2[11337] = 32'b11111111111111101011101010011000;
assign LUT_2[11338] = 32'b11111111111111110101101010111011;
assign LUT_2[11339] = 32'b11111111111111110010100011010100;
assign LUT_2[11340] = 32'b11111111111111101011001111100111;
assign LUT_2[11341] = 32'b11111111111111101000001000000000;
assign LUT_2[11342] = 32'b11111111111111110010001000100011;
assign LUT_2[11343] = 32'b11111111111111101111000000111100;
assign LUT_2[11344] = 32'b11111111111111101110100100101100;
assign LUT_2[11345] = 32'b11111111111111101011011101000101;
assign LUT_2[11346] = 32'b11111111111111110101011101101000;
assign LUT_2[11347] = 32'b11111111111111110010010110000001;
assign LUT_2[11348] = 32'b11111111111111101011000010010100;
assign LUT_2[11349] = 32'b11111111111111100111111010101101;
assign LUT_2[11350] = 32'b11111111111111110001111011010000;
assign LUT_2[11351] = 32'b11111111111111101110110011101001;
assign LUT_2[11352] = 32'b11111111111111101001010110001001;
assign LUT_2[11353] = 32'b11111111111111100110001110100010;
assign LUT_2[11354] = 32'b11111111111111110000001111000101;
assign LUT_2[11355] = 32'b11111111111111101101000111011110;
assign LUT_2[11356] = 32'b11111111111111100101110011110001;
assign LUT_2[11357] = 32'b11111111111111100010101100001010;
assign LUT_2[11358] = 32'b11111111111111101100101100101101;
assign LUT_2[11359] = 32'b11111111111111101001100101000110;
assign LUT_2[11360] = 32'b11111111111111110100011100001011;
assign LUT_2[11361] = 32'b11111111111111110001010100100100;
assign LUT_2[11362] = 32'b11111111111111111011010101000111;
assign LUT_2[11363] = 32'b11111111111111111000001101100000;
assign LUT_2[11364] = 32'b11111111111111110000111001110011;
assign LUT_2[11365] = 32'b11111111111111101101110010001100;
assign LUT_2[11366] = 32'b11111111111111110111110010101111;
assign LUT_2[11367] = 32'b11111111111111110100101011001000;
assign LUT_2[11368] = 32'b11111111111111101111001101101000;
assign LUT_2[11369] = 32'b11111111111111101100000110000001;
assign LUT_2[11370] = 32'b11111111111111110110000110100100;
assign LUT_2[11371] = 32'b11111111111111110010111110111101;
assign LUT_2[11372] = 32'b11111111111111101011101011010000;
assign LUT_2[11373] = 32'b11111111111111101000100011101001;
assign LUT_2[11374] = 32'b11111111111111110010100100001100;
assign LUT_2[11375] = 32'b11111111111111101111011100100101;
assign LUT_2[11376] = 32'b11111111111111101111000000010101;
assign LUT_2[11377] = 32'b11111111111111101011111000101110;
assign LUT_2[11378] = 32'b11111111111111110101111001010001;
assign LUT_2[11379] = 32'b11111111111111110010110001101010;
assign LUT_2[11380] = 32'b11111111111111101011011101111101;
assign LUT_2[11381] = 32'b11111111111111101000010110010110;
assign LUT_2[11382] = 32'b11111111111111110010010110111001;
assign LUT_2[11383] = 32'b11111111111111101111001111010010;
assign LUT_2[11384] = 32'b11111111111111101001110001110010;
assign LUT_2[11385] = 32'b11111111111111100110101010001011;
assign LUT_2[11386] = 32'b11111111111111110000101010101110;
assign LUT_2[11387] = 32'b11111111111111101101100011000111;
assign LUT_2[11388] = 32'b11111111111111100110001111011010;
assign LUT_2[11389] = 32'b11111111111111100011000111110011;
assign LUT_2[11390] = 32'b11111111111111101101001000010110;
assign LUT_2[11391] = 32'b11111111111111101010000000101111;
assign LUT_2[11392] = 32'b00000000000000000000001100001110;
assign LUT_2[11393] = 32'b11111111111111111101000100100111;
assign LUT_2[11394] = 32'b00000000000000000111000101001010;
assign LUT_2[11395] = 32'b00000000000000000011111101100011;
assign LUT_2[11396] = 32'b11111111111111111100101001110110;
assign LUT_2[11397] = 32'b11111111111111111001100010001111;
assign LUT_2[11398] = 32'b00000000000000000011100010110010;
assign LUT_2[11399] = 32'b00000000000000000000011011001011;
assign LUT_2[11400] = 32'b11111111111111111010111101101011;
assign LUT_2[11401] = 32'b11111111111111110111110110000100;
assign LUT_2[11402] = 32'b00000000000000000001110110100111;
assign LUT_2[11403] = 32'b11111111111111111110101111000000;
assign LUT_2[11404] = 32'b11111111111111110111011011010011;
assign LUT_2[11405] = 32'b11111111111111110100010011101100;
assign LUT_2[11406] = 32'b11111111111111111110010100001111;
assign LUT_2[11407] = 32'b11111111111111111011001100101000;
assign LUT_2[11408] = 32'b11111111111111111010110000011000;
assign LUT_2[11409] = 32'b11111111111111110111101000110001;
assign LUT_2[11410] = 32'b00000000000000000001101001010100;
assign LUT_2[11411] = 32'b11111111111111111110100001101101;
assign LUT_2[11412] = 32'b11111111111111110111001110000000;
assign LUT_2[11413] = 32'b11111111111111110100000110011001;
assign LUT_2[11414] = 32'b11111111111111111110000110111100;
assign LUT_2[11415] = 32'b11111111111111111010111111010101;
assign LUT_2[11416] = 32'b11111111111111110101100001110101;
assign LUT_2[11417] = 32'b11111111111111110010011010001110;
assign LUT_2[11418] = 32'b11111111111111111100011010110001;
assign LUT_2[11419] = 32'b11111111111111111001010011001010;
assign LUT_2[11420] = 32'b11111111111111110001111111011101;
assign LUT_2[11421] = 32'b11111111111111101110110111110110;
assign LUT_2[11422] = 32'b11111111111111111000111000011001;
assign LUT_2[11423] = 32'b11111111111111110101110000110010;
assign LUT_2[11424] = 32'b00000000000000000000100111110111;
assign LUT_2[11425] = 32'b11111111111111111101100000010000;
assign LUT_2[11426] = 32'b00000000000000000111100000110011;
assign LUT_2[11427] = 32'b00000000000000000100011001001100;
assign LUT_2[11428] = 32'b11111111111111111101000101011111;
assign LUT_2[11429] = 32'b11111111111111111001111101111000;
assign LUT_2[11430] = 32'b00000000000000000011111110011011;
assign LUT_2[11431] = 32'b00000000000000000000110110110100;
assign LUT_2[11432] = 32'b11111111111111111011011001010100;
assign LUT_2[11433] = 32'b11111111111111111000010001101101;
assign LUT_2[11434] = 32'b00000000000000000010010010010000;
assign LUT_2[11435] = 32'b11111111111111111111001010101001;
assign LUT_2[11436] = 32'b11111111111111110111110110111100;
assign LUT_2[11437] = 32'b11111111111111110100101111010101;
assign LUT_2[11438] = 32'b11111111111111111110101111111000;
assign LUT_2[11439] = 32'b11111111111111111011101000010001;
assign LUT_2[11440] = 32'b11111111111111111011001100000001;
assign LUT_2[11441] = 32'b11111111111111111000000100011010;
assign LUT_2[11442] = 32'b00000000000000000010000100111101;
assign LUT_2[11443] = 32'b11111111111111111110111101010110;
assign LUT_2[11444] = 32'b11111111111111110111101001101001;
assign LUT_2[11445] = 32'b11111111111111110100100010000010;
assign LUT_2[11446] = 32'b11111111111111111110100010100101;
assign LUT_2[11447] = 32'b11111111111111111011011010111110;
assign LUT_2[11448] = 32'b11111111111111110101111101011110;
assign LUT_2[11449] = 32'b11111111111111110010110101110111;
assign LUT_2[11450] = 32'b11111111111111111100110110011010;
assign LUT_2[11451] = 32'b11111111111111111001101110110011;
assign LUT_2[11452] = 32'b11111111111111110010011011000110;
assign LUT_2[11453] = 32'b11111111111111101111010011011111;
assign LUT_2[11454] = 32'b11111111111111111001010100000010;
assign LUT_2[11455] = 32'b11111111111111110110001100011011;
assign LUT_2[11456] = 32'b11111111111111111000010100110001;
assign LUT_2[11457] = 32'b11111111111111110101001101001010;
assign LUT_2[11458] = 32'b11111111111111111111001101101101;
assign LUT_2[11459] = 32'b11111111111111111100000110000110;
assign LUT_2[11460] = 32'b11111111111111110100110010011001;
assign LUT_2[11461] = 32'b11111111111111110001101010110010;
assign LUT_2[11462] = 32'b11111111111111111011101011010101;
assign LUT_2[11463] = 32'b11111111111111111000100011101110;
assign LUT_2[11464] = 32'b11111111111111110011000110001110;
assign LUT_2[11465] = 32'b11111111111111101111111110100111;
assign LUT_2[11466] = 32'b11111111111111111001111111001010;
assign LUT_2[11467] = 32'b11111111111111110110110111100011;
assign LUT_2[11468] = 32'b11111111111111101111100011110110;
assign LUT_2[11469] = 32'b11111111111111101100011100001111;
assign LUT_2[11470] = 32'b11111111111111110110011100110010;
assign LUT_2[11471] = 32'b11111111111111110011010101001011;
assign LUT_2[11472] = 32'b11111111111111110010111000111011;
assign LUT_2[11473] = 32'b11111111111111101111110001010100;
assign LUT_2[11474] = 32'b11111111111111111001110001110111;
assign LUT_2[11475] = 32'b11111111111111110110101010010000;
assign LUT_2[11476] = 32'b11111111111111101111010110100011;
assign LUT_2[11477] = 32'b11111111111111101100001110111100;
assign LUT_2[11478] = 32'b11111111111111110110001111011111;
assign LUT_2[11479] = 32'b11111111111111110011000111111000;
assign LUT_2[11480] = 32'b11111111111111101101101010011000;
assign LUT_2[11481] = 32'b11111111111111101010100010110001;
assign LUT_2[11482] = 32'b11111111111111110100100011010100;
assign LUT_2[11483] = 32'b11111111111111110001011011101101;
assign LUT_2[11484] = 32'b11111111111111101010001000000000;
assign LUT_2[11485] = 32'b11111111111111100111000000011001;
assign LUT_2[11486] = 32'b11111111111111110001000000111100;
assign LUT_2[11487] = 32'b11111111111111101101111001010101;
assign LUT_2[11488] = 32'b11111111111111111000110000011010;
assign LUT_2[11489] = 32'b11111111111111110101101000110011;
assign LUT_2[11490] = 32'b11111111111111111111101001010110;
assign LUT_2[11491] = 32'b11111111111111111100100001101111;
assign LUT_2[11492] = 32'b11111111111111110101001110000010;
assign LUT_2[11493] = 32'b11111111111111110010000110011011;
assign LUT_2[11494] = 32'b11111111111111111100000110111110;
assign LUT_2[11495] = 32'b11111111111111111000111111010111;
assign LUT_2[11496] = 32'b11111111111111110011100001110111;
assign LUT_2[11497] = 32'b11111111111111110000011010010000;
assign LUT_2[11498] = 32'b11111111111111111010011010110011;
assign LUT_2[11499] = 32'b11111111111111110111010011001100;
assign LUT_2[11500] = 32'b11111111111111101111111111011111;
assign LUT_2[11501] = 32'b11111111111111101100110111111000;
assign LUT_2[11502] = 32'b11111111111111110110111000011011;
assign LUT_2[11503] = 32'b11111111111111110011110000110100;
assign LUT_2[11504] = 32'b11111111111111110011010100100100;
assign LUT_2[11505] = 32'b11111111111111110000001100111101;
assign LUT_2[11506] = 32'b11111111111111111010001101100000;
assign LUT_2[11507] = 32'b11111111111111110111000101111001;
assign LUT_2[11508] = 32'b11111111111111101111110010001100;
assign LUT_2[11509] = 32'b11111111111111101100101010100101;
assign LUT_2[11510] = 32'b11111111111111110110101011001000;
assign LUT_2[11511] = 32'b11111111111111110011100011100001;
assign LUT_2[11512] = 32'b11111111111111101110000110000001;
assign LUT_2[11513] = 32'b11111111111111101010111110011010;
assign LUT_2[11514] = 32'b11111111111111110100111110111101;
assign LUT_2[11515] = 32'b11111111111111110001110111010110;
assign LUT_2[11516] = 32'b11111111111111101010100011101001;
assign LUT_2[11517] = 32'b11111111111111100111011100000010;
assign LUT_2[11518] = 32'b11111111111111110001011100100101;
assign LUT_2[11519] = 32'b11111111111111101110010100111110;
assign LUT_2[11520] = 32'b11111111111111111111110110100101;
assign LUT_2[11521] = 32'b11111111111111111100101110111110;
assign LUT_2[11522] = 32'b00000000000000000110101111100001;
assign LUT_2[11523] = 32'b00000000000000000011100111111010;
assign LUT_2[11524] = 32'b11111111111111111100010100001101;
assign LUT_2[11525] = 32'b11111111111111111001001100100110;
assign LUT_2[11526] = 32'b00000000000000000011001101001001;
assign LUT_2[11527] = 32'b00000000000000000000000101100010;
assign LUT_2[11528] = 32'b11111111111111111010101000000010;
assign LUT_2[11529] = 32'b11111111111111110111100000011011;
assign LUT_2[11530] = 32'b00000000000000000001100000111110;
assign LUT_2[11531] = 32'b11111111111111111110011001010111;
assign LUT_2[11532] = 32'b11111111111111110111000101101010;
assign LUT_2[11533] = 32'b11111111111111110011111110000011;
assign LUT_2[11534] = 32'b11111111111111111101111110100110;
assign LUT_2[11535] = 32'b11111111111111111010110110111111;
assign LUT_2[11536] = 32'b11111111111111111010011010101111;
assign LUT_2[11537] = 32'b11111111111111110111010011001000;
assign LUT_2[11538] = 32'b00000000000000000001010011101011;
assign LUT_2[11539] = 32'b11111111111111111110001100000100;
assign LUT_2[11540] = 32'b11111111111111110110111000010111;
assign LUT_2[11541] = 32'b11111111111111110011110000110000;
assign LUT_2[11542] = 32'b11111111111111111101110001010011;
assign LUT_2[11543] = 32'b11111111111111111010101001101100;
assign LUT_2[11544] = 32'b11111111111111110101001100001100;
assign LUT_2[11545] = 32'b11111111111111110010000100100101;
assign LUT_2[11546] = 32'b11111111111111111100000101001000;
assign LUT_2[11547] = 32'b11111111111111111000111101100001;
assign LUT_2[11548] = 32'b11111111111111110001101001110100;
assign LUT_2[11549] = 32'b11111111111111101110100010001101;
assign LUT_2[11550] = 32'b11111111111111111000100010110000;
assign LUT_2[11551] = 32'b11111111111111110101011011001001;
assign LUT_2[11552] = 32'b00000000000000000000010010001110;
assign LUT_2[11553] = 32'b11111111111111111101001010100111;
assign LUT_2[11554] = 32'b00000000000000000111001011001010;
assign LUT_2[11555] = 32'b00000000000000000100000011100011;
assign LUT_2[11556] = 32'b11111111111111111100101111110110;
assign LUT_2[11557] = 32'b11111111111111111001101000001111;
assign LUT_2[11558] = 32'b00000000000000000011101000110010;
assign LUT_2[11559] = 32'b00000000000000000000100001001011;
assign LUT_2[11560] = 32'b11111111111111111011000011101011;
assign LUT_2[11561] = 32'b11111111111111110111111100000100;
assign LUT_2[11562] = 32'b00000000000000000001111100100111;
assign LUT_2[11563] = 32'b11111111111111111110110101000000;
assign LUT_2[11564] = 32'b11111111111111110111100001010011;
assign LUT_2[11565] = 32'b11111111111111110100011001101100;
assign LUT_2[11566] = 32'b11111111111111111110011010001111;
assign LUT_2[11567] = 32'b11111111111111111011010010101000;
assign LUT_2[11568] = 32'b11111111111111111010110110011000;
assign LUT_2[11569] = 32'b11111111111111110111101110110001;
assign LUT_2[11570] = 32'b00000000000000000001101111010100;
assign LUT_2[11571] = 32'b11111111111111111110100111101101;
assign LUT_2[11572] = 32'b11111111111111110111010100000000;
assign LUT_2[11573] = 32'b11111111111111110100001100011001;
assign LUT_2[11574] = 32'b11111111111111111110001100111100;
assign LUT_2[11575] = 32'b11111111111111111011000101010101;
assign LUT_2[11576] = 32'b11111111111111110101100111110101;
assign LUT_2[11577] = 32'b11111111111111110010100000001110;
assign LUT_2[11578] = 32'b11111111111111111100100000110001;
assign LUT_2[11579] = 32'b11111111111111111001011001001010;
assign LUT_2[11580] = 32'b11111111111111110010000101011101;
assign LUT_2[11581] = 32'b11111111111111101110111101110110;
assign LUT_2[11582] = 32'b11111111111111111000111110011001;
assign LUT_2[11583] = 32'b11111111111111110101110110110010;
assign LUT_2[11584] = 32'b11111111111111110111111111001000;
assign LUT_2[11585] = 32'b11111111111111110100110111100001;
assign LUT_2[11586] = 32'b11111111111111111110111000000100;
assign LUT_2[11587] = 32'b11111111111111111011110000011101;
assign LUT_2[11588] = 32'b11111111111111110100011100110000;
assign LUT_2[11589] = 32'b11111111111111110001010101001001;
assign LUT_2[11590] = 32'b11111111111111111011010101101100;
assign LUT_2[11591] = 32'b11111111111111111000001110000101;
assign LUT_2[11592] = 32'b11111111111111110010110000100101;
assign LUT_2[11593] = 32'b11111111111111101111101000111110;
assign LUT_2[11594] = 32'b11111111111111111001101001100001;
assign LUT_2[11595] = 32'b11111111111111110110100001111010;
assign LUT_2[11596] = 32'b11111111111111101111001110001101;
assign LUT_2[11597] = 32'b11111111111111101100000110100110;
assign LUT_2[11598] = 32'b11111111111111110110000111001001;
assign LUT_2[11599] = 32'b11111111111111110010111111100010;
assign LUT_2[11600] = 32'b11111111111111110010100011010010;
assign LUT_2[11601] = 32'b11111111111111101111011011101011;
assign LUT_2[11602] = 32'b11111111111111111001011100001110;
assign LUT_2[11603] = 32'b11111111111111110110010100100111;
assign LUT_2[11604] = 32'b11111111111111101111000000111010;
assign LUT_2[11605] = 32'b11111111111111101011111001010011;
assign LUT_2[11606] = 32'b11111111111111110101111001110110;
assign LUT_2[11607] = 32'b11111111111111110010110010001111;
assign LUT_2[11608] = 32'b11111111111111101101010100101111;
assign LUT_2[11609] = 32'b11111111111111101010001101001000;
assign LUT_2[11610] = 32'b11111111111111110100001101101011;
assign LUT_2[11611] = 32'b11111111111111110001000110000100;
assign LUT_2[11612] = 32'b11111111111111101001110010010111;
assign LUT_2[11613] = 32'b11111111111111100110101010110000;
assign LUT_2[11614] = 32'b11111111111111110000101011010011;
assign LUT_2[11615] = 32'b11111111111111101101100011101100;
assign LUT_2[11616] = 32'b11111111111111111000011010110001;
assign LUT_2[11617] = 32'b11111111111111110101010011001010;
assign LUT_2[11618] = 32'b11111111111111111111010011101101;
assign LUT_2[11619] = 32'b11111111111111111100001100000110;
assign LUT_2[11620] = 32'b11111111111111110100111000011001;
assign LUT_2[11621] = 32'b11111111111111110001110000110010;
assign LUT_2[11622] = 32'b11111111111111111011110001010101;
assign LUT_2[11623] = 32'b11111111111111111000101001101110;
assign LUT_2[11624] = 32'b11111111111111110011001100001110;
assign LUT_2[11625] = 32'b11111111111111110000000100100111;
assign LUT_2[11626] = 32'b11111111111111111010000101001010;
assign LUT_2[11627] = 32'b11111111111111110110111101100011;
assign LUT_2[11628] = 32'b11111111111111101111101001110110;
assign LUT_2[11629] = 32'b11111111111111101100100010001111;
assign LUT_2[11630] = 32'b11111111111111110110100010110010;
assign LUT_2[11631] = 32'b11111111111111110011011011001011;
assign LUT_2[11632] = 32'b11111111111111110010111110111011;
assign LUT_2[11633] = 32'b11111111111111101111110111010100;
assign LUT_2[11634] = 32'b11111111111111111001110111110111;
assign LUT_2[11635] = 32'b11111111111111110110110000010000;
assign LUT_2[11636] = 32'b11111111111111101111011100100011;
assign LUT_2[11637] = 32'b11111111111111101100010100111100;
assign LUT_2[11638] = 32'b11111111111111110110010101011111;
assign LUT_2[11639] = 32'b11111111111111110011001101111000;
assign LUT_2[11640] = 32'b11111111111111101101110000011000;
assign LUT_2[11641] = 32'b11111111111111101010101000110001;
assign LUT_2[11642] = 32'b11111111111111110100101001010100;
assign LUT_2[11643] = 32'b11111111111111110001100001101101;
assign LUT_2[11644] = 32'b11111111111111101010001110000000;
assign LUT_2[11645] = 32'b11111111111111100111000110011001;
assign LUT_2[11646] = 32'b11111111111111110001000110111100;
assign LUT_2[11647] = 32'b11111111111111101101111111010101;
assign LUT_2[11648] = 32'b00000000000000000100001010110100;
assign LUT_2[11649] = 32'b00000000000000000001000011001101;
assign LUT_2[11650] = 32'b00000000000000001011000011110000;
assign LUT_2[11651] = 32'b00000000000000000111111100001001;
assign LUT_2[11652] = 32'b00000000000000000000101000011100;
assign LUT_2[11653] = 32'b11111111111111111101100000110101;
assign LUT_2[11654] = 32'b00000000000000000111100001011000;
assign LUT_2[11655] = 32'b00000000000000000100011001110001;
assign LUT_2[11656] = 32'b11111111111111111110111100010001;
assign LUT_2[11657] = 32'b11111111111111111011110100101010;
assign LUT_2[11658] = 32'b00000000000000000101110101001101;
assign LUT_2[11659] = 32'b00000000000000000010101101100110;
assign LUT_2[11660] = 32'b11111111111111111011011001111001;
assign LUT_2[11661] = 32'b11111111111111111000010010010010;
assign LUT_2[11662] = 32'b00000000000000000010010010110101;
assign LUT_2[11663] = 32'b11111111111111111111001011001110;
assign LUT_2[11664] = 32'b11111111111111111110101110111110;
assign LUT_2[11665] = 32'b11111111111111111011100111010111;
assign LUT_2[11666] = 32'b00000000000000000101100111111010;
assign LUT_2[11667] = 32'b00000000000000000010100000010011;
assign LUT_2[11668] = 32'b11111111111111111011001100100110;
assign LUT_2[11669] = 32'b11111111111111111000000100111111;
assign LUT_2[11670] = 32'b00000000000000000010000101100010;
assign LUT_2[11671] = 32'b11111111111111111110111101111011;
assign LUT_2[11672] = 32'b11111111111111111001100000011011;
assign LUT_2[11673] = 32'b11111111111111110110011000110100;
assign LUT_2[11674] = 32'b00000000000000000000011001010111;
assign LUT_2[11675] = 32'b11111111111111111101010001110000;
assign LUT_2[11676] = 32'b11111111111111110101111110000011;
assign LUT_2[11677] = 32'b11111111111111110010110110011100;
assign LUT_2[11678] = 32'b11111111111111111100110110111111;
assign LUT_2[11679] = 32'b11111111111111111001101111011000;
assign LUT_2[11680] = 32'b00000000000000000100100110011101;
assign LUT_2[11681] = 32'b00000000000000000001011110110110;
assign LUT_2[11682] = 32'b00000000000000001011011111011001;
assign LUT_2[11683] = 32'b00000000000000001000010111110010;
assign LUT_2[11684] = 32'b00000000000000000001000100000101;
assign LUT_2[11685] = 32'b11111111111111111101111100011110;
assign LUT_2[11686] = 32'b00000000000000000111111101000001;
assign LUT_2[11687] = 32'b00000000000000000100110101011010;
assign LUT_2[11688] = 32'b11111111111111111111010111111010;
assign LUT_2[11689] = 32'b11111111111111111100010000010011;
assign LUT_2[11690] = 32'b00000000000000000110010000110110;
assign LUT_2[11691] = 32'b00000000000000000011001001001111;
assign LUT_2[11692] = 32'b11111111111111111011110101100010;
assign LUT_2[11693] = 32'b11111111111111111000101101111011;
assign LUT_2[11694] = 32'b00000000000000000010101110011110;
assign LUT_2[11695] = 32'b11111111111111111111100110110111;
assign LUT_2[11696] = 32'b11111111111111111111001010100111;
assign LUT_2[11697] = 32'b11111111111111111100000011000000;
assign LUT_2[11698] = 32'b00000000000000000110000011100011;
assign LUT_2[11699] = 32'b00000000000000000010111011111100;
assign LUT_2[11700] = 32'b11111111111111111011101000001111;
assign LUT_2[11701] = 32'b11111111111111111000100000101000;
assign LUT_2[11702] = 32'b00000000000000000010100001001011;
assign LUT_2[11703] = 32'b11111111111111111111011001100100;
assign LUT_2[11704] = 32'b11111111111111111001111100000100;
assign LUT_2[11705] = 32'b11111111111111110110110100011101;
assign LUT_2[11706] = 32'b00000000000000000000110101000000;
assign LUT_2[11707] = 32'b11111111111111111101101101011001;
assign LUT_2[11708] = 32'b11111111111111110110011001101100;
assign LUT_2[11709] = 32'b11111111111111110011010010000101;
assign LUT_2[11710] = 32'b11111111111111111101010010101000;
assign LUT_2[11711] = 32'b11111111111111111010001011000001;
assign LUT_2[11712] = 32'b11111111111111111100010011010111;
assign LUT_2[11713] = 32'b11111111111111111001001011110000;
assign LUT_2[11714] = 32'b00000000000000000011001100010011;
assign LUT_2[11715] = 32'b00000000000000000000000100101100;
assign LUT_2[11716] = 32'b11111111111111111000110000111111;
assign LUT_2[11717] = 32'b11111111111111110101101001011000;
assign LUT_2[11718] = 32'b11111111111111111111101001111011;
assign LUT_2[11719] = 32'b11111111111111111100100010010100;
assign LUT_2[11720] = 32'b11111111111111110111000100110100;
assign LUT_2[11721] = 32'b11111111111111110011111101001101;
assign LUT_2[11722] = 32'b11111111111111111101111101110000;
assign LUT_2[11723] = 32'b11111111111111111010110110001001;
assign LUT_2[11724] = 32'b11111111111111110011100010011100;
assign LUT_2[11725] = 32'b11111111111111110000011010110101;
assign LUT_2[11726] = 32'b11111111111111111010011011011000;
assign LUT_2[11727] = 32'b11111111111111110111010011110001;
assign LUT_2[11728] = 32'b11111111111111110110110111100001;
assign LUT_2[11729] = 32'b11111111111111110011101111111010;
assign LUT_2[11730] = 32'b11111111111111111101110000011101;
assign LUT_2[11731] = 32'b11111111111111111010101000110110;
assign LUT_2[11732] = 32'b11111111111111110011010101001001;
assign LUT_2[11733] = 32'b11111111111111110000001101100010;
assign LUT_2[11734] = 32'b11111111111111111010001110000101;
assign LUT_2[11735] = 32'b11111111111111110111000110011110;
assign LUT_2[11736] = 32'b11111111111111110001101000111110;
assign LUT_2[11737] = 32'b11111111111111101110100001010111;
assign LUT_2[11738] = 32'b11111111111111111000100001111010;
assign LUT_2[11739] = 32'b11111111111111110101011010010011;
assign LUT_2[11740] = 32'b11111111111111101110000110100110;
assign LUT_2[11741] = 32'b11111111111111101010111110111111;
assign LUT_2[11742] = 32'b11111111111111110100111111100010;
assign LUT_2[11743] = 32'b11111111111111110001110111111011;
assign LUT_2[11744] = 32'b11111111111111111100101111000000;
assign LUT_2[11745] = 32'b11111111111111111001100111011001;
assign LUT_2[11746] = 32'b00000000000000000011100111111100;
assign LUT_2[11747] = 32'b00000000000000000000100000010101;
assign LUT_2[11748] = 32'b11111111111111111001001100101000;
assign LUT_2[11749] = 32'b11111111111111110110000101000001;
assign LUT_2[11750] = 32'b00000000000000000000000101100100;
assign LUT_2[11751] = 32'b11111111111111111100111101111101;
assign LUT_2[11752] = 32'b11111111111111110111100000011101;
assign LUT_2[11753] = 32'b11111111111111110100011000110110;
assign LUT_2[11754] = 32'b11111111111111111110011001011001;
assign LUT_2[11755] = 32'b11111111111111111011010001110010;
assign LUT_2[11756] = 32'b11111111111111110011111110000101;
assign LUT_2[11757] = 32'b11111111111111110000110110011110;
assign LUT_2[11758] = 32'b11111111111111111010110111000001;
assign LUT_2[11759] = 32'b11111111111111110111101111011010;
assign LUT_2[11760] = 32'b11111111111111110111010011001010;
assign LUT_2[11761] = 32'b11111111111111110100001011100011;
assign LUT_2[11762] = 32'b11111111111111111110001100000110;
assign LUT_2[11763] = 32'b11111111111111111011000100011111;
assign LUT_2[11764] = 32'b11111111111111110011110000110010;
assign LUT_2[11765] = 32'b11111111111111110000101001001011;
assign LUT_2[11766] = 32'b11111111111111111010101001101110;
assign LUT_2[11767] = 32'b11111111111111110111100010000111;
assign LUT_2[11768] = 32'b11111111111111110010000100100111;
assign LUT_2[11769] = 32'b11111111111111101110111101000000;
assign LUT_2[11770] = 32'b11111111111111111000111101100011;
assign LUT_2[11771] = 32'b11111111111111110101110101111100;
assign LUT_2[11772] = 32'b11111111111111101110100010001111;
assign LUT_2[11773] = 32'b11111111111111101011011010101000;
assign LUT_2[11774] = 32'b11111111111111110101011011001011;
assign LUT_2[11775] = 32'b11111111111111110010010011100100;
assign LUT_2[11776] = 32'b00000000000000000000101001110001;
assign LUT_2[11777] = 32'b11111111111111111101100010001010;
assign LUT_2[11778] = 32'b00000000000000000111100010101101;
assign LUT_2[11779] = 32'b00000000000000000100011011000110;
assign LUT_2[11780] = 32'b11111111111111111101000111011001;
assign LUT_2[11781] = 32'b11111111111111111001111111110010;
assign LUT_2[11782] = 32'b00000000000000000100000000010101;
assign LUT_2[11783] = 32'b00000000000000000000111000101110;
assign LUT_2[11784] = 32'b11111111111111111011011011001110;
assign LUT_2[11785] = 32'b11111111111111111000010011100111;
assign LUT_2[11786] = 32'b00000000000000000010010100001010;
assign LUT_2[11787] = 32'b11111111111111111111001100100011;
assign LUT_2[11788] = 32'b11111111111111110111111000110110;
assign LUT_2[11789] = 32'b11111111111111110100110001001111;
assign LUT_2[11790] = 32'b11111111111111111110110001110010;
assign LUT_2[11791] = 32'b11111111111111111011101010001011;
assign LUT_2[11792] = 32'b11111111111111111011001101111011;
assign LUT_2[11793] = 32'b11111111111111111000000110010100;
assign LUT_2[11794] = 32'b00000000000000000010000110110111;
assign LUT_2[11795] = 32'b11111111111111111110111111010000;
assign LUT_2[11796] = 32'b11111111111111110111101011100011;
assign LUT_2[11797] = 32'b11111111111111110100100011111100;
assign LUT_2[11798] = 32'b11111111111111111110100100011111;
assign LUT_2[11799] = 32'b11111111111111111011011100111000;
assign LUT_2[11800] = 32'b11111111111111110101111111011000;
assign LUT_2[11801] = 32'b11111111111111110010110111110001;
assign LUT_2[11802] = 32'b11111111111111111100111000010100;
assign LUT_2[11803] = 32'b11111111111111111001110000101101;
assign LUT_2[11804] = 32'b11111111111111110010011101000000;
assign LUT_2[11805] = 32'b11111111111111101111010101011001;
assign LUT_2[11806] = 32'b11111111111111111001010101111100;
assign LUT_2[11807] = 32'b11111111111111110110001110010101;
assign LUT_2[11808] = 32'b00000000000000000001000101011010;
assign LUT_2[11809] = 32'b11111111111111111101111101110011;
assign LUT_2[11810] = 32'b00000000000000000111111110010110;
assign LUT_2[11811] = 32'b00000000000000000100110110101111;
assign LUT_2[11812] = 32'b11111111111111111101100011000010;
assign LUT_2[11813] = 32'b11111111111111111010011011011011;
assign LUT_2[11814] = 32'b00000000000000000100011011111110;
assign LUT_2[11815] = 32'b00000000000000000001010100010111;
assign LUT_2[11816] = 32'b11111111111111111011110110110111;
assign LUT_2[11817] = 32'b11111111111111111000101111010000;
assign LUT_2[11818] = 32'b00000000000000000010101111110011;
assign LUT_2[11819] = 32'b11111111111111111111101000001100;
assign LUT_2[11820] = 32'b11111111111111111000010100011111;
assign LUT_2[11821] = 32'b11111111111111110101001100111000;
assign LUT_2[11822] = 32'b11111111111111111111001101011011;
assign LUT_2[11823] = 32'b11111111111111111100000101110100;
assign LUT_2[11824] = 32'b11111111111111111011101001100100;
assign LUT_2[11825] = 32'b11111111111111111000100001111101;
assign LUT_2[11826] = 32'b00000000000000000010100010100000;
assign LUT_2[11827] = 32'b11111111111111111111011010111001;
assign LUT_2[11828] = 32'b11111111111111111000000111001100;
assign LUT_2[11829] = 32'b11111111111111110100111111100101;
assign LUT_2[11830] = 32'b11111111111111111111000000001000;
assign LUT_2[11831] = 32'b11111111111111111011111000100001;
assign LUT_2[11832] = 32'b11111111111111110110011011000001;
assign LUT_2[11833] = 32'b11111111111111110011010011011010;
assign LUT_2[11834] = 32'b11111111111111111101010011111101;
assign LUT_2[11835] = 32'b11111111111111111010001100010110;
assign LUT_2[11836] = 32'b11111111111111110010111000101001;
assign LUT_2[11837] = 32'b11111111111111101111110001000010;
assign LUT_2[11838] = 32'b11111111111111111001110001100101;
assign LUT_2[11839] = 32'b11111111111111110110101001111110;
assign LUT_2[11840] = 32'b11111111111111111000110010010100;
assign LUT_2[11841] = 32'b11111111111111110101101010101101;
assign LUT_2[11842] = 32'b11111111111111111111101011010000;
assign LUT_2[11843] = 32'b11111111111111111100100011101001;
assign LUT_2[11844] = 32'b11111111111111110101001111111100;
assign LUT_2[11845] = 32'b11111111111111110010001000010101;
assign LUT_2[11846] = 32'b11111111111111111100001000111000;
assign LUT_2[11847] = 32'b11111111111111111001000001010001;
assign LUT_2[11848] = 32'b11111111111111110011100011110001;
assign LUT_2[11849] = 32'b11111111111111110000011100001010;
assign LUT_2[11850] = 32'b11111111111111111010011100101101;
assign LUT_2[11851] = 32'b11111111111111110111010101000110;
assign LUT_2[11852] = 32'b11111111111111110000000001011001;
assign LUT_2[11853] = 32'b11111111111111101100111001110010;
assign LUT_2[11854] = 32'b11111111111111110110111010010101;
assign LUT_2[11855] = 32'b11111111111111110011110010101110;
assign LUT_2[11856] = 32'b11111111111111110011010110011110;
assign LUT_2[11857] = 32'b11111111111111110000001110110111;
assign LUT_2[11858] = 32'b11111111111111111010001111011010;
assign LUT_2[11859] = 32'b11111111111111110111000111110011;
assign LUT_2[11860] = 32'b11111111111111101111110100000110;
assign LUT_2[11861] = 32'b11111111111111101100101100011111;
assign LUT_2[11862] = 32'b11111111111111110110101101000010;
assign LUT_2[11863] = 32'b11111111111111110011100101011011;
assign LUT_2[11864] = 32'b11111111111111101110000111111011;
assign LUT_2[11865] = 32'b11111111111111101011000000010100;
assign LUT_2[11866] = 32'b11111111111111110101000000110111;
assign LUT_2[11867] = 32'b11111111111111110001111001010000;
assign LUT_2[11868] = 32'b11111111111111101010100101100011;
assign LUT_2[11869] = 32'b11111111111111100111011101111100;
assign LUT_2[11870] = 32'b11111111111111110001011110011111;
assign LUT_2[11871] = 32'b11111111111111101110010110111000;
assign LUT_2[11872] = 32'b11111111111111111001001101111101;
assign LUT_2[11873] = 32'b11111111111111110110000110010110;
assign LUT_2[11874] = 32'b00000000000000000000000110111001;
assign LUT_2[11875] = 32'b11111111111111111100111111010010;
assign LUT_2[11876] = 32'b11111111111111110101101011100101;
assign LUT_2[11877] = 32'b11111111111111110010100011111110;
assign LUT_2[11878] = 32'b11111111111111111100100100100001;
assign LUT_2[11879] = 32'b11111111111111111001011100111010;
assign LUT_2[11880] = 32'b11111111111111110011111111011010;
assign LUT_2[11881] = 32'b11111111111111110000110111110011;
assign LUT_2[11882] = 32'b11111111111111111010111000010110;
assign LUT_2[11883] = 32'b11111111111111110111110000101111;
assign LUT_2[11884] = 32'b11111111111111110000011101000010;
assign LUT_2[11885] = 32'b11111111111111101101010101011011;
assign LUT_2[11886] = 32'b11111111111111110111010101111110;
assign LUT_2[11887] = 32'b11111111111111110100001110010111;
assign LUT_2[11888] = 32'b11111111111111110011110010000111;
assign LUT_2[11889] = 32'b11111111111111110000101010100000;
assign LUT_2[11890] = 32'b11111111111111111010101011000011;
assign LUT_2[11891] = 32'b11111111111111110111100011011100;
assign LUT_2[11892] = 32'b11111111111111110000001111101111;
assign LUT_2[11893] = 32'b11111111111111101101001000001000;
assign LUT_2[11894] = 32'b11111111111111110111001000101011;
assign LUT_2[11895] = 32'b11111111111111110100000001000100;
assign LUT_2[11896] = 32'b11111111111111101110100011100100;
assign LUT_2[11897] = 32'b11111111111111101011011011111101;
assign LUT_2[11898] = 32'b11111111111111110101011100100000;
assign LUT_2[11899] = 32'b11111111111111110010010100111001;
assign LUT_2[11900] = 32'b11111111111111101011000001001100;
assign LUT_2[11901] = 32'b11111111111111100111111001100101;
assign LUT_2[11902] = 32'b11111111111111110001111010001000;
assign LUT_2[11903] = 32'b11111111111111101110110010100001;
assign LUT_2[11904] = 32'b00000000000000000100111110000000;
assign LUT_2[11905] = 32'b00000000000000000001110110011001;
assign LUT_2[11906] = 32'b00000000000000001011110110111100;
assign LUT_2[11907] = 32'b00000000000000001000101111010101;
assign LUT_2[11908] = 32'b00000000000000000001011011101000;
assign LUT_2[11909] = 32'b11111111111111111110010100000001;
assign LUT_2[11910] = 32'b00000000000000001000010100100100;
assign LUT_2[11911] = 32'b00000000000000000101001100111101;
assign LUT_2[11912] = 32'b11111111111111111111101111011101;
assign LUT_2[11913] = 32'b11111111111111111100100111110110;
assign LUT_2[11914] = 32'b00000000000000000110101000011001;
assign LUT_2[11915] = 32'b00000000000000000011100000110010;
assign LUT_2[11916] = 32'b11111111111111111100001101000101;
assign LUT_2[11917] = 32'b11111111111111111001000101011110;
assign LUT_2[11918] = 32'b00000000000000000011000110000001;
assign LUT_2[11919] = 32'b11111111111111111111111110011010;
assign LUT_2[11920] = 32'b11111111111111111111100010001010;
assign LUT_2[11921] = 32'b11111111111111111100011010100011;
assign LUT_2[11922] = 32'b00000000000000000110011011000110;
assign LUT_2[11923] = 32'b00000000000000000011010011011111;
assign LUT_2[11924] = 32'b11111111111111111011111111110010;
assign LUT_2[11925] = 32'b11111111111111111000111000001011;
assign LUT_2[11926] = 32'b00000000000000000010111000101110;
assign LUT_2[11927] = 32'b11111111111111111111110001000111;
assign LUT_2[11928] = 32'b11111111111111111010010011100111;
assign LUT_2[11929] = 32'b11111111111111110111001100000000;
assign LUT_2[11930] = 32'b00000000000000000001001100100011;
assign LUT_2[11931] = 32'b11111111111111111110000100111100;
assign LUT_2[11932] = 32'b11111111111111110110110001001111;
assign LUT_2[11933] = 32'b11111111111111110011101001101000;
assign LUT_2[11934] = 32'b11111111111111111101101010001011;
assign LUT_2[11935] = 32'b11111111111111111010100010100100;
assign LUT_2[11936] = 32'b00000000000000000101011001101001;
assign LUT_2[11937] = 32'b00000000000000000010010010000010;
assign LUT_2[11938] = 32'b00000000000000001100010010100101;
assign LUT_2[11939] = 32'b00000000000000001001001010111110;
assign LUT_2[11940] = 32'b00000000000000000001110111010001;
assign LUT_2[11941] = 32'b11111111111111111110101111101010;
assign LUT_2[11942] = 32'b00000000000000001000110000001101;
assign LUT_2[11943] = 32'b00000000000000000101101000100110;
assign LUT_2[11944] = 32'b00000000000000000000001011000110;
assign LUT_2[11945] = 32'b11111111111111111101000011011111;
assign LUT_2[11946] = 32'b00000000000000000111000100000010;
assign LUT_2[11947] = 32'b00000000000000000011111100011011;
assign LUT_2[11948] = 32'b11111111111111111100101000101110;
assign LUT_2[11949] = 32'b11111111111111111001100001000111;
assign LUT_2[11950] = 32'b00000000000000000011100001101010;
assign LUT_2[11951] = 32'b00000000000000000000011010000011;
assign LUT_2[11952] = 32'b11111111111111111111111101110011;
assign LUT_2[11953] = 32'b11111111111111111100110110001100;
assign LUT_2[11954] = 32'b00000000000000000110110110101111;
assign LUT_2[11955] = 32'b00000000000000000011101111001000;
assign LUT_2[11956] = 32'b11111111111111111100011011011011;
assign LUT_2[11957] = 32'b11111111111111111001010011110100;
assign LUT_2[11958] = 32'b00000000000000000011010100010111;
assign LUT_2[11959] = 32'b00000000000000000000001100110000;
assign LUT_2[11960] = 32'b11111111111111111010101111010000;
assign LUT_2[11961] = 32'b11111111111111110111100111101001;
assign LUT_2[11962] = 32'b00000000000000000001101000001100;
assign LUT_2[11963] = 32'b11111111111111111110100000100101;
assign LUT_2[11964] = 32'b11111111111111110111001100111000;
assign LUT_2[11965] = 32'b11111111111111110100000101010001;
assign LUT_2[11966] = 32'b11111111111111111110000101110100;
assign LUT_2[11967] = 32'b11111111111111111010111110001101;
assign LUT_2[11968] = 32'b11111111111111111101000110100011;
assign LUT_2[11969] = 32'b11111111111111111001111110111100;
assign LUT_2[11970] = 32'b00000000000000000011111111011111;
assign LUT_2[11971] = 32'b00000000000000000000110111111000;
assign LUT_2[11972] = 32'b11111111111111111001100100001011;
assign LUT_2[11973] = 32'b11111111111111110110011100100100;
assign LUT_2[11974] = 32'b00000000000000000000011101000111;
assign LUT_2[11975] = 32'b11111111111111111101010101100000;
assign LUT_2[11976] = 32'b11111111111111110111111000000000;
assign LUT_2[11977] = 32'b11111111111111110100110000011001;
assign LUT_2[11978] = 32'b11111111111111111110110000111100;
assign LUT_2[11979] = 32'b11111111111111111011101001010101;
assign LUT_2[11980] = 32'b11111111111111110100010101101000;
assign LUT_2[11981] = 32'b11111111111111110001001110000001;
assign LUT_2[11982] = 32'b11111111111111111011001110100100;
assign LUT_2[11983] = 32'b11111111111111111000000110111101;
assign LUT_2[11984] = 32'b11111111111111110111101010101101;
assign LUT_2[11985] = 32'b11111111111111110100100011000110;
assign LUT_2[11986] = 32'b11111111111111111110100011101001;
assign LUT_2[11987] = 32'b11111111111111111011011100000010;
assign LUT_2[11988] = 32'b11111111111111110100001000010101;
assign LUT_2[11989] = 32'b11111111111111110001000000101110;
assign LUT_2[11990] = 32'b11111111111111111011000001010001;
assign LUT_2[11991] = 32'b11111111111111110111111001101010;
assign LUT_2[11992] = 32'b11111111111111110010011100001010;
assign LUT_2[11993] = 32'b11111111111111101111010100100011;
assign LUT_2[11994] = 32'b11111111111111111001010101000110;
assign LUT_2[11995] = 32'b11111111111111110110001101011111;
assign LUT_2[11996] = 32'b11111111111111101110111001110010;
assign LUT_2[11997] = 32'b11111111111111101011110010001011;
assign LUT_2[11998] = 32'b11111111111111110101110010101110;
assign LUT_2[11999] = 32'b11111111111111110010101011000111;
assign LUT_2[12000] = 32'b11111111111111111101100010001100;
assign LUT_2[12001] = 32'b11111111111111111010011010100101;
assign LUT_2[12002] = 32'b00000000000000000100011011001000;
assign LUT_2[12003] = 32'b00000000000000000001010011100001;
assign LUT_2[12004] = 32'b11111111111111111001111111110100;
assign LUT_2[12005] = 32'b11111111111111110110111000001101;
assign LUT_2[12006] = 32'b00000000000000000000111000110000;
assign LUT_2[12007] = 32'b11111111111111111101110001001001;
assign LUT_2[12008] = 32'b11111111111111111000010011101001;
assign LUT_2[12009] = 32'b11111111111111110101001100000010;
assign LUT_2[12010] = 32'b11111111111111111111001100100101;
assign LUT_2[12011] = 32'b11111111111111111100000100111110;
assign LUT_2[12012] = 32'b11111111111111110100110001010001;
assign LUT_2[12013] = 32'b11111111111111110001101001101010;
assign LUT_2[12014] = 32'b11111111111111111011101010001101;
assign LUT_2[12015] = 32'b11111111111111111000100010100110;
assign LUT_2[12016] = 32'b11111111111111111000000110010110;
assign LUT_2[12017] = 32'b11111111111111110100111110101111;
assign LUT_2[12018] = 32'b11111111111111111110111111010010;
assign LUT_2[12019] = 32'b11111111111111111011110111101011;
assign LUT_2[12020] = 32'b11111111111111110100100011111110;
assign LUT_2[12021] = 32'b11111111111111110001011100010111;
assign LUT_2[12022] = 32'b11111111111111111011011100111010;
assign LUT_2[12023] = 32'b11111111111111111000010101010011;
assign LUT_2[12024] = 32'b11111111111111110010110111110011;
assign LUT_2[12025] = 32'b11111111111111101111110000001100;
assign LUT_2[12026] = 32'b11111111111111111001110000101111;
assign LUT_2[12027] = 32'b11111111111111110110101001001000;
assign LUT_2[12028] = 32'b11111111111111101111010101011011;
assign LUT_2[12029] = 32'b11111111111111101100001101110100;
assign LUT_2[12030] = 32'b11111111111111110110001110010111;
assign LUT_2[12031] = 32'b11111111111111110011000110110000;
assign LUT_2[12032] = 32'b00000000000000000100101000010111;
assign LUT_2[12033] = 32'b00000000000000000001100000110000;
assign LUT_2[12034] = 32'b00000000000000001011100001010011;
assign LUT_2[12035] = 32'b00000000000000001000011001101100;
assign LUT_2[12036] = 32'b00000000000000000001000101111111;
assign LUT_2[12037] = 32'b11111111111111111101111110011000;
assign LUT_2[12038] = 32'b00000000000000000111111110111011;
assign LUT_2[12039] = 32'b00000000000000000100110111010100;
assign LUT_2[12040] = 32'b11111111111111111111011001110100;
assign LUT_2[12041] = 32'b11111111111111111100010010001101;
assign LUT_2[12042] = 32'b00000000000000000110010010110000;
assign LUT_2[12043] = 32'b00000000000000000011001011001001;
assign LUT_2[12044] = 32'b11111111111111111011110111011100;
assign LUT_2[12045] = 32'b11111111111111111000101111110101;
assign LUT_2[12046] = 32'b00000000000000000010110000011000;
assign LUT_2[12047] = 32'b11111111111111111111101000110001;
assign LUT_2[12048] = 32'b11111111111111111111001100100001;
assign LUT_2[12049] = 32'b11111111111111111100000100111010;
assign LUT_2[12050] = 32'b00000000000000000110000101011101;
assign LUT_2[12051] = 32'b00000000000000000010111101110110;
assign LUT_2[12052] = 32'b11111111111111111011101010001001;
assign LUT_2[12053] = 32'b11111111111111111000100010100010;
assign LUT_2[12054] = 32'b00000000000000000010100011000101;
assign LUT_2[12055] = 32'b11111111111111111111011011011110;
assign LUT_2[12056] = 32'b11111111111111111001111101111110;
assign LUT_2[12057] = 32'b11111111111111110110110110010111;
assign LUT_2[12058] = 32'b00000000000000000000110110111010;
assign LUT_2[12059] = 32'b11111111111111111101101111010011;
assign LUT_2[12060] = 32'b11111111111111110110011011100110;
assign LUT_2[12061] = 32'b11111111111111110011010011111111;
assign LUT_2[12062] = 32'b11111111111111111101010100100010;
assign LUT_2[12063] = 32'b11111111111111111010001100111011;
assign LUT_2[12064] = 32'b00000000000000000101000100000000;
assign LUT_2[12065] = 32'b00000000000000000001111100011001;
assign LUT_2[12066] = 32'b00000000000000001011111100111100;
assign LUT_2[12067] = 32'b00000000000000001000110101010101;
assign LUT_2[12068] = 32'b00000000000000000001100001101000;
assign LUT_2[12069] = 32'b11111111111111111110011010000001;
assign LUT_2[12070] = 32'b00000000000000001000011010100100;
assign LUT_2[12071] = 32'b00000000000000000101010010111101;
assign LUT_2[12072] = 32'b11111111111111111111110101011101;
assign LUT_2[12073] = 32'b11111111111111111100101101110110;
assign LUT_2[12074] = 32'b00000000000000000110101110011001;
assign LUT_2[12075] = 32'b00000000000000000011100110110010;
assign LUT_2[12076] = 32'b11111111111111111100010011000101;
assign LUT_2[12077] = 32'b11111111111111111001001011011110;
assign LUT_2[12078] = 32'b00000000000000000011001100000001;
assign LUT_2[12079] = 32'b00000000000000000000000100011010;
assign LUT_2[12080] = 32'b11111111111111111111101000001010;
assign LUT_2[12081] = 32'b11111111111111111100100000100011;
assign LUT_2[12082] = 32'b00000000000000000110100001000110;
assign LUT_2[12083] = 32'b00000000000000000011011001011111;
assign LUT_2[12084] = 32'b11111111111111111100000101110010;
assign LUT_2[12085] = 32'b11111111111111111000111110001011;
assign LUT_2[12086] = 32'b00000000000000000010111110101110;
assign LUT_2[12087] = 32'b11111111111111111111110111000111;
assign LUT_2[12088] = 32'b11111111111111111010011001100111;
assign LUT_2[12089] = 32'b11111111111111110111010010000000;
assign LUT_2[12090] = 32'b00000000000000000001010010100011;
assign LUT_2[12091] = 32'b11111111111111111110001010111100;
assign LUT_2[12092] = 32'b11111111111111110110110111001111;
assign LUT_2[12093] = 32'b11111111111111110011101111101000;
assign LUT_2[12094] = 32'b11111111111111111101110000001011;
assign LUT_2[12095] = 32'b11111111111111111010101000100100;
assign LUT_2[12096] = 32'b11111111111111111100110000111010;
assign LUT_2[12097] = 32'b11111111111111111001101001010011;
assign LUT_2[12098] = 32'b00000000000000000011101001110110;
assign LUT_2[12099] = 32'b00000000000000000000100010001111;
assign LUT_2[12100] = 32'b11111111111111111001001110100010;
assign LUT_2[12101] = 32'b11111111111111110110000110111011;
assign LUT_2[12102] = 32'b00000000000000000000000111011110;
assign LUT_2[12103] = 32'b11111111111111111100111111110111;
assign LUT_2[12104] = 32'b11111111111111110111100010010111;
assign LUT_2[12105] = 32'b11111111111111110100011010110000;
assign LUT_2[12106] = 32'b11111111111111111110011011010011;
assign LUT_2[12107] = 32'b11111111111111111011010011101100;
assign LUT_2[12108] = 32'b11111111111111110011111111111111;
assign LUT_2[12109] = 32'b11111111111111110000111000011000;
assign LUT_2[12110] = 32'b11111111111111111010111000111011;
assign LUT_2[12111] = 32'b11111111111111110111110001010100;
assign LUT_2[12112] = 32'b11111111111111110111010101000100;
assign LUT_2[12113] = 32'b11111111111111110100001101011101;
assign LUT_2[12114] = 32'b11111111111111111110001110000000;
assign LUT_2[12115] = 32'b11111111111111111011000110011001;
assign LUT_2[12116] = 32'b11111111111111110011110010101100;
assign LUT_2[12117] = 32'b11111111111111110000101011000101;
assign LUT_2[12118] = 32'b11111111111111111010101011101000;
assign LUT_2[12119] = 32'b11111111111111110111100100000001;
assign LUT_2[12120] = 32'b11111111111111110010000110100001;
assign LUT_2[12121] = 32'b11111111111111101110111110111010;
assign LUT_2[12122] = 32'b11111111111111111000111111011101;
assign LUT_2[12123] = 32'b11111111111111110101110111110110;
assign LUT_2[12124] = 32'b11111111111111101110100100001001;
assign LUT_2[12125] = 32'b11111111111111101011011100100010;
assign LUT_2[12126] = 32'b11111111111111110101011101000101;
assign LUT_2[12127] = 32'b11111111111111110010010101011110;
assign LUT_2[12128] = 32'b11111111111111111101001100100011;
assign LUT_2[12129] = 32'b11111111111111111010000100111100;
assign LUT_2[12130] = 32'b00000000000000000100000101011111;
assign LUT_2[12131] = 32'b00000000000000000000111101111000;
assign LUT_2[12132] = 32'b11111111111111111001101010001011;
assign LUT_2[12133] = 32'b11111111111111110110100010100100;
assign LUT_2[12134] = 32'b00000000000000000000100011000111;
assign LUT_2[12135] = 32'b11111111111111111101011011100000;
assign LUT_2[12136] = 32'b11111111111111110111111110000000;
assign LUT_2[12137] = 32'b11111111111111110100110110011001;
assign LUT_2[12138] = 32'b11111111111111111110110110111100;
assign LUT_2[12139] = 32'b11111111111111111011101111010101;
assign LUT_2[12140] = 32'b11111111111111110100011011101000;
assign LUT_2[12141] = 32'b11111111111111110001010100000001;
assign LUT_2[12142] = 32'b11111111111111111011010100100100;
assign LUT_2[12143] = 32'b11111111111111111000001100111101;
assign LUT_2[12144] = 32'b11111111111111110111110000101101;
assign LUT_2[12145] = 32'b11111111111111110100101001000110;
assign LUT_2[12146] = 32'b11111111111111111110101001101001;
assign LUT_2[12147] = 32'b11111111111111111011100010000010;
assign LUT_2[12148] = 32'b11111111111111110100001110010101;
assign LUT_2[12149] = 32'b11111111111111110001000110101110;
assign LUT_2[12150] = 32'b11111111111111111011000111010001;
assign LUT_2[12151] = 32'b11111111111111110111111111101010;
assign LUT_2[12152] = 32'b11111111111111110010100010001010;
assign LUT_2[12153] = 32'b11111111111111101111011010100011;
assign LUT_2[12154] = 32'b11111111111111111001011011000110;
assign LUT_2[12155] = 32'b11111111111111110110010011011111;
assign LUT_2[12156] = 32'b11111111111111101110111111110010;
assign LUT_2[12157] = 32'b11111111111111101011111000001011;
assign LUT_2[12158] = 32'b11111111111111110101111000101110;
assign LUT_2[12159] = 32'b11111111111111110010110001000111;
assign LUT_2[12160] = 32'b00000000000000001000111100100110;
assign LUT_2[12161] = 32'b00000000000000000101110100111111;
assign LUT_2[12162] = 32'b00000000000000001111110101100010;
assign LUT_2[12163] = 32'b00000000000000001100101101111011;
assign LUT_2[12164] = 32'b00000000000000000101011010001110;
assign LUT_2[12165] = 32'b00000000000000000010010010100111;
assign LUT_2[12166] = 32'b00000000000000001100010011001010;
assign LUT_2[12167] = 32'b00000000000000001001001011100011;
assign LUT_2[12168] = 32'b00000000000000000011101110000011;
assign LUT_2[12169] = 32'b00000000000000000000100110011100;
assign LUT_2[12170] = 32'b00000000000000001010100110111111;
assign LUT_2[12171] = 32'b00000000000000000111011111011000;
assign LUT_2[12172] = 32'b00000000000000000000001011101011;
assign LUT_2[12173] = 32'b11111111111111111101000100000100;
assign LUT_2[12174] = 32'b00000000000000000111000100100111;
assign LUT_2[12175] = 32'b00000000000000000011111101000000;
assign LUT_2[12176] = 32'b00000000000000000011100000110000;
assign LUT_2[12177] = 32'b00000000000000000000011001001001;
assign LUT_2[12178] = 32'b00000000000000001010011001101100;
assign LUT_2[12179] = 32'b00000000000000000111010010000101;
assign LUT_2[12180] = 32'b11111111111111111111111110011000;
assign LUT_2[12181] = 32'b11111111111111111100110110110001;
assign LUT_2[12182] = 32'b00000000000000000110110111010100;
assign LUT_2[12183] = 32'b00000000000000000011101111101101;
assign LUT_2[12184] = 32'b11111111111111111110010010001101;
assign LUT_2[12185] = 32'b11111111111111111011001010100110;
assign LUT_2[12186] = 32'b00000000000000000101001011001001;
assign LUT_2[12187] = 32'b00000000000000000010000011100010;
assign LUT_2[12188] = 32'b11111111111111111010101111110101;
assign LUT_2[12189] = 32'b11111111111111110111101000001110;
assign LUT_2[12190] = 32'b00000000000000000001101000110001;
assign LUT_2[12191] = 32'b11111111111111111110100001001010;
assign LUT_2[12192] = 32'b00000000000000001001011000001111;
assign LUT_2[12193] = 32'b00000000000000000110010000101000;
assign LUT_2[12194] = 32'b00000000000000010000010001001011;
assign LUT_2[12195] = 32'b00000000000000001101001001100100;
assign LUT_2[12196] = 32'b00000000000000000101110101110111;
assign LUT_2[12197] = 32'b00000000000000000010101110010000;
assign LUT_2[12198] = 32'b00000000000000001100101110110011;
assign LUT_2[12199] = 32'b00000000000000001001100111001100;
assign LUT_2[12200] = 32'b00000000000000000100001001101100;
assign LUT_2[12201] = 32'b00000000000000000001000010000101;
assign LUT_2[12202] = 32'b00000000000000001011000010101000;
assign LUT_2[12203] = 32'b00000000000000000111111011000001;
assign LUT_2[12204] = 32'b00000000000000000000100111010100;
assign LUT_2[12205] = 32'b11111111111111111101011111101101;
assign LUT_2[12206] = 32'b00000000000000000111100000010000;
assign LUT_2[12207] = 32'b00000000000000000100011000101001;
assign LUT_2[12208] = 32'b00000000000000000011111100011001;
assign LUT_2[12209] = 32'b00000000000000000000110100110010;
assign LUT_2[12210] = 32'b00000000000000001010110101010101;
assign LUT_2[12211] = 32'b00000000000000000111101101101110;
assign LUT_2[12212] = 32'b00000000000000000000011010000001;
assign LUT_2[12213] = 32'b11111111111111111101010010011010;
assign LUT_2[12214] = 32'b00000000000000000111010010111101;
assign LUT_2[12215] = 32'b00000000000000000100001011010110;
assign LUT_2[12216] = 32'b11111111111111111110101101110110;
assign LUT_2[12217] = 32'b11111111111111111011100110001111;
assign LUT_2[12218] = 32'b00000000000000000101100110110010;
assign LUT_2[12219] = 32'b00000000000000000010011111001011;
assign LUT_2[12220] = 32'b11111111111111111011001011011110;
assign LUT_2[12221] = 32'b11111111111111111000000011110111;
assign LUT_2[12222] = 32'b00000000000000000010000100011010;
assign LUT_2[12223] = 32'b11111111111111111110111100110011;
assign LUT_2[12224] = 32'b00000000000000000001000101001001;
assign LUT_2[12225] = 32'b11111111111111111101111101100010;
assign LUT_2[12226] = 32'b00000000000000000111111110000101;
assign LUT_2[12227] = 32'b00000000000000000100110110011110;
assign LUT_2[12228] = 32'b11111111111111111101100010110001;
assign LUT_2[12229] = 32'b11111111111111111010011011001010;
assign LUT_2[12230] = 32'b00000000000000000100011011101101;
assign LUT_2[12231] = 32'b00000000000000000001010100000110;
assign LUT_2[12232] = 32'b11111111111111111011110110100110;
assign LUT_2[12233] = 32'b11111111111111111000101110111111;
assign LUT_2[12234] = 32'b00000000000000000010101111100010;
assign LUT_2[12235] = 32'b11111111111111111111100111111011;
assign LUT_2[12236] = 32'b11111111111111111000010100001110;
assign LUT_2[12237] = 32'b11111111111111110101001100100111;
assign LUT_2[12238] = 32'b11111111111111111111001101001010;
assign LUT_2[12239] = 32'b11111111111111111100000101100011;
assign LUT_2[12240] = 32'b11111111111111111011101001010011;
assign LUT_2[12241] = 32'b11111111111111111000100001101100;
assign LUT_2[12242] = 32'b00000000000000000010100010001111;
assign LUT_2[12243] = 32'b11111111111111111111011010101000;
assign LUT_2[12244] = 32'b11111111111111111000000110111011;
assign LUT_2[12245] = 32'b11111111111111110100111111010100;
assign LUT_2[12246] = 32'b11111111111111111110111111110111;
assign LUT_2[12247] = 32'b11111111111111111011111000010000;
assign LUT_2[12248] = 32'b11111111111111110110011010110000;
assign LUT_2[12249] = 32'b11111111111111110011010011001001;
assign LUT_2[12250] = 32'b11111111111111111101010011101100;
assign LUT_2[12251] = 32'b11111111111111111010001100000101;
assign LUT_2[12252] = 32'b11111111111111110010111000011000;
assign LUT_2[12253] = 32'b11111111111111101111110000110001;
assign LUT_2[12254] = 32'b11111111111111111001110001010100;
assign LUT_2[12255] = 32'b11111111111111110110101001101101;
assign LUT_2[12256] = 32'b00000000000000000001100000110010;
assign LUT_2[12257] = 32'b11111111111111111110011001001011;
assign LUT_2[12258] = 32'b00000000000000001000011001101110;
assign LUT_2[12259] = 32'b00000000000000000101010010000111;
assign LUT_2[12260] = 32'b11111111111111111101111110011010;
assign LUT_2[12261] = 32'b11111111111111111010110110110011;
assign LUT_2[12262] = 32'b00000000000000000100110111010110;
assign LUT_2[12263] = 32'b00000000000000000001101111101111;
assign LUT_2[12264] = 32'b11111111111111111100010010001111;
assign LUT_2[12265] = 32'b11111111111111111001001010101000;
assign LUT_2[12266] = 32'b00000000000000000011001011001011;
assign LUT_2[12267] = 32'b00000000000000000000000011100100;
assign LUT_2[12268] = 32'b11111111111111111000101111110111;
assign LUT_2[12269] = 32'b11111111111111110101101000010000;
assign LUT_2[12270] = 32'b11111111111111111111101000110011;
assign LUT_2[12271] = 32'b11111111111111111100100001001100;
assign LUT_2[12272] = 32'b11111111111111111100000100111100;
assign LUT_2[12273] = 32'b11111111111111111000111101010101;
assign LUT_2[12274] = 32'b00000000000000000010111101111000;
assign LUT_2[12275] = 32'b11111111111111111111110110010001;
assign LUT_2[12276] = 32'b11111111111111111000100010100100;
assign LUT_2[12277] = 32'b11111111111111110101011010111101;
assign LUT_2[12278] = 32'b11111111111111111111011011100000;
assign LUT_2[12279] = 32'b11111111111111111100010011111001;
assign LUT_2[12280] = 32'b11111111111111110110110110011001;
assign LUT_2[12281] = 32'b11111111111111110011101110110010;
assign LUT_2[12282] = 32'b11111111111111111101101111010101;
assign LUT_2[12283] = 32'b11111111111111111010100111101110;
assign LUT_2[12284] = 32'b11111111111111110011010100000001;
assign LUT_2[12285] = 32'b11111111111111110000001100011010;
assign LUT_2[12286] = 32'b11111111111111111010001100111101;
assign LUT_2[12287] = 32'b11111111111111110111000101010110;
assign LUT_2[12288] = 32'b11111111111111111000011010001001;
assign LUT_2[12289] = 32'b11111111111111110101010010100010;
assign LUT_2[12290] = 32'b11111111111111111111010011000101;
assign LUT_2[12291] = 32'b11111111111111111100001011011110;
assign LUT_2[12292] = 32'b11111111111111110100110111110001;
assign LUT_2[12293] = 32'b11111111111111110001110000001010;
assign LUT_2[12294] = 32'b11111111111111111011110000101101;
assign LUT_2[12295] = 32'b11111111111111111000101001000110;
assign LUT_2[12296] = 32'b11111111111111110011001011100110;
assign LUT_2[12297] = 32'b11111111111111110000000011111111;
assign LUT_2[12298] = 32'b11111111111111111010000100100010;
assign LUT_2[12299] = 32'b11111111111111110110111100111011;
assign LUT_2[12300] = 32'b11111111111111101111101001001110;
assign LUT_2[12301] = 32'b11111111111111101100100001100111;
assign LUT_2[12302] = 32'b11111111111111110110100010001010;
assign LUT_2[12303] = 32'b11111111111111110011011010100011;
assign LUT_2[12304] = 32'b11111111111111110010111110010011;
assign LUT_2[12305] = 32'b11111111111111101111110110101100;
assign LUT_2[12306] = 32'b11111111111111111001110111001111;
assign LUT_2[12307] = 32'b11111111111111110110101111101000;
assign LUT_2[12308] = 32'b11111111111111101111011011111011;
assign LUT_2[12309] = 32'b11111111111111101100010100010100;
assign LUT_2[12310] = 32'b11111111111111110110010100110111;
assign LUT_2[12311] = 32'b11111111111111110011001101010000;
assign LUT_2[12312] = 32'b11111111111111101101101111110000;
assign LUT_2[12313] = 32'b11111111111111101010101000001001;
assign LUT_2[12314] = 32'b11111111111111110100101000101100;
assign LUT_2[12315] = 32'b11111111111111110001100001000101;
assign LUT_2[12316] = 32'b11111111111111101010001101011000;
assign LUT_2[12317] = 32'b11111111111111100111000101110001;
assign LUT_2[12318] = 32'b11111111111111110001000110010100;
assign LUT_2[12319] = 32'b11111111111111101101111110101101;
assign LUT_2[12320] = 32'b11111111111111111000110101110010;
assign LUT_2[12321] = 32'b11111111111111110101101110001011;
assign LUT_2[12322] = 32'b11111111111111111111101110101110;
assign LUT_2[12323] = 32'b11111111111111111100100111000111;
assign LUT_2[12324] = 32'b11111111111111110101010011011010;
assign LUT_2[12325] = 32'b11111111111111110010001011110011;
assign LUT_2[12326] = 32'b11111111111111111100001100010110;
assign LUT_2[12327] = 32'b11111111111111111001000100101111;
assign LUT_2[12328] = 32'b11111111111111110011100111001111;
assign LUT_2[12329] = 32'b11111111111111110000011111101000;
assign LUT_2[12330] = 32'b11111111111111111010100000001011;
assign LUT_2[12331] = 32'b11111111111111110111011000100100;
assign LUT_2[12332] = 32'b11111111111111110000000100110111;
assign LUT_2[12333] = 32'b11111111111111101100111101010000;
assign LUT_2[12334] = 32'b11111111111111110110111101110011;
assign LUT_2[12335] = 32'b11111111111111110011110110001100;
assign LUT_2[12336] = 32'b11111111111111110011011001111100;
assign LUT_2[12337] = 32'b11111111111111110000010010010101;
assign LUT_2[12338] = 32'b11111111111111111010010010111000;
assign LUT_2[12339] = 32'b11111111111111110111001011010001;
assign LUT_2[12340] = 32'b11111111111111101111110111100100;
assign LUT_2[12341] = 32'b11111111111111101100101111111101;
assign LUT_2[12342] = 32'b11111111111111110110110000100000;
assign LUT_2[12343] = 32'b11111111111111110011101000111001;
assign LUT_2[12344] = 32'b11111111111111101110001011011001;
assign LUT_2[12345] = 32'b11111111111111101011000011110010;
assign LUT_2[12346] = 32'b11111111111111110101000100010101;
assign LUT_2[12347] = 32'b11111111111111110001111100101110;
assign LUT_2[12348] = 32'b11111111111111101010101001000001;
assign LUT_2[12349] = 32'b11111111111111100111100001011010;
assign LUT_2[12350] = 32'b11111111111111110001100001111101;
assign LUT_2[12351] = 32'b11111111111111101110011010010110;
assign LUT_2[12352] = 32'b11111111111111110000100010101100;
assign LUT_2[12353] = 32'b11111111111111101101011011000101;
assign LUT_2[12354] = 32'b11111111111111110111011011101000;
assign LUT_2[12355] = 32'b11111111111111110100010100000001;
assign LUT_2[12356] = 32'b11111111111111101101000000010100;
assign LUT_2[12357] = 32'b11111111111111101001111000101101;
assign LUT_2[12358] = 32'b11111111111111110011111001010000;
assign LUT_2[12359] = 32'b11111111111111110000110001101001;
assign LUT_2[12360] = 32'b11111111111111101011010100001001;
assign LUT_2[12361] = 32'b11111111111111101000001100100010;
assign LUT_2[12362] = 32'b11111111111111110010001101000101;
assign LUT_2[12363] = 32'b11111111111111101111000101011110;
assign LUT_2[12364] = 32'b11111111111111100111110001110001;
assign LUT_2[12365] = 32'b11111111111111100100101010001010;
assign LUT_2[12366] = 32'b11111111111111101110101010101101;
assign LUT_2[12367] = 32'b11111111111111101011100011000110;
assign LUT_2[12368] = 32'b11111111111111101011000110110110;
assign LUT_2[12369] = 32'b11111111111111100111111111001111;
assign LUT_2[12370] = 32'b11111111111111110001111111110010;
assign LUT_2[12371] = 32'b11111111111111101110111000001011;
assign LUT_2[12372] = 32'b11111111111111100111100100011110;
assign LUT_2[12373] = 32'b11111111111111100100011100110111;
assign LUT_2[12374] = 32'b11111111111111101110011101011010;
assign LUT_2[12375] = 32'b11111111111111101011010101110011;
assign LUT_2[12376] = 32'b11111111111111100101111000010011;
assign LUT_2[12377] = 32'b11111111111111100010110000101100;
assign LUT_2[12378] = 32'b11111111111111101100110001001111;
assign LUT_2[12379] = 32'b11111111111111101001101001101000;
assign LUT_2[12380] = 32'b11111111111111100010010101111011;
assign LUT_2[12381] = 32'b11111111111111011111001110010100;
assign LUT_2[12382] = 32'b11111111111111101001001110110111;
assign LUT_2[12383] = 32'b11111111111111100110000111010000;
assign LUT_2[12384] = 32'b11111111111111110000111110010101;
assign LUT_2[12385] = 32'b11111111111111101101110110101110;
assign LUT_2[12386] = 32'b11111111111111110111110111010001;
assign LUT_2[12387] = 32'b11111111111111110100101111101010;
assign LUT_2[12388] = 32'b11111111111111101101011011111101;
assign LUT_2[12389] = 32'b11111111111111101010010100010110;
assign LUT_2[12390] = 32'b11111111111111110100010100111001;
assign LUT_2[12391] = 32'b11111111111111110001001101010010;
assign LUT_2[12392] = 32'b11111111111111101011101111110010;
assign LUT_2[12393] = 32'b11111111111111101000101000001011;
assign LUT_2[12394] = 32'b11111111111111110010101000101110;
assign LUT_2[12395] = 32'b11111111111111101111100001000111;
assign LUT_2[12396] = 32'b11111111111111101000001101011010;
assign LUT_2[12397] = 32'b11111111111111100101000101110011;
assign LUT_2[12398] = 32'b11111111111111101111000110010110;
assign LUT_2[12399] = 32'b11111111111111101011111110101111;
assign LUT_2[12400] = 32'b11111111111111101011100010011111;
assign LUT_2[12401] = 32'b11111111111111101000011010111000;
assign LUT_2[12402] = 32'b11111111111111110010011011011011;
assign LUT_2[12403] = 32'b11111111111111101111010011110100;
assign LUT_2[12404] = 32'b11111111111111101000000000000111;
assign LUT_2[12405] = 32'b11111111111111100100111000100000;
assign LUT_2[12406] = 32'b11111111111111101110111001000011;
assign LUT_2[12407] = 32'b11111111111111101011110001011100;
assign LUT_2[12408] = 32'b11111111111111100110010011111100;
assign LUT_2[12409] = 32'b11111111111111100011001100010101;
assign LUT_2[12410] = 32'b11111111111111101101001100111000;
assign LUT_2[12411] = 32'b11111111111111101010000101010001;
assign LUT_2[12412] = 32'b11111111111111100010110001100100;
assign LUT_2[12413] = 32'b11111111111111011111101001111101;
assign LUT_2[12414] = 32'b11111111111111101001101010100000;
assign LUT_2[12415] = 32'b11111111111111100110100010111001;
assign LUT_2[12416] = 32'b11111111111111111100101110011000;
assign LUT_2[12417] = 32'b11111111111111111001100110110001;
assign LUT_2[12418] = 32'b00000000000000000011100111010100;
assign LUT_2[12419] = 32'b00000000000000000000011111101101;
assign LUT_2[12420] = 32'b11111111111111111001001100000000;
assign LUT_2[12421] = 32'b11111111111111110110000100011001;
assign LUT_2[12422] = 32'b00000000000000000000000100111100;
assign LUT_2[12423] = 32'b11111111111111111100111101010101;
assign LUT_2[12424] = 32'b11111111111111110111011111110101;
assign LUT_2[12425] = 32'b11111111111111110100011000001110;
assign LUT_2[12426] = 32'b11111111111111111110011000110001;
assign LUT_2[12427] = 32'b11111111111111111011010001001010;
assign LUT_2[12428] = 32'b11111111111111110011111101011101;
assign LUT_2[12429] = 32'b11111111111111110000110101110110;
assign LUT_2[12430] = 32'b11111111111111111010110110011001;
assign LUT_2[12431] = 32'b11111111111111110111101110110010;
assign LUT_2[12432] = 32'b11111111111111110111010010100010;
assign LUT_2[12433] = 32'b11111111111111110100001010111011;
assign LUT_2[12434] = 32'b11111111111111111110001011011110;
assign LUT_2[12435] = 32'b11111111111111111011000011110111;
assign LUT_2[12436] = 32'b11111111111111110011110000001010;
assign LUT_2[12437] = 32'b11111111111111110000101000100011;
assign LUT_2[12438] = 32'b11111111111111111010101001000110;
assign LUT_2[12439] = 32'b11111111111111110111100001011111;
assign LUT_2[12440] = 32'b11111111111111110010000011111111;
assign LUT_2[12441] = 32'b11111111111111101110111100011000;
assign LUT_2[12442] = 32'b11111111111111111000111100111011;
assign LUT_2[12443] = 32'b11111111111111110101110101010100;
assign LUT_2[12444] = 32'b11111111111111101110100001100111;
assign LUT_2[12445] = 32'b11111111111111101011011010000000;
assign LUT_2[12446] = 32'b11111111111111110101011010100011;
assign LUT_2[12447] = 32'b11111111111111110010010010111100;
assign LUT_2[12448] = 32'b11111111111111111101001010000001;
assign LUT_2[12449] = 32'b11111111111111111010000010011010;
assign LUT_2[12450] = 32'b00000000000000000100000010111101;
assign LUT_2[12451] = 32'b00000000000000000000111011010110;
assign LUT_2[12452] = 32'b11111111111111111001100111101001;
assign LUT_2[12453] = 32'b11111111111111110110100000000010;
assign LUT_2[12454] = 32'b00000000000000000000100000100101;
assign LUT_2[12455] = 32'b11111111111111111101011000111110;
assign LUT_2[12456] = 32'b11111111111111110111111011011110;
assign LUT_2[12457] = 32'b11111111111111110100110011110111;
assign LUT_2[12458] = 32'b11111111111111111110110100011010;
assign LUT_2[12459] = 32'b11111111111111111011101100110011;
assign LUT_2[12460] = 32'b11111111111111110100011001000110;
assign LUT_2[12461] = 32'b11111111111111110001010001011111;
assign LUT_2[12462] = 32'b11111111111111111011010010000010;
assign LUT_2[12463] = 32'b11111111111111111000001010011011;
assign LUT_2[12464] = 32'b11111111111111110111101110001011;
assign LUT_2[12465] = 32'b11111111111111110100100110100100;
assign LUT_2[12466] = 32'b11111111111111111110100111000111;
assign LUT_2[12467] = 32'b11111111111111111011011111100000;
assign LUT_2[12468] = 32'b11111111111111110100001011110011;
assign LUT_2[12469] = 32'b11111111111111110001000100001100;
assign LUT_2[12470] = 32'b11111111111111111011000100101111;
assign LUT_2[12471] = 32'b11111111111111110111111101001000;
assign LUT_2[12472] = 32'b11111111111111110010011111101000;
assign LUT_2[12473] = 32'b11111111111111101111011000000001;
assign LUT_2[12474] = 32'b11111111111111111001011000100100;
assign LUT_2[12475] = 32'b11111111111111110110010000111101;
assign LUT_2[12476] = 32'b11111111111111101110111101010000;
assign LUT_2[12477] = 32'b11111111111111101011110101101001;
assign LUT_2[12478] = 32'b11111111111111110101110110001100;
assign LUT_2[12479] = 32'b11111111111111110010101110100101;
assign LUT_2[12480] = 32'b11111111111111110100110110111011;
assign LUT_2[12481] = 32'b11111111111111110001101111010100;
assign LUT_2[12482] = 32'b11111111111111111011101111110111;
assign LUT_2[12483] = 32'b11111111111111111000101000010000;
assign LUT_2[12484] = 32'b11111111111111110001010100100011;
assign LUT_2[12485] = 32'b11111111111111101110001100111100;
assign LUT_2[12486] = 32'b11111111111111111000001101011111;
assign LUT_2[12487] = 32'b11111111111111110101000101111000;
assign LUT_2[12488] = 32'b11111111111111101111101000011000;
assign LUT_2[12489] = 32'b11111111111111101100100000110001;
assign LUT_2[12490] = 32'b11111111111111110110100001010100;
assign LUT_2[12491] = 32'b11111111111111110011011001101101;
assign LUT_2[12492] = 32'b11111111111111101100000110000000;
assign LUT_2[12493] = 32'b11111111111111101000111110011001;
assign LUT_2[12494] = 32'b11111111111111110010111110111100;
assign LUT_2[12495] = 32'b11111111111111101111110111010101;
assign LUT_2[12496] = 32'b11111111111111101111011011000101;
assign LUT_2[12497] = 32'b11111111111111101100010011011110;
assign LUT_2[12498] = 32'b11111111111111110110010100000001;
assign LUT_2[12499] = 32'b11111111111111110011001100011010;
assign LUT_2[12500] = 32'b11111111111111101011111000101101;
assign LUT_2[12501] = 32'b11111111111111101000110001000110;
assign LUT_2[12502] = 32'b11111111111111110010110001101001;
assign LUT_2[12503] = 32'b11111111111111101111101010000010;
assign LUT_2[12504] = 32'b11111111111111101010001100100010;
assign LUT_2[12505] = 32'b11111111111111100111000100111011;
assign LUT_2[12506] = 32'b11111111111111110001000101011110;
assign LUT_2[12507] = 32'b11111111111111101101111101110111;
assign LUT_2[12508] = 32'b11111111111111100110101010001010;
assign LUT_2[12509] = 32'b11111111111111100011100010100011;
assign LUT_2[12510] = 32'b11111111111111101101100011000110;
assign LUT_2[12511] = 32'b11111111111111101010011011011111;
assign LUT_2[12512] = 32'b11111111111111110101010010100100;
assign LUT_2[12513] = 32'b11111111111111110010001010111101;
assign LUT_2[12514] = 32'b11111111111111111100001011100000;
assign LUT_2[12515] = 32'b11111111111111111001000011111001;
assign LUT_2[12516] = 32'b11111111111111110001110000001100;
assign LUT_2[12517] = 32'b11111111111111101110101000100101;
assign LUT_2[12518] = 32'b11111111111111111000101001001000;
assign LUT_2[12519] = 32'b11111111111111110101100001100001;
assign LUT_2[12520] = 32'b11111111111111110000000100000001;
assign LUT_2[12521] = 32'b11111111111111101100111100011010;
assign LUT_2[12522] = 32'b11111111111111110110111100111101;
assign LUT_2[12523] = 32'b11111111111111110011110101010110;
assign LUT_2[12524] = 32'b11111111111111101100100001101001;
assign LUT_2[12525] = 32'b11111111111111101001011010000010;
assign LUT_2[12526] = 32'b11111111111111110011011010100101;
assign LUT_2[12527] = 32'b11111111111111110000010010111110;
assign LUT_2[12528] = 32'b11111111111111101111110110101110;
assign LUT_2[12529] = 32'b11111111111111101100101111000111;
assign LUT_2[12530] = 32'b11111111111111110110101111101010;
assign LUT_2[12531] = 32'b11111111111111110011101000000011;
assign LUT_2[12532] = 32'b11111111111111101100010100010110;
assign LUT_2[12533] = 32'b11111111111111101001001100101111;
assign LUT_2[12534] = 32'b11111111111111110011001101010010;
assign LUT_2[12535] = 32'b11111111111111110000000101101011;
assign LUT_2[12536] = 32'b11111111111111101010101000001011;
assign LUT_2[12537] = 32'b11111111111111100111100000100100;
assign LUT_2[12538] = 32'b11111111111111110001100001000111;
assign LUT_2[12539] = 32'b11111111111111101110011001100000;
assign LUT_2[12540] = 32'b11111111111111100111000101110011;
assign LUT_2[12541] = 32'b11111111111111100011111110001100;
assign LUT_2[12542] = 32'b11111111111111101101111110101111;
assign LUT_2[12543] = 32'b11111111111111101010110111001000;
assign LUT_2[12544] = 32'b11111111111111111100011000101111;
assign LUT_2[12545] = 32'b11111111111111111001010001001000;
assign LUT_2[12546] = 32'b00000000000000000011010001101011;
assign LUT_2[12547] = 32'b00000000000000000000001010000100;
assign LUT_2[12548] = 32'b11111111111111111000110110010111;
assign LUT_2[12549] = 32'b11111111111111110101101110110000;
assign LUT_2[12550] = 32'b11111111111111111111101111010011;
assign LUT_2[12551] = 32'b11111111111111111100100111101100;
assign LUT_2[12552] = 32'b11111111111111110111001010001100;
assign LUT_2[12553] = 32'b11111111111111110100000010100101;
assign LUT_2[12554] = 32'b11111111111111111110000011001000;
assign LUT_2[12555] = 32'b11111111111111111010111011100001;
assign LUT_2[12556] = 32'b11111111111111110011100111110100;
assign LUT_2[12557] = 32'b11111111111111110000100000001101;
assign LUT_2[12558] = 32'b11111111111111111010100000110000;
assign LUT_2[12559] = 32'b11111111111111110111011001001001;
assign LUT_2[12560] = 32'b11111111111111110110111100111001;
assign LUT_2[12561] = 32'b11111111111111110011110101010010;
assign LUT_2[12562] = 32'b11111111111111111101110101110101;
assign LUT_2[12563] = 32'b11111111111111111010101110001110;
assign LUT_2[12564] = 32'b11111111111111110011011010100001;
assign LUT_2[12565] = 32'b11111111111111110000010010111010;
assign LUT_2[12566] = 32'b11111111111111111010010011011101;
assign LUT_2[12567] = 32'b11111111111111110111001011110110;
assign LUT_2[12568] = 32'b11111111111111110001101110010110;
assign LUT_2[12569] = 32'b11111111111111101110100110101111;
assign LUT_2[12570] = 32'b11111111111111111000100111010010;
assign LUT_2[12571] = 32'b11111111111111110101011111101011;
assign LUT_2[12572] = 32'b11111111111111101110001011111110;
assign LUT_2[12573] = 32'b11111111111111101011000100010111;
assign LUT_2[12574] = 32'b11111111111111110101000100111010;
assign LUT_2[12575] = 32'b11111111111111110001111101010011;
assign LUT_2[12576] = 32'b11111111111111111100110100011000;
assign LUT_2[12577] = 32'b11111111111111111001101100110001;
assign LUT_2[12578] = 32'b00000000000000000011101101010100;
assign LUT_2[12579] = 32'b00000000000000000000100101101101;
assign LUT_2[12580] = 32'b11111111111111111001010010000000;
assign LUT_2[12581] = 32'b11111111111111110110001010011001;
assign LUT_2[12582] = 32'b00000000000000000000001010111100;
assign LUT_2[12583] = 32'b11111111111111111101000011010101;
assign LUT_2[12584] = 32'b11111111111111110111100101110101;
assign LUT_2[12585] = 32'b11111111111111110100011110001110;
assign LUT_2[12586] = 32'b11111111111111111110011110110001;
assign LUT_2[12587] = 32'b11111111111111111011010111001010;
assign LUT_2[12588] = 32'b11111111111111110100000011011101;
assign LUT_2[12589] = 32'b11111111111111110000111011110110;
assign LUT_2[12590] = 32'b11111111111111111010111100011001;
assign LUT_2[12591] = 32'b11111111111111110111110100110010;
assign LUT_2[12592] = 32'b11111111111111110111011000100010;
assign LUT_2[12593] = 32'b11111111111111110100010000111011;
assign LUT_2[12594] = 32'b11111111111111111110010001011110;
assign LUT_2[12595] = 32'b11111111111111111011001001110111;
assign LUT_2[12596] = 32'b11111111111111110011110110001010;
assign LUT_2[12597] = 32'b11111111111111110000101110100011;
assign LUT_2[12598] = 32'b11111111111111111010101111000110;
assign LUT_2[12599] = 32'b11111111111111110111100111011111;
assign LUT_2[12600] = 32'b11111111111111110010001001111111;
assign LUT_2[12601] = 32'b11111111111111101111000010011000;
assign LUT_2[12602] = 32'b11111111111111111001000010111011;
assign LUT_2[12603] = 32'b11111111111111110101111011010100;
assign LUT_2[12604] = 32'b11111111111111101110100111100111;
assign LUT_2[12605] = 32'b11111111111111101011100000000000;
assign LUT_2[12606] = 32'b11111111111111110101100000100011;
assign LUT_2[12607] = 32'b11111111111111110010011000111100;
assign LUT_2[12608] = 32'b11111111111111110100100001010010;
assign LUT_2[12609] = 32'b11111111111111110001011001101011;
assign LUT_2[12610] = 32'b11111111111111111011011010001110;
assign LUT_2[12611] = 32'b11111111111111111000010010100111;
assign LUT_2[12612] = 32'b11111111111111110000111110111010;
assign LUT_2[12613] = 32'b11111111111111101101110111010011;
assign LUT_2[12614] = 32'b11111111111111110111110111110110;
assign LUT_2[12615] = 32'b11111111111111110100110000001111;
assign LUT_2[12616] = 32'b11111111111111101111010010101111;
assign LUT_2[12617] = 32'b11111111111111101100001011001000;
assign LUT_2[12618] = 32'b11111111111111110110001011101011;
assign LUT_2[12619] = 32'b11111111111111110011000100000100;
assign LUT_2[12620] = 32'b11111111111111101011110000010111;
assign LUT_2[12621] = 32'b11111111111111101000101000110000;
assign LUT_2[12622] = 32'b11111111111111110010101001010011;
assign LUT_2[12623] = 32'b11111111111111101111100001101100;
assign LUT_2[12624] = 32'b11111111111111101111000101011100;
assign LUT_2[12625] = 32'b11111111111111101011111101110101;
assign LUT_2[12626] = 32'b11111111111111110101111110011000;
assign LUT_2[12627] = 32'b11111111111111110010110110110001;
assign LUT_2[12628] = 32'b11111111111111101011100011000100;
assign LUT_2[12629] = 32'b11111111111111101000011011011101;
assign LUT_2[12630] = 32'b11111111111111110010011100000000;
assign LUT_2[12631] = 32'b11111111111111101111010100011001;
assign LUT_2[12632] = 32'b11111111111111101001110110111001;
assign LUT_2[12633] = 32'b11111111111111100110101111010010;
assign LUT_2[12634] = 32'b11111111111111110000101111110101;
assign LUT_2[12635] = 32'b11111111111111101101101000001110;
assign LUT_2[12636] = 32'b11111111111111100110010100100001;
assign LUT_2[12637] = 32'b11111111111111100011001100111010;
assign LUT_2[12638] = 32'b11111111111111101101001101011101;
assign LUT_2[12639] = 32'b11111111111111101010000101110110;
assign LUT_2[12640] = 32'b11111111111111110100111100111011;
assign LUT_2[12641] = 32'b11111111111111110001110101010100;
assign LUT_2[12642] = 32'b11111111111111111011110101110111;
assign LUT_2[12643] = 32'b11111111111111111000101110010000;
assign LUT_2[12644] = 32'b11111111111111110001011010100011;
assign LUT_2[12645] = 32'b11111111111111101110010010111100;
assign LUT_2[12646] = 32'b11111111111111111000010011011111;
assign LUT_2[12647] = 32'b11111111111111110101001011111000;
assign LUT_2[12648] = 32'b11111111111111101111101110011000;
assign LUT_2[12649] = 32'b11111111111111101100100110110001;
assign LUT_2[12650] = 32'b11111111111111110110100111010100;
assign LUT_2[12651] = 32'b11111111111111110011011111101101;
assign LUT_2[12652] = 32'b11111111111111101100001100000000;
assign LUT_2[12653] = 32'b11111111111111101001000100011001;
assign LUT_2[12654] = 32'b11111111111111110011000100111100;
assign LUT_2[12655] = 32'b11111111111111101111111101010101;
assign LUT_2[12656] = 32'b11111111111111101111100001000101;
assign LUT_2[12657] = 32'b11111111111111101100011001011110;
assign LUT_2[12658] = 32'b11111111111111110110011010000001;
assign LUT_2[12659] = 32'b11111111111111110011010010011010;
assign LUT_2[12660] = 32'b11111111111111101011111110101101;
assign LUT_2[12661] = 32'b11111111111111101000110111000110;
assign LUT_2[12662] = 32'b11111111111111110010110111101001;
assign LUT_2[12663] = 32'b11111111111111101111110000000010;
assign LUT_2[12664] = 32'b11111111111111101010010010100010;
assign LUT_2[12665] = 32'b11111111111111100111001010111011;
assign LUT_2[12666] = 32'b11111111111111110001001011011110;
assign LUT_2[12667] = 32'b11111111111111101110000011110111;
assign LUT_2[12668] = 32'b11111111111111100110110000001010;
assign LUT_2[12669] = 32'b11111111111111100011101000100011;
assign LUT_2[12670] = 32'b11111111111111101101101001000110;
assign LUT_2[12671] = 32'b11111111111111101010100001011111;
assign LUT_2[12672] = 32'b00000000000000000000101100111110;
assign LUT_2[12673] = 32'b11111111111111111101100101010111;
assign LUT_2[12674] = 32'b00000000000000000111100101111010;
assign LUT_2[12675] = 32'b00000000000000000100011110010011;
assign LUT_2[12676] = 32'b11111111111111111101001010100110;
assign LUT_2[12677] = 32'b11111111111111111010000010111111;
assign LUT_2[12678] = 32'b00000000000000000100000011100010;
assign LUT_2[12679] = 32'b00000000000000000000111011111011;
assign LUT_2[12680] = 32'b11111111111111111011011110011011;
assign LUT_2[12681] = 32'b11111111111111111000010110110100;
assign LUT_2[12682] = 32'b00000000000000000010010111010111;
assign LUT_2[12683] = 32'b11111111111111111111001111110000;
assign LUT_2[12684] = 32'b11111111111111110111111100000011;
assign LUT_2[12685] = 32'b11111111111111110100110100011100;
assign LUT_2[12686] = 32'b11111111111111111110110100111111;
assign LUT_2[12687] = 32'b11111111111111111011101101011000;
assign LUT_2[12688] = 32'b11111111111111111011010001001000;
assign LUT_2[12689] = 32'b11111111111111111000001001100001;
assign LUT_2[12690] = 32'b00000000000000000010001010000100;
assign LUT_2[12691] = 32'b11111111111111111111000010011101;
assign LUT_2[12692] = 32'b11111111111111110111101110110000;
assign LUT_2[12693] = 32'b11111111111111110100100111001001;
assign LUT_2[12694] = 32'b11111111111111111110100111101100;
assign LUT_2[12695] = 32'b11111111111111111011100000000101;
assign LUT_2[12696] = 32'b11111111111111110110000010100101;
assign LUT_2[12697] = 32'b11111111111111110010111010111110;
assign LUT_2[12698] = 32'b11111111111111111100111011100001;
assign LUT_2[12699] = 32'b11111111111111111001110011111010;
assign LUT_2[12700] = 32'b11111111111111110010100000001101;
assign LUT_2[12701] = 32'b11111111111111101111011000100110;
assign LUT_2[12702] = 32'b11111111111111111001011001001001;
assign LUT_2[12703] = 32'b11111111111111110110010001100010;
assign LUT_2[12704] = 32'b00000000000000000001001000100111;
assign LUT_2[12705] = 32'b11111111111111111110000001000000;
assign LUT_2[12706] = 32'b00000000000000001000000001100011;
assign LUT_2[12707] = 32'b00000000000000000100111001111100;
assign LUT_2[12708] = 32'b11111111111111111101100110001111;
assign LUT_2[12709] = 32'b11111111111111111010011110101000;
assign LUT_2[12710] = 32'b00000000000000000100011111001011;
assign LUT_2[12711] = 32'b00000000000000000001010111100100;
assign LUT_2[12712] = 32'b11111111111111111011111010000100;
assign LUT_2[12713] = 32'b11111111111111111000110010011101;
assign LUT_2[12714] = 32'b00000000000000000010110011000000;
assign LUT_2[12715] = 32'b11111111111111111111101011011001;
assign LUT_2[12716] = 32'b11111111111111111000010111101100;
assign LUT_2[12717] = 32'b11111111111111110101010000000101;
assign LUT_2[12718] = 32'b11111111111111111111010000101000;
assign LUT_2[12719] = 32'b11111111111111111100001001000001;
assign LUT_2[12720] = 32'b11111111111111111011101100110001;
assign LUT_2[12721] = 32'b11111111111111111000100101001010;
assign LUT_2[12722] = 32'b00000000000000000010100101101101;
assign LUT_2[12723] = 32'b11111111111111111111011110000110;
assign LUT_2[12724] = 32'b11111111111111111000001010011001;
assign LUT_2[12725] = 32'b11111111111111110101000010110010;
assign LUT_2[12726] = 32'b11111111111111111111000011010101;
assign LUT_2[12727] = 32'b11111111111111111011111011101110;
assign LUT_2[12728] = 32'b11111111111111110110011110001110;
assign LUT_2[12729] = 32'b11111111111111110011010110100111;
assign LUT_2[12730] = 32'b11111111111111111101010111001010;
assign LUT_2[12731] = 32'b11111111111111111010001111100011;
assign LUT_2[12732] = 32'b11111111111111110010111011110110;
assign LUT_2[12733] = 32'b11111111111111101111110100001111;
assign LUT_2[12734] = 32'b11111111111111111001110100110010;
assign LUT_2[12735] = 32'b11111111111111110110101101001011;
assign LUT_2[12736] = 32'b11111111111111111000110101100001;
assign LUT_2[12737] = 32'b11111111111111110101101101111010;
assign LUT_2[12738] = 32'b11111111111111111111101110011101;
assign LUT_2[12739] = 32'b11111111111111111100100110110110;
assign LUT_2[12740] = 32'b11111111111111110101010011001001;
assign LUT_2[12741] = 32'b11111111111111110010001011100010;
assign LUT_2[12742] = 32'b11111111111111111100001100000101;
assign LUT_2[12743] = 32'b11111111111111111001000100011110;
assign LUT_2[12744] = 32'b11111111111111110011100110111110;
assign LUT_2[12745] = 32'b11111111111111110000011111010111;
assign LUT_2[12746] = 32'b11111111111111111010011111111010;
assign LUT_2[12747] = 32'b11111111111111110111011000010011;
assign LUT_2[12748] = 32'b11111111111111110000000100100110;
assign LUT_2[12749] = 32'b11111111111111101100111100111111;
assign LUT_2[12750] = 32'b11111111111111110110111101100010;
assign LUT_2[12751] = 32'b11111111111111110011110101111011;
assign LUT_2[12752] = 32'b11111111111111110011011001101011;
assign LUT_2[12753] = 32'b11111111111111110000010010000100;
assign LUT_2[12754] = 32'b11111111111111111010010010100111;
assign LUT_2[12755] = 32'b11111111111111110111001011000000;
assign LUT_2[12756] = 32'b11111111111111101111110111010011;
assign LUT_2[12757] = 32'b11111111111111101100101111101100;
assign LUT_2[12758] = 32'b11111111111111110110110000001111;
assign LUT_2[12759] = 32'b11111111111111110011101000101000;
assign LUT_2[12760] = 32'b11111111111111101110001011001000;
assign LUT_2[12761] = 32'b11111111111111101011000011100001;
assign LUT_2[12762] = 32'b11111111111111110101000100000100;
assign LUT_2[12763] = 32'b11111111111111110001111100011101;
assign LUT_2[12764] = 32'b11111111111111101010101000110000;
assign LUT_2[12765] = 32'b11111111111111100111100001001001;
assign LUT_2[12766] = 32'b11111111111111110001100001101100;
assign LUT_2[12767] = 32'b11111111111111101110011010000101;
assign LUT_2[12768] = 32'b11111111111111111001010001001010;
assign LUT_2[12769] = 32'b11111111111111110110001001100011;
assign LUT_2[12770] = 32'b00000000000000000000001010000110;
assign LUT_2[12771] = 32'b11111111111111111101000010011111;
assign LUT_2[12772] = 32'b11111111111111110101101110110010;
assign LUT_2[12773] = 32'b11111111111111110010100111001011;
assign LUT_2[12774] = 32'b11111111111111111100100111101110;
assign LUT_2[12775] = 32'b11111111111111111001100000000111;
assign LUT_2[12776] = 32'b11111111111111110100000010100111;
assign LUT_2[12777] = 32'b11111111111111110000111011000000;
assign LUT_2[12778] = 32'b11111111111111111010111011100011;
assign LUT_2[12779] = 32'b11111111111111110111110011111100;
assign LUT_2[12780] = 32'b11111111111111110000100000001111;
assign LUT_2[12781] = 32'b11111111111111101101011000101000;
assign LUT_2[12782] = 32'b11111111111111110111011001001011;
assign LUT_2[12783] = 32'b11111111111111110100010001100100;
assign LUT_2[12784] = 32'b11111111111111110011110101010100;
assign LUT_2[12785] = 32'b11111111111111110000101101101101;
assign LUT_2[12786] = 32'b11111111111111111010101110010000;
assign LUT_2[12787] = 32'b11111111111111110111100110101001;
assign LUT_2[12788] = 32'b11111111111111110000010010111100;
assign LUT_2[12789] = 32'b11111111111111101101001011010101;
assign LUT_2[12790] = 32'b11111111111111110111001011111000;
assign LUT_2[12791] = 32'b11111111111111110100000100010001;
assign LUT_2[12792] = 32'b11111111111111101110100110110001;
assign LUT_2[12793] = 32'b11111111111111101011011111001010;
assign LUT_2[12794] = 32'b11111111111111110101011111101101;
assign LUT_2[12795] = 32'b11111111111111110010011000000110;
assign LUT_2[12796] = 32'b11111111111111101011000100011001;
assign LUT_2[12797] = 32'b11111111111111100111111100110010;
assign LUT_2[12798] = 32'b11111111111111110001111101010101;
assign LUT_2[12799] = 32'b11111111111111101110110101101110;
assign LUT_2[12800] = 32'b11111111111111111101001011111011;
assign LUT_2[12801] = 32'b11111111111111111010000100010100;
assign LUT_2[12802] = 32'b00000000000000000100000100110111;
assign LUT_2[12803] = 32'b00000000000000000000111101010000;
assign LUT_2[12804] = 32'b11111111111111111001101001100011;
assign LUT_2[12805] = 32'b11111111111111110110100001111100;
assign LUT_2[12806] = 32'b00000000000000000000100010011111;
assign LUT_2[12807] = 32'b11111111111111111101011010111000;
assign LUT_2[12808] = 32'b11111111111111110111111101011000;
assign LUT_2[12809] = 32'b11111111111111110100110101110001;
assign LUT_2[12810] = 32'b11111111111111111110110110010100;
assign LUT_2[12811] = 32'b11111111111111111011101110101101;
assign LUT_2[12812] = 32'b11111111111111110100011011000000;
assign LUT_2[12813] = 32'b11111111111111110001010011011001;
assign LUT_2[12814] = 32'b11111111111111111011010011111100;
assign LUT_2[12815] = 32'b11111111111111111000001100010101;
assign LUT_2[12816] = 32'b11111111111111110111110000000101;
assign LUT_2[12817] = 32'b11111111111111110100101000011110;
assign LUT_2[12818] = 32'b11111111111111111110101001000001;
assign LUT_2[12819] = 32'b11111111111111111011100001011010;
assign LUT_2[12820] = 32'b11111111111111110100001101101101;
assign LUT_2[12821] = 32'b11111111111111110001000110000110;
assign LUT_2[12822] = 32'b11111111111111111011000110101001;
assign LUT_2[12823] = 32'b11111111111111110111111111000010;
assign LUT_2[12824] = 32'b11111111111111110010100001100010;
assign LUT_2[12825] = 32'b11111111111111101111011001111011;
assign LUT_2[12826] = 32'b11111111111111111001011010011110;
assign LUT_2[12827] = 32'b11111111111111110110010010110111;
assign LUT_2[12828] = 32'b11111111111111101110111111001010;
assign LUT_2[12829] = 32'b11111111111111101011110111100011;
assign LUT_2[12830] = 32'b11111111111111110101111000000110;
assign LUT_2[12831] = 32'b11111111111111110010110000011111;
assign LUT_2[12832] = 32'b11111111111111111101100111100100;
assign LUT_2[12833] = 32'b11111111111111111010011111111101;
assign LUT_2[12834] = 32'b00000000000000000100100000100000;
assign LUT_2[12835] = 32'b00000000000000000001011000111001;
assign LUT_2[12836] = 32'b11111111111111111010000101001100;
assign LUT_2[12837] = 32'b11111111111111110110111101100101;
assign LUT_2[12838] = 32'b00000000000000000000111110001000;
assign LUT_2[12839] = 32'b11111111111111111101110110100001;
assign LUT_2[12840] = 32'b11111111111111111000011001000001;
assign LUT_2[12841] = 32'b11111111111111110101010001011010;
assign LUT_2[12842] = 32'b11111111111111111111010001111101;
assign LUT_2[12843] = 32'b11111111111111111100001010010110;
assign LUT_2[12844] = 32'b11111111111111110100110110101001;
assign LUT_2[12845] = 32'b11111111111111110001101111000010;
assign LUT_2[12846] = 32'b11111111111111111011101111100101;
assign LUT_2[12847] = 32'b11111111111111111000100111111110;
assign LUT_2[12848] = 32'b11111111111111111000001011101110;
assign LUT_2[12849] = 32'b11111111111111110101000100000111;
assign LUT_2[12850] = 32'b11111111111111111111000100101010;
assign LUT_2[12851] = 32'b11111111111111111011111101000011;
assign LUT_2[12852] = 32'b11111111111111110100101001010110;
assign LUT_2[12853] = 32'b11111111111111110001100001101111;
assign LUT_2[12854] = 32'b11111111111111111011100010010010;
assign LUT_2[12855] = 32'b11111111111111111000011010101011;
assign LUT_2[12856] = 32'b11111111111111110010111101001011;
assign LUT_2[12857] = 32'b11111111111111101111110101100100;
assign LUT_2[12858] = 32'b11111111111111111001110110000111;
assign LUT_2[12859] = 32'b11111111111111110110101110100000;
assign LUT_2[12860] = 32'b11111111111111101111011010110011;
assign LUT_2[12861] = 32'b11111111111111101100010011001100;
assign LUT_2[12862] = 32'b11111111111111110110010011101111;
assign LUT_2[12863] = 32'b11111111111111110011001100001000;
assign LUT_2[12864] = 32'b11111111111111110101010100011110;
assign LUT_2[12865] = 32'b11111111111111110010001100110111;
assign LUT_2[12866] = 32'b11111111111111111100001101011010;
assign LUT_2[12867] = 32'b11111111111111111001000101110011;
assign LUT_2[12868] = 32'b11111111111111110001110010000110;
assign LUT_2[12869] = 32'b11111111111111101110101010011111;
assign LUT_2[12870] = 32'b11111111111111111000101011000010;
assign LUT_2[12871] = 32'b11111111111111110101100011011011;
assign LUT_2[12872] = 32'b11111111111111110000000101111011;
assign LUT_2[12873] = 32'b11111111111111101100111110010100;
assign LUT_2[12874] = 32'b11111111111111110110111110110111;
assign LUT_2[12875] = 32'b11111111111111110011110111010000;
assign LUT_2[12876] = 32'b11111111111111101100100011100011;
assign LUT_2[12877] = 32'b11111111111111101001011011111100;
assign LUT_2[12878] = 32'b11111111111111110011011100011111;
assign LUT_2[12879] = 32'b11111111111111110000010100111000;
assign LUT_2[12880] = 32'b11111111111111101111111000101000;
assign LUT_2[12881] = 32'b11111111111111101100110001000001;
assign LUT_2[12882] = 32'b11111111111111110110110001100100;
assign LUT_2[12883] = 32'b11111111111111110011101001111101;
assign LUT_2[12884] = 32'b11111111111111101100010110010000;
assign LUT_2[12885] = 32'b11111111111111101001001110101001;
assign LUT_2[12886] = 32'b11111111111111110011001111001100;
assign LUT_2[12887] = 32'b11111111111111110000000111100101;
assign LUT_2[12888] = 32'b11111111111111101010101010000101;
assign LUT_2[12889] = 32'b11111111111111100111100010011110;
assign LUT_2[12890] = 32'b11111111111111110001100011000001;
assign LUT_2[12891] = 32'b11111111111111101110011011011010;
assign LUT_2[12892] = 32'b11111111111111100111000111101101;
assign LUT_2[12893] = 32'b11111111111111100100000000000110;
assign LUT_2[12894] = 32'b11111111111111101110000000101001;
assign LUT_2[12895] = 32'b11111111111111101010111001000010;
assign LUT_2[12896] = 32'b11111111111111110101110000000111;
assign LUT_2[12897] = 32'b11111111111111110010101000100000;
assign LUT_2[12898] = 32'b11111111111111111100101001000011;
assign LUT_2[12899] = 32'b11111111111111111001100001011100;
assign LUT_2[12900] = 32'b11111111111111110010001101101111;
assign LUT_2[12901] = 32'b11111111111111101111000110001000;
assign LUT_2[12902] = 32'b11111111111111111001000110101011;
assign LUT_2[12903] = 32'b11111111111111110101111111000100;
assign LUT_2[12904] = 32'b11111111111111110000100001100100;
assign LUT_2[12905] = 32'b11111111111111101101011001111101;
assign LUT_2[12906] = 32'b11111111111111110111011010100000;
assign LUT_2[12907] = 32'b11111111111111110100010010111001;
assign LUT_2[12908] = 32'b11111111111111101100111111001100;
assign LUT_2[12909] = 32'b11111111111111101001110111100101;
assign LUT_2[12910] = 32'b11111111111111110011111000001000;
assign LUT_2[12911] = 32'b11111111111111110000110000100001;
assign LUT_2[12912] = 32'b11111111111111110000010100010001;
assign LUT_2[12913] = 32'b11111111111111101101001100101010;
assign LUT_2[12914] = 32'b11111111111111110111001101001101;
assign LUT_2[12915] = 32'b11111111111111110100000101100110;
assign LUT_2[12916] = 32'b11111111111111101100110001111001;
assign LUT_2[12917] = 32'b11111111111111101001101010010010;
assign LUT_2[12918] = 32'b11111111111111110011101010110101;
assign LUT_2[12919] = 32'b11111111111111110000100011001110;
assign LUT_2[12920] = 32'b11111111111111101011000101101110;
assign LUT_2[12921] = 32'b11111111111111100111111110000111;
assign LUT_2[12922] = 32'b11111111111111110001111110101010;
assign LUT_2[12923] = 32'b11111111111111101110110111000011;
assign LUT_2[12924] = 32'b11111111111111100111100011010110;
assign LUT_2[12925] = 32'b11111111111111100100011011101111;
assign LUT_2[12926] = 32'b11111111111111101110011100010010;
assign LUT_2[12927] = 32'b11111111111111101011010100101011;
assign LUT_2[12928] = 32'b00000000000000000001100000001010;
assign LUT_2[12929] = 32'b11111111111111111110011000100011;
assign LUT_2[12930] = 32'b00000000000000001000011001000110;
assign LUT_2[12931] = 32'b00000000000000000101010001011111;
assign LUT_2[12932] = 32'b11111111111111111101111101110010;
assign LUT_2[12933] = 32'b11111111111111111010110110001011;
assign LUT_2[12934] = 32'b00000000000000000100110110101110;
assign LUT_2[12935] = 32'b00000000000000000001101111000111;
assign LUT_2[12936] = 32'b11111111111111111100010001100111;
assign LUT_2[12937] = 32'b11111111111111111001001010000000;
assign LUT_2[12938] = 32'b00000000000000000011001010100011;
assign LUT_2[12939] = 32'b00000000000000000000000010111100;
assign LUT_2[12940] = 32'b11111111111111111000101111001111;
assign LUT_2[12941] = 32'b11111111111111110101100111101000;
assign LUT_2[12942] = 32'b11111111111111111111101000001011;
assign LUT_2[12943] = 32'b11111111111111111100100000100100;
assign LUT_2[12944] = 32'b11111111111111111100000100010100;
assign LUT_2[12945] = 32'b11111111111111111000111100101101;
assign LUT_2[12946] = 32'b00000000000000000010111101010000;
assign LUT_2[12947] = 32'b11111111111111111111110101101001;
assign LUT_2[12948] = 32'b11111111111111111000100001111100;
assign LUT_2[12949] = 32'b11111111111111110101011010010101;
assign LUT_2[12950] = 32'b11111111111111111111011010111000;
assign LUT_2[12951] = 32'b11111111111111111100010011010001;
assign LUT_2[12952] = 32'b11111111111111110110110101110001;
assign LUT_2[12953] = 32'b11111111111111110011101110001010;
assign LUT_2[12954] = 32'b11111111111111111101101110101101;
assign LUT_2[12955] = 32'b11111111111111111010100111000110;
assign LUT_2[12956] = 32'b11111111111111110011010011011001;
assign LUT_2[12957] = 32'b11111111111111110000001011110010;
assign LUT_2[12958] = 32'b11111111111111111010001100010101;
assign LUT_2[12959] = 32'b11111111111111110111000100101110;
assign LUT_2[12960] = 32'b00000000000000000001111011110011;
assign LUT_2[12961] = 32'b11111111111111111110110100001100;
assign LUT_2[12962] = 32'b00000000000000001000110100101111;
assign LUT_2[12963] = 32'b00000000000000000101101101001000;
assign LUT_2[12964] = 32'b11111111111111111110011001011011;
assign LUT_2[12965] = 32'b11111111111111111011010001110100;
assign LUT_2[12966] = 32'b00000000000000000101010010010111;
assign LUT_2[12967] = 32'b00000000000000000010001010110000;
assign LUT_2[12968] = 32'b11111111111111111100101101010000;
assign LUT_2[12969] = 32'b11111111111111111001100101101001;
assign LUT_2[12970] = 32'b00000000000000000011100110001100;
assign LUT_2[12971] = 32'b00000000000000000000011110100101;
assign LUT_2[12972] = 32'b11111111111111111001001010111000;
assign LUT_2[12973] = 32'b11111111111111110110000011010001;
assign LUT_2[12974] = 32'b00000000000000000000000011110100;
assign LUT_2[12975] = 32'b11111111111111111100111100001101;
assign LUT_2[12976] = 32'b11111111111111111100011111111101;
assign LUT_2[12977] = 32'b11111111111111111001011000010110;
assign LUT_2[12978] = 32'b00000000000000000011011000111001;
assign LUT_2[12979] = 32'b00000000000000000000010001010010;
assign LUT_2[12980] = 32'b11111111111111111000111101100101;
assign LUT_2[12981] = 32'b11111111111111110101110101111110;
assign LUT_2[12982] = 32'b11111111111111111111110110100001;
assign LUT_2[12983] = 32'b11111111111111111100101110111010;
assign LUT_2[12984] = 32'b11111111111111110111010001011010;
assign LUT_2[12985] = 32'b11111111111111110100001001110011;
assign LUT_2[12986] = 32'b11111111111111111110001010010110;
assign LUT_2[12987] = 32'b11111111111111111011000010101111;
assign LUT_2[12988] = 32'b11111111111111110011101111000010;
assign LUT_2[12989] = 32'b11111111111111110000100111011011;
assign LUT_2[12990] = 32'b11111111111111111010100111111110;
assign LUT_2[12991] = 32'b11111111111111110111100000010111;
assign LUT_2[12992] = 32'b11111111111111111001101000101101;
assign LUT_2[12993] = 32'b11111111111111110110100001000110;
assign LUT_2[12994] = 32'b00000000000000000000100001101001;
assign LUT_2[12995] = 32'b11111111111111111101011010000010;
assign LUT_2[12996] = 32'b11111111111111110110000110010101;
assign LUT_2[12997] = 32'b11111111111111110010111110101110;
assign LUT_2[12998] = 32'b11111111111111111100111111010001;
assign LUT_2[12999] = 32'b11111111111111111001110111101010;
assign LUT_2[13000] = 32'b11111111111111110100011010001010;
assign LUT_2[13001] = 32'b11111111111111110001010010100011;
assign LUT_2[13002] = 32'b11111111111111111011010011000110;
assign LUT_2[13003] = 32'b11111111111111111000001011011111;
assign LUT_2[13004] = 32'b11111111111111110000110111110010;
assign LUT_2[13005] = 32'b11111111111111101101110000001011;
assign LUT_2[13006] = 32'b11111111111111110111110000101110;
assign LUT_2[13007] = 32'b11111111111111110100101001000111;
assign LUT_2[13008] = 32'b11111111111111110100001100110111;
assign LUT_2[13009] = 32'b11111111111111110001000101010000;
assign LUT_2[13010] = 32'b11111111111111111011000101110011;
assign LUT_2[13011] = 32'b11111111111111110111111110001100;
assign LUT_2[13012] = 32'b11111111111111110000101010011111;
assign LUT_2[13013] = 32'b11111111111111101101100010111000;
assign LUT_2[13014] = 32'b11111111111111110111100011011011;
assign LUT_2[13015] = 32'b11111111111111110100011011110100;
assign LUT_2[13016] = 32'b11111111111111101110111110010100;
assign LUT_2[13017] = 32'b11111111111111101011110110101101;
assign LUT_2[13018] = 32'b11111111111111110101110111010000;
assign LUT_2[13019] = 32'b11111111111111110010101111101001;
assign LUT_2[13020] = 32'b11111111111111101011011011111100;
assign LUT_2[13021] = 32'b11111111111111101000010100010101;
assign LUT_2[13022] = 32'b11111111111111110010010100111000;
assign LUT_2[13023] = 32'b11111111111111101111001101010001;
assign LUT_2[13024] = 32'b11111111111111111010000100010110;
assign LUT_2[13025] = 32'b11111111111111110110111100101111;
assign LUT_2[13026] = 32'b00000000000000000000111101010010;
assign LUT_2[13027] = 32'b11111111111111111101110101101011;
assign LUT_2[13028] = 32'b11111111111111110110100001111110;
assign LUT_2[13029] = 32'b11111111111111110011011010010111;
assign LUT_2[13030] = 32'b11111111111111111101011010111010;
assign LUT_2[13031] = 32'b11111111111111111010010011010011;
assign LUT_2[13032] = 32'b11111111111111110100110101110011;
assign LUT_2[13033] = 32'b11111111111111110001101110001100;
assign LUT_2[13034] = 32'b11111111111111111011101110101111;
assign LUT_2[13035] = 32'b11111111111111111000100111001000;
assign LUT_2[13036] = 32'b11111111111111110001010011011011;
assign LUT_2[13037] = 32'b11111111111111101110001011110100;
assign LUT_2[13038] = 32'b11111111111111111000001100010111;
assign LUT_2[13039] = 32'b11111111111111110101000100110000;
assign LUT_2[13040] = 32'b11111111111111110100101000100000;
assign LUT_2[13041] = 32'b11111111111111110001100000111001;
assign LUT_2[13042] = 32'b11111111111111111011100001011100;
assign LUT_2[13043] = 32'b11111111111111111000011001110101;
assign LUT_2[13044] = 32'b11111111111111110001000110001000;
assign LUT_2[13045] = 32'b11111111111111101101111110100001;
assign LUT_2[13046] = 32'b11111111111111110111111111000100;
assign LUT_2[13047] = 32'b11111111111111110100110111011101;
assign LUT_2[13048] = 32'b11111111111111101111011001111101;
assign LUT_2[13049] = 32'b11111111111111101100010010010110;
assign LUT_2[13050] = 32'b11111111111111110110010010111001;
assign LUT_2[13051] = 32'b11111111111111110011001011010010;
assign LUT_2[13052] = 32'b11111111111111101011110111100101;
assign LUT_2[13053] = 32'b11111111111111101000101111111110;
assign LUT_2[13054] = 32'b11111111111111110010110000100001;
assign LUT_2[13055] = 32'b11111111111111101111101000111010;
assign LUT_2[13056] = 32'b00000000000000000001001010100001;
assign LUT_2[13057] = 32'b11111111111111111110000010111010;
assign LUT_2[13058] = 32'b00000000000000001000000011011101;
assign LUT_2[13059] = 32'b00000000000000000100111011110110;
assign LUT_2[13060] = 32'b11111111111111111101101000001001;
assign LUT_2[13061] = 32'b11111111111111111010100000100010;
assign LUT_2[13062] = 32'b00000000000000000100100001000101;
assign LUT_2[13063] = 32'b00000000000000000001011001011110;
assign LUT_2[13064] = 32'b11111111111111111011111011111110;
assign LUT_2[13065] = 32'b11111111111111111000110100010111;
assign LUT_2[13066] = 32'b00000000000000000010110100111010;
assign LUT_2[13067] = 32'b11111111111111111111101101010011;
assign LUT_2[13068] = 32'b11111111111111111000011001100110;
assign LUT_2[13069] = 32'b11111111111111110101010001111111;
assign LUT_2[13070] = 32'b11111111111111111111010010100010;
assign LUT_2[13071] = 32'b11111111111111111100001010111011;
assign LUT_2[13072] = 32'b11111111111111111011101110101011;
assign LUT_2[13073] = 32'b11111111111111111000100111000100;
assign LUT_2[13074] = 32'b00000000000000000010100111100111;
assign LUT_2[13075] = 32'b11111111111111111111100000000000;
assign LUT_2[13076] = 32'b11111111111111111000001100010011;
assign LUT_2[13077] = 32'b11111111111111110101000100101100;
assign LUT_2[13078] = 32'b11111111111111111111000101001111;
assign LUT_2[13079] = 32'b11111111111111111011111101101000;
assign LUT_2[13080] = 32'b11111111111111110110100000001000;
assign LUT_2[13081] = 32'b11111111111111110011011000100001;
assign LUT_2[13082] = 32'b11111111111111111101011001000100;
assign LUT_2[13083] = 32'b11111111111111111010010001011101;
assign LUT_2[13084] = 32'b11111111111111110010111101110000;
assign LUT_2[13085] = 32'b11111111111111101111110110001001;
assign LUT_2[13086] = 32'b11111111111111111001110110101100;
assign LUT_2[13087] = 32'b11111111111111110110101111000101;
assign LUT_2[13088] = 32'b00000000000000000001100110001010;
assign LUT_2[13089] = 32'b11111111111111111110011110100011;
assign LUT_2[13090] = 32'b00000000000000001000011111000110;
assign LUT_2[13091] = 32'b00000000000000000101010111011111;
assign LUT_2[13092] = 32'b11111111111111111110000011110010;
assign LUT_2[13093] = 32'b11111111111111111010111100001011;
assign LUT_2[13094] = 32'b00000000000000000100111100101110;
assign LUT_2[13095] = 32'b00000000000000000001110101000111;
assign LUT_2[13096] = 32'b11111111111111111100010111100111;
assign LUT_2[13097] = 32'b11111111111111111001010000000000;
assign LUT_2[13098] = 32'b00000000000000000011010000100011;
assign LUT_2[13099] = 32'b00000000000000000000001000111100;
assign LUT_2[13100] = 32'b11111111111111111000110101001111;
assign LUT_2[13101] = 32'b11111111111111110101101101101000;
assign LUT_2[13102] = 32'b11111111111111111111101110001011;
assign LUT_2[13103] = 32'b11111111111111111100100110100100;
assign LUT_2[13104] = 32'b11111111111111111100001010010100;
assign LUT_2[13105] = 32'b11111111111111111001000010101101;
assign LUT_2[13106] = 32'b00000000000000000011000011010000;
assign LUT_2[13107] = 32'b11111111111111111111111011101001;
assign LUT_2[13108] = 32'b11111111111111111000100111111100;
assign LUT_2[13109] = 32'b11111111111111110101100000010101;
assign LUT_2[13110] = 32'b11111111111111111111100000111000;
assign LUT_2[13111] = 32'b11111111111111111100011001010001;
assign LUT_2[13112] = 32'b11111111111111110110111011110001;
assign LUT_2[13113] = 32'b11111111111111110011110100001010;
assign LUT_2[13114] = 32'b11111111111111111101110100101101;
assign LUT_2[13115] = 32'b11111111111111111010101101000110;
assign LUT_2[13116] = 32'b11111111111111110011011001011001;
assign LUT_2[13117] = 32'b11111111111111110000010001110010;
assign LUT_2[13118] = 32'b11111111111111111010010010010101;
assign LUT_2[13119] = 32'b11111111111111110111001010101110;
assign LUT_2[13120] = 32'b11111111111111111001010011000100;
assign LUT_2[13121] = 32'b11111111111111110110001011011101;
assign LUT_2[13122] = 32'b00000000000000000000001100000000;
assign LUT_2[13123] = 32'b11111111111111111101000100011001;
assign LUT_2[13124] = 32'b11111111111111110101110000101100;
assign LUT_2[13125] = 32'b11111111111111110010101001000101;
assign LUT_2[13126] = 32'b11111111111111111100101001101000;
assign LUT_2[13127] = 32'b11111111111111111001100010000001;
assign LUT_2[13128] = 32'b11111111111111110100000100100001;
assign LUT_2[13129] = 32'b11111111111111110000111100111010;
assign LUT_2[13130] = 32'b11111111111111111010111101011101;
assign LUT_2[13131] = 32'b11111111111111110111110101110110;
assign LUT_2[13132] = 32'b11111111111111110000100010001001;
assign LUT_2[13133] = 32'b11111111111111101101011010100010;
assign LUT_2[13134] = 32'b11111111111111110111011011000101;
assign LUT_2[13135] = 32'b11111111111111110100010011011110;
assign LUT_2[13136] = 32'b11111111111111110011110111001110;
assign LUT_2[13137] = 32'b11111111111111110000101111100111;
assign LUT_2[13138] = 32'b11111111111111111010110000001010;
assign LUT_2[13139] = 32'b11111111111111110111101000100011;
assign LUT_2[13140] = 32'b11111111111111110000010100110110;
assign LUT_2[13141] = 32'b11111111111111101101001101001111;
assign LUT_2[13142] = 32'b11111111111111110111001101110010;
assign LUT_2[13143] = 32'b11111111111111110100000110001011;
assign LUT_2[13144] = 32'b11111111111111101110101000101011;
assign LUT_2[13145] = 32'b11111111111111101011100001000100;
assign LUT_2[13146] = 32'b11111111111111110101100001100111;
assign LUT_2[13147] = 32'b11111111111111110010011010000000;
assign LUT_2[13148] = 32'b11111111111111101011000110010011;
assign LUT_2[13149] = 32'b11111111111111100111111110101100;
assign LUT_2[13150] = 32'b11111111111111110001111111001111;
assign LUT_2[13151] = 32'b11111111111111101110110111101000;
assign LUT_2[13152] = 32'b11111111111111111001101110101101;
assign LUT_2[13153] = 32'b11111111111111110110100111000110;
assign LUT_2[13154] = 32'b00000000000000000000100111101001;
assign LUT_2[13155] = 32'b11111111111111111101100000000010;
assign LUT_2[13156] = 32'b11111111111111110110001100010101;
assign LUT_2[13157] = 32'b11111111111111110011000100101110;
assign LUT_2[13158] = 32'b11111111111111111101000101010001;
assign LUT_2[13159] = 32'b11111111111111111001111101101010;
assign LUT_2[13160] = 32'b11111111111111110100100000001010;
assign LUT_2[13161] = 32'b11111111111111110001011000100011;
assign LUT_2[13162] = 32'b11111111111111111011011001000110;
assign LUT_2[13163] = 32'b11111111111111111000010001011111;
assign LUT_2[13164] = 32'b11111111111111110000111101110010;
assign LUT_2[13165] = 32'b11111111111111101101110110001011;
assign LUT_2[13166] = 32'b11111111111111110111110110101110;
assign LUT_2[13167] = 32'b11111111111111110100101111000111;
assign LUT_2[13168] = 32'b11111111111111110100010010110111;
assign LUT_2[13169] = 32'b11111111111111110001001011010000;
assign LUT_2[13170] = 32'b11111111111111111011001011110011;
assign LUT_2[13171] = 32'b11111111111111111000000100001100;
assign LUT_2[13172] = 32'b11111111111111110000110000011111;
assign LUT_2[13173] = 32'b11111111111111101101101000111000;
assign LUT_2[13174] = 32'b11111111111111110111101001011011;
assign LUT_2[13175] = 32'b11111111111111110100100001110100;
assign LUT_2[13176] = 32'b11111111111111101111000100010100;
assign LUT_2[13177] = 32'b11111111111111101011111100101101;
assign LUT_2[13178] = 32'b11111111111111110101111101010000;
assign LUT_2[13179] = 32'b11111111111111110010110101101001;
assign LUT_2[13180] = 32'b11111111111111101011100001111100;
assign LUT_2[13181] = 32'b11111111111111101000011010010101;
assign LUT_2[13182] = 32'b11111111111111110010011010111000;
assign LUT_2[13183] = 32'b11111111111111101111010011010001;
assign LUT_2[13184] = 32'b00000000000000000101011110110000;
assign LUT_2[13185] = 32'b00000000000000000010010111001001;
assign LUT_2[13186] = 32'b00000000000000001100010111101100;
assign LUT_2[13187] = 32'b00000000000000001001010000000101;
assign LUT_2[13188] = 32'b00000000000000000001111100011000;
assign LUT_2[13189] = 32'b11111111111111111110110100110001;
assign LUT_2[13190] = 32'b00000000000000001000110101010100;
assign LUT_2[13191] = 32'b00000000000000000101101101101101;
assign LUT_2[13192] = 32'b00000000000000000000010000001101;
assign LUT_2[13193] = 32'b11111111111111111101001000100110;
assign LUT_2[13194] = 32'b00000000000000000111001001001001;
assign LUT_2[13195] = 32'b00000000000000000100000001100010;
assign LUT_2[13196] = 32'b11111111111111111100101101110101;
assign LUT_2[13197] = 32'b11111111111111111001100110001110;
assign LUT_2[13198] = 32'b00000000000000000011100110110001;
assign LUT_2[13199] = 32'b00000000000000000000011111001010;
assign LUT_2[13200] = 32'b00000000000000000000000010111010;
assign LUT_2[13201] = 32'b11111111111111111100111011010011;
assign LUT_2[13202] = 32'b00000000000000000110111011110110;
assign LUT_2[13203] = 32'b00000000000000000011110100001111;
assign LUT_2[13204] = 32'b11111111111111111100100000100010;
assign LUT_2[13205] = 32'b11111111111111111001011000111011;
assign LUT_2[13206] = 32'b00000000000000000011011001011110;
assign LUT_2[13207] = 32'b00000000000000000000010001110111;
assign LUT_2[13208] = 32'b11111111111111111010110100010111;
assign LUT_2[13209] = 32'b11111111111111110111101100110000;
assign LUT_2[13210] = 32'b00000000000000000001101101010011;
assign LUT_2[13211] = 32'b11111111111111111110100101101100;
assign LUT_2[13212] = 32'b11111111111111110111010001111111;
assign LUT_2[13213] = 32'b11111111111111110100001010011000;
assign LUT_2[13214] = 32'b11111111111111111110001010111011;
assign LUT_2[13215] = 32'b11111111111111111011000011010100;
assign LUT_2[13216] = 32'b00000000000000000101111010011001;
assign LUT_2[13217] = 32'b00000000000000000010110010110010;
assign LUT_2[13218] = 32'b00000000000000001100110011010101;
assign LUT_2[13219] = 32'b00000000000000001001101011101110;
assign LUT_2[13220] = 32'b00000000000000000010011000000001;
assign LUT_2[13221] = 32'b11111111111111111111010000011010;
assign LUT_2[13222] = 32'b00000000000000001001010000111101;
assign LUT_2[13223] = 32'b00000000000000000110001001010110;
assign LUT_2[13224] = 32'b00000000000000000000101011110110;
assign LUT_2[13225] = 32'b11111111111111111101100100001111;
assign LUT_2[13226] = 32'b00000000000000000111100100110010;
assign LUT_2[13227] = 32'b00000000000000000100011101001011;
assign LUT_2[13228] = 32'b11111111111111111101001001011110;
assign LUT_2[13229] = 32'b11111111111111111010000001110111;
assign LUT_2[13230] = 32'b00000000000000000100000010011010;
assign LUT_2[13231] = 32'b00000000000000000000111010110011;
assign LUT_2[13232] = 32'b00000000000000000000011110100011;
assign LUT_2[13233] = 32'b11111111111111111101010110111100;
assign LUT_2[13234] = 32'b00000000000000000111010111011111;
assign LUT_2[13235] = 32'b00000000000000000100001111111000;
assign LUT_2[13236] = 32'b11111111111111111100111100001011;
assign LUT_2[13237] = 32'b11111111111111111001110100100100;
assign LUT_2[13238] = 32'b00000000000000000011110101000111;
assign LUT_2[13239] = 32'b00000000000000000000101101100000;
assign LUT_2[13240] = 32'b11111111111111111011010000000000;
assign LUT_2[13241] = 32'b11111111111111111000001000011001;
assign LUT_2[13242] = 32'b00000000000000000010001000111100;
assign LUT_2[13243] = 32'b11111111111111111111000001010101;
assign LUT_2[13244] = 32'b11111111111111110111101101101000;
assign LUT_2[13245] = 32'b11111111111111110100100110000001;
assign LUT_2[13246] = 32'b11111111111111111110100110100100;
assign LUT_2[13247] = 32'b11111111111111111011011110111101;
assign LUT_2[13248] = 32'b11111111111111111101100111010011;
assign LUT_2[13249] = 32'b11111111111111111010011111101100;
assign LUT_2[13250] = 32'b00000000000000000100100000001111;
assign LUT_2[13251] = 32'b00000000000000000001011000101000;
assign LUT_2[13252] = 32'b11111111111111111010000100111011;
assign LUT_2[13253] = 32'b11111111111111110110111101010100;
assign LUT_2[13254] = 32'b00000000000000000000111101110111;
assign LUT_2[13255] = 32'b11111111111111111101110110010000;
assign LUT_2[13256] = 32'b11111111111111111000011000110000;
assign LUT_2[13257] = 32'b11111111111111110101010001001001;
assign LUT_2[13258] = 32'b11111111111111111111010001101100;
assign LUT_2[13259] = 32'b11111111111111111100001010000101;
assign LUT_2[13260] = 32'b11111111111111110100110110011000;
assign LUT_2[13261] = 32'b11111111111111110001101110110001;
assign LUT_2[13262] = 32'b11111111111111111011101111010100;
assign LUT_2[13263] = 32'b11111111111111111000100111101101;
assign LUT_2[13264] = 32'b11111111111111111000001011011101;
assign LUT_2[13265] = 32'b11111111111111110101000011110110;
assign LUT_2[13266] = 32'b11111111111111111111000100011001;
assign LUT_2[13267] = 32'b11111111111111111011111100110010;
assign LUT_2[13268] = 32'b11111111111111110100101001000101;
assign LUT_2[13269] = 32'b11111111111111110001100001011110;
assign LUT_2[13270] = 32'b11111111111111111011100010000001;
assign LUT_2[13271] = 32'b11111111111111111000011010011010;
assign LUT_2[13272] = 32'b11111111111111110010111100111010;
assign LUT_2[13273] = 32'b11111111111111101111110101010011;
assign LUT_2[13274] = 32'b11111111111111111001110101110110;
assign LUT_2[13275] = 32'b11111111111111110110101110001111;
assign LUT_2[13276] = 32'b11111111111111101111011010100010;
assign LUT_2[13277] = 32'b11111111111111101100010010111011;
assign LUT_2[13278] = 32'b11111111111111110110010011011110;
assign LUT_2[13279] = 32'b11111111111111110011001011110111;
assign LUT_2[13280] = 32'b11111111111111111110000010111100;
assign LUT_2[13281] = 32'b11111111111111111010111011010101;
assign LUT_2[13282] = 32'b00000000000000000100111011111000;
assign LUT_2[13283] = 32'b00000000000000000001110100010001;
assign LUT_2[13284] = 32'b11111111111111111010100000100100;
assign LUT_2[13285] = 32'b11111111111111110111011000111101;
assign LUT_2[13286] = 32'b00000000000000000001011001100000;
assign LUT_2[13287] = 32'b11111111111111111110010001111001;
assign LUT_2[13288] = 32'b11111111111111111000110100011001;
assign LUT_2[13289] = 32'b11111111111111110101101100110010;
assign LUT_2[13290] = 32'b11111111111111111111101101010101;
assign LUT_2[13291] = 32'b11111111111111111100100101101110;
assign LUT_2[13292] = 32'b11111111111111110101010010000001;
assign LUT_2[13293] = 32'b11111111111111110010001010011010;
assign LUT_2[13294] = 32'b11111111111111111100001010111101;
assign LUT_2[13295] = 32'b11111111111111111001000011010110;
assign LUT_2[13296] = 32'b11111111111111111000100111000110;
assign LUT_2[13297] = 32'b11111111111111110101011111011111;
assign LUT_2[13298] = 32'b11111111111111111111100000000010;
assign LUT_2[13299] = 32'b11111111111111111100011000011011;
assign LUT_2[13300] = 32'b11111111111111110101000100101110;
assign LUT_2[13301] = 32'b11111111111111110001111101000111;
assign LUT_2[13302] = 32'b11111111111111111011111101101010;
assign LUT_2[13303] = 32'b11111111111111111000110110000011;
assign LUT_2[13304] = 32'b11111111111111110011011000100011;
assign LUT_2[13305] = 32'b11111111111111110000010000111100;
assign LUT_2[13306] = 32'b11111111111111111010010001011111;
assign LUT_2[13307] = 32'b11111111111111110111001001111000;
assign LUT_2[13308] = 32'b11111111111111101111110110001011;
assign LUT_2[13309] = 32'b11111111111111101100101110100100;
assign LUT_2[13310] = 32'b11111111111111110110101111000111;
assign LUT_2[13311] = 32'b11111111111111110011100111100000;
assign LUT_2[13312] = 32'b11111111111111111111000110001110;
assign LUT_2[13313] = 32'b11111111111111111011111110100111;
assign LUT_2[13314] = 32'b00000000000000000101111111001010;
assign LUT_2[13315] = 32'b00000000000000000010110111100011;
assign LUT_2[13316] = 32'b11111111111111111011100011110110;
assign LUT_2[13317] = 32'b11111111111111111000011100001111;
assign LUT_2[13318] = 32'b00000000000000000010011100110010;
assign LUT_2[13319] = 32'b11111111111111111111010101001011;
assign LUT_2[13320] = 32'b11111111111111111001110111101011;
assign LUT_2[13321] = 32'b11111111111111110110110000000100;
assign LUT_2[13322] = 32'b00000000000000000000110000100111;
assign LUT_2[13323] = 32'b11111111111111111101101001000000;
assign LUT_2[13324] = 32'b11111111111111110110010101010011;
assign LUT_2[13325] = 32'b11111111111111110011001101101100;
assign LUT_2[13326] = 32'b11111111111111111101001110001111;
assign LUT_2[13327] = 32'b11111111111111111010000110101000;
assign LUT_2[13328] = 32'b11111111111111111001101010011000;
assign LUT_2[13329] = 32'b11111111111111110110100010110001;
assign LUT_2[13330] = 32'b00000000000000000000100011010100;
assign LUT_2[13331] = 32'b11111111111111111101011011101101;
assign LUT_2[13332] = 32'b11111111111111110110001000000000;
assign LUT_2[13333] = 32'b11111111111111110011000000011001;
assign LUT_2[13334] = 32'b11111111111111111101000000111100;
assign LUT_2[13335] = 32'b11111111111111111001111001010101;
assign LUT_2[13336] = 32'b11111111111111110100011011110101;
assign LUT_2[13337] = 32'b11111111111111110001010100001110;
assign LUT_2[13338] = 32'b11111111111111111011010100110001;
assign LUT_2[13339] = 32'b11111111111111111000001101001010;
assign LUT_2[13340] = 32'b11111111111111110000111001011101;
assign LUT_2[13341] = 32'b11111111111111101101110001110110;
assign LUT_2[13342] = 32'b11111111111111110111110010011001;
assign LUT_2[13343] = 32'b11111111111111110100101010110010;
assign LUT_2[13344] = 32'b11111111111111111111100001110111;
assign LUT_2[13345] = 32'b11111111111111111100011010010000;
assign LUT_2[13346] = 32'b00000000000000000110011010110011;
assign LUT_2[13347] = 32'b00000000000000000011010011001100;
assign LUT_2[13348] = 32'b11111111111111111011111111011111;
assign LUT_2[13349] = 32'b11111111111111111000110111111000;
assign LUT_2[13350] = 32'b00000000000000000010111000011011;
assign LUT_2[13351] = 32'b11111111111111111111110000110100;
assign LUT_2[13352] = 32'b11111111111111111010010011010100;
assign LUT_2[13353] = 32'b11111111111111110111001011101101;
assign LUT_2[13354] = 32'b00000000000000000001001100010000;
assign LUT_2[13355] = 32'b11111111111111111110000100101001;
assign LUT_2[13356] = 32'b11111111111111110110110000111100;
assign LUT_2[13357] = 32'b11111111111111110011101001010101;
assign LUT_2[13358] = 32'b11111111111111111101101001111000;
assign LUT_2[13359] = 32'b11111111111111111010100010010001;
assign LUT_2[13360] = 32'b11111111111111111010000110000001;
assign LUT_2[13361] = 32'b11111111111111110110111110011010;
assign LUT_2[13362] = 32'b00000000000000000000111110111101;
assign LUT_2[13363] = 32'b11111111111111111101110111010110;
assign LUT_2[13364] = 32'b11111111111111110110100011101001;
assign LUT_2[13365] = 32'b11111111111111110011011100000010;
assign LUT_2[13366] = 32'b11111111111111111101011100100101;
assign LUT_2[13367] = 32'b11111111111111111010010100111110;
assign LUT_2[13368] = 32'b11111111111111110100110111011110;
assign LUT_2[13369] = 32'b11111111111111110001101111110111;
assign LUT_2[13370] = 32'b11111111111111111011110000011010;
assign LUT_2[13371] = 32'b11111111111111111000101000110011;
assign LUT_2[13372] = 32'b11111111111111110001010101000110;
assign LUT_2[13373] = 32'b11111111111111101110001101011111;
assign LUT_2[13374] = 32'b11111111111111111000001110000010;
assign LUT_2[13375] = 32'b11111111111111110101000110011011;
assign LUT_2[13376] = 32'b11111111111111110111001110110001;
assign LUT_2[13377] = 32'b11111111111111110100000111001010;
assign LUT_2[13378] = 32'b11111111111111111110000111101101;
assign LUT_2[13379] = 32'b11111111111111111011000000000110;
assign LUT_2[13380] = 32'b11111111111111110011101100011001;
assign LUT_2[13381] = 32'b11111111111111110000100100110010;
assign LUT_2[13382] = 32'b11111111111111111010100101010101;
assign LUT_2[13383] = 32'b11111111111111110111011101101110;
assign LUT_2[13384] = 32'b11111111111111110010000000001110;
assign LUT_2[13385] = 32'b11111111111111101110111000100111;
assign LUT_2[13386] = 32'b11111111111111111000111001001010;
assign LUT_2[13387] = 32'b11111111111111110101110001100011;
assign LUT_2[13388] = 32'b11111111111111101110011101110110;
assign LUT_2[13389] = 32'b11111111111111101011010110001111;
assign LUT_2[13390] = 32'b11111111111111110101010110110010;
assign LUT_2[13391] = 32'b11111111111111110010001111001011;
assign LUT_2[13392] = 32'b11111111111111110001110010111011;
assign LUT_2[13393] = 32'b11111111111111101110101011010100;
assign LUT_2[13394] = 32'b11111111111111111000101011110111;
assign LUT_2[13395] = 32'b11111111111111110101100100010000;
assign LUT_2[13396] = 32'b11111111111111101110010000100011;
assign LUT_2[13397] = 32'b11111111111111101011001000111100;
assign LUT_2[13398] = 32'b11111111111111110101001001011111;
assign LUT_2[13399] = 32'b11111111111111110010000001111000;
assign LUT_2[13400] = 32'b11111111111111101100100100011000;
assign LUT_2[13401] = 32'b11111111111111101001011100110001;
assign LUT_2[13402] = 32'b11111111111111110011011101010100;
assign LUT_2[13403] = 32'b11111111111111110000010101101101;
assign LUT_2[13404] = 32'b11111111111111101001000010000000;
assign LUT_2[13405] = 32'b11111111111111100101111010011001;
assign LUT_2[13406] = 32'b11111111111111101111111010111100;
assign LUT_2[13407] = 32'b11111111111111101100110011010101;
assign LUT_2[13408] = 32'b11111111111111110111101010011010;
assign LUT_2[13409] = 32'b11111111111111110100100010110011;
assign LUT_2[13410] = 32'b11111111111111111110100011010110;
assign LUT_2[13411] = 32'b11111111111111111011011011101111;
assign LUT_2[13412] = 32'b11111111111111110100001000000010;
assign LUT_2[13413] = 32'b11111111111111110001000000011011;
assign LUT_2[13414] = 32'b11111111111111111011000000111110;
assign LUT_2[13415] = 32'b11111111111111110111111001010111;
assign LUT_2[13416] = 32'b11111111111111110010011011110111;
assign LUT_2[13417] = 32'b11111111111111101111010100010000;
assign LUT_2[13418] = 32'b11111111111111111001010100110011;
assign LUT_2[13419] = 32'b11111111111111110110001101001100;
assign LUT_2[13420] = 32'b11111111111111101110111001011111;
assign LUT_2[13421] = 32'b11111111111111101011110001111000;
assign LUT_2[13422] = 32'b11111111111111110101110010011011;
assign LUT_2[13423] = 32'b11111111111111110010101010110100;
assign LUT_2[13424] = 32'b11111111111111110010001110100100;
assign LUT_2[13425] = 32'b11111111111111101111000110111101;
assign LUT_2[13426] = 32'b11111111111111111001000111100000;
assign LUT_2[13427] = 32'b11111111111111110101111111111001;
assign LUT_2[13428] = 32'b11111111111111101110101100001100;
assign LUT_2[13429] = 32'b11111111111111101011100100100101;
assign LUT_2[13430] = 32'b11111111111111110101100101001000;
assign LUT_2[13431] = 32'b11111111111111110010011101100001;
assign LUT_2[13432] = 32'b11111111111111101101000000000001;
assign LUT_2[13433] = 32'b11111111111111101001111000011010;
assign LUT_2[13434] = 32'b11111111111111110011111000111101;
assign LUT_2[13435] = 32'b11111111111111110000110001010110;
assign LUT_2[13436] = 32'b11111111111111101001011101101001;
assign LUT_2[13437] = 32'b11111111111111100110010110000010;
assign LUT_2[13438] = 32'b11111111111111110000010110100101;
assign LUT_2[13439] = 32'b11111111111111101101001110111110;
assign LUT_2[13440] = 32'b00000000000000000011011010011101;
assign LUT_2[13441] = 32'b00000000000000000000010010110110;
assign LUT_2[13442] = 32'b00000000000000001010010011011001;
assign LUT_2[13443] = 32'b00000000000000000111001011110010;
assign LUT_2[13444] = 32'b11111111111111111111111000000101;
assign LUT_2[13445] = 32'b11111111111111111100110000011110;
assign LUT_2[13446] = 32'b00000000000000000110110001000001;
assign LUT_2[13447] = 32'b00000000000000000011101001011010;
assign LUT_2[13448] = 32'b11111111111111111110001011111010;
assign LUT_2[13449] = 32'b11111111111111111011000100010011;
assign LUT_2[13450] = 32'b00000000000000000101000100110110;
assign LUT_2[13451] = 32'b00000000000000000001111101001111;
assign LUT_2[13452] = 32'b11111111111111111010101001100010;
assign LUT_2[13453] = 32'b11111111111111110111100001111011;
assign LUT_2[13454] = 32'b00000000000000000001100010011110;
assign LUT_2[13455] = 32'b11111111111111111110011010110111;
assign LUT_2[13456] = 32'b11111111111111111101111110100111;
assign LUT_2[13457] = 32'b11111111111111111010110111000000;
assign LUT_2[13458] = 32'b00000000000000000100110111100011;
assign LUT_2[13459] = 32'b00000000000000000001101111111100;
assign LUT_2[13460] = 32'b11111111111111111010011100001111;
assign LUT_2[13461] = 32'b11111111111111110111010100101000;
assign LUT_2[13462] = 32'b00000000000000000001010101001011;
assign LUT_2[13463] = 32'b11111111111111111110001101100100;
assign LUT_2[13464] = 32'b11111111111111111000110000000100;
assign LUT_2[13465] = 32'b11111111111111110101101000011101;
assign LUT_2[13466] = 32'b11111111111111111111101001000000;
assign LUT_2[13467] = 32'b11111111111111111100100001011001;
assign LUT_2[13468] = 32'b11111111111111110101001101101100;
assign LUT_2[13469] = 32'b11111111111111110010000110000101;
assign LUT_2[13470] = 32'b11111111111111111100000110101000;
assign LUT_2[13471] = 32'b11111111111111111000111111000001;
assign LUT_2[13472] = 32'b00000000000000000011110110000110;
assign LUT_2[13473] = 32'b00000000000000000000101110011111;
assign LUT_2[13474] = 32'b00000000000000001010101111000010;
assign LUT_2[13475] = 32'b00000000000000000111100111011011;
assign LUT_2[13476] = 32'b00000000000000000000010011101110;
assign LUT_2[13477] = 32'b11111111111111111101001100000111;
assign LUT_2[13478] = 32'b00000000000000000111001100101010;
assign LUT_2[13479] = 32'b00000000000000000100000101000011;
assign LUT_2[13480] = 32'b11111111111111111110100111100011;
assign LUT_2[13481] = 32'b11111111111111111011011111111100;
assign LUT_2[13482] = 32'b00000000000000000101100000011111;
assign LUT_2[13483] = 32'b00000000000000000010011000111000;
assign LUT_2[13484] = 32'b11111111111111111011000101001011;
assign LUT_2[13485] = 32'b11111111111111110111111101100100;
assign LUT_2[13486] = 32'b00000000000000000001111110000111;
assign LUT_2[13487] = 32'b11111111111111111110110110100000;
assign LUT_2[13488] = 32'b11111111111111111110011010010000;
assign LUT_2[13489] = 32'b11111111111111111011010010101001;
assign LUT_2[13490] = 32'b00000000000000000101010011001100;
assign LUT_2[13491] = 32'b00000000000000000010001011100101;
assign LUT_2[13492] = 32'b11111111111111111010110111111000;
assign LUT_2[13493] = 32'b11111111111111110111110000010001;
assign LUT_2[13494] = 32'b00000000000000000001110000110100;
assign LUT_2[13495] = 32'b11111111111111111110101001001101;
assign LUT_2[13496] = 32'b11111111111111111001001011101101;
assign LUT_2[13497] = 32'b11111111111111110110000100000110;
assign LUT_2[13498] = 32'b00000000000000000000000100101001;
assign LUT_2[13499] = 32'b11111111111111111100111101000010;
assign LUT_2[13500] = 32'b11111111111111110101101001010101;
assign LUT_2[13501] = 32'b11111111111111110010100001101110;
assign LUT_2[13502] = 32'b11111111111111111100100010010001;
assign LUT_2[13503] = 32'b11111111111111111001011010101010;
assign LUT_2[13504] = 32'b11111111111111111011100011000000;
assign LUT_2[13505] = 32'b11111111111111111000011011011001;
assign LUT_2[13506] = 32'b00000000000000000010011011111100;
assign LUT_2[13507] = 32'b11111111111111111111010100010101;
assign LUT_2[13508] = 32'b11111111111111111000000000101000;
assign LUT_2[13509] = 32'b11111111111111110100111001000001;
assign LUT_2[13510] = 32'b11111111111111111110111001100100;
assign LUT_2[13511] = 32'b11111111111111111011110001111101;
assign LUT_2[13512] = 32'b11111111111111110110010100011101;
assign LUT_2[13513] = 32'b11111111111111110011001100110110;
assign LUT_2[13514] = 32'b11111111111111111101001101011001;
assign LUT_2[13515] = 32'b11111111111111111010000101110010;
assign LUT_2[13516] = 32'b11111111111111110010110010000101;
assign LUT_2[13517] = 32'b11111111111111101111101010011110;
assign LUT_2[13518] = 32'b11111111111111111001101011000001;
assign LUT_2[13519] = 32'b11111111111111110110100011011010;
assign LUT_2[13520] = 32'b11111111111111110110000111001010;
assign LUT_2[13521] = 32'b11111111111111110010111111100011;
assign LUT_2[13522] = 32'b11111111111111111101000000000110;
assign LUT_2[13523] = 32'b11111111111111111001111000011111;
assign LUT_2[13524] = 32'b11111111111111110010100100110010;
assign LUT_2[13525] = 32'b11111111111111101111011101001011;
assign LUT_2[13526] = 32'b11111111111111111001011101101110;
assign LUT_2[13527] = 32'b11111111111111110110010110000111;
assign LUT_2[13528] = 32'b11111111111111110000111000100111;
assign LUT_2[13529] = 32'b11111111111111101101110001000000;
assign LUT_2[13530] = 32'b11111111111111110111110001100011;
assign LUT_2[13531] = 32'b11111111111111110100101001111100;
assign LUT_2[13532] = 32'b11111111111111101101010110001111;
assign LUT_2[13533] = 32'b11111111111111101010001110101000;
assign LUT_2[13534] = 32'b11111111111111110100001111001011;
assign LUT_2[13535] = 32'b11111111111111110001000111100100;
assign LUT_2[13536] = 32'b11111111111111111011111110101001;
assign LUT_2[13537] = 32'b11111111111111111000110111000010;
assign LUT_2[13538] = 32'b00000000000000000010110111100101;
assign LUT_2[13539] = 32'b11111111111111111111101111111110;
assign LUT_2[13540] = 32'b11111111111111111000011100010001;
assign LUT_2[13541] = 32'b11111111111111110101010100101010;
assign LUT_2[13542] = 32'b11111111111111111111010101001101;
assign LUT_2[13543] = 32'b11111111111111111100001101100110;
assign LUT_2[13544] = 32'b11111111111111110110110000000110;
assign LUT_2[13545] = 32'b11111111111111110011101000011111;
assign LUT_2[13546] = 32'b11111111111111111101101001000010;
assign LUT_2[13547] = 32'b11111111111111111010100001011011;
assign LUT_2[13548] = 32'b11111111111111110011001101101110;
assign LUT_2[13549] = 32'b11111111111111110000000110000111;
assign LUT_2[13550] = 32'b11111111111111111010000110101010;
assign LUT_2[13551] = 32'b11111111111111110110111111000011;
assign LUT_2[13552] = 32'b11111111111111110110100010110011;
assign LUT_2[13553] = 32'b11111111111111110011011011001100;
assign LUT_2[13554] = 32'b11111111111111111101011011101111;
assign LUT_2[13555] = 32'b11111111111111111010010100001000;
assign LUT_2[13556] = 32'b11111111111111110011000000011011;
assign LUT_2[13557] = 32'b11111111111111101111111000110100;
assign LUT_2[13558] = 32'b11111111111111111001111001010111;
assign LUT_2[13559] = 32'b11111111111111110110110001110000;
assign LUT_2[13560] = 32'b11111111111111110001010100010000;
assign LUT_2[13561] = 32'b11111111111111101110001100101001;
assign LUT_2[13562] = 32'b11111111111111111000001101001100;
assign LUT_2[13563] = 32'b11111111111111110101000101100101;
assign LUT_2[13564] = 32'b11111111111111101101110001111000;
assign LUT_2[13565] = 32'b11111111111111101010101010010001;
assign LUT_2[13566] = 32'b11111111111111110100101010110100;
assign LUT_2[13567] = 32'b11111111111111110001100011001101;
assign LUT_2[13568] = 32'b00000000000000000011000100110100;
assign LUT_2[13569] = 32'b11111111111111111111111101001101;
assign LUT_2[13570] = 32'b00000000000000001001111101110000;
assign LUT_2[13571] = 32'b00000000000000000110110110001001;
assign LUT_2[13572] = 32'b11111111111111111111100010011100;
assign LUT_2[13573] = 32'b11111111111111111100011010110101;
assign LUT_2[13574] = 32'b00000000000000000110011011011000;
assign LUT_2[13575] = 32'b00000000000000000011010011110001;
assign LUT_2[13576] = 32'b11111111111111111101110110010001;
assign LUT_2[13577] = 32'b11111111111111111010101110101010;
assign LUT_2[13578] = 32'b00000000000000000100101111001101;
assign LUT_2[13579] = 32'b00000000000000000001100111100110;
assign LUT_2[13580] = 32'b11111111111111111010010011111001;
assign LUT_2[13581] = 32'b11111111111111110111001100010010;
assign LUT_2[13582] = 32'b00000000000000000001001100110101;
assign LUT_2[13583] = 32'b11111111111111111110000101001110;
assign LUT_2[13584] = 32'b11111111111111111101101000111110;
assign LUT_2[13585] = 32'b11111111111111111010100001010111;
assign LUT_2[13586] = 32'b00000000000000000100100001111010;
assign LUT_2[13587] = 32'b00000000000000000001011010010011;
assign LUT_2[13588] = 32'b11111111111111111010000110100110;
assign LUT_2[13589] = 32'b11111111111111110110111110111111;
assign LUT_2[13590] = 32'b00000000000000000000111111100010;
assign LUT_2[13591] = 32'b11111111111111111101110111111011;
assign LUT_2[13592] = 32'b11111111111111111000011010011011;
assign LUT_2[13593] = 32'b11111111111111110101010010110100;
assign LUT_2[13594] = 32'b11111111111111111111010011010111;
assign LUT_2[13595] = 32'b11111111111111111100001011110000;
assign LUT_2[13596] = 32'b11111111111111110100111000000011;
assign LUT_2[13597] = 32'b11111111111111110001110000011100;
assign LUT_2[13598] = 32'b11111111111111111011110000111111;
assign LUT_2[13599] = 32'b11111111111111111000101001011000;
assign LUT_2[13600] = 32'b00000000000000000011100000011101;
assign LUT_2[13601] = 32'b00000000000000000000011000110110;
assign LUT_2[13602] = 32'b00000000000000001010011001011001;
assign LUT_2[13603] = 32'b00000000000000000111010001110010;
assign LUT_2[13604] = 32'b11111111111111111111111110000101;
assign LUT_2[13605] = 32'b11111111111111111100110110011110;
assign LUT_2[13606] = 32'b00000000000000000110110111000001;
assign LUT_2[13607] = 32'b00000000000000000011101111011010;
assign LUT_2[13608] = 32'b11111111111111111110010001111010;
assign LUT_2[13609] = 32'b11111111111111111011001010010011;
assign LUT_2[13610] = 32'b00000000000000000101001010110110;
assign LUT_2[13611] = 32'b00000000000000000010000011001111;
assign LUT_2[13612] = 32'b11111111111111111010101111100010;
assign LUT_2[13613] = 32'b11111111111111110111100111111011;
assign LUT_2[13614] = 32'b00000000000000000001101000011110;
assign LUT_2[13615] = 32'b11111111111111111110100000110111;
assign LUT_2[13616] = 32'b11111111111111111110000100100111;
assign LUT_2[13617] = 32'b11111111111111111010111101000000;
assign LUT_2[13618] = 32'b00000000000000000100111101100011;
assign LUT_2[13619] = 32'b00000000000000000001110101111100;
assign LUT_2[13620] = 32'b11111111111111111010100010001111;
assign LUT_2[13621] = 32'b11111111111111110111011010101000;
assign LUT_2[13622] = 32'b00000000000000000001011011001011;
assign LUT_2[13623] = 32'b11111111111111111110010011100100;
assign LUT_2[13624] = 32'b11111111111111111000110110000100;
assign LUT_2[13625] = 32'b11111111111111110101101110011101;
assign LUT_2[13626] = 32'b11111111111111111111101111000000;
assign LUT_2[13627] = 32'b11111111111111111100100111011001;
assign LUT_2[13628] = 32'b11111111111111110101010011101100;
assign LUT_2[13629] = 32'b11111111111111110010001100000101;
assign LUT_2[13630] = 32'b11111111111111111100001100101000;
assign LUT_2[13631] = 32'b11111111111111111001000101000001;
assign LUT_2[13632] = 32'b11111111111111111011001101010111;
assign LUT_2[13633] = 32'b11111111111111111000000101110000;
assign LUT_2[13634] = 32'b00000000000000000010000110010011;
assign LUT_2[13635] = 32'b11111111111111111110111110101100;
assign LUT_2[13636] = 32'b11111111111111110111101010111111;
assign LUT_2[13637] = 32'b11111111111111110100100011011000;
assign LUT_2[13638] = 32'b11111111111111111110100011111011;
assign LUT_2[13639] = 32'b11111111111111111011011100010100;
assign LUT_2[13640] = 32'b11111111111111110101111110110100;
assign LUT_2[13641] = 32'b11111111111111110010110111001101;
assign LUT_2[13642] = 32'b11111111111111111100110111110000;
assign LUT_2[13643] = 32'b11111111111111111001110000001001;
assign LUT_2[13644] = 32'b11111111111111110010011100011100;
assign LUT_2[13645] = 32'b11111111111111101111010100110101;
assign LUT_2[13646] = 32'b11111111111111111001010101011000;
assign LUT_2[13647] = 32'b11111111111111110110001101110001;
assign LUT_2[13648] = 32'b11111111111111110101110001100001;
assign LUT_2[13649] = 32'b11111111111111110010101001111010;
assign LUT_2[13650] = 32'b11111111111111111100101010011101;
assign LUT_2[13651] = 32'b11111111111111111001100010110110;
assign LUT_2[13652] = 32'b11111111111111110010001111001001;
assign LUT_2[13653] = 32'b11111111111111101111000111100010;
assign LUT_2[13654] = 32'b11111111111111111001001000000101;
assign LUT_2[13655] = 32'b11111111111111110110000000011110;
assign LUT_2[13656] = 32'b11111111111111110000100010111110;
assign LUT_2[13657] = 32'b11111111111111101101011011010111;
assign LUT_2[13658] = 32'b11111111111111110111011011111010;
assign LUT_2[13659] = 32'b11111111111111110100010100010011;
assign LUT_2[13660] = 32'b11111111111111101101000000100110;
assign LUT_2[13661] = 32'b11111111111111101001111000111111;
assign LUT_2[13662] = 32'b11111111111111110011111001100010;
assign LUT_2[13663] = 32'b11111111111111110000110001111011;
assign LUT_2[13664] = 32'b11111111111111111011101001000000;
assign LUT_2[13665] = 32'b11111111111111111000100001011001;
assign LUT_2[13666] = 32'b00000000000000000010100001111100;
assign LUT_2[13667] = 32'b11111111111111111111011010010101;
assign LUT_2[13668] = 32'b11111111111111111000000110101000;
assign LUT_2[13669] = 32'b11111111111111110100111111000001;
assign LUT_2[13670] = 32'b11111111111111111110111111100100;
assign LUT_2[13671] = 32'b11111111111111111011110111111101;
assign LUT_2[13672] = 32'b11111111111111110110011010011101;
assign LUT_2[13673] = 32'b11111111111111110011010010110110;
assign LUT_2[13674] = 32'b11111111111111111101010011011001;
assign LUT_2[13675] = 32'b11111111111111111010001011110010;
assign LUT_2[13676] = 32'b11111111111111110010111000000101;
assign LUT_2[13677] = 32'b11111111111111101111110000011110;
assign LUT_2[13678] = 32'b11111111111111111001110001000001;
assign LUT_2[13679] = 32'b11111111111111110110101001011010;
assign LUT_2[13680] = 32'b11111111111111110110001101001010;
assign LUT_2[13681] = 32'b11111111111111110011000101100011;
assign LUT_2[13682] = 32'b11111111111111111101000110000110;
assign LUT_2[13683] = 32'b11111111111111111001111110011111;
assign LUT_2[13684] = 32'b11111111111111110010101010110010;
assign LUT_2[13685] = 32'b11111111111111101111100011001011;
assign LUT_2[13686] = 32'b11111111111111111001100011101110;
assign LUT_2[13687] = 32'b11111111111111110110011100000111;
assign LUT_2[13688] = 32'b11111111111111110000111110100111;
assign LUT_2[13689] = 32'b11111111111111101101110111000000;
assign LUT_2[13690] = 32'b11111111111111110111110111100011;
assign LUT_2[13691] = 32'b11111111111111110100101111111100;
assign LUT_2[13692] = 32'b11111111111111101101011100001111;
assign LUT_2[13693] = 32'b11111111111111101010010100101000;
assign LUT_2[13694] = 32'b11111111111111110100010101001011;
assign LUT_2[13695] = 32'b11111111111111110001001101100100;
assign LUT_2[13696] = 32'b00000000000000000111011001000011;
assign LUT_2[13697] = 32'b00000000000000000100010001011100;
assign LUT_2[13698] = 32'b00000000000000001110010001111111;
assign LUT_2[13699] = 32'b00000000000000001011001010011000;
assign LUT_2[13700] = 32'b00000000000000000011110110101011;
assign LUT_2[13701] = 32'b00000000000000000000101111000100;
assign LUT_2[13702] = 32'b00000000000000001010101111100111;
assign LUT_2[13703] = 32'b00000000000000000111101000000000;
assign LUT_2[13704] = 32'b00000000000000000010001010100000;
assign LUT_2[13705] = 32'b11111111111111111111000010111001;
assign LUT_2[13706] = 32'b00000000000000001001000011011100;
assign LUT_2[13707] = 32'b00000000000000000101111011110101;
assign LUT_2[13708] = 32'b11111111111111111110101000001000;
assign LUT_2[13709] = 32'b11111111111111111011100000100001;
assign LUT_2[13710] = 32'b00000000000000000101100001000100;
assign LUT_2[13711] = 32'b00000000000000000010011001011101;
assign LUT_2[13712] = 32'b00000000000000000001111101001101;
assign LUT_2[13713] = 32'b11111111111111111110110101100110;
assign LUT_2[13714] = 32'b00000000000000001000110110001001;
assign LUT_2[13715] = 32'b00000000000000000101101110100010;
assign LUT_2[13716] = 32'b11111111111111111110011010110101;
assign LUT_2[13717] = 32'b11111111111111111011010011001110;
assign LUT_2[13718] = 32'b00000000000000000101010011110001;
assign LUT_2[13719] = 32'b00000000000000000010001100001010;
assign LUT_2[13720] = 32'b11111111111111111100101110101010;
assign LUT_2[13721] = 32'b11111111111111111001100111000011;
assign LUT_2[13722] = 32'b00000000000000000011100111100110;
assign LUT_2[13723] = 32'b00000000000000000000011111111111;
assign LUT_2[13724] = 32'b11111111111111111001001100010010;
assign LUT_2[13725] = 32'b11111111111111110110000100101011;
assign LUT_2[13726] = 32'b00000000000000000000000101001110;
assign LUT_2[13727] = 32'b11111111111111111100111101100111;
assign LUT_2[13728] = 32'b00000000000000000111110100101100;
assign LUT_2[13729] = 32'b00000000000000000100101101000101;
assign LUT_2[13730] = 32'b00000000000000001110101101101000;
assign LUT_2[13731] = 32'b00000000000000001011100110000001;
assign LUT_2[13732] = 32'b00000000000000000100010010010100;
assign LUT_2[13733] = 32'b00000000000000000001001010101101;
assign LUT_2[13734] = 32'b00000000000000001011001011010000;
assign LUT_2[13735] = 32'b00000000000000001000000011101001;
assign LUT_2[13736] = 32'b00000000000000000010100110001001;
assign LUT_2[13737] = 32'b11111111111111111111011110100010;
assign LUT_2[13738] = 32'b00000000000000001001011111000101;
assign LUT_2[13739] = 32'b00000000000000000110010111011110;
assign LUT_2[13740] = 32'b11111111111111111111000011110001;
assign LUT_2[13741] = 32'b11111111111111111011111100001010;
assign LUT_2[13742] = 32'b00000000000000000101111100101101;
assign LUT_2[13743] = 32'b00000000000000000010110101000110;
assign LUT_2[13744] = 32'b00000000000000000010011000110110;
assign LUT_2[13745] = 32'b11111111111111111111010001001111;
assign LUT_2[13746] = 32'b00000000000000001001010001110010;
assign LUT_2[13747] = 32'b00000000000000000110001010001011;
assign LUT_2[13748] = 32'b11111111111111111110110110011110;
assign LUT_2[13749] = 32'b11111111111111111011101110110111;
assign LUT_2[13750] = 32'b00000000000000000101101111011010;
assign LUT_2[13751] = 32'b00000000000000000010100111110011;
assign LUT_2[13752] = 32'b11111111111111111101001010010011;
assign LUT_2[13753] = 32'b11111111111111111010000010101100;
assign LUT_2[13754] = 32'b00000000000000000100000011001111;
assign LUT_2[13755] = 32'b00000000000000000000111011101000;
assign LUT_2[13756] = 32'b11111111111111111001100111111011;
assign LUT_2[13757] = 32'b11111111111111110110100000010100;
assign LUT_2[13758] = 32'b00000000000000000000100000110111;
assign LUT_2[13759] = 32'b11111111111111111101011001010000;
assign LUT_2[13760] = 32'b11111111111111111111100001100110;
assign LUT_2[13761] = 32'b11111111111111111100011001111111;
assign LUT_2[13762] = 32'b00000000000000000110011010100010;
assign LUT_2[13763] = 32'b00000000000000000011010010111011;
assign LUT_2[13764] = 32'b11111111111111111011111111001110;
assign LUT_2[13765] = 32'b11111111111111111000110111100111;
assign LUT_2[13766] = 32'b00000000000000000010111000001010;
assign LUT_2[13767] = 32'b11111111111111111111110000100011;
assign LUT_2[13768] = 32'b11111111111111111010010011000011;
assign LUT_2[13769] = 32'b11111111111111110111001011011100;
assign LUT_2[13770] = 32'b00000000000000000001001011111111;
assign LUT_2[13771] = 32'b11111111111111111110000100011000;
assign LUT_2[13772] = 32'b11111111111111110110110000101011;
assign LUT_2[13773] = 32'b11111111111111110011101001000100;
assign LUT_2[13774] = 32'b11111111111111111101101001100111;
assign LUT_2[13775] = 32'b11111111111111111010100010000000;
assign LUT_2[13776] = 32'b11111111111111111010000101110000;
assign LUT_2[13777] = 32'b11111111111111110110111110001001;
assign LUT_2[13778] = 32'b00000000000000000000111110101100;
assign LUT_2[13779] = 32'b11111111111111111101110111000101;
assign LUT_2[13780] = 32'b11111111111111110110100011011000;
assign LUT_2[13781] = 32'b11111111111111110011011011110001;
assign LUT_2[13782] = 32'b11111111111111111101011100010100;
assign LUT_2[13783] = 32'b11111111111111111010010100101101;
assign LUT_2[13784] = 32'b11111111111111110100110111001101;
assign LUT_2[13785] = 32'b11111111111111110001101111100110;
assign LUT_2[13786] = 32'b11111111111111111011110000001001;
assign LUT_2[13787] = 32'b11111111111111111000101000100010;
assign LUT_2[13788] = 32'b11111111111111110001010100110101;
assign LUT_2[13789] = 32'b11111111111111101110001101001110;
assign LUT_2[13790] = 32'b11111111111111111000001101110001;
assign LUT_2[13791] = 32'b11111111111111110101000110001010;
assign LUT_2[13792] = 32'b11111111111111111111111101001111;
assign LUT_2[13793] = 32'b11111111111111111100110101101000;
assign LUT_2[13794] = 32'b00000000000000000110110110001011;
assign LUT_2[13795] = 32'b00000000000000000011101110100100;
assign LUT_2[13796] = 32'b11111111111111111100011010110111;
assign LUT_2[13797] = 32'b11111111111111111001010011010000;
assign LUT_2[13798] = 32'b00000000000000000011010011110011;
assign LUT_2[13799] = 32'b00000000000000000000001100001100;
assign LUT_2[13800] = 32'b11111111111111111010101110101100;
assign LUT_2[13801] = 32'b11111111111111110111100111000101;
assign LUT_2[13802] = 32'b00000000000000000001100111101000;
assign LUT_2[13803] = 32'b11111111111111111110100000000001;
assign LUT_2[13804] = 32'b11111111111111110111001100010100;
assign LUT_2[13805] = 32'b11111111111111110100000100101101;
assign LUT_2[13806] = 32'b11111111111111111110000101010000;
assign LUT_2[13807] = 32'b11111111111111111010111101101001;
assign LUT_2[13808] = 32'b11111111111111111010100001011001;
assign LUT_2[13809] = 32'b11111111111111110111011001110010;
assign LUT_2[13810] = 32'b00000000000000000001011010010101;
assign LUT_2[13811] = 32'b11111111111111111110010010101110;
assign LUT_2[13812] = 32'b11111111111111110110111111000001;
assign LUT_2[13813] = 32'b11111111111111110011110111011010;
assign LUT_2[13814] = 32'b11111111111111111101110111111101;
assign LUT_2[13815] = 32'b11111111111111111010110000010110;
assign LUT_2[13816] = 32'b11111111111111110101010010110110;
assign LUT_2[13817] = 32'b11111111111111110010001011001111;
assign LUT_2[13818] = 32'b11111111111111111100001011110010;
assign LUT_2[13819] = 32'b11111111111111111001000100001011;
assign LUT_2[13820] = 32'b11111111111111110001110000011110;
assign LUT_2[13821] = 32'b11111111111111101110101000110111;
assign LUT_2[13822] = 32'b11111111111111111000101001011010;
assign LUT_2[13823] = 32'b11111111111111110101100001110011;
assign LUT_2[13824] = 32'b00000000000000000011111000000000;
assign LUT_2[13825] = 32'b00000000000000000000110000011001;
assign LUT_2[13826] = 32'b00000000000000001010110000111100;
assign LUT_2[13827] = 32'b00000000000000000111101001010101;
assign LUT_2[13828] = 32'b00000000000000000000010101101000;
assign LUT_2[13829] = 32'b11111111111111111101001110000001;
assign LUT_2[13830] = 32'b00000000000000000111001110100100;
assign LUT_2[13831] = 32'b00000000000000000100000110111101;
assign LUT_2[13832] = 32'b11111111111111111110101001011101;
assign LUT_2[13833] = 32'b11111111111111111011100001110110;
assign LUT_2[13834] = 32'b00000000000000000101100010011001;
assign LUT_2[13835] = 32'b00000000000000000010011010110010;
assign LUT_2[13836] = 32'b11111111111111111011000111000101;
assign LUT_2[13837] = 32'b11111111111111110111111111011110;
assign LUT_2[13838] = 32'b00000000000000000010000000000001;
assign LUT_2[13839] = 32'b11111111111111111110111000011010;
assign LUT_2[13840] = 32'b11111111111111111110011100001010;
assign LUT_2[13841] = 32'b11111111111111111011010100100011;
assign LUT_2[13842] = 32'b00000000000000000101010101000110;
assign LUT_2[13843] = 32'b00000000000000000010001101011111;
assign LUT_2[13844] = 32'b11111111111111111010111001110010;
assign LUT_2[13845] = 32'b11111111111111110111110010001011;
assign LUT_2[13846] = 32'b00000000000000000001110010101110;
assign LUT_2[13847] = 32'b11111111111111111110101011000111;
assign LUT_2[13848] = 32'b11111111111111111001001101100111;
assign LUT_2[13849] = 32'b11111111111111110110000110000000;
assign LUT_2[13850] = 32'b00000000000000000000000110100011;
assign LUT_2[13851] = 32'b11111111111111111100111110111100;
assign LUT_2[13852] = 32'b11111111111111110101101011001111;
assign LUT_2[13853] = 32'b11111111111111110010100011101000;
assign LUT_2[13854] = 32'b11111111111111111100100100001011;
assign LUT_2[13855] = 32'b11111111111111111001011100100100;
assign LUT_2[13856] = 32'b00000000000000000100010011101001;
assign LUT_2[13857] = 32'b00000000000000000001001100000010;
assign LUT_2[13858] = 32'b00000000000000001011001100100101;
assign LUT_2[13859] = 32'b00000000000000001000000100111110;
assign LUT_2[13860] = 32'b00000000000000000000110001010001;
assign LUT_2[13861] = 32'b11111111111111111101101001101010;
assign LUT_2[13862] = 32'b00000000000000000111101010001101;
assign LUT_2[13863] = 32'b00000000000000000100100010100110;
assign LUT_2[13864] = 32'b11111111111111111111000101000110;
assign LUT_2[13865] = 32'b11111111111111111011111101011111;
assign LUT_2[13866] = 32'b00000000000000000101111110000010;
assign LUT_2[13867] = 32'b00000000000000000010110110011011;
assign LUT_2[13868] = 32'b11111111111111111011100010101110;
assign LUT_2[13869] = 32'b11111111111111111000011011000111;
assign LUT_2[13870] = 32'b00000000000000000010011011101010;
assign LUT_2[13871] = 32'b11111111111111111111010100000011;
assign LUT_2[13872] = 32'b11111111111111111110110111110011;
assign LUT_2[13873] = 32'b11111111111111111011110000001100;
assign LUT_2[13874] = 32'b00000000000000000101110000101111;
assign LUT_2[13875] = 32'b00000000000000000010101001001000;
assign LUT_2[13876] = 32'b11111111111111111011010101011011;
assign LUT_2[13877] = 32'b11111111111111111000001101110100;
assign LUT_2[13878] = 32'b00000000000000000010001110010111;
assign LUT_2[13879] = 32'b11111111111111111111000110110000;
assign LUT_2[13880] = 32'b11111111111111111001101001010000;
assign LUT_2[13881] = 32'b11111111111111110110100001101001;
assign LUT_2[13882] = 32'b00000000000000000000100010001100;
assign LUT_2[13883] = 32'b11111111111111111101011010100101;
assign LUT_2[13884] = 32'b11111111111111110110000110111000;
assign LUT_2[13885] = 32'b11111111111111110010111111010001;
assign LUT_2[13886] = 32'b11111111111111111100111111110100;
assign LUT_2[13887] = 32'b11111111111111111001111000001101;
assign LUT_2[13888] = 32'b11111111111111111100000000100011;
assign LUT_2[13889] = 32'b11111111111111111000111000111100;
assign LUT_2[13890] = 32'b00000000000000000010111001011111;
assign LUT_2[13891] = 32'b11111111111111111111110001111000;
assign LUT_2[13892] = 32'b11111111111111111000011110001011;
assign LUT_2[13893] = 32'b11111111111111110101010110100100;
assign LUT_2[13894] = 32'b11111111111111111111010111000111;
assign LUT_2[13895] = 32'b11111111111111111100001111100000;
assign LUT_2[13896] = 32'b11111111111111110110110010000000;
assign LUT_2[13897] = 32'b11111111111111110011101010011001;
assign LUT_2[13898] = 32'b11111111111111111101101010111100;
assign LUT_2[13899] = 32'b11111111111111111010100011010101;
assign LUT_2[13900] = 32'b11111111111111110011001111101000;
assign LUT_2[13901] = 32'b11111111111111110000001000000001;
assign LUT_2[13902] = 32'b11111111111111111010001000100100;
assign LUT_2[13903] = 32'b11111111111111110111000000111101;
assign LUT_2[13904] = 32'b11111111111111110110100100101101;
assign LUT_2[13905] = 32'b11111111111111110011011101000110;
assign LUT_2[13906] = 32'b11111111111111111101011101101001;
assign LUT_2[13907] = 32'b11111111111111111010010110000010;
assign LUT_2[13908] = 32'b11111111111111110011000010010101;
assign LUT_2[13909] = 32'b11111111111111101111111010101110;
assign LUT_2[13910] = 32'b11111111111111111001111011010001;
assign LUT_2[13911] = 32'b11111111111111110110110011101010;
assign LUT_2[13912] = 32'b11111111111111110001010110001010;
assign LUT_2[13913] = 32'b11111111111111101110001110100011;
assign LUT_2[13914] = 32'b11111111111111111000001111000110;
assign LUT_2[13915] = 32'b11111111111111110101000111011111;
assign LUT_2[13916] = 32'b11111111111111101101110011110010;
assign LUT_2[13917] = 32'b11111111111111101010101100001011;
assign LUT_2[13918] = 32'b11111111111111110100101100101110;
assign LUT_2[13919] = 32'b11111111111111110001100101000111;
assign LUT_2[13920] = 32'b11111111111111111100011100001100;
assign LUT_2[13921] = 32'b11111111111111111001010100100101;
assign LUT_2[13922] = 32'b00000000000000000011010101001000;
assign LUT_2[13923] = 32'b00000000000000000000001101100001;
assign LUT_2[13924] = 32'b11111111111111111000111001110100;
assign LUT_2[13925] = 32'b11111111111111110101110010001101;
assign LUT_2[13926] = 32'b11111111111111111111110010110000;
assign LUT_2[13927] = 32'b11111111111111111100101011001001;
assign LUT_2[13928] = 32'b11111111111111110111001101101001;
assign LUT_2[13929] = 32'b11111111111111110100000110000010;
assign LUT_2[13930] = 32'b11111111111111111110000110100101;
assign LUT_2[13931] = 32'b11111111111111111010111110111110;
assign LUT_2[13932] = 32'b11111111111111110011101011010001;
assign LUT_2[13933] = 32'b11111111111111110000100011101010;
assign LUT_2[13934] = 32'b11111111111111111010100100001101;
assign LUT_2[13935] = 32'b11111111111111110111011100100110;
assign LUT_2[13936] = 32'b11111111111111110111000000010110;
assign LUT_2[13937] = 32'b11111111111111110011111000101111;
assign LUT_2[13938] = 32'b11111111111111111101111001010010;
assign LUT_2[13939] = 32'b11111111111111111010110001101011;
assign LUT_2[13940] = 32'b11111111111111110011011101111110;
assign LUT_2[13941] = 32'b11111111111111110000010110010111;
assign LUT_2[13942] = 32'b11111111111111111010010110111010;
assign LUT_2[13943] = 32'b11111111111111110111001111010011;
assign LUT_2[13944] = 32'b11111111111111110001110001110011;
assign LUT_2[13945] = 32'b11111111111111101110101010001100;
assign LUT_2[13946] = 32'b11111111111111111000101010101111;
assign LUT_2[13947] = 32'b11111111111111110101100011001000;
assign LUT_2[13948] = 32'b11111111111111101110001111011011;
assign LUT_2[13949] = 32'b11111111111111101011000111110100;
assign LUT_2[13950] = 32'b11111111111111110101001000010111;
assign LUT_2[13951] = 32'b11111111111111110010000000110000;
assign LUT_2[13952] = 32'b00000000000000001000001100001111;
assign LUT_2[13953] = 32'b00000000000000000101000100101000;
assign LUT_2[13954] = 32'b00000000000000001111000101001011;
assign LUT_2[13955] = 32'b00000000000000001011111101100100;
assign LUT_2[13956] = 32'b00000000000000000100101001110111;
assign LUT_2[13957] = 32'b00000000000000000001100010010000;
assign LUT_2[13958] = 32'b00000000000000001011100010110011;
assign LUT_2[13959] = 32'b00000000000000001000011011001100;
assign LUT_2[13960] = 32'b00000000000000000010111101101100;
assign LUT_2[13961] = 32'b11111111111111111111110110000101;
assign LUT_2[13962] = 32'b00000000000000001001110110101000;
assign LUT_2[13963] = 32'b00000000000000000110101111000001;
assign LUT_2[13964] = 32'b11111111111111111111011011010100;
assign LUT_2[13965] = 32'b11111111111111111100010011101101;
assign LUT_2[13966] = 32'b00000000000000000110010100010000;
assign LUT_2[13967] = 32'b00000000000000000011001100101001;
assign LUT_2[13968] = 32'b00000000000000000010110000011001;
assign LUT_2[13969] = 32'b11111111111111111111101000110010;
assign LUT_2[13970] = 32'b00000000000000001001101001010101;
assign LUT_2[13971] = 32'b00000000000000000110100001101110;
assign LUT_2[13972] = 32'b11111111111111111111001110000001;
assign LUT_2[13973] = 32'b11111111111111111100000110011010;
assign LUT_2[13974] = 32'b00000000000000000110000110111101;
assign LUT_2[13975] = 32'b00000000000000000010111111010110;
assign LUT_2[13976] = 32'b11111111111111111101100001110110;
assign LUT_2[13977] = 32'b11111111111111111010011010001111;
assign LUT_2[13978] = 32'b00000000000000000100011010110010;
assign LUT_2[13979] = 32'b00000000000000000001010011001011;
assign LUT_2[13980] = 32'b11111111111111111001111111011110;
assign LUT_2[13981] = 32'b11111111111111110110110111110111;
assign LUT_2[13982] = 32'b00000000000000000000111000011010;
assign LUT_2[13983] = 32'b11111111111111111101110000110011;
assign LUT_2[13984] = 32'b00000000000000001000100111111000;
assign LUT_2[13985] = 32'b00000000000000000101100000010001;
assign LUT_2[13986] = 32'b00000000000000001111100000110100;
assign LUT_2[13987] = 32'b00000000000000001100011001001101;
assign LUT_2[13988] = 32'b00000000000000000101000101100000;
assign LUT_2[13989] = 32'b00000000000000000001111101111001;
assign LUT_2[13990] = 32'b00000000000000001011111110011100;
assign LUT_2[13991] = 32'b00000000000000001000110110110101;
assign LUT_2[13992] = 32'b00000000000000000011011001010101;
assign LUT_2[13993] = 32'b00000000000000000000010001101110;
assign LUT_2[13994] = 32'b00000000000000001010010010010001;
assign LUT_2[13995] = 32'b00000000000000000111001010101010;
assign LUT_2[13996] = 32'b11111111111111111111110110111101;
assign LUT_2[13997] = 32'b11111111111111111100101111010110;
assign LUT_2[13998] = 32'b00000000000000000110101111111001;
assign LUT_2[13999] = 32'b00000000000000000011101000010010;
assign LUT_2[14000] = 32'b00000000000000000011001100000010;
assign LUT_2[14001] = 32'b00000000000000000000000100011011;
assign LUT_2[14002] = 32'b00000000000000001010000100111110;
assign LUT_2[14003] = 32'b00000000000000000110111101010111;
assign LUT_2[14004] = 32'b11111111111111111111101001101010;
assign LUT_2[14005] = 32'b11111111111111111100100010000011;
assign LUT_2[14006] = 32'b00000000000000000110100010100110;
assign LUT_2[14007] = 32'b00000000000000000011011010111111;
assign LUT_2[14008] = 32'b11111111111111111101111101011111;
assign LUT_2[14009] = 32'b11111111111111111010110101111000;
assign LUT_2[14010] = 32'b00000000000000000100110110011011;
assign LUT_2[14011] = 32'b00000000000000000001101110110100;
assign LUT_2[14012] = 32'b11111111111111111010011011000111;
assign LUT_2[14013] = 32'b11111111111111110111010011100000;
assign LUT_2[14014] = 32'b00000000000000000001010100000011;
assign LUT_2[14015] = 32'b11111111111111111110001100011100;
assign LUT_2[14016] = 32'b00000000000000000000010100110010;
assign LUT_2[14017] = 32'b11111111111111111101001101001011;
assign LUT_2[14018] = 32'b00000000000000000111001101101110;
assign LUT_2[14019] = 32'b00000000000000000100000110000111;
assign LUT_2[14020] = 32'b11111111111111111100110010011010;
assign LUT_2[14021] = 32'b11111111111111111001101010110011;
assign LUT_2[14022] = 32'b00000000000000000011101011010110;
assign LUT_2[14023] = 32'b00000000000000000000100011101111;
assign LUT_2[14024] = 32'b11111111111111111011000110001111;
assign LUT_2[14025] = 32'b11111111111111110111111110101000;
assign LUT_2[14026] = 32'b00000000000000000001111111001011;
assign LUT_2[14027] = 32'b11111111111111111110110111100100;
assign LUT_2[14028] = 32'b11111111111111110111100011110111;
assign LUT_2[14029] = 32'b11111111111111110100011100010000;
assign LUT_2[14030] = 32'b11111111111111111110011100110011;
assign LUT_2[14031] = 32'b11111111111111111011010101001100;
assign LUT_2[14032] = 32'b11111111111111111010111000111100;
assign LUT_2[14033] = 32'b11111111111111110111110001010101;
assign LUT_2[14034] = 32'b00000000000000000001110001111000;
assign LUT_2[14035] = 32'b11111111111111111110101010010001;
assign LUT_2[14036] = 32'b11111111111111110111010110100100;
assign LUT_2[14037] = 32'b11111111111111110100001110111101;
assign LUT_2[14038] = 32'b11111111111111111110001111100000;
assign LUT_2[14039] = 32'b11111111111111111011000111111001;
assign LUT_2[14040] = 32'b11111111111111110101101010011001;
assign LUT_2[14041] = 32'b11111111111111110010100010110010;
assign LUT_2[14042] = 32'b11111111111111111100100011010101;
assign LUT_2[14043] = 32'b11111111111111111001011011101110;
assign LUT_2[14044] = 32'b11111111111111110010001000000001;
assign LUT_2[14045] = 32'b11111111111111101111000000011010;
assign LUT_2[14046] = 32'b11111111111111111001000000111101;
assign LUT_2[14047] = 32'b11111111111111110101111001010110;
assign LUT_2[14048] = 32'b00000000000000000000110000011011;
assign LUT_2[14049] = 32'b11111111111111111101101000110100;
assign LUT_2[14050] = 32'b00000000000000000111101001010111;
assign LUT_2[14051] = 32'b00000000000000000100100001110000;
assign LUT_2[14052] = 32'b11111111111111111101001110000011;
assign LUT_2[14053] = 32'b11111111111111111010000110011100;
assign LUT_2[14054] = 32'b00000000000000000100000110111111;
assign LUT_2[14055] = 32'b00000000000000000000111111011000;
assign LUT_2[14056] = 32'b11111111111111111011100001111000;
assign LUT_2[14057] = 32'b11111111111111111000011010010001;
assign LUT_2[14058] = 32'b00000000000000000010011010110100;
assign LUT_2[14059] = 32'b11111111111111111111010011001101;
assign LUT_2[14060] = 32'b11111111111111110111111111100000;
assign LUT_2[14061] = 32'b11111111111111110100110111111001;
assign LUT_2[14062] = 32'b11111111111111111110111000011100;
assign LUT_2[14063] = 32'b11111111111111111011110000110101;
assign LUT_2[14064] = 32'b11111111111111111011010100100101;
assign LUT_2[14065] = 32'b11111111111111111000001100111110;
assign LUT_2[14066] = 32'b00000000000000000010001101100001;
assign LUT_2[14067] = 32'b11111111111111111111000101111010;
assign LUT_2[14068] = 32'b11111111111111110111110010001101;
assign LUT_2[14069] = 32'b11111111111111110100101010100110;
assign LUT_2[14070] = 32'b11111111111111111110101011001001;
assign LUT_2[14071] = 32'b11111111111111111011100011100010;
assign LUT_2[14072] = 32'b11111111111111110110000110000010;
assign LUT_2[14073] = 32'b11111111111111110010111110011011;
assign LUT_2[14074] = 32'b11111111111111111100111110111110;
assign LUT_2[14075] = 32'b11111111111111111001110111010111;
assign LUT_2[14076] = 32'b11111111111111110010100011101010;
assign LUT_2[14077] = 32'b11111111111111101111011100000011;
assign LUT_2[14078] = 32'b11111111111111111001011100100110;
assign LUT_2[14079] = 32'b11111111111111110110010100111111;
assign LUT_2[14080] = 32'b00000000000000000111110110100110;
assign LUT_2[14081] = 32'b00000000000000000100101110111111;
assign LUT_2[14082] = 32'b00000000000000001110101111100010;
assign LUT_2[14083] = 32'b00000000000000001011100111111011;
assign LUT_2[14084] = 32'b00000000000000000100010100001110;
assign LUT_2[14085] = 32'b00000000000000000001001100100111;
assign LUT_2[14086] = 32'b00000000000000001011001101001010;
assign LUT_2[14087] = 32'b00000000000000001000000101100011;
assign LUT_2[14088] = 32'b00000000000000000010101000000011;
assign LUT_2[14089] = 32'b11111111111111111111100000011100;
assign LUT_2[14090] = 32'b00000000000000001001100000111111;
assign LUT_2[14091] = 32'b00000000000000000110011001011000;
assign LUT_2[14092] = 32'b11111111111111111111000101101011;
assign LUT_2[14093] = 32'b11111111111111111011111110000100;
assign LUT_2[14094] = 32'b00000000000000000101111110100111;
assign LUT_2[14095] = 32'b00000000000000000010110111000000;
assign LUT_2[14096] = 32'b00000000000000000010011010110000;
assign LUT_2[14097] = 32'b11111111111111111111010011001001;
assign LUT_2[14098] = 32'b00000000000000001001010011101100;
assign LUT_2[14099] = 32'b00000000000000000110001100000101;
assign LUT_2[14100] = 32'b11111111111111111110111000011000;
assign LUT_2[14101] = 32'b11111111111111111011110000110001;
assign LUT_2[14102] = 32'b00000000000000000101110001010100;
assign LUT_2[14103] = 32'b00000000000000000010101001101101;
assign LUT_2[14104] = 32'b11111111111111111101001100001101;
assign LUT_2[14105] = 32'b11111111111111111010000100100110;
assign LUT_2[14106] = 32'b00000000000000000100000101001001;
assign LUT_2[14107] = 32'b00000000000000000000111101100010;
assign LUT_2[14108] = 32'b11111111111111111001101001110101;
assign LUT_2[14109] = 32'b11111111111111110110100010001110;
assign LUT_2[14110] = 32'b00000000000000000000100010110001;
assign LUT_2[14111] = 32'b11111111111111111101011011001010;
assign LUT_2[14112] = 32'b00000000000000001000010010001111;
assign LUT_2[14113] = 32'b00000000000000000101001010101000;
assign LUT_2[14114] = 32'b00000000000000001111001011001011;
assign LUT_2[14115] = 32'b00000000000000001100000011100100;
assign LUT_2[14116] = 32'b00000000000000000100101111110111;
assign LUT_2[14117] = 32'b00000000000000000001101000010000;
assign LUT_2[14118] = 32'b00000000000000001011101000110011;
assign LUT_2[14119] = 32'b00000000000000001000100001001100;
assign LUT_2[14120] = 32'b00000000000000000011000011101100;
assign LUT_2[14121] = 32'b11111111111111111111111100000101;
assign LUT_2[14122] = 32'b00000000000000001001111100101000;
assign LUT_2[14123] = 32'b00000000000000000110110101000001;
assign LUT_2[14124] = 32'b11111111111111111111100001010100;
assign LUT_2[14125] = 32'b11111111111111111100011001101101;
assign LUT_2[14126] = 32'b00000000000000000110011010010000;
assign LUT_2[14127] = 32'b00000000000000000011010010101001;
assign LUT_2[14128] = 32'b00000000000000000010110110011001;
assign LUT_2[14129] = 32'b11111111111111111111101110110010;
assign LUT_2[14130] = 32'b00000000000000001001101111010101;
assign LUT_2[14131] = 32'b00000000000000000110100111101110;
assign LUT_2[14132] = 32'b11111111111111111111010100000001;
assign LUT_2[14133] = 32'b11111111111111111100001100011010;
assign LUT_2[14134] = 32'b00000000000000000110001100111101;
assign LUT_2[14135] = 32'b00000000000000000011000101010110;
assign LUT_2[14136] = 32'b11111111111111111101100111110110;
assign LUT_2[14137] = 32'b11111111111111111010100000001111;
assign LUT_2[14138] = 32'b00000000000000000100100000110010;
assign LUT_2[14139] = 32'b00000000000000000001011001001011;
assign LUT_2[14140] = 32'b11111111111111111010000101011110;
assign LUT_2[14141] = 32'b11111111111111110110111101110111;
assign LUT_2[14142] = 32'b00000000000000000000111110011010;
assign LUT_2[14143] = 32'b11111111111111111101110110110011;
assign LUT_2[14144] = 32'b11111111111111111111111111001001;
assign LUT_2[14145] = 32'b11111111111111111100110111100010;
assign LUT_2[14146] = 32'b00000000000000000110111000000101;
assign LUT_2[14147] = 32'b00000000000000000011110000011110;
assign LUT_2[14148] = 32'b11111111111111111100011100110001;
assign LUT_2[14149] = 32'b11111111111111111001010101001010;
assign LUT_2[14150] = 32'b00000000000000000011010101101101;
assign LUT_2[14151] = 32'b00000000000000000000001110000110;
assign LUT_2[14152] = 32'b11111111111111111010110000100110;
assign LUT_2[14153] = 32'b11111111111111110111101000111111;
assign LUT_2[14154] = 32'b00000000000000000001101001100010;
assign LUT_2[14155] = 32'b11111111111111111110100001111011;
assign LUT_2[14156] = 32'b11111111111111110111001110001110;
assign LUT_2[14157] = 32'b11111111111111110100000110100111;
assign LUT_2[14158] = 32'b11111111111111111110000111001010;
assign LUT_2[14159] = 32'b11111111111111111010111111100011;
assign LUT_2[14160] = 32'b11111111111111111010100011010011;
assign LUT_2[14161] = 32'b11111111111111110111011011101100;
assign LUT_2[14162] = 32'b00000000000000000001011100001111;
assign LUT_2[14163] = 32'b11111111111111111110010100101000;
assign LUT_2[14164] = 32'b11111111111111110111000000111011;
assign LUT_2[14165] = 32'b11111111111111110011111001010100;
assign LUT_2[14166] = 32'b11111111111111111101111001110111;
assign LUT_2[14167] = 32'b11111111111111111010110010010000;
assign LUT_2[14168] = 32'b11111111111111110101010100110000;
assign LUT_2[14169] = 32'b11111111111111110010001101001001;
assign LUT_2[14170] = 32'b11111111111111111100001101101100;
assign LUT_2[14171] = 32'b11111111111111111001000110000101;
assign LUT_2[14172] = 32'b11111111111111110001110010011000;
assign LUT_2[14173] = 32'b11111111111111101110101010110001;
assign LUT_2[14174] = 32'b11111111111111111000101011010100;
assign LUT_2[14175] = 32'b11111111111111110101100011101101;
assign LUT_2[14176] = 32'b00000000000000000000011010110010;
assign LUT_2[14177] = 32'b11111111111111111101010011001011;
assign LUT_2[14178] = 32'b00000000000000000111010011101110;
assign LUT_2[14179] = 32'b00000000000000000100001100000111;
assign LUT_2[14180] = 32'b11111111111111111100111000011010;
assign LUT_2[14181] = 32'b11111111111111111001110000110011;
assign LUT_2[14182] = 32'b00000000000000000011110001010110;
assign LUT_2[14183] = 32'b00000000000000000000101001101111;
assign LUT_2[14184] = 32'b11111111111111111011001100001111;
assign LUT_2[14185] = 32'b11111111111111111000000100101000;
assign LUT_2[14186] = 32'b00000000000000000010000101001011;
assign LUT_2[14187] = 32'b11111111111111111110111101100100;
assign LUT_2[14188] = 32'b11111111111111110111101001110111;
assign LUT_2[14189] = 32'b11111111111111110100100010010000;
assign LUT_2[14190] = 32'b11111111111111111110100010110011;
assign LUT_2[14191] = 32'b11111111111111111011011011001100;
assign LUT_2[14192] = 32'b11111111111111111010111110111100;
assign LUT_2[14193] = 32'b11111111111111110111110111010101;
assign LUT_2[14194] = 32'b00000000000000000001110111111000;
assign LUT_2[14195] = 32'b11111111111111111110110000010001;
assign LUT_2[14196] = 32'b11111111111111110111011100100100;
assign LUT_2[14197] = 32'b11111111111111110100010100111101;
assign LUT_2[14198] = 32'b11111111111111111110010101100000;
assign LUT_2[14199] = 32'b11111111111111111011001101111001;
assign LUT_2[14200] = 32'b11111111111111110101110000011001;
assign LUT_2[14201] = 32'b11111111111111110010101000110010;
assign LUT_2[14202] = 32'b11111111111111111100101001010101;
assign LUT_2[14203] = 32'b11111111111111111001100001101110;
assign LUT_2[14204] = 32'b11111111111111110010001110000001;
assign LUT_2[14205] = 32'b11111111111111101111000110011010;
assign LUT_2[14206] = 32'b11111111111111111001000110111101;
assign LUT_2[14207] = 32'b11111111111111110101111111010110;
assign LUT_2[14208] = 32'b00000000000000001100001010110101;
assign LUT_2[14209] = 32'b00000000000000001001000011001110;
assign LUT_2[14210] = 32'b00000000000000010011000011110001;
assign LUT_2[14211] = 32'b00000000000000001111111100001010;
assign LUT_2[14212] = 32'b00000000000000001000101000011101;
assign LUT_2[14213] = 32'b00000000000000000101100000110110;
assign LUT_2[14214] = 32'b00000000000000001111100001011001;
assign LUT_2[14215] = 32'b00000000000000001100011001110010;
assign LUT_2[14216] = 32'b00000000000000000110111100010010;
assign LUT_2[14217] = 32'b00000000000000000011110100101011;
assign LUT_2[14218] = 32'b00000000000000001101110101001110;
assign LUT_2[14219] = 32'b00000000000000001010101101100111;
assign LUT_2[14220] = 32'b00000000000000000011011001111010;
assign LUT_2[14221] = 32'b00000000000000000000010010010011;
assign LUT_2[14222] = 32'b00000000000000001010010010110110;
assign LUT_2[14223] = 32'b00000000000000000111001011001111;
assign LUT_2[14224] = 32'b00000000000000000110101110111111;
assign LUT_2[14225] = 32'b00000000000000000011100111011000;
assign LUT_2[14226] = 32'b00000000000000001101100111111011;
assign LUT_2[14227] = 32'b00000000000000001010100000010100;
assign LUT_2[14228] = 32'b00000000000000000011001100100111;
assign LUT_2[14229] = 32'b00000000000000000000000101000000;
assign LUT_2[14230] = 32'b00000000000000001010000101100011;
assign LUT_2[14231] = 32'b00000000000000000110111101111100;
assign LUT_2[14232] = 32'b00000000000000000001100000011100;
assign LUT_2[14233] = 32'b11111111111111111110011000110101;
assign LUT_2[14234] = 32'b00000000000000001000011001011000;
assign LUT_2[14235] = 32'b00000000000000000101010001110001;
assign LUT_2[14236] = 32'b11111111111111111101111110000100;
assign LUT_2[14237] = 32'b11111111111111111010110110011101;
assign LUT_2[14238] = 32'b00000000000000000100110111000000;
assign LUT_2[14239] = 32'b00000000000000000001101111011001;
assign LUT_2[14240] = 32'b00000000000000001100100110011110;
assign LUT_2[14241] = 32'b00000000000000001001011110110111;
assign LUT_2[14242] = 32'b00000000000000010011011111011010;
assign LUT_2[14243] = 32'b00000000000000010000010111110011;
assign LUT_2[14244] = 32'b00000000000000001001000100000110;
assign LUT_2[14245] = 32'b00000000000000000101111100011111;
assign LUT_2[14246] = 32'b00000000000000001111111101000010;
assign LUT_2[14247] = 32'b00000000000000001100110101011011;
assign LUT_2[14248] = 32'b00000000000000000111010111111011;
assign LUT_2[14249] = 32'b00000000000000000100010000010100;
assign LUT_2[14250] = 32'b00000000000000001110010000110111;
assign LUT_2[14251] = 32'b00000000000000001011001001010000;
assign LUT_2[14252] = 32'b00000000000000000011110101100011;
assign LUT_2[14253] = 32'b00000000000000000000101101111100;
assign LUT_2[14254] = 32'b00000000000000001010101110011111;
assign LUT_2[14255] = 32'b00000000000000000111100110111000;
assign LUT_2[14256] = 32'b00000000000000000111001010101000;
assign LUT_2[14257] = 32'b00000000000000000100000011000001;
assign LUT_2[14258] = 32'b00000000000000001110000011100100;
assign LUT_2[14259] = 32'b00000000000000001010111011111101;
assign LUT_2[14260] = 32'b00000000000000000011101000010000;
assign LUT_2[14261] = 32'b00000000000000000000100000101001;
assign LUT_2[14262] = 32'b00000000000000001010100001001100;
assign LUT_2[14263] = 32'b00000000000000000111011001100101;
assign LUT_2[14264] = 32'b00000000000000000001111100000101;
assign LUT_2[14265] = 32'b11111111111111111110110100011110;
assign LUT_2[14266] = 32'b00000000000000001000110101000001;
assign LUT_2[14267] = 32'b00000000000000000101101101011010;
assign LUT_2[14268] = 32'b11111111111111111110011001101101;
assign LUT_2[14269] = 32'b11111111111111111011010010000110;
assign LUT_2[14270] = 32'b00000000000000000101010010101001;
assign LUT_2[14271] = 32'b00000000000000000010001011000010;
assign LUT_2[14272] = 32'b00000000000000000100010011011000;
assign LUT_2[14273] = 32'b00000000000000000001001011110001;
assign LUT_2[14274] = 32'b00000000000000001011001100010100;
assign LUT_2[14275] = 32'b00000000000000001000000100101101;
assign LUT_2[14276] = 32'b00000000000000000000110001000000;
assign LUT_2[14277] = 32'b11111111111111111101101001011001;
assign LUT_2[14278] = 32'b00000000000000000111101001111100;
assign LUT_2[14279] = 32'b00000000000000000100100010010101;
assign LUT_2[14280] = 32'b11111111111111111111000100110101;
assign LUT_2[14281] = 32'b11111111111111111011111101001110;
assign LUT_2[14282] = 32'b00000000000000000101111101110001;
assign LUT_2[14283] = 32'b00000000000000000010110110001010;
assign LUT_2[14284] = 32'b11111111111111111011100010011101;
assign LUT_2[14285] = 32'b11111111111111111000011010110110;
assign LUT_2[14286] = 32'b00000000000000000010011011011001;
assign LUT_2[14287] = 32'b11111111111111111111010011110010;
assign LUT_2[14288] = 32'b11111111111111111110110111100010;
assign LUT_2[14289] = 32'b11111111111111111011101111111011;
assign LUT_2[14290] = 32'b00000000000000000101110000011110;
assign LUT_2[14291] = 32'b00000000000000000010101000110111;
assign LUT_2[14292] = 32'b11111111111111111011010101001010;
assign LUT_2[14293] = 32'b11111111111111111000001101100011;
assign LUT_2[14294] = 32'b00000000000000000010001110000110;
assign LUT_2[14295] = 32'b11111111111111111111000110011111;
assign LUT_2[14296] = 32'b11111111111111111001101000111111;
assign LUT_2[14297] = 32'b11111111111111110110100001011000;
assign LUT_2[14298] = 32'b00000000000000000000100001111011;
assign LUT_2[14299] = 32'b11111111111111111101011010010100;
assign LUT_2[14300] = 32'b11111111111111110110000110100111;
assign LUT_2[14301] = 32'b11111111111111110010111111000000;
assign LUT_2[14302] = 32'b11111111111111111100111111100011;
assign LUT_2[14303] = 32'b11111111111111111001110111111100;
assign LUT_2[14304] = 32'b00000000000000000100101111000001;
assign LUT_2[14305] = 32'b00000000000000000001100111011010;
assign LUT_2[14306] = 32'b00000000000000001011100111111101;
assign LUT_2[14307] = 32'b00000000000000001000100000010110;
assign LUT_2[14308] = 32'b00000000000000000001001100101001;
assign LUT_2[14309] = 32'b11111111111111111110000101000010;
assign LUT_2[14310] = 32'b00000000000000001000000101100101;
assign LUT_2[14311] = 32'b00000000000000000100111101111110;
assign LUT_2[14312] = 32'b11111111111111111111100000011110;
assign LUT_2[14313] = 32'b11111111111111111100011000110111;
assign LUT_2[14314] = 32'b00000000000000000110011001011010;
assign LUT_2[14315] = 32'b00000000000000000011010001110011;
assign LUT_2[14316] = 32'b11111111111111111011111110000110;
assign LUT_2[14317] = 32'b11111111111111111000110110011111;
assign LUT_2[14318] = 32'b00000000000000000010110111000010;
assign LUT_2[14319] = 32'b11111111111111111111101111011011;
assign LUT_2[14320] = 32'b11111111111111111111010011001011;
assign LUT_2[14321] = 32'b11111111111111111100001011100100;
assign LUT_2[14322] = 32'b00000000000000000110001100000111;
assign LUT_2[14323] = 32'b00000000000000000011000100100000;
assign LUT_2[14324] = 32'b11111111111111111011110000110011;
assign LUT_2[14325] = 32'b11111111111111111000101001001100;
assign LUT_2[14326] = 32'b00000000000000000010101001101111;
assign LUT_2[14327] = 32'b11111111111111111111100010001000;
assign LUT_2[14328] = 32'b11111111111111111010000100101000;
assign LUT_2[14329] = 32'b11111111111111110110111101000001;
assign LUT_2[14330] = 32'b00000000000000000000111101100100;
assign LUT_2[14331] = 32'b11111111111111111101110101111101;
assign LUT_2[14332] = 32'b11111111111111110110100010010000;
assign LUT_2[14333] = 32'b11111111111111110011011010101001;
assign LUT_2[14334] = 32'b11111111111111111101011011001100;
assign LUT_2[14335] = 32'b11111111111111111010010011100101;
assign LUT_2[14336] = 32'b11111111111111110100010000000101;
assign LUT_2[14337] = 32'b11111111111111110001001000011110;
assign LUT_2[14338] = 32'b11111111111111111011001001000001;
assign LUT_2[14339] = 32'b11111111111111111000000001011010;
assign LUT_2[14340] = 32'b11111111111111110000101101101101;
assign LUT_2[14341] = 32'b11111111111111101101100110000110;
assign LUT_2[14342] = 32'b11111111111111110111100110101001;
assign LUT_2[14343] = 32'b11111111111111110100011111000010;
assign LUT_2[14344] = 32'b11111111111111101111000001100010;
assign LUT_2[14345] = 32'b11111111111111101011111001111011;
assign LUT_2[14346] = 32'b11111111111111110101111010011110;
assign LUT_2[14347] = 32'b11111111111111110010110010110111;
assign LUT_2[14348] = 32'b11111111111111101011011111001010;
assign LUT_2[14349] = 32'b11111111111111101000010111100011;
assign LUT_2[14350] = 32'b11111111111111110010011000000110;
assign LUT_2[14351] = 32'b11111111111111101111010000011111;
assign LUT_2[14352] = 32'b11111111111111101110110100001111;
assign LUT_2[14353] = 32'b11111111111111101011101100101000;
assign LUT_2[14354] = 32'b11111111111111110101101101001011;
assign LUT_2[14355] = 32'b11111111111111110010100101100100;
assign LUT_2[14356] = 32'b11111111111111101011010001110111;
assign LUT_2[14357] = 32'b11111111111111101000001010010000;
assign LUT_2[14358] = 32'b11111111111111110010001010110011;
assign LUT_2[14359] = 32'b11111111111111101111000011001100;
assign LUT_2[14360] = 32'b11111111111111101001100101101100;
assign LUT_2[14361] = 32'b11111111111111100110011110000101;
assign LUT_2[14362] = 32'b11111111111111110000011110101000;
assign LUT_2[14363] = 32'b11111111111111101101010111000001;
assign LUT_2[14364] = 32'b11111111111111100110000011010100;
assign LUT_2[14365] = 32'b11111111111111100010111011101101;
assign LUT_2[14366] = 32'b11111111111111101100111100010000;
assign LUT_2[14367] = 32'b11111111111111101001110100101001;
assign LUT_2[14368] = 32'b11111111111111110100101011101110;
assign LUT_2[14369] = 32'b11111111111111110001100100000111;
assign LUT_2[14370] = 32'b11111111111111111011100100101010;
assign LUT_2[14371] = 32'b11111111111111111000011101000011;
assign LUT_2[14372] = 32'b11111111111111110001001001010110;
assign LUT_2[14373] = 32'b11111111111111101110000001101111;
assign LUT_2[14374] = 32'b11111111111111111000000010010010;
assign LUT_2[14375] = 32'b11111111111111110100111010101011;
assign LUT_2[14376] = 32'b11111111111111101111011101001011;
assign LUT_2[14377] = 32'b11111111111111101100010101100100;
assign LUT_2[14378] = 32'b11111111111111110110010110000111;
assign LUT_2[14379] = 32'b11111111111111110011001110100000;
assign LUT_2[14380] = 32'b11111111111111101011111010110011;
assign LUT_2[14381] = 32'b11111111111111101000110011001100;
assign LUT_2[14382] = 32'b11111111111111110010110011101111;
assign LUT_2[14383] = 32'b11111111111111101111101100001000;
assign LUT_2[14384] = 32'b11111111111111101111001111111000;
assign LUT_2[14385] = 32'b11111111111111101100001000010001;
assign LUT_2[14386] = 32'b11111111111111110110001000110100;
assign LUT_2[14387] = 32'b11111111111111110011000001001101;
assign LUT_2[14388] = 32'b11111111111111101011101101100000;
assign LUT_2[14389] = 32'b11111111111111101000100101111001;
assign LUT_2[14390] = 32'b11111111111111110010100110011100;
assign LUT_2[14391] = 32'b11111111111111101111011110110101;
assign LUT_2[14392] = 32'b11111111111111101010000001010101;
assign LUT_2[14393] = 32'b11111111111111100110111001101110;
assign LUT_2[14394] = 32'b11111111111111110000111010010001;
assign LUT_2[14395] = 32'b11111111111111101101110010101010;
assign LUT_2[14396] = 32'b11111111111111100110011110111101;
assign LUT_2[14397] = 32'b11111111111111100011010111010110;
assign LUT_2[14398] = 32'b11111111111111101101010111111001;
assign LUT_2[14399] = 32'b11111111111111101010010000010010;
assign LUT_2[14400] = 32'b11111111111111101100011000101000;
assign LUT_2[14401] = 32'b11111111111111101001010001000001;
assign LUT_2[14402] = 32'b11111111111111110011010001100100;
assign LUT_2[14403] = 32'b11111111111111110000001001111101;
assign LUT_2[14404] = 32'b11111111111111101000110110010000;
assign LUT_2[14405] = 32'b11111111111111100101101110101001;
assign LUT_2[14406] = 32'b11111111111111101111101111001100;
assign LUT_2[14407] = 32'b11111111111111101100100111100101;
assign LUT_2[14408] = 32'b11111111111111100111001010000101;
assign LUT_2[14409] = 32'b11111111111111100100000010011110;
assign LUT_2[14410] = 32'b11111111111111101110000011000001;
assign LUT_2[14411] = 32'b11111111111111101010111011011010;
assign LUT_2[14412] = 32'b11111111111111100011100111101101;
assign LUT_2[14413] = 32'b11111111111111100000100000000110;
assign LUT_2[14414] = 32'b11111111111111101010100000101001;
assign LUT_2[14415] = 32'b11111111111111100111011001000010;
assign LUT_2[14416] = 32'b11111111111111100110111100110010;
assign LUT_2[14417] = 32'b11111111111111100011110101001011;
assign LUT_2[14418] = 32'b11111111111111101101110101101110;
assign LUT_2[14419] = 32'b11111111111111101010101110000111;
assign LUT_2[14420] = 32'b11111111111111100011011010011010;
assign LUT_2[14421] = 32'b11111111111111100000010010110011;
assign LUT_2[14422] = 32'b11111111111111101010010011010110;
assign LUT_2[14423] = 32'b11111111111111100111001011101111;
assign LUT_2[14424] = 32'b11111111111111100001101110001111;
assign LUT_2[14425] = 32'b11111111111111011110100110101000;
assign LUT_2[14426] = 32'b11111111111111101000100111001011;
assign LUT_2[14427] = 32'b11111111111111100101011111100100;
assign LUT_2[14428] = 32'b11111111111111011110001011110111;
assign LUT_2[14429] = 32'b11111111111111011011000100010000;
assign LUT_2[14430] = 32'b11111111111111100101000100110011;
assign LUT_2[14431] = 32'b11111111111111100001111101001100;
assign LUT_2[14432] = 32'b11111111111111101100110100010001;
assign LUT_2[14433] = 32'b11111111111111101001101100101010;
assign LUT_2[14434] = 32'b11111111111111110011101101001101;
assign LUT_2[14435] = 32'b11111111111111110000100101100110;
assign LUT_2[14436] = 32'b11111111111111101001010001111001;
assign LUT_2[14437] = 32'b11111111111111100110001010010010;
assign LUT_2[14438] = 32'b11111111111111110000001010110101;
assign LUT_2[14439] = 32'b11111111111111101101000011001110;
assign LUT_2[14440] = 32'b11111111111111100111100101101110;
assign LUT_2[14441] = 32'b11111111111111100100011110000111;
assign LUT_2[14442] = 32'b11111111111111101110011110101010;
assign LUT_2[14443] = 32'b11111111111111101011010111000011;
assign LUT_2[14444] = 32'b11111111111111100100000011010110;
assign LUT_2[14445] = 32'b11111111111111100000111011101111;
assign LUT_2[14446] = 32'b11111111111111101010111100010010;
assign LUT_2[14447] = 32'b11111111111111100111110100101011;
assign LUT_2[14448] = 32'b11111111111111100111011000011011;
assign LUT_2[14449] = 32'b11111111111111100100010000110100;
assign LUT_2[14450] = 32'b11111111111111101110010001010111;
assign LUT_2[14451] = 32'b11111111111111101011001001110000;
assign LUT_2[14452] = 32'b11111111111111100011110110000011;
assign LUT_2[14453] = 32'b11111111111111100000101110011100;
assign LUT_2[14454] = 32'b11111111111111101010101110111111;
assign LUT_2[14455] = 32'b11111111111111100111100111011000;
assign LUT_2[14456] = 32'b11111111111111100010001001111000;
assign LUT_2[14457] = 32'b11111111111111011111000010010001;
assign LUT_2[14458] = 32'b11111111111111101001000010110100;
assign LUT_2[14459] = 32'b11111111111111100101111011001101;
assign LUT_2[14460] = 32'b11111111111111011110100111100000;
assign LUT_2[14461] = 32'b11111111111111011011011111111001;
assign LUT_2[14462] = 32'b11111111111111100101100000011100;
assign LUT_2[14463] = 32'b11111111111111100010011000110101;
assign LUT_2[14464] = 32'b11111111111111111000100100010100;
assign LUT_2[14465] = 32'b11111111111111110101011100101101;
assign LUT_2[14466] = 32'b11111111111111111111011101010000;
assign LUT_2[14467] = 32'b11111111111111111100010101101001;
assign LUT_2[14468] = 32'b11111111111111110101000001111100;
assign LUT_2[14469] = 32'b11111111111111110001111010010101;
assign LUT_2[14470] = 32'b11111111111111111011111010111000;
assign LUT_2[14471] = 32'b11111111111111111000110011010001;
assign LUT_2[14472] = 32'b11111111111111110011010101110001;
assign LUT_2[14473] = 32'b11111111111111110000001110001010;
assign LUT_2[14474] = 32'b11111111111111111010001110101101;
assign LUT_2[14475] = 32'b11111111111111110111000111000110;
assign LUT_2[14476] = 32'b11111111111111101111110011011001;
assign LUT_2[14477] = 32'b11111111111111101100101011110010;
assign LUT_2[14478] = 32'b11111111111111110110101100010101;
assign LUT_2[14479] = 32'b11111111111111110011100100101110;
assign LUT_2[14480] = 32'b11111111111111110011001000011110;
assign LUT_2[14481] = 32'b11111111111111110000000000110111;
assign LUT_2[14482] = 32'b11111111111111111010000001011010;
assign LUT_2[14483] = 32'b11111111111111110110111001110011;
assign LUT_2[14484] = 32'b11111111111111101111100110000110;
assign LUT_2[14485] = 32'b11111111111111101100011110011111;
assign LUT_2[14486] = 32'b11111111111111110110011111000010;
assign LUT_2[14487] = 32'b11111111111111110011010111011011;
assign LUT_2[14488] = 32'b11111111111111101101111001111011;
assign LUT_2[14489] = 32'b11111111111111101010110010010100;
assign LUT_2[14490] = 32'b11111111111111110100110010110111;
assign LUT_2[14491] = 32'b11111111111111110001101011010000;
assign LUT_2[14492] = 32'b11111111111111101010010111100011;
assign LUT_2[14493] = 32'b11111111111111100111001111111100;
assign LUT_2[14494] = 32'b11111111111111110001010000011111;
assign LUT_2[14495] = 32'b11111111111111101110001000111000;
assign LUT_2[14496] = 32'b11111111111111111000111111111101;
assign LUT_2[14497] = 32'b11111111111111110101111000010110;
assign LUT_2[14498] = 32'b11111111111111111111111000111001;
assign LUT_2[14499] = 32'b11111111111111111100110001010010;
assign LUT_2[14500] = 32'b11111111111111110101011101100101;
assign LUT_2[14501] = 32'b11111111111111110010010101111110;
assign LUT_2[14502] = 32'b11111111111111111100010110100001;
assign LUT_2[14503] = 32'b11111111111111111001001110111010;
assign LUT_2[14504] = 32'b11111111111111110011110001011010;
assign LUT_2[14505] = 32'b11111111111111110000101001110011;
assign LUT_2[14506] = 32'b11111111111111111010101010010110;
assign LUT_2[14507] = 32'b11111111111111110111100010101111;
assign LUT_2[14508] = 32'b11111111111111110000001111000010;
assign LUT_2[14509] = 32'b11111111111111101101000111011011;
assign LUT_2[14510] = 32'b11111111111111110111000111111110;
assign LUT_2[14511] = 32'b11111111111111110100000000010111;
assign LUT_2[14512] = 32'b11111111111111110011100100000111;
assign LUT_2[14513] = 32'b11111111111111110000011100100000;
assign LUT_2[14514] = 32'b11111111111111111010011101000011;
assign LUT_2[14515] = 32'b11111111111111110111010101011100;
assign LUT_2[14516] = 32'b11111111111111110000000001101111;
assign LUT_2[14517] = 32'b11111111111111101100111010001000;
assign LUT_2[14518] = 32'b11111111111111110110111010101011;
assign LUT_2[14519] = 32'b11111111111111110011110011000100;
assign LUT_2[14520] = 32'b11111111111111101110010101100100;
assign LUT_2[14521] = 32'b11111111111111101011001101111101;
assign LUT_2[14522] = 32'b11111111111111110101001110100000;
assign LUT_2[14523] = 32'b11111111111111110010000110111001;
assign LUT_2[14524] = 32'b11111111111111101010110011001100;
assign LUT_2[14525] = 32'b11111111111111100111101011100101;
assign LUT_2[14526] = 32'b11111111111111110001101100001000;
assign LUT_2[14527] = 32'b11111111111111101110100100100001;
assign LUT_2[14528] = 32'b11111111111111110000101100110111;
assign LUT_2[14529] = 32'b11111111111111101101100101010000;
assign LUT_2[14530] = 32'b11111111111111110111100101110011;
assign LUT_2[14531] = 32'b11111111111111110100011110001100;
assign LUT_2[14532] = 32'b11111111111111101101001010011111;
assign LUT_2[14533] = 32'b11111111111111101010000010111000;
assign LUT_2[14534] = 32'b11111111111111110100000011011011;
assign LUT_2[14535] = 32'b11111111111111110000111011110100;
assign LUT_2[14536] = 32'b11111111111111101011011110010100;
assign LUT_2[14537] = 32'b11111111111111101000010110101101;
assign LUT_2[14538] = 32'b11111111111111110010010111010000;
assign LUT_2[14539] = 32'b11111111111111101111001111101001;
assign LUT_2[14540] = 32'b11111111111111100111111011111100;
assign LUT_2[14541] = 32'b11111111111111100100110100010101;
assign LUT_2[14542] = 32'b11111111111111101110110100111000;
assign LUT_2[14543] = 32'b11111111111111101011101101010001;
assign LUT_2[14544] = 32'b11111111111111101011010001000001;
assign LUT_2[14545] = 32'b11111111111111101000001001011010;
assign LUT_2[14546] = 32'b11111111111111110010001001111101;
assign LUT_2[14547] = 32'b11111111111111101111000010010110;
assign LUT_2[14548] = 32'b11111111111111100111101110101001;
assign LUT_2[14549] = 32'b11111111111111100100100111000010;
assign LUT_2[14550] = 32'b11111111111111101110100111100101;
assign LUT_2[14551] = 32'b11111111111111101011011111111110;
assign LUT_2[14552] = 32'b11111111111111100110000010011110;
assign LUT_2[14553] = 32'b11111111111111100010111010110111;
assign LUT_2[14554] = 32'b11111111111111101100111011011010;
assign LUT_2[14555] = 32'b11111111111111101001110011110011;
assign LUT_2[14556] = 32'b11111111111111100010100000000110;
assign LUT_2[14557] = 32'b11111111111111011111011000011111;
assign LUT_2[14558] = 32'b11111111111111101001011001000010;
assign LUT_2[14559] = 32'b11111111111111100110010001011011;
assign LUT_2[14560] = 32'b11111111111111110001001000100000;
assign LUT_2[14561] = 32'b11111111111111101110000000111001;
assign LUT_2[14562] = 32'b11111111111111111000000001011100;
assign LUT_2[14563] = 32'b11111111111111110100111001110101;
assign LUT_2[14564] = 32'b11111111111111101101100110001000;
assign LUT_2[14565] = 32'b11111111111111101010011110100001;
assign LUT_2[14566] = 32'b11111111111111110100011111000100;
assign LUT_2[14567] = 32'b11111111111111110001010111011101;
assign LUT_2[14568] = 32'b11111111111111101011111001111101;
assign LUT_2[14569] = 32'b11111111111111101000110010010110;
assign LUT_2[14570] = 32'b11111111111111110010110010111001;
assign LUT_2[14571] = 32'b11111111111111101111101011010010;
assign LUT_2[14572] = 32'b11111111111111101000010111100101;
assign LUT_2[14573] = 32'b11111111111111100101001111111110;
assign LUT_2[14574] = 32'b11111111111111101111010000100001;
assign LUT_2[14575] = 32'b11111111111111101100001000111010;
assign LUT_2[14576] = 32'b11111111111111101011101100101010;
assign LUT_2[14577] = 32'b11111111111111101000100101000011;
assign LUT_2[14578] = 32'b11111111111111110010100101100110;
assign LUT_2[14579] = 32'b11111111111111101111011101111111;
assign LUT_2[14580] = 32'b11111111111111101000001010010010;
assign LUT_2[14581] = 32'b11111111111111100101000010101011;
assign LUT_2[14582] = 32'b11111111111111101111000011001110;
assign LUT_2[14583] = 32'b11111111111111101011111011100111;
assign LUT_2[14584] = 32'b11111111111111100110011110000111;
assign LUT_2[14585] = 32'b11111111111111100011010110100000;
assign LUT_2[14586] = 32'b11111111111111101101010111000011;
assign LUT_2[14587] = 32'b11111111111111101010001111011100;
assign LUT_2[14588] = 32'b11111111111111100010111011101111;
assign LUT_2[14589] = 32'b11111111111111011111110100001000;
assign LUT_2[14590] = 32'b11111111111111101001110100101011;
assign LUT_2[14591] = 32'b11111111111111100110101101000100;
assign LUT_2[14592] = 32'b11111111111111111000001110101011;
assign LUT_2[14593] = 32'b11111111111111110101000111000100;
assign LUT_2[14594] = 32'b11111111111111111111000111100111;
assign LUT_2[14595] = 32'b11111111111111111100000000000000;
assign LUT_2[14596] = 32'b11111111111111110100101100010011;
assign LUT_2[14597] = 32'b11111111111111110001100100101100;
assign LUT_2[14598] = 32'b11111111111111111011100101001111;
assign LUT_2[14599] = 32'b11111111111111111000011101101000;
assign LUT_2[14600] = 32'b11111111111111110011000000001000;
assign LUT_2[14601] = 32'b11111111111111101111111000100001;
assign LUT_2[14602] = 32'b11111111111111111001111001000100;
assign LUT_2[14603] = 32'b11111111111111110110110001011101;
assign LUT_2[14604] = 32'b11111111111111101111011101110000;
assign LUT_2[14605] = 32'b11111111111111101100010110001001;
assign LUT_2[14606] = 32'b11111111111111110110010110101100;
assign LUT_2[14607] = 32'b11111111111111110011001111000101;
assign LUT_2[14608] = 32'b11111111111111110010110010110101;
assign LUT_2[14609] = 32'b11111111111111101111101011001110;
assign LUT_2[14610] = 32'b11111111111111111001101011110001;
assign LUT_2[14611] = 32'b11111111111111110110100100001010;
assign LUT_2[14612] = 32'b11111111111111101111010000011101;
assign LUT_2[14613] = 32'b11111111111111101100001000110110;
assign LUT_2[14614] = 32'b11111111111111110110001001011001;
assign LUT_2[14615] = 32'b11111111111111110011000001110010;
assign LUT_2[14616] = 32'b11111111111111101101100100010010;
assign LUT_2[14617] = 32'b11111111111111101010011100101011;
assign LUT_2[14618] = 32'b11111111111111110100011101001110;
assign LUT_2[14619] = 32'b11111111111111110001010101100111;
assign LUT_2[14620] = 32'b11111111111111101010000001111010;
assign LUT_2[14621] = 32'b11111111111111100110111010010011;
assign LUT_2[14622] = 32'b11111111111111110000111010110110;
assign LUT_2[14623] = 32'b11111111111111101101110011001111;
assign LUT_2[14624] = 32'b11111111111111111000101010010100;
assign LUT_2[14625] = 32'b11111111111111110101100010101101;
assign LUT_2[14626] = 32'b11111111111111111111100011010000;
assign LUT_2[14627] = 32'b11111111111111111100011011101001;
assign LUT_2[14628] = 32'b11111111111111110101000111111100;
assign LUT_2[14629] = 32'b11111111111111110010000000010101;
assign LUT_2[14630] = 32'b11111111111111111100000000111000;
assign LUT_2[14631] = 32'b11111111111111111000111001010001;
assign LUT_2[14632] = 32'b11111111111111110011011011110001;
assign LUT_2[14633] = 32'b11111111111111110000010100001010;
assign LUT_2[14634] = 32'b11111111111111111010010100101101;
assign LUT_2[14635] = 32'b11111111111111110111001101000110;
assign LUT_2[14636] = 32'b11111111111111101111111001011001;
assign LUT_2[14637] = 32'b11111111111111101100110001110010;
assign LUT_2[14638] = 32'b11111111111111110110110010010101;
assign LUT_2[14639] = 32'b11111111111111110011101010101110;
assign LUT_2[14640] = 32'b11111111111111110011001110011110;
assign LUT_2[14641] = 32'b11111111111111110000000110110111;
assign LUT_2[14642] = 32'b11111111111111111010000111011010;
assign LUT_2[14643] = 32'b11111111111111110110111111110011;
assign LUT_2[14644] = 32'b11111111111111101111101100000110;
assign LUT_2[14645] = 32'b11111111111111101100100100011111;
assign LUT_2[14646] = 32'b11111111111111110110100101000010;
assign LUT_2[14647] = 32'b11111111111111110011011101011011;
assign LUT_2[14648] = 32'b11111111111111101101111111111011;
assign LUT_2[14649] = 32'b11111111111111101010111000010100;
assign LUT_2[14650] = 32'b11111111111111110100111000110111;
assign LUT_2[14651] = 32'b11111111111111110001110001010000;
assign LUT_2[14652] = 32'b11111111111111101010011101100011;
assign LUT_2[14653] = 32'b11111111111111100111010101111100;
assign LUT_2[14654] = 32'b11111111111111110001010110011111;
assign LUT_2[14655] = 32'b11111111111111101110001110111000;
assign LUT_2[14656] = 32'b11111111111111110000010111001110;
assign LUT_2[14657] = 32'b11111111111111101101001111100111;
assign LUT_2[14658] = 32'b11111111111111110111010000001010;
assign LUT_2[14659] = 32'b11111111111111110100001000100011;
assign LUT_2[14660] = 32'b11111111111111101100110100110110;
assign LUT_2[14661] = 32'b11111111111111101001101101001111;
assign LUT_2[14662] = 32'b11111111111111110011101101110010;
assign LUT_2[14663] = 32'b11111111111111110000100110001011;
assign LUT_2[14664] = 32'b11111111111111101011001000101011;
assign LUT_2[14665] = 32'b11111111111111101000000001000100;
assign LUT_2[14666] = 32'b11111111111111110010000001100111;
assign LUT_2[14667] = 32'b11111111111111101110111010000000;
assign LUT_2[14668] = 32'b11111111111111100111100110010011;
assign LUT_2[14669] = 32'b11111111111111100100011110101100;
assign LUT_2[14670] = 32'b11111111111111101110011111001111;
assign LUT_2[14671] = 32'b11111111111111101011010111101000;
assign LUT_2[14672] = 32'b11111111111111101010111011011000;
assign LUT_2[14673] = 32'b11111111111111100111110011110001;
assign LUT_2[14674] = 32'b11111111111111110001110100010100;
assign LUT_2[14675] = 32'b11111111111111101110101100101101;
assign LUT_2[14676] = 32'b11111111111111100111011001000000;
assign LUT_2[14677] = 32'b11111111111111100100010001011001;
assign LUT_2[14678] = 32'b11111111111111101110010001111100;
assign LUT_2[14679] = 32'b11111111111111101011001010010101;
assign LUT_2[14680] = 32'b11111111111111100101101100110101;
assign LUT_2[14681] = 32'b11111111111111100010100101001110;
assign LUT_2[14682] = 32'b11111111111111101100100101110001;
assign LUT_2[14683] = 32'b11111111111111101001011110001010;
assign LUT_2[14684] = 32'b11111111111111100010001010011101;
assign LUT_2[14685] = 32'b11111111111111011111000010110110;
assign LUT_2[14686] = 32'b11111111111111101001000011011001;
assign LUT_2[14687] = 32'b11111111111111100101111011110010;
assign LUT_2[14688] = 32'b11111111111111110000110010110111;
assign LUT_2[14689] = 32'b11111111111111101101101011010000;
assign LUT_2[14690] = 32'b11111111111111110111101011110011;
assign LUT_2[14691] = 32'b11111111111111110100100100001100;
assign LUT_2[14692] = 32'b11111111111111101101010000011111;
assign LUT_2[14693] = 32'b11111111111111101010001000111000;
assign LUT_2[14694] = 32'b11111111111111110100001001011011;
assign LUT_2[14695] = 32'b11111111111111110001000001110100;
assign LUT_2[14696] = 32'b11111111111111101011100100010100;
assign LUT_2[14697] = 32'b11111111111111101000011100101101;
assign LUT_2[14698] = 32'b11111111111111110010011101010000;
assign LUT_2[14699] = 32'b11111111111111101111010101101001;
assign LUT_2[14700] = 32'b11111111111111101000000001111100;
assign LUT_2[14701] = 32'b11111111111111100100111010010101;
assign LUT_2[14702] = 32'b11111111111111101110111010111000;
assign LUT_2[14703] = 32'b11111111111111101011110011010001;
assign LUT_2[14704] = 32'b11111111111111101011010111000001;
assign LUT_2[14705] = 32'b11111111111111101000001111011010;
assign LUT_2[14706] = 32'b11111111111111110010001111111101;
assign LUT_2[14707] = 32'b11111111111111101111001000010110;
assign LUT_2[14708] = 32'b11111111111111100111110100101001;
assign LUT_2[14709] = 32'b11111111111111100100101101000010;
assign LUT_2[14710] = 32'b11111111111111101110101101100101;
assign LUT_2[14711] = 32'b11111111111111101011100101111110;
assign LUT_2[14712] = 32'b11111111111111100110001000011110;
assign LUT_2[14713] = 32'b11111111111111100011000000110111;
assign LUT_2[14714] = 32'b11111111111111101101000001011010;
assign LUT_2[14715] = 32'b11111111111111101001111001110011;
assign LUT_2[14716] = 32'b11111111111111100010100110000110;
assign LUT_2[14717] = 32'b11111111111111011111011110011111;
assign LUT_2[14718] = 32'b11111111111111101001011111000010;
assign LUT_2[14719] = 32'b11111111111111100110010111011011;
assign LUT_2[14720] = 32'b11111111111111111100100010111010;
assign LUT_2[14721] = 32'b11111111111111111001011011010011;
assign LUT_2[14722] = 32'b00000000000000000011011011110110;
assign LUT_2[14723] = 32'b00000000000000000000010100001111;
assign LUT_2[14724] = 32'b11111111111111111001000000100010;
assign LUT_2[14725] = 32'b11111111111111110101111000111011;
assign LUT_2[14726] = 32'b11111111111111111111111001011110;
assign LUT_2[14727] = 32'b11111111111111111100110001110111;
assign LUT_2[14728] = 32'b11111111111111110111010100010111;
assign LUT_2[14729] = 32'b11111111111111110100001100110000;
assign LUT_2[14730] = 32'b11111111111111111110001101010011;
assign LUT_2[14731] = 32'b11111111111111111011000101101100;
assign LUT_2[14732] = 32'b11111111111111110011110001111111;
assign LUT_2[14733] = 32'b11111111111111110000101010011000;
assign LUT_2[14734] = 32'b11111111111111111010101010111011;
assign LUT_2[14735] = 32'b11111111111111110111100011010100;
assign LUT_2[14736] = 32'b11111111111111110111000111000100;
assign LUT_2[14737] = 32'b11111111111111110011111111011101;
assign LUT_2[14738] = 32'b11111111111111111110000000000000;
assign LUT_2[14739] = 32'b11111111111111111010111000011001;
assign LUT_2[14740] = 32'b11111111111111110011100100101100;
assign LUT_2[14741] = 32'b11111111111111110000011101000101;
assign LUT_2[14742] = 32'b11111111111111111010011101101000;
assign LUT_2[14743] = 32'b11111111111111110111010110000001;
assign LUT_2[14744] = 32'b11111111111111110001111000100001;
assign LUT_2[14745] = 32'b11111111111111101110110000111010;
assign LUT_2[14746] = 32'b11111111111111111000110001011101;
assign LUT_2[14747] = 32'b11111111111111110101101001110110;
assign LUT_2[14748] = 32'b11111111111111101110010110001001;
assign LUT_2[14749] = 32'b11111111111111101011001110100010;
assign LUT_2[14750] = 32'b11111111111111110101001111000101;
assign LUT_2[14751] = 32'b11111111111111110010000111011110;
assign LUT_2[14752] = 32'b11111111111111111100111110100011;
assign LUT_2[14753] = 32'b11111111111111111001110110111100;
assign LUT_2[14754] = 32'b00000000000000000011110111011111;
assign LUT_2[14755] = 32'b00000000000000000000101111111000;
assign LUT_2[14756] = 32'b11111111111111111001011100001011;
assign LUT_2[14757] = 32'b11111111111111110110010100100100;
assign LUT_2[14758] = 32'b00000000000000000000010101000111;
assign LUT_2[14759] = 32'b11111111111111111101001101100000;
assign LUT_2[14760] = 32'b11111111111111110111110000000000;
assign LUT_2[14761] = 32'b11111111111111110100101000011001;
assign LUT_2[14762] = 32'b11111111111111111110101000111100;
assign LUT_2[14763] = 32'b11111111111111111011100001010101;
assign LUT_2[14764] = 32'b11111111111111110100001101101000;
assign LUT_2[14765] = 32'b11111111111111110001000110000001;
assign LUT_2[14766] = 32'b11111111111111111011000110100100;
assign LUT_2[14767] = 32'b11111111111111110111111110111101;
assign LUT_2[14768] = 32'b11111111111111110111100010101101;
assign LUT_2[14769] = 32'b11111111111111110100011011000110;
assign LUT_2[14770] = 32'b11111111111111111110011011101001;
assign LUT_2[14771] = 32'b11111111111111111011010100000010;
assign LUT_2[14772] = 32'b11111111111111110100000000010101;
assign LUT_2[14773] = 32'b11111111111111110000111000101110;
assign LUT_2[14774] = 32'b11111111111111111010111001010001;
assign LUT_2[14775] = 32'b11111111111111110111110001101010;
assign LUT_2[14776] = 32'b11111111111111110010010100001010;
assign LUT_2[14777] = 32'b11111111111111101111001100100011;
assign LUT_2[14778] = 32'b11111111111111111001001101000110;
assign LUT_2[14779] = 32'b11111111111111110110000101011111;
assign LUT_2[14780] = 32'b11111111111111101110110001110010;
assign LUT_2[14781] = 32'b11111111111111101011101010001011;
assign LUT_2[14782] = 32'b11111111111111110101101010101110;
assign LUT_2[14783] = 32'b11111111111111110010100011000111;
assign LUT_2[14784] = 32'b11111111111111110100101011011101;
assign LUT_2[14785] = 32'b11111111111111110001100011110110;
assign LUT_2[14786] = 32'b11111111111111111011100100011001;
assign LUT_2[14787] = 32'b11111111111111111000011100110010;
assign LUT_2[14788] = 32'b11111111111111110001001001000101;
assign LUT_2[14789] = 32'b11111111111111101110000001011110;
assign LUT_2[14790] = 32'b11111111111111111000000010000001;
assign LUT_2[14791] = 32'b11111111111111110100111010011010;
assign LUT_2[14792] = 32'b11111111111111101111011100111010;
assign LUT_2[14793] = 32'b11111111111111101100010101010011;
assign LUT_2[14794] = 32'b11111111111111110110010101110110;
assign LUT_2[14795] = 32'b11111111111111110011001110001111;
assign LUT_2[14796] = 32'b11111111111111101011111010100010;
assign LUT_2[14797] = 32'b11111111111111101000110010111011;
assign LUT_2[14798] = 32'b11111111111111110010110011011110;
assign LUT_2[14799] = 32'b11111111111111101111101011110111;
assign LUT_2[14800] = 32'b11111111111111101111001111100111;
assign LUT_2[14801] = 32'b11111111111111101100001000000000;
assign LUT_2[14802] = 32'b11111111111111110110001000100011;
assign LUT_2[14803] = 32'b11111111111111110011000000111100;
assign LUT_2[14804] = 32'b11111111111111101011101101001111;
assign LUT_2[14805] = 32'b11111111111111101000100101101000;
assign LUT_2[14806] = 32'b11111111111111110010100110001011;
assign LUT_2[14807] = 32'b11111111111111101111011110100100;
assign LUT_2[14808] = 32'b11111111111111101010000001000100;
assign LUT_2[14809] = 32'b11111111111111100110111001011101;
assign LUT_2[14810] = 32'b11111111111111110000111010000000;
assign LUT_2[14811] = 32'b11111111111111101101110010011001;
assign LUT_2[14812] = 32'b11111111111111100110011110101100;
assign LUT_2[14813] = 32'b11111111111111100011010111000101;
assign LUT_2[14814] = 32'b11111111111111101101010111101000;
assign LUT_2[14815] = 32'b11111111111111101010010000000001;
assign LUT_2[14816] = 32'b11111111111111110101000111000110;
assign LUT_2[14817] = 32'b11111111111111110001111111011111;
assign LUT_2[14818] = 32'b11111111111111111100000000000010;
assign LUT_2[14819] = 32'b11111111111111111000111000011011;
assign LUT_2[14820] = 32'b11111111111111110001100100101110;
assign LUT_2[14821] = 32'b11111111111111101110011101000111;
assign LUT_2[14822] = 32'b11111111111111111000011101101010;
assign LUT_2[14823] = 32'b11111111111111110101010110000011;
assign LUT_2[14824] = 32'b11111111111111101111111000100011;
assign LUT_2[14825] = 32'b11111111111111101100110000111100;
assign LUT_2[14826] = 32'b11111111111111110110110001011111;
assign LUT_2[14827] = 32'b11111111111111110011101001111000;
assign LUT_2[14828] = 32'b11111111111111101100010110001011;
assign LUT_2[14829] = 32'b11111111111111101001001110100100;
assign LUT_2[14830] = 32'b11111111111111110011001111000111;
assign LUT_2[14831] = 32'b11111111111111110000000111100000;
assign LUT_2[14832] = 32'b11111111111111101111101011010000;
assign LUT_2[14833] = 32'b11111111111111101100100011101001;
assign LUT_2[14834] = 32'b11111111111111110110100100001100;
assign LUT_2[14835] = 32'b11111111111111110011011100100101;
assign LUT_2[14836] = 32'b11111111111111101100001000111000;
assign LUT_2[14837] = 32'b11111111111111101001000001010001;
assign LUT_2[14838] = 32'b11111111111111110011000001110100;
assign LUT_2[14839] = 32'b11111111111111101111111010001101;
assign LUT_2[14840] = 32'b11111111111111101010011100101101;
assign LUT_2[14841] = 32'b11111111111111100111010101000110;
assign LUT_2[14842] = 32'b11111111111111110001010101101001;
assign LUT_2[14843] = 32'b11111111111111101110001110000010;
assign LUT_2[14844] = 32'b11111111111111100110111010010101;
assign LUT_2[14845] = 32'b11111111111111100011110010101110;
assign LUT_2[14846] = 32'b11111111111111101101110011010001;
assign LUT_2[14847] = 32'b11111111111111101010101011101010;
assign LUT_2[14848] = 32'b11111111111111111001000001110111;
assign LUT_2[14849] = 32'b11111111111111110101111010010000;
assign LUT_2[14850] = 32'b11111111111111111111111010110011;
assign LUT_2[14851] = 32'b11111111111111111100110011001100;
assign LUT_2[14852] = 32'b11111111111111110101011111011111;
assign LUT_2[14853] = 32'b11111111111111110010010111111000;
assign LUT_2[14854] = 32'b11111111111111111100011000011011;
assign LUT_2[14855] = 32'b11111111111111111001010000110100;
assign LUT_2[14856] = 32'b11111111111111110011110011010100;
assign LUT_2[14857] = 32'b11111111111111110000101011101101;
assign LUT_2[14858] = 32'b11111111111111111010101100010000;
assign LUT_2[14859] = 32'b11111111111111110111100100101001;
assign LUT_2[14860] = 32'b11111111111111110000010000111100;
assign LUT_2[14861] = 32'b11111111111111101101001001010101;
assign LUT_2[14862] = 32'b11111111111111110111001001111000;
assign LUT_2[14863] = 32'b11111111111111110100000010010001;
assign LUT_2[14864] = 32'b11111111111111110011100110000001;
assign LUT_2[14865] = 32'b11111111111111110000011110011010;
assign LUT_2[14866] = 32'b11111111111111111010011110111101;
assign LUT_2[14867] = 32'b11111111111111110111010111010110;
assign LUT_2[14868] = 32'b11111111111111110000000011101001;
assign LUT_2[14869] = 32'b11111111111111101100111100000010;
assign LUT_2[14870] = 32'b11111111111111110110111100100101;
assign LUT_2[14871] = 32'b11111111111111110011110100111110;
assign LUT_2[14872] = 32'b11111111111111101110010111011110;
assign LUT_2[14873] = 32'b11111111111111101011001111110111;
assign LUT_2[14874] = 32'b11111111111111110101010000011010;
assign LUT_2[14875] = 32'b11111111111111110010001000110011;
assign LUT_2[14876] = 32'b11111111111111101010110101000110;
assign LUT_2[14877] = 32'b11111111111111100111101101011111;
assign LUT_2[14878] = 32'b11111111111111110001101110000010;
assign LUT_2[14879] = 32'b11111111111111101110100110011011;
assign LUT_2[14880] = 32'b11111111111111111001011101100000;
assign LUT_2[14881] = 32'b11111111111111110110010101111001;
assign LUT_2[14882] = 32'b00000000000000000000010110011100;
assign LUT_2[14883] = 32'b11111111111111111101001110110101;
assign LUT_2[14884] = 32'b11111111111111110101111011001000;
assign LUT_2[14885] = 32'b11111111111111110010110011100001;
assign LUT_2[14886] = 32'b11111111111111111100110100000100;
assign LUT_2[14887] = 32'b11111111111111111001101100011101;
assign LUT_2[14888] = 32'b11111111111111110100001110111101;
assign LUT_2[14889] = 32'b11111111111111110001000111010110;
assign LUT_2[14890] = 32'b11111111111111111011000111111001;
assign LUT_2[14891] = 32'b11111111111111111000000000010010;
assign LUT_2[14892] = 32'b11111111111111110000101100100101;
assign LUT_2[14893] = 32'b11111111111111101101100100111110;
assign LUT_2[14894] = 32'b11111111111111110111100101100001;
assign LUT_2[14895] = 32'b11111111111111110100011101111010;
assign LUT_2[14896] = 32'b11111111111111110100000001101010;
assign LUT_2[14897] = 32'b11111111111111110000111010000011;
assign LUT_2[14898] = 32'b11111111111111111010111010100110;
assign LUT_2[14899] = 32'b11111111111111110111110010111111;
assign LUT_2[14900] = 32'b11111111111111110000011111010010;
assign LUT_2[14901] = 32'b11111111111111101101010111101011;
assign LUT_2[14902] = 32'b11111111111111110111011000001110;
assign LUT_2[14903] = 32'b11111111111111110100010000100111;
assign LUT_2[14904] = 32'b11111111111111101110110011000111;
assign LUT_2[14905] = 32'b11111111111111101011101011100000;
assign LUT_2[14906] = 32'b11111111111111110101101100000011;
assign LUT_2[14907] = 32'b11111111111111110010100100011100;
assign LUT_2[14908] = 32'b11111111111111101011010000101111;
assign LUT_2[14909] = 32'b11111111111111101000001001001000;
assign LUT_2[14910] = 32'b11111111111111110010001001101011;
assign LUT_2[14911] = 32'b11111111111111101111000010000100;
assign LUT_2[14912] = 32'b11111111111111110001001010011010;
assign LUT_2[14913] = 32'b11111111111111101110000010110011;
assign LUT_2[14914] = 32'b11111111111111111000000011010110;
assign LUT_2[14915] = 32'b11111111111111110100111011101111;
assign LUT_2[14916] = 32'b11111111111111101101101000000010;
assign LUT_2[14917] = 32'b11111111111111101010100000011011;
assign LUT_2[14918] = 32'b11111111111111110100100000111110;
assign LUT_2[14919] = 32'b11111111111111110001011001010111;
assign LUT_2[14920] = 32'b11111111111111101011111011110111;
assign LUT_2[14921] = 32'b11111111111111101000110100010000;
assign LUT_2[14922] = 32'b11111111111111110010110100110011;
assign LUT_2[14923] = 32'b11111111111111101111101101001100;
assign LUT_2[14924] = 32'b11111111111111101000011001011111;
assign LUT_2[14925] = 32'b11111111111111100101010001111000;
assign LUT_2[14926] = 32'b11111111111111101111010010011011;
assign LUT_2[14927] = 32'b11111111111111101100001010110100;
assign LUT_2[14928] = 32'b11111111111111101011101110100100;
assign LUT_2[14929] = 32'b11111111111111101000100110111101;
assign LUT_2[14930] = 32'b11111111111111110010100111100000;
assign LUT_2[14931] = 32'b11111111111111101111011111111001;
assign LUT_2[14932] = 32'b11111111111111101000001100001100;
assign LUT_2[14933] = 32'b11111111111111100101000100100101;
assign LUT_2[14934] = 32'b11111111111111101111000101001000;
assign LUT_2[14935] = 32'b11111111111111101011111101100001;
assign LUT_2[14936] = 32'b11111111111111100110100000000001;
assign LUT_2[14937] = 32'b11111111111111100011011000011010;
assign LUT_2[14938] = 32'b11111111111111101101011000111101;
assign LUT_2[14939] = 32'b11111111111111101010010001010110;
assign LUT_2[14940] = 32'b11111111111111100010111101101001;
assign LUT_2[14941] = 32'b11111111111111011111110110000010;
assign LUT_2[14942] = 32'b11111111111111101001110110100101;
assign LUT_2[14943] = 32'b11111111111111100110101110111110;
assign LUT_2[14944] = 32'b11111111111111110001100110000011;
assign LUT_2[14945] = 32'b11111111111111101110011110011100;
assign LUT_2[14946] = 32'b11111111111111111000011110111111;
assign LUT_2[14947] = 32'b11111111111111110101010111011000;
assign LUT_2[14948] = 32'b11111111111111101110000011101011;
assign LUT_2[14949] = 32'b11111111111111101010111100000100;
assign LUT_2[14950] = 32'b11111111111111110100111100100111;
assign LUT_2[14951] = 32'b11111111111111110001110101000000;
assign LUT_2[14952] = 32'b11111111111111101100010111100000;
assign LUT_2[14953] = 32'b11111111111111101001001111111001;
assign LUT_2[14954] = 32'b11111111111111110011010000011100;
assign LUT_2[14955] = 32'b11111111111111110000001000110101;
assign LUT_2[14956] = 32'b11111111111111101000110101001000;
assign LUT_2[14957] = 32'b11111111111111100101101101100001;
assign LUT_2[14958] = 32'b11111111111111101111101110000100;
assign LUT_2[14959] = 32'b11111111111111101100100110011101;
assign LUT_2[14960] = 32'b11111111111111101100001010001101;
assign LUT_2[14961] = 32'b11111111111111101001000010100110;
assign LUT_2[14962] = 32'b11111111111111110011000011001001;
assign LUT_2[14963] = 32'b11111111111111101111111011100010;
assign LUT_2[14964] = 32'b11111111111111101000100111110101;
assign LUT_2[14965] = 32'b11111111111111100101100000001110;
assign LUT_2[14966] = 32'b11111111111111101111100000110001;
assign LUT_2[14967] = 32'b11111111111111101100011001001010;
assign LUT_2[14968] = 32'b11111111111111100110111011101010;
assign LUT_2[14969] = 32'b11111111111111100011110100000011;
assign LUT_2[14970] = 32'b11111111111111101101110100100110;
assign LUT_2[14971] = 32'b11111111111111101010101100111111;
assign LUT_2[14972] = 32'b11111111111111100011011001010010;
assign LUT_2[14973] = 32'b11111111111111100000010001101011;
assign LUT_2[14974] = 32'b11111111111111101010010010001110;
assign LUT_2[14975] = 32'b11111111111111100111001010100111;
assign LUT_2[14976] = 32'b11111111111111111101010110000110;
assign LUT_2[14977] = 32'b11111111111111111010001110011111;
assign LUT_2[14978] = 32'b00000000000000000100001111000010;
assign LUT_2[14979] = 32'b00000000000000000001000111011011;
assign LUT_2[14980] = 32'b11111111111111111001110011101110;
assign LUT_2[14981] = 32'b11111111111111110110101100000111;
assign LUT_2[14982] = 32'b00000000000000000000101100101010;
assign LUT_2[14983] = 32'b11111111111111111101100101000011;
assign LUT_2[14984] = 32'b11111111111111111000000111100011;
assign LUT_2[14985] = 32'b11111111111111110100111111111100;
assign LUT_2[14986] = 32'b11111111111111111111000000011111;
assign LUT_2[14987] = 32'b11111111111111111011111000111000;
assign LUT_2[14988] = 32'b11111111111111110100100101001011;
assign LUT_2[14989] = 32'b11111111111111110001011101100100;
assign LUT_2[14990] = 32'b11111111111111111011011110000111;
assign LUT_2[14991] = 32'b11111111111111111000010110100000;
assign LUT_2[14992] = 32'b11111111111111110111111010010000;
assign LUT_2[14993] = 32'b11111111111111110100110010101001;
assign LUT_2[14994] = 32'b11111111111111111110110011001100;
assign LUT_2[14995] = 32'b11111111111111111011101011100101;
assign LUT_2[14996] = 32'b11111111111111110100010111111000;
assign LUT_2[14997] = 32'b11111111111111110001010000010001;
assign LUT_2[14998] = 32'b11111111111111111011010000110100;
assign LUT_2[14999] = 32'b11111111111111111000001001001101;
assign LUT_2[15000] = 32'b11111111111111110010101011101101;
assign LUT_2[15001] = 32'b11111111111111101111100100000110;
assign LUT_2[15002] = 32'b11111111111111111001100100101001;
assign LUT_2[15003] = 32'b11111111111111110110011101000010;
assign LUT_2[15004] = 32'b11111111111111101111001001010101;
assign LUT_2[15005] = 32'b11111111111111101100000001101110;
assign LUT_2[15006] = 32'b11111111111111110110000010010001;
assign LUT_2[15007] = 32'b11111111111111110010111010101010;
assign LUT_2[15008] = 32'b11111111111111111101110001101111;
assign LUT_2[15009] = 32'b11111111111111111010101010001000;
assign LUT_2[15010] = 32'b00000000000000000100101010101011;
assign LUT_2[15011] = 32'b00000000000000000001100011000100;
assign LUT_2[15012] = 32'b11111111111111111010001111010111;
assign LUT_2[15013] = 32'b11111111111111110111000111110000;
assign LUT_2[15014] = 32'b00000000000000000001001000010011;
assign LUT_2[15015] = 32'b11111111111111111110000000101100;
assign LUT_2[15016] = 32'b11111111111111111000100011001100;
assign LUT_2[15017] = 32'b11111111111111110101011011100101;
assign LUT_2[15018] = 32'b11111111111111111111011100001000;
assign LUT_2[15019] = 32'b11111111111111111100010100100001;
assign LUT_2[15020] = 32'b11111111111111110101000000110100;
assign LUT_2[15021] = 32'b11111111111111110001111001001101;
assign LUT_2[15022] = 32'b11111111111111111011111001110000;
assign LUT_2[15023] = 32'b11111111111111111000110010001001;
assign LUT_2[15024] = 32'b11111111111111111000010101111001;
assign LUT_2[15025] = 32'b11111111111111110101001110010010;
assign LUT_2[15026] = 32'b11111111111111111111001110110101;
assign LUT_2[15027] = 32'b11111111111111111100000111001110;
assign LUT_2[15028] = 32'b11111111111111110100110011100001;
assign LUT_2[15029] = 32'b11111111111111110001101011111010;
assign LUT_2[15030] = 32'b11111111111111111011101100011101;
assign LUT_2[15031] = 32'b11111111111111111000100100110110;
assign LUT_2[15032] = 32'b11111111111111110011000111010110;
assign LUT_2[15033] = 32'b11111111111111101111111111101111;
assign LUT_2[15034] = 32'b11111111111111111010000000010010;
assign LUT_2[15035] = 32'b11111111111111110110111000101011;
assign LUT_2[15036] = 32'b11111111111111101111100100111110;
assign LUT_2[15037] = 32'b11111111111111101100011101010111;
assign LUT_2[15038] = 32'b11111111111111110110011101111010;
assign LUT_2[15039] = 32'b11111111111111110011010110010011;
assign LUT_2[15040] = 32'b11111111111111110101011110101001;
assign LUT_2[15041] = 32'b11111111111111110010010111000010;
assign LUT_2[15042] = 32'b11111111111111111100010111100101;
assign LUT_2[15043] = 32'b11111111111111111001001111111110;
assign LUT_2[15044] = 32'b11111111111111110001111100010001;
assign LUT_2[15045] = 32'b11111111111111101110110100101010;
assign LUT_2[15046] = 32'b11111111111111111000110101001101;
assign LUT_2[15047] = 32'b11111111111111110101101101100110;
assign LUT_2[15048] = 32'b11111111111111110000010000000110;
assign LUT_2[15049] = 32'b11111111111111101101001000011111;
assign LUT_2[15050] = 32'b11111111111111110111001001000010;
assign LUT_2[15051] = 32'b11111111111111110100000001011011;
assign LUT_2[15052] = 32'b11111111111111101100101101101110;
assign LUT_2[15053] = 32'b11111111111111101001100110000111;
assign LUT_2[15054] = 32'b11111111111111110011100110101010;
assign LUT_2[15055] = 32'b11111111111111110000011111000011;
assign LUT_2[15056] = 32'b11111111111111110000000010110011;
assign LUT_2[15057] = 32'b11111111111111101100111011001100;
assign LUT_2[15058] = 32'b11111111111111110110111011101111;
assign LUT_2[15059] = 32'b11111111111111110011110100001000;
assign LUT_2[15060] = 32'b11111111111111101100100000011011;
assign LUT_2[15061] = 32'b11111111111111101001011000110100;
assign LUT_2[15062] = 32'b11111111111111110011011001010111;
assign LUT_2[15063] = 32'b11111111111111110000010001110000;
assign LUT_2[15064] = 32'b11111111111111101010110100010000;
assign LUT_2[15065] = 32'b11111111111111100111101100101001;
assign LUT_2[15066] = 32'b11111111111111110001101101001100;
assign LUT_2[15067] = 32'b11111111111111101110100101100101;
assign LUT_2[15068] = 32'b11111111111111100111010001111000;
assign LUT_2[15069] = 32'b11111111111111100100001010010001;
assign LUT_2[15070] = 32'b11111111111111101110001010110100;
assign LUT_2[15071] = 32'b11111111111111101011000011001101;
assign LUT_2[15072] = 32'b11111111111111110101111010010010;
assign LUT_2[15073] = 32'b11111111111111110010110010101011;
assign LUT_2[15074] = 32'b11111111111111111100110011001110;
assign LUT_2[15075] = 32'b11111111111111111001101011100111;
assign LUT_2[15076] = 32'b11111111111111110010010111111010;
assign LUT_2[15077] = 32'b11111111111111101111010000010011;
assign LUT_2[15078] = 32'b11111111111111111001010000110110;
assign LUT_2[15079] = 32'b11111111111111110110001001001111;
assign LUT_2[15080] = 32'b11111111111111110000101011101111;
assign LUT_2[15081] = 32'b11111111111111101101100100001000;
assign LUT_2[15082] = 32'b11111111111111110111100100101011;
assign LUT_2[15083] = 32'b11111111111111110100011101000100;
assign LUT_2[15084] = 32'b11111111111111101101001001010111;
assign LUT_2[15085] = 32'b11111111111111101010000001110000;
assign LUT_2[15086] = 32'b11111111111111110100000010010011;
assign LUT_2[15087] = 32'b11111111111111110000111010101100;
assign LUT_2[15088] = 32'b11111111111111110000011110011100;
assign LUT_2[15089] = 32'b11111111111111101101010110110101;
assign LUT_2[15090] = 32'b11111111111111110111010111011000;
assign LUT_2[15091] = 32'b11111111111111110100001111110001;
assign LUT_2[15092] = 32'b11111111111111101100111100000100;
assign LUT_2[15093] = 32'b11111111111111101001110100011101;
assign LUT_2[15094] = 32'b11111111111111110011110101000000;
assign LUT_2[15095] = 32'b11111111111111110000101101011001;
assign LUT_2[15096] = 32'b11111111111111101011001111111001;
assign LUT_2[15097] = 32'b11111111111111101000001000010010;
assign LUT_2[15098] = 32'b11111111111111110010001000110101;
assign LUT_2[15099] = 32'b11111111111111101111000001001110;
assign LUT_2[15100] = 32'b11111111111111100111101101100001;
assign LUT_2[15101] = 32'b11111111111111100100100101111010;
assign LUT_2[15102] = 32'b11111111111111101110100110011101;
assign LUT_2[15103] = 32'b11111111111111101011011110110110;
assign LUT_2[15104] = 32'b11111111111111111101000000011101;
assign LUT_2[15105] = 32'b11111111111111111001111000110110;
assign LUT_2[15106] = 32'b00000000000000000011111001011001;
assign LUT_2[15107] = 32'b00000000000000000000110001110010;
assign LUT_2[15108] = 32'b11111111111111111001011110000101;
assign LUT_2[15109] = 32'b11111111111111110110010110011110;
assign LUT_2[15110] = 32'b00000000000000000000010111000001;
assign LUT_2[15111] = 32'b11111111111111111101001111011010;
assign LUT_2[15112] = 32'b11111111111111110111110001111010;
assign LUT_2[15113] = 32'b11111111111111110100101010010011;
assign LUT_2[15114] = 32'b11111111111111111110101010110110;
assign LUT_2[15115] = 32'b11111111111111111011100011001111;
assign LUT_2[15116] = 32'b11111111111111110100001111100010;
assign LUT_2[15117] = 32'b11111111111111110001000111111011;
assign LUT_2[15118] = 32'b11111111111111111011001000011110;
assign LUT_2[15119] = 32'b11111111111111111000000000110111;
assign LUT_2[15120] = 32'b11111111111111110111100100100111;
assign LUT_2[15121] = 32'b11111111111111110100011101000000;
assign LUT_2[15122] = 32'b11111111111111111110011101100011;
assign LUT_2[15123] = 32'b11111111111111111011010101111100;
assign LUT_2[15124] = 32'b11111111111111110100000010001111;
assign LUT_2[15125] = 32'b11111111111111110000111010101000;
assign LUT_2[15126] = 32'b11111111111111111010111011001011;
assign LUT_2[15127] = 32'b11111111111111110111110011100100;
assign LUT_2[15128] = 32'b11111111111111110010010110000100;
assign LUT_2[15129] = 32'b11111111111111101111001110011101;
assign LUT_2[15130] = 32'b11111111111111111001001111000000;
assign LUT_2[15131] = 32'b11111111111111110110000111011001;
assign LUT_2[15132] = 32'b11111111111111101110110011101100;
assign LUT_2[15133] = 32'b11111111111111101011101100000101;
assign LUT_2[15134] = 32'b11111111111111110101101100101000;
assign LUT_2[15135] = 32'b11111111111111110010100101000001;
assign LUT_2[15136] = 32'b11111111111111111101011100000110;
assign LUT_2[15137] = 32'b11111111111111111010010100011111;
assign LUT_2[15138] = 32'b00000000000000000100010101000010;
assign LUT_2[15139] = 32'b00000000000000000001001101011011;
assign LUT_2[15140] = 32'b11111111111111111001111001101110;
assign LUT_2[15141] = 32'b11111111111111110110110010000111;
assign LUT_2[15142] = 32'b00000000000000000000110010101010;
assign LUT_2[15143] = 32'b11111111111111111101101011000011;
assign LUT_2[15144] = 32'b11111111111111111000001101100011;
assign LUT_2[15145] = 32'b11111111111111110101000101111100;
assign LUT_2[15146] = 32'b11111111111111111111000110011111;
assign LUT_2[15147] = 32'b11111111111111111011111110111000;
assign LUT_2[15148] = 32'b11111111111111110100101011001011;
assign LUT_2[15149] = 32'b11111111111111110001100011100100;
assign LUT_2[15150] = 32'b11111111111111111011100100000111;
assign LUT_2[15151] = 32'b11111111111111111000011100100000;
assign LUT_2[15152] = 32'b11111111111111111000000000010000;
assign LUT_2[15153] = 32'b11111111111111110100111000101001;
assign LUT_2[15154] = 32'b11111111111111111110111001001100;
assign LUT_2[15155] = 32'b11111111111111111011110001100101;
assign LUT_2[15156] = 32'b11111111111111110100011101111000;
assign LUT_2[15157] = 32'b11111111111111110001010110010001;
assign LUT_2[15158] = 32'b11111111111111111011010110110100;
assign LUT_2[15159] = 32'b11111111111111111000001111001101;
assign LUT_2[15160] = 32'b11111111111111110010110001101101;
assign LUT_2[15161] = 32'b11111111111111101111101010000110;
assign LUT_2[15162] = 32'b11111111111111111001101010101001;
assign LUT_2[15163] = 32'b11111111111111110110100011000010;
assign LUT_2[15164] = 32'b11111111111111101111001111010101;
assign LUT_2[15165] = 32'b11111111111111101100000111101110;
assign LUT_2[15166] = 32'b11111111111111110110001000010001;
assign LUT_2[15167] = 32'b11111111111111110011000000101010;
assign LUT_2[15168] = 32'b11111111111111110101001001000000;
assign LUT_2[15169] = 32'b11111111111111110010000001011001;
assign LUT_2[15170] = 32'b11111111111111111100000001111100;
assign LUT_2[15171] = 32'b11111111111111111000111010010101;
assign LUT_2[15172] = 32'b11111111111111110001100110101000;
assign LUT_2[15173] = 32'b11111111111111101110011111000001;
assign LUT_2[15174] = 32'b11111111111111111000011111100100;
assign LUT_2[15175] = 32'b11111111111111110101010111111101;
assign LUT_2[15176] = 32'b11111111111111101111111010011101;
assign LUT_2[15177] = 32'b11111111111111101100110010110110;
assign LUT_2[15178] = 32'b11111111111111110110110011011001;
assign LUT_2[15179] = 32'b11111111111111110011101011110010;
assign LUT_2[15180] = 32'b11111111111111101100011000000101;
assign LUT_2[15181] = 32'b11111111111111101001010000011110;
assign LUT_2[15182] = 32'b11111111111111110011010001000001;
assign LUT_2[15183] = 32'b11111111111111110000001001011010;
assign LUT_2[15184] = 32'b11111111111111101111101101001010;
assign LUT_2[15185] = 32'b11111111111111101100100101100011;
assign LUT_2[15186] = 32'b11111111111111110110100110000110;
assign LUT_2[15187] = 32'b11111111111111110011011110011111;
assign LUT_2[15188] = 32'b11111111111111101100001010110010;
assign LUT_2[15189] = 32'b11111111111111101001000011001011;
assign LUT_2[15190] = 32'b11111111111111110011000011101110;
assign LUT_2[15191] = 32'b11111111111111101111111100000111;
assign LUT_2[15192] = 32'b11111111111111101010011110100111;
assign LUT_2[15193] = 32'b11111111111111100111010111000000;
assign LUT_2[15194] = 32'b11111111111111110001010111100011;
assign LUT_2[15195] = 32'b11111111111111101110001111111100;
assign LUT_2[15196] = 32'b11111111111111100110111100001111;
assign LUT_2[15197] = 32'b11111111111111100011110100101000;
assign LUT_2[15198] = 32'b11111111111111101101110101001011;
assign LUT_2[15199] = 32'b11111111111111101010101101100100;
assign LUT_2[15200] = 32'b11111111111111110101100100101001;
assign LUT_2[15201] = 32'b11111111111111110010011101000010;
assign LUT_2[15202] = 32'b11111111111111111100011101100101;
assign LUT_2[15203] = 32'b11111111111111111001010101111110;
assign LUT_2[15204] = 32'b11111111111111110010000010010001;
assign LUT_2[15205] = 32'b11111111111111101110111010101010;
assign LUT_2[15206] = 32'b11111111111111111000111011001101;
assign LUT_2[15207] = 32'b11111111111111110101110011100110;
assign LUT_2[15208] = 32'b11111111111111110000010110000110;
assign LUT_2[15209] = 32'b11111111111111101101001110011111;
assign LUT_2[15210] = 32'b11111111111111110111001111000010;
assign LUT_2[15211] = 32'b11111111111111110100000111011011;
assign LUT_2[15212] = 32'b11111111111111101100110011101110;
assign LUT_2[15213] = 32'b11111111111111101001101100000111;
assign LUT_2[15214] = 32'b11111111111111110011101100101010;
assign LUT_2[15215] = 32'b11111111111111110000100101000011;
assign LUT_2[15216] = 32'b11111111111111110000001000110011;
assign LUT_2[15217] = 32'b11111111111111101101000001001100;
assign LUT_2[15218] = 32'b11111111111111110111000001101111;
assign LUT_2[15219] = 32'b11111111111111110011111010001000;
assign LUT_2[15220] = 32'b11111111111111101100100110011011;
assign LUT_2[15221] = 32'b11111111111111101001011110110100;
assign LUT_2[15222] = 32'b11111111111111110011011111010111;
assign LUT_2[15223] = 32'b11111111111111110000010111110000;
assign LUT_2[15224] = 32'b11111111111111101010111010010000;
assign LUT_2[15225] = 32'b11111111111111100111110010101001;
assign LUT_2[15226] = 32'b11111111111111110001110011001100;
assign LUT_2[15227] = 32'b11111111111111101110101011100101;
assign LUT_2[15228] = 32'b11111111111111100111010111111000;
assign LUT_2[15229] = 32'b11111111111111100100010000010001;
assign LUT_2[15230] = 32'b11111111111111101110010000110100;
assign LUT_2[15231] = 32'b11111111111111101011001001001101;
assign LUT_2[15232] = 32'b00000000000000000001010100101100;
assign LUT_2[15233] = 32'b11111111111111111110001101000101;
assign LUT_2[15234] = 32'b00000000000000001000001101101000;
assign LUT_2[15235] = 32'b00000000000000000101000110000001;
assign LUT_2[15236] = 32'b11111111111111111101110010010100;
assign LUT_2[15237] = 32'b11111111111111111010101010101101;
assign LUT_2[15238] = 32'b00000000000000000100101011010000;
assign LUT_2[15239] = 32'b00000000000000000001100011101001;
assign LUT_2[15240] = 32'b11111111111111111100000110001001;
assign LUT_2[15241] = 32'b11111111111111111000111110100010;
assign LUT_2[15242] = 32'b00000000000000000010111111000101;
assign LUT_2[15243] = 32'b11111111111111111111110111011110;
assign LUT_2[15244] = 32'b11111111111111111000100011110001;
assign LUT_2[15245] = 32'b11111111111111110101011100001010;
assign LUT_2[15246] = 32'b11111111111111111111011100101101;
assign LUT_2[15247] = 32'b11111111111111111100010101000110;
assign LUT_2[15248] = 32'b11111111111111111011111000110110;
assign LUT_2[15249] = 32'b11111111111111111000110001001111;
assign LUT_2[15250] = 32'b00000000000000000010110001110010;
assign LUT_2[15251] = 32'b11111111111111111111101010001011;
assign LUT_2[15252] = 32'b11111111111111111000010110011110;
assign LUT_2[15253] = 32'b11111111111111110101001110110111;
assign LUT_2[15254] = 32'b11111111111111111111001111011010;
assign LUT_2[15255] = 32'b11111111111111111100000111110011;
assign LUT_2[15256] = 32'b11111111111111110110101010010011;
assign LUT_2[15257] = 32'b11111111111111110011100010101100;
assign LUT_2[15258] = 32'b11111111111111111101100011001111;
assign LUT_2[15259] = 32'b11111111111111111010011011101000;
assign LUT_2[15260] = 32'b11111111111111110011000111111011;
assign LUT_2[15261] = 32'b11111111111111110000000000010100;
assign LUT_2[15262] = 32'b11111111111111111010000000110111;
assign LUT_2[15263] = 32'b11111111111111110110111001010000;
assign LUT_2[15264] = 32'b00000000000000000001110000010101;
assign LUT_2[15265] = 32'b11111111111111111110101000101110;
assign LUT_2[15266] = 32'b00000000000000001000101001010001;
assign LUT_2[15267] = 32'b00000000000000000101100001101010;
assign LUT_2[15268] = 32'b11111111111111111110001101111101;
assign LUT_2[15269] = 32'b11111111111111111011000110010110;
assign LUT_2[15270] = 32'b00000000000000000101000110111001;
assign LUT_2[15271] = 32'b00000000000000000001111111010010;
assign LUT_2[15272] = 32'b11111111111111111100100001110010;
assign LUT_2[15273] = 32'b11111111111111111001011010001011;
assign LUT_2[15274] = 32'b00000000000000000011011010101110;
assign LUT_2[15275] = 32'b00000000000000000000010011000111;
assign LUT_2[15276] = 32'b11111111111111111000111111011010;
assign LUT_2[15277] = 32'b11111111111111110101110111110011;
assign LUT_2[15278] = 32'b11111111111111111111111000010110;
assign LUT_2[15279] = 32'b11111111111111111100110000101111;
assign LUT_2[15280] = 32'b11111111111111111100010100011111;
assign LUT_2[15281] = 32'b11111111111111111001001100111000;
assign LUT_2[15282] = 32'b00000000000000000011001101011011;
assign LUT_2[15283] = 32'b00000000000000000000000101110100;
assign LUT_2[15284] = 32'b11111111111111111000110010000111;
assign LUT_2[15285] = 32'b11111111111111110101101010100000;
assign LUT_2[15286] = 32'b11111111111111111111101011000011;
assign LUT_2[15287] = 32'b11111111111111111100100011011100;
assign LUT_2[15288] = 32'b11111111111111110111000101111100;
assign LUT_2[15289] = 32'b11111111111111110011111110010101;
assign LUT_2[15290] = 32'b11111111111111111101111110111000;
assign LUT_2[15291] = 32'b11111111111111111010110111010001;
assign LUT_2[15292] = 32'b11111111111111110011100011100100;
assign LUT_2[15293] = 32'b11111111111111110000011011111101;
assign LUT_2[15294] = 32'b11111111111111111010011100100000;
assign LUT_2[15295] = 32'b11111111111111110111010100111001;
assign LUT_2[15296] = 32'b11111111111111111001011101001111;
assign LUT_2[15297] = 32'b11111111111111110110010101101000;
assign LUT_2[15298] = 32'b00000000000000000000010110001011;
assign LUT_2[15299] = 32'b11111111111111111101001110100100;
assign LUT_2[15300] = 32'b11111111111111110101111010110111;
assign LUT_2[15301] = 32'b11111111111111110010110011010000;
assign LUT_2[15302] = 32'b11111111111111111100110011110011;
assign LUT_2[15303] = 32'b11111111111111111001101100001100;
assign LUT_2[15304] = 32'b11111111111111110100001110101100;
assign LUT_2[15305] = 32'b11111111111111110001000111000101;
assign LUT_2[15306] = 32'b11111111111111111011000111101000;
assign LUT_2[15307] = 32'b11111111111111111000000000000001;
assign LUT_2[15308] = 32'b11111111111111110000101100010100;
assign LUT_2[15309] = 32'b11111111111111101101100100101101;
assign LUT_2[15310] = 32'b11111111111111110111100101010000;
assign LUT_2[15311] = 32'b11111111111111110100011101101001;
assign LUT_2[15312] = 32'b11111111111111110100000001011001;
assign LUT_2[15313] = 32'b11111111111111110000111001110010;
assign LUT_2[15314] = 32'b11111111111111111010111010010101;
assign LUT_2[15315] = 32'b11111111111111110111110010101110;
assign LUT_2[15316] = 32'b11111111111111110000011111000001;
assign LUT_2[15317] = 32'b11111111111111101101010111011010;
assign LUT_2[15318] = 32'b11111111111111110111010111111101;
assign LUT_2[15319] = 32'b11111111111111110100010000010110;
assign LUT_2[15320] = 32'b11111111111111101110110010110110;
assign LUT_2[15321] = 32'b11111111111111101011101011001111;
assign LUT_2[15322] = 32'b11111111111111110101101011110010;
assign LUT_2[15323] = 32'b11111111111111110010100100001011;
assign LUT_2[15324] = 32'b11111111111111101011010000011110;
assign LUT_2[15325] = 32'b11111111111111101000001000110111;
assign LUT_2[15326] = 32'b11111111111111110010001001011010;
assign LUT_2[15327] = 32'b11111111111111101111000001110011;
assign LUT_2[15328] = 32'b11111111111111111001111000111000;
assign LUT_2[15329] = 32'b11111111111111110110110001010001;
assign LUT_2[15330] = 32'b00000000000000000000110001110100;
assign LUT_2[15331] = 32'b11111111111111111101101010001101;
assign LUT_2[15332] = 32'b11111111111111110110010110100000;
assign LUT_2[15333] = 32'b11111111111111110011001110111001;
assign LUT_2[15334] = 32'b11111111111111111101001111011100;
assign LUT_2[15335] = 32'b11111111111111111010000111110101;
assign LUT_2[15336] = 32'b11111111111111110100101010010101;
assign LUT_2[15337] = 32'b11111111111111110001100010101110;
assign LUT_2[15338] = 32'b11111111111111111011100011010001;
assign LUT_2[15339] = 32'b11111111111111111000011011101010;
assign LUT_2[15340] = 32'b11111111111111110001000111111101;
assign LUT_2[15341] = 32'b11111111111111101110000000010110;
assign LUT_2[15342] = 32'b11111111111111111000000000111001;
assign LUT_2[15343] = 32'b11111111111111110100111001010010;
assign LUT_2[15344] = 32'b11111111111111110100011101000010;
assign LUT_2[15345] = 32'b11111111111111110001010101011011;
assign LUT_2[15346] = 32'b11111111111111111011010101111110;
assign LUT_2[15347] = 32'b11111111111111111000001110010111;
assign LUT_2[15348] = 32'b11111111111111110000111010101010;
assign LUT_2[15349] = 32'b11111111111111101101110011000011;
assign LUT_2[15350] = 32'b11111111111111110111110011100110;
assign LUT_2[15351] = 32'b11111111111111110100101011111111;
assign LUT_2[15352] = 32'b11111111111111101111001110011111;
assign LUT_2[15353] = 32'b11111111111111101100000110111000;
assign LUT_2[15354] = 32'b11111111111111110110000111011011;
assign LUT_2[15355] = 32'b11111111111111110010111111110100;
assign LUT_2[15356] = 32'b11111111111111101011101100000111;
assign LUT_2[15357] = 32'b11111111111111101000100100100000;
assign LUT_2[15358] = 32'b11111111111111110010100101000011;
assign LUT_2[15359] = 32'b11111111111111101111011101011100;
assign LUT_2[15360] = 32'b11111111111111111010111100001010;
assign LUT_2[15361] = 32'b11111111111111110111110100100011;
assign LUT_2[15362] = 32'b00000000000000000001110101000110;
assign LUT_2[15363] = 32'b11111111111111111110101101011111;
assign LUT_2[15364] = 32'b11111111111111110111011001110010;
assign LUT_2[15365] = 32'b11111111111111110100010010001011;
assign LUT_2[15366] = 32'b11111111111111111110010010101110;
assign LUT_2[15367] = 32'b11111111111111111011001011000111;
assign LUT_2[15368] = 32'b11111111111111110101101101100111;
assign LUT_2[15369] = 32'b11111111111111110010100110000000;
assign LUT_2[15370] = 32'b11111111111111111100100110100011;
assign LUT_2[15371] = 32'b11111111111111111001011110111100;
assign LUT_2[15372] = 32'b11111111111111110010001011001111;
assign LUT_2[15373] = 32'b11111111111111101111000011101000;
assign LUT_2[15374] = 32'b11111111111111111001000100001011;
assign LUT_2[15375] = 32'b11111111111111110101111100100100;
assign LUT_2[15376] = 32'b11111111111111110101100000010100;
assign LUT_2[15377] = 32'b11111111111111110010011000101101;
assign LUT_2[15378] = 32'b11111111111111111100011001010000;
assign LUT_2[15379] = 32'b11111111111111111001010001101001;
assign LUT_2[15380] = 32'b11111111111111110001111101111100;
assign LUT_2[15381] = 32'b11111111111111101110110110010101;
assign LUT_2[15382] = 32'b11111111111111111000110110111000;
assign LUT_2[15383] = 32'b11111111111111110101101111010001;
assign LUT_2[15384] = 32'b11111111111111110000010001110001;
assign LUT_2[15385] = 32'b11111111111111101101001010001010;
assign LUT_2[15386] = 32'b11111111111111110111001010101101;
assign LUT_2[15387] = 32'b11111111111111110100000011000110;
assign LUT_2[15388] = 32'b11111111111111101100101111011001;
assign LUT_2[15389] = 32'b11111111111111101001100111110010;
assign LUT_2[15390] = 32'b11111111111111110011101000010101;
assign LUT_2[15391] = 32'b11111111111111110000100000101110;
assign LUT_2[15392] = 32'b11111111111111111011010111110011;
assign LUT_2[15393] = 32'b11111111111111111000010000001100;
assign LUT_2[15394] = 32'b00000000000000000010010000101111;
assign LUT_2[15395] = 32'b11111111111111111111001001001000;
assign LUT_2[15396] = 32'b11111111111111110111110101011011;
assign LUT_2[15397] = 32'b11111111111111110100101101110100;
assign LUT_2[15398] = 32'b11111111111111111110101110010111;
assign LUT_2[15399] = 32'b11111111111111111011100110110000;
assign LUT_2[15400] = 32'b11111111111111110110001001010000;
assign LUT_2[15401] = 32'b11111111111111110011000001101001;
assign LUT_2[15402] = 32'b11111111111111111101000010001100;
assign LUT_2[15403] = 32'b11111111111111111001111010100101;
assign LUT_2[15404] = 32'b11111111111111110010100110111000;
assign LUT_2[15405] = 32'b11111111111111101111011111010001;
assign LUT_2[15406] = 32'b11111111111111111001011111110100;
assign LUT_2[15407] = 32'b11111111111111110110011000001101;
assign LUT_2[15408] = 32'b11111111111111110101111011111101;
assign LUT_2[15409] = 32'b11111111111111110010110100010110;
assign LUT_2[15410] = 32'b11111111111111111100110100111001;
assign LUT_2[15411] = 32'b11111111111111111001101101010010;
assign LUT_2[15412] = 32'b11111111111111110010011001100101;
assign LUT_2[15413] = 32'b11111111111111101111010001111110;
assign LUT_2[15414] = 32'b11111111111111111001010010100001;
assign LUT_2[15415] = 32'b11111111111111110110001010111010;
assign LUT_2[15416] = 32'b11111111111111110000101101011010;
assign LUT_2[15417] = 32'b11111111111111101101100101110011;
assign LUT_2[15418] = 32'b11111111111111110111100110010110;
assign LUT_2[15419] = 32'b11111111111111110100011110101111;
assign LUT_2[15420] = 32'b11111111111111101101001011000010;
assign LUT_2[15421] = 32'b11111111111111101010000011011011;
assign LUT_2[15422] = 32'b11111111111111110100000011111110;
assign LUT_2[15423] = 32'b11111111111111110000111100010111;
assign LUT_2[15424] = 32'b11111111111111110011000100101101;
assign LUT_2[15425] = 32'b11111111111111101111111101000110;
assign LUT_2[15426] = 32'b11111111111111111001111101101001;
assign LUT_2[15427] = 32'b11111111111111110110110110000010;
assign LUT_2[15428] = 32'b11111111111111101111100010010101;
assign LUT_2[15429] = 32'b11111111111111101100011010101110;
assign LUT_2[15430] = 32'b11111111111111110110011011010001;
assign LUT_2[15431] = 32'b11111111111111110011010011101010;
assign LUT_2[15432] = 32'b11111111111111101101110110001010;
assign LUT_2[15433] = 32'b11111111111111101010101110100011;
assign LUT_2[15434] = 32'b11111111111111110100101111000110;
assign LUT_2[15435] = 32'b11111111111111110001100111011111;
assign LUT_2[15436] = 32'b11111111111111101010010011110010;
assign LUT_2[15437] = 32'b11111111111111100111001100001011;
assign LUT_2[15438] = 32'b11111111111111110001001100101110;
assign LUT_2[15439] = 32'b11111111111111101110000101000111;
assign LUT_2[15440] = 32'b11111111111111101101101000110111;
assign LUT_2[15441] = 32'b11111111111111101010100001010000;
assign LUT_2[15442] = 32'b11111111111111110100100001110011;
assign LUT_2[15443] = 32'b11111111111111110001011010001100;
assign LUT_2[15444] = 32'b11111111111111101010000110011111;
assign LUT_2[15445] = 32'b11111111111111100110111110111000;
assign LUT_2[15446] = 32'b11111111111111110000111111011011;
assign LUT_2[15447] = 32'b11111111111111101101110111110100;
assign LUT_2[15448] = 32'b11111111111111101000011010010100;
assign LUT_2[15449] = 32'b11111111111111100101010010101101;
assign LUT_2[15450] = 32'b11111111111111101111010011010000;
assign LUT_2[15451] = 32'b11111111111111101100001011101001;
assign LUT_2[15452] = 32'b11111111111111100100110111111100;
assign LUT_2[15453] = 32'b11111111111111100001110000010101;
assign LUT_2[15454] = 32'b11111111111111101011110000111000;
assign LUT_2[15455] = 32'b11111111111111101000101001010001;
assign LUT_2[15456] = 32'b11111111111111110011100000010110;
assign LUT_2[15457] = 32'b11111111111111110000011000101111;
assign LUT_2[15458] = 32'b11111111111111111010011001010010;
assign LUT_2[15459] = 32'b11111111111111110111010001101011;
assign LUT_2[15460] = 32'b11111111111111101111111101111110;
assign LUT_2[15461] = 32'b11111111111111101100110110010111;
assign LUT_2[15462] = 32'b11111111111111110110110110111010;
assign LUT_2[15463] = 32'b11111111111111110011101111010011;
assign LUT_2[15464] = 32'b11111111111111101110010001110011;
assign LUT_2[15465] = 32'b11111111111111101011001010001100;
assign LUT_2[15466] = 32'b11111111111111110101001010101111;
assign LUT_2[15467] = 32'b11111111111111110010000011001000;
assign LUT_2[15468] = 32'b11111111111111101010101111011011;
assign LUT_2[15469] = 32'b11111111111111100111100111110100;
assign LUT_2[15470] = 32'b11111111111111110001101000010111;
assign LUT_2[15471] = 32'b11111111111111101110100000110000;
assign LUT_2[15472] = 32'b11111111111111101110000100100000;
assign LUT_2[15473] = 32'b11111111111111101010111100111001;
assign LUT_2[15474] = 32'b11111111111111110100111101011100;
assign LUT_2[15475] = 32'b11111111111111110001110101110101;
assign LUT_2[15476] = 32'b11111111111111101010100010001000;
assign LUT_2[15477] = 32'b11111111111111100111011010100001;
assign LUT_2[15478] = 32'b11111111111111110001011011000100;
assign LUT_2[15479] = 32'b11111111111111101110010011011101;
assign LUT_2[15480] = 32'b11111111111111101000110101111101;
assign LUT_2[15481] = 32'b11111111111111100101101110010110;
assign LUT_2[15482] = 32'b11111111111111101111101110111001;
assign LUT_2[15483] = 32'b11111111111111101100100111010010;
assign LUT_2[15484] = 32'b11111111111111100101010011100101;
assign LUT_2[15485] = 32'b11111111111111100010001011111110;
assign LUT_2[15486] = 32'b11111111111111101100001100100001;
assign LUT_2[15487] = 32'b11111111111111101001000100111010;
assign LUT_2[15488] = 32'b11111111111111111111010000011001;
assign LUT_2[15489] = 32'b11111111111111111100001000110010;
assign LUT_2[15490] = 32'b00000000000000000110001001010101;
assign LUT_2[15491] = 32'b00000000000000000011000001101110;
assign LUT_2[15492] = 32'b11111111111111111011101110000001;
assign LUT_2[15493] = 32'b11111111111111111000100110011010;
assign LUT_2[15494] = 32'b00000000000000000010100110111101;
assign LUT_2[15495] = 32'b11111111111111111111011111010110;
assign LUT_2[15496] = 32'b11111111111111111010000001110110;
assign LUT_2[15497] = 32'b11111111111111110110111010001111;
assign LUT_2[15498] = 32'b00000000000000000000111010110010;
assign LUT_2[15499] = 32'b11111111111111111101110011001011;
assign LUT_2[15500] = 32'b11111111111111110110011111011110;
assign LUT_2[15501] = 32'b11111111111111110011010111110111;
assign LUT_2[15502] = 32'b11111111111111111101011000011010;
assign LUT_2[15503] = 32'b11111111111111111010010000110011;
assign LUT_2[15504] = 32'b11111111111111111001110100100011;
assign LUT_2[15505] = 32'b11111111111111110110101100111100;
assign LUT_2[15506] = 32'b00000000000000000000101101011111;
assign LUT_2[15507] = 32'b11111111111111111101100101111000;
assign LUT_2[15508] = 32'b11111111111111110110010010001011;
assign LUT_2[15509] = 32'b11111111111111110011001010100100;
assign LUT_2[15510] = 32'b11111111111111111101001011000111;
assign LUT_2[15511] = 32'b11111111111111111010000011100000;
assign LUT_2[15512] = 32'b11111111111111110100100110000000;
assign LUT_2[15513] = 32'b11111111111111110001011110011001;
assign LUT_2[15514] = 32'b11111111111111111011011110111100;
assign LUT_2[15515] = 32'b11111111111111111000010111010101;
assign LUT_2[15516] = 32'b11111111111111110001000011101000;
assign LUT_2[15517] = 32'b11111111111111101101111100000001;
assign LUT_2[15518] = 32'b11111111111111110111111100100100;
assign LUT_2[15519] = 32'b11111111111111110100110100111101;
assign LUT_2[15520] = 32'b11111111111111111111101100000010;
assign LUT_2[15521] = 32'b11111111111111111100100100011011;
assign LUT_2[15522] = 32'b00000000000000000110100100111110;
assign LUT_2[15523] = 32'b00000000000000000011011101010111;
assign LUT_2[15524] = 32'b11111111111111111100001001101010;
assign LUT_2[15525] = 32'b11111111111111111001000010000011;
assign LUT_2[15526] = 32'b00000000000000000011000010100110;
assign LUT_2[15527] = 32'b11111111111111111111111010111111;
assign LUT_2[15528] = 32'b11111111111111111010011101011111;
assign LUT_2[15529] = 32'b11111111111111110111010101111000;
assign LUT_2[15530] = 32'b00000000000000000001010110011011;
assign LUT_2[15531] = 32'b11111111111111111110001110110100;
assign LUT_2[15532] = 32'b11111111111111110110111011000111;
assign LUT_2[15533] = 32'b11111111111111110011110011100000;
assign LUT_2[15534] = 32'b11111111111111111101110100000011;
assign LUT_2[15535] = 32'b11111111111111111010101100011100;
assign LUT_2[15536] = 32'b11111111111111111010010000001100;
assign LUT_2[15537] = 32'b11111111111111110111001000100101;
assign LUT_2[15538] = 32'b00000000000000000001001001001000;
assign LUT_2[15539] = 32'b11111111111111111110000001100001;
assign LUT_2[15540] = 32'b11111111111111110110101101110100;
assign LUT_2[15541] = 32'b11111111111111110011100110001101;
assign LUT_2[15542] = 32'b11111111111111111101100110110000;
assign LUT_2[15543] = 32'b11111111111111111010011111001001;
assign LUT_2[15544] = 32'b11111111111111110101000001101001;
assign LUT_2[15545] = 32'b11111111111111110001111010000010;
assign LUT_2[15546] = 32'b11111111111111111011111010100101;
assign LUT_2[15547] = 32'b11111111111111111000110010111110;
assign LUT_2[15548] = 32'b11111111111111110001011111010001;
assign LUT_2[15549] = 32'b11111111111111101110010111101010;
assign LUT_2[15550] = 32'b11111111111111111000011000001101;
assign LUT_2[15551] = 32'b11111111111111110101010000100110;
assign LUT_2[15552] = 32'b11111111111111110111011000111100;
assign LUT_2[15553] = 32'b11111111111111110100010001010101;
assign LUT_2[15554] = 32'b11111111111111111110010001111000;
assign LUT_2[15555] = 32'b11111111111111111011001010010001;
assign LUT_2[15556] = 32'b11111111111111110011110110100100;
assign LUT_2[15557] = 32'b11111111111111110000101110111101;
assign LUT_2[15558] = 32'b11111111111111111010101111100000;
assign LUT_2[15559] = 32'b11111111111111110111100111111001;
assign LUT_2[15560] = 32'b11111111111111110010001010011001;
assign LUT_2[15561] = 32'b11111111111111101111000010110010;
assign LUT_2[15562] = 32'b11111111111111111001000011010101;
assign LUT_2[15563] = 32'b11111111111111110101111011101110;
assign LUT_2[15564] = 32'b11111111111111101110101000000001;
assign LUT_2[15565] = 32'b11111111111111101011100000011010;
assign LUT_2[15566] = 32'b11111111111111110101100000111101;
assign LUT_2[15567] = 32'b11111111111111110010011001010110;
assign LUT_2[15568] = 32'b11111111111111110001111101000110;
assign LUT_2[15569] = 32'b11111111111111101110110101011111;
assign LUT_2[15570] = 32'b11111111111111111000110110000010;
assign LUT_2[15571] = 32'b11111111111111110101101110011011;
assign LUT_2[15572] = 32'b11111111111111101110011010101110;
assign LUT_2[15573] = 32'b11111111111111101011010011000111;
assign LUT_2[15574] = 32'b11111111111111110101010011101010;
assign LUT_2[15575] = 32'b11111111111111110010001100000011;
assign LUT_2[15576] = 32'b11111111111111101100101110100011;
assign LUT_2[15577] = 32'b11111111111111101001100110111100;
assign LUT_2[15578] = 32'b11111111111111110011100111011111;
assign LUT_2[15579] = 32'b11111111111111110000011111111000;
assign LUT_2[15580] = 32'b11111111111111101001001100001011;
assign LUT_2[15581] = 32'b11111111111111100110000100100100;
assign LUT_2[15582] = 32'b11111111111111110000000101000111;
assign LUT_2[15583] = 32'b11111111111111101100111101100000;
assign LUT_2[15584] = 32'b11111111111111110111110100100101;
assign LUT_2[15585] = 32'b11111111111111110100101100111110;
assign LUT_2[15586] = 32'b11111111111111111110101101100001;
assign LUT_2[15587] = 32'b11111111111111111011100101111010;
assign LUT_2[15588] = 32'b11111111111111110100010010001101;
assign LUT_2[15589] = 32'b11111111111111110001001010100110;
assign LUT_2[15590] = 32'b11111111111111111011001011001001;
assign LUT_2[15591] = 32'b11111111111111111000000011100010;
assign LUT_2[15592] = 32'b11111111111111110010100110000010;
assign LUT_2[15593] = 32'b11111111111111101111011110011011;
assign LUT_2[15594] = 32'b11111111111111111001011110111110;
assign LUT_2[15595] = 32'b11111111111111110110010111010111;
assign LUT_2[15596] = 32'b11111111111111101111000011101010;
assign LUT_2[15597] = 32'b11111111111111101011111100000011;
assign LUT_2[15598] = 32'b11111111111111110101111100100110;
assign LUT_2[15599] = 32'b11111111111111110010110100111111;
assign LUT_2[15600] = 32'b11111111111111110010011000101111;
assign LUT_2[15601] = 32'b11111111111111101111010001001000;
assign LUT_2[15602] = 32'b11111111111111111001010001101011;
assign LUT_2[15603] = 32'b11111111111111110110001010000100;
assign LUT_2[15604] = 32'b11111111111111101110110110010111;
assign LUT_2[15605] = 32'b11111111111111101011101110110000;
assign LUT_2[15606] = 32'b11111111111111110101101111010011;
assign LUT_2[15607] = 32'b11111111111111110010100111101100;
assign LUT_2[15608] = 32'b11111111111111101101001010001100;
assign LUT_2[15609] = 32'b11111111111111101010000010100101;
assign LUT_2[15610] = 32'b11111111111111110100000011001000;
assign LUT_2[15611] = 32'b11111111111111110000111011100001;
assign LUT_2[15612] = 32'b11111111111111101001100111110100;
assign LUT_2[15613] = 32'b11111111111111100110100000001101;
assign LUT_2[15614] = 32'b11111111111111110000100000110000;
assign LUT_2[15615] = 32'b11111111111111101101011001001001;
assign LUT_2[15616] = 32'b11111111111111111110111010110000;
assign LUT_2[15617] = 32'b11111111111111111011110011001001;
assign LUT_2[15618] = 32'b00000000000000000101110011101100;
assign LUT_2[15619] = 32'b00000000000000000010101100000101;
assign LUT_2[15620] = 32'b11111111111111111011011000011000;
assign LUT_2[15621] = 32'b11111111111111111000010000110001;
assign LUT_2[15622] = 32'b00000000000000000010010001010100;
assign LUT_2[15623] = 32'b11111111111111111111001001101101;
assign LUT_2[15624] = 32'b11111111111111111001101100001101;
assign LUT_2[15625] = 32'b11111111111111110110100100100110;
assign LUT_2[15626] = 32'b00000000000000000000100101001001;
assign LUT_2[15627] = 32'b11111111111111111101011101100010;
assign LUT_2[15628] = 32'b11111111111111110110001001110101;
assign LUT_2[15629] = 32'b11111111111111110011000010001110;
assign LUT_2[15630] = 32'b11111111111111111101000010110001;
assign LUT_2[15631] = 32'b11111111111111111001111011001010;
assign LUT_2[15632] = 32'b11111111111111111001011110111010;
assign LUT_2[15633] = 32'b11111111111111110110010111010011;
assign LUT_2[15634] = 32'b00000000000000000000010111110110;
assign LUT_2[15635] = 32'b11111111111111111101010000001111;
assign LUT_2[15636] = 32'b11111111111111110101111100100010;
assign LUT_2[15637] = 32'b11111111111111110010110100111011;
assign LUT_2[15638] = 32'b11111111111111111100110101011110;
assign LUT_2[15639] = 32'b11111111111111111001101101110111;
assign LUT_2[15640] = 32'b11111111111111110100010000010111;
assign LUT_2[15641] = 32'b11111111111111110001001000110000;
assign LUT_2[15642] = 32'b11111111111111111011001001010011;
assign LUT_2[15643] = 32'b11111111111111111000000001101100;
assign LUT_2[15644] = 32'b11111111111111110000101101111111;
assign LUT_2[15645] = 32'b11111111111111101101100110011000;
assign LUT_2[15646] = 32'b11111111111111110111100110111011;
assign LUT_2[15647] = 32'b11111111111111110100011111010100;
assign LUT_2[15648] = 32'b11111111111111111111010110011001;
assign LUT_2[15649] = 32'b11111111111111111100001110110010;
assign LUT_2[15650] = 32'b00000000000000000110001111010101;
assign LUT_2[15651] = 32'b00000000000000000011000111101110;
assign LUT_2[15652] = 32'b11111111111111111011110100000001;
assign LUT_2[15653] = 32'b11111111111111111000101100011010;
assign LUT_2[15654] = 32'b00000000000000000010101100111101;
assign LUT_2[15655] = 32'b11111111111111111111100101010110;
assign LUT_2[15656] = 32'b11111111111111111010000111110110;
assign LUT_2[15657] = 32'b11111111111111110111000000001111;
assign LUT_2[15658] = 32'b00000000000000000001000000110010;
assign LUT_2[15659] = 32'b11111111111111111101111001001011;
assign LUT_2[15660] = 32'b11111111111111110110100101011110;
assign LUT_2[15661] = 32'b11111111111111110011011101110111;
assign LUT_2[15662] = 32'b11111111111111111101011110011010;
assign LUT_2[15663] = 32'b11111111111111111010010110110011;
assign LUT_2[15664] = 32'b11111111111111111001111010100011;
assign LUT_2[15665] = 32'b11111111111111110110110010111100;
assign LUT_2[15666] = 32'b00000000000000000000110011011111;
assign LUT_2[15667] = 32'b11111111111111111101101011111000;
assign LUT_2[15668] = 32'b11111111111111110110011000001011;
assign LUT_2[15669] = 32'b11111111111111110011010000100100;
assign LUT_2[15670] = 32'b11111111111111111101010001000111;
assign LUT_2[15671] = 32'b11111111111111111010001001100000;
assign LUT_2[15672] = 32'b11111111111111110100101100000000;
assign LUT_2[15673] = 32'b11111111111111110001100100011001;
assign LUT_2[15674] = 32'b11111111111111111011100100111100;
assign LUT_2[15675] = 32'b11111111111111111000011101010101;
assign LUT_2[15676] = 32'b11111111111111110001001001101000;
assign LUT_2[15677] = 32'b11111111111111101110000010000001;
assign LUT_2[15678] = 32'b11111111111111111000000010100100;
assign LUT_2[15679] = 32'b11111111111111110100111010111101;
assign LUT_2[15680] = 32'b11111111111111110111000011010011;
assign LUT_2[15681] = 32'b11111111111111110011111011101100;
assign LUT_2[15682] = 32'b11111111111111111101111100001111;
assign LUT_2[15683] = 32'b11111111111111111010110100101000;
assign LUT_2[15684] = 32'b11111111111111110011100000111011;
assign LUT_2[15685] = 32'b11111111111111110000011001010100;
assign LUT_2[15686] = 32'b11111111111111111010011001110111;
assign LUT_2[15687] = 32'b11111111111111110111010010010000;
assign LUT_2[15688] = 32'b11111111111111110001110100110000;
assign LUT_2[15689] = 32'b11111111111111101110101101001001;
assign LUT_2[15690] = 32'b11111111111111111000101101101100;
assign LUT_2[15691] = 32'b11111111111111110101100110000101;
assign LUT_2[15692] = 32'b11111111111111101110010010011000;
assign LUT_2[15693] = 32'b11111111111111101011001010110001;
assign LUT_2[15694] = 32'b11111111111111110101001011010100;
assign LUT_2[15695] = 32'b11111111111111110010000011101101;
assign LUT_2[15696] = 32'b11111111111111110001100111011101;
assign LUT_2[15697] = 32'b11111111111111101110011111110110;
assign LUT_2[15698] = 32'b11111111111111111000100000011001;
assign LUT_2[15699] = 32'b11111111111111110101011000110010;
assign LUT_2[15700] = 32'b11111111111111101110000101000101;
assign LUT_2[15701] = 32'b11111111111111101010111101011110;
assign LUT_2[15702] = 32'b11111111111111110100111110000001;
assign LUT_2[15703] = 32'b11111111111111110001110110011010;
assign LUT_2[15704] = 32'b11111111111111101100011000111010;
assign LUT_2[15705] = 32'b11111111111111101001010001010011;
assign LUT_2[15706] = 32'b11111111111111110011010001110110;
assign LUT_2[15707] = 32'b11111111111111110000001010001111;
assign LUT_2[15708] = 32'b11111111111111101000110110100010;
assign LUT_2[15709] = 32'b11111111111111100101101110111011;
assign LUT_2[15710] = 32'b11111111111111101111101111011110;
assign LUT_2[15711] = 32'b11111111111111101100100111110111;
assign LUT_2[15712] = 32'b11111111111111110111011110111100;
assign LUT_2[15713] = 32'b11111111111111110100010111010101;
assign LUT_2[15714] = 32'b11111111111111111110010111111000;
assign LUT_2[15715] = 32'b11111111111111111011010000010001;
assign LUT_2[15716] = 32'b11111111111111110011111100100100;
assign LUT_2[15717] = 32'b11111111111111110000110100111101;
assign LUT_2[15718] = 32'b11111111111111111010110101100000;
assign LUT_2[15719] = 32'b11111111111111110111101101111001;
assign LUT_2[15720] = 32'b11111111111111110010010000011001;
assign LUT_2[15721] = 32'b11111111111111101111001000110010;
assign LUT_2[15722] = 32'b11111111111111111001001001010101;
assign LUT_2[15723] = 32'b11111111111111110110000001101110;
assign LUT_2[15724] = 32'b11111111111111101110101110000001;
assign LUT_2[15725] = 32'b11111111111111101011100110011010;
assign LUT_2[15726] = 32'b11111111111111110101100110111101;
assign LUT_2[15727] = 32'b11111111111111110010011111010110;
assign LUT_2[15728] = 32'b11111111111111110010000011000110;
assign LUT_2[15729] = 32'b11111111111111101110111011011111;
assign LUT_2[15730] = 32'b11111111111111111000111100000010;
assign LUT_2[15731] = 32'b11111111111111110101110100011011;
assign LUT_2[15732] = 32'b11111111111111101110100000101110;
assign LUT_2[15733] = 32'b11111111111111101011011001000111;
assign LUT_2[15734] = 32'b11111111111111110101011001101010;
assign LUT_2[15735] = 32'b11111111111111110010010010000011;
assign LUT_2[15736] = 32'b11111111111111101100110100100011;
assign LUT_2[15737] = 32'b11111111111111101001101100111100;
assign LUT_2[15738] = 32'b11111111111111110011101101011111;
assign LUT_2[15739] = 32'b11111111111111110000100101111000;
assign LUT_2[15740] = 32'b11111111111111101001010010001011;
assign LUT_2[15741] = 32'b11111111111111100110001010100100;
assign LUT_2[15742] = 32'b11111111111111110000001011000111;
assign LUT_2[15743] = 32'b11111111111111101101000011100000;
assign LUT_2[15744] = 32'b00000000000000000011001110111111;
assign LUT_2[15745] = 32'b00000000000000000000000111011000;
assign LUT_2[15746] = 32'b00000000000000001010000111111011;
assign LUT_2[15747] = 32'b00000000000000000111000000010100;
assign LUT_2[15748] = 32'b11111111111111111111101100100111;
assign LUT_2[15749] = 32'b11111111111111111100100101000000;
assign LUT_2[15750] = 32'b00000000000000000110100101100011;
assign LUT_2[15751] = 32'b00000000000000000011011101111100;
assign LUT_2[15752] = 32'b11111111111111111110000000011100;
assign LUT_2[15753] = 32'b11111111111111111010111000110101;
assign LUT_2[15754] = 32'b00000000000000000100111001011000;
assign LUT_2[15755] = 32'b00000000000000000001110001110001;
assign LUT_2[15756] = 32'b11111111111111111010011110000100;
assign LUT_2[15757] = 32'b11111111111111110111010110011101;
assign LUT_2[15758] = 32'b00000000000000000001010111000000;
assign LUT_2[15759] = 32'b11111111111111111110001111011001;
assign LUT_2[15760] = 32'b11111111111111111101110011001001;
assign LUT_2[15761] = 32'b11111111111111111010101011100010;
assign LUT_2[15762] = 32'b00000000000000000100101100000101;
assign LUT_2[15763] = 32'b00000000000000000001100100011110;
assign LUT_2[15764] = 32'b11111111111111111010010000110001;
assign LUT_2[15765] = 32'b11111111111111110111001001001010;
assign LUT_2[15766] = 32'b00000000000000000001001001101101;
assign LUT_2[15767] = 32'b11111111111111111110000010000110;
assign LUT_2[15768] = 32'b11111111111111111000100100100110;
assign LUT_2[15769] = 32'b11111111111111110101011100111111;
assign LUT_2[15770] = 32'b11111111111111111111011101100010;
assign LUT_2[15771] = 32'b11111111111111111100010101111011;
assign LUT_2[15772] = 32'b11111111111111110101000010001110;
assign LUT_2[15773] = 32'b11111111111111110001111010100111;
assign LUT_2[15774] = 32'b11111111111111111011111011001010;
assign LUT_2[15775] = 32'b11111111111111111000110011100011;
assign LUT_2[15776] = 32'b00000000000000000011101010101000;
assign LUT_2[15777] = 32'b00000000000000000000100011000001;
assign LUT_2[15778] = 32'b00000000000000001010100011100100;
assign LUT_2[15779] = 32'b00000000000000000111011011111101;
assign LUT_2[15780] = 32'b00000000000000000000001000010000;
assign LUT_2[15781] = 32'b11111111111111111101000000101001;
assign LUT_2[15782] = 32'b00000000000000000111000001001100;
assign LUT_2[15783] = 32'b00000000000000000011111001100101;
assign LUT_2[15784] = 32'b11111111111111111110011100000101;
assign LUT_2[15785] = 32'b11111111111111111011010100011110;
assign LUT_2[15786] = 32'b00000000000000000101010101000001;
assign LUT_2[15787] = 32'b00000000000000000010001101011010;
assign LUT_2[15788] = 32'b11111111111111111010111001101101;
assign LUT_2[15789] = 32'b11111111111111110111110010000110;
assign LUT_2[15790] = 32'b00000000000000000001110010101001;
assign LUT_2[15791] = 32'b11111111111111111110101011000010;
assign LUT_2[15792] = 32'b11111111111111111110001110110010;
assign LUT_2[15793] = 32'b11111111111111111011000111001011;
assign LUT_2[15794] = 32'b00000000000000000101000111101110;
assign LUT_2[15795] = 32'b00000000000000000010000000000111;
assign LUT_2[15796] = 32'b11111111111111111010101100011010;
assign LUT_2[15797] = 32'b11111111111111110111100100110011;
assign LUT_2[15798] = 32'b00000000000000000001100101010110;
assign LUT_2[15799] = 32'b11111111111111111110011101101111;
assign LUT_2[15800] = 32'b11111111111111111001000000001111;
assign LUT_2[15801] = 32'b11111111111111110101111000101000;
assign LUT_2[15802] = 32'b11111111111111111111111001001011;
assign LUT_2[15803] = 32'b11111111111111111100110001100100;
assign LUT_2[15804] = 32'b11111111111111110101011101110111;
assign LUT_2[15805] = 32'b11111111111111110010010110010000;
assign LUT_2[15806] = 32'b11111111111111111100010110110011;
assign LUT_2[15807] = 32'b11111111111111111001001111001100;
assign LUT_2[15808] = 32'b11111111111111111011010111100010;
assign LUT_2[15809] = 32'b11111111111111111000001111111011;
assign LUT_2[15810] = 32'b00000000000000000010010000011110;
assign LUT_2[15811] = 32'b11111111111111111111001000110111;
assign LUT_2[15812] = 32'b11111111111111110111110101001010;
assign LUT_2[15813] = 32'b11111111111111110100101101100011;
assign LUT_2[15814] = 32'b11111111111111111110101110000110;
assign LUT_2[15815] = 32'b11111111111111111011100110011111;
assign LUT_2[15816] = 32'b11111111111111110110001000111111;
assign LUT_2[15817] = 32'b11111111111111110011000001011000;
assign LUT_2[15818] = 32'b11111111111111111101000001111011;
assign LUT_2[15819] = 32'b11111111111111111001111010010100;
assign LUT_2[15820] = 32'b11111111111111110010100110100111;
assign LUT_2[15821] = 32'b11111111111111101111011111000000;
assign LUT_2[15822] = 32'b11111111111111111001011111100011;
assign LUT_2[15823] = 32'b11111111111111110110010111111100;
assign LUT_2[15824] = 32'b11111111111111110101111011101100;
assign LUT_2[15825] = 32'b11111111111111110010110100000101;
assign LUT_2[15826] = 32'b11111111111111111100110100101000;
assign LUT_2[15827] = 32'b11111111111111111001101101000001;
assign LUT_2[15828] = 32'b11111111111111110010011001010100;
assign LUT_2[15829] = 32'b11111111111111101111010001101101;
assign LUT_2[15830] = 32'b11111111111111111001010010010000;
assign LUT_2[15831] = 32'b11111111111111110110001010101001;
assign LUT_2[15832] = 32'b11111111111111110000101101001001;
assign LUT_2[15833] = 32'b11111111111111101101100101100010;
assign LUT_2[15834] = 32'b11111111111111110111100110000101;
assign LUT_2[15835] = 32'b11111111111111110100011110011110;
assign LUT_2[15836] = 32'b11111111111111101101001010110001;
assign LUT_2[15837] = 32'b11111111111111101010000011001010;
assign LUT_2[15838] = 32'b11111111111111110100000011101101;
assign LUT_2[15839] = 32'b11111111111111110000111100000110;
assign LUT_2[15840] = 32'b11111111111111111011110011001011;
assign LUT_2[15841] = 32'b11111111111111111000101011100100;
assign LUT_2[15842] = 32'b00000000000000000010101100000111;
assign LUT_2[15843] = 32'b11111111111111111111100100100000;
assign LUT_2[15844] = 32'b11111111111111111000010000110011;
assign LUT_2[15845] = 32'b11111111111111110101001001001100;
assign LUT_2[15846] = 32'b11111111111111111111001001101111;
assign LUT_2[15847] = 32'b11111111111111111100000010001000;
assign LUT_2[15848] = 32'b11111111111111110110100100101000;
assign LUT_2[15849] = 32'b11111111111111110011011101000001;
assign LUT_2[15850] = 32'b11111111111111111101011101100100;
assign LUT_2[15851] = 32'b11111111111111111010010101111101;
assign LUT_2[15852] = 32'b11111111111111110011000010010000;
assign LUT_2[15853] = 32'b11111111111111101111111010101001;
assign LUT_2[15854] = 32'b11111111111111111001111011001100;
assign LUT_2[15855] = 32'b11111111111111110110110011100101;
assign LUT_2[15856] = 32'b11111111111111110110010111010101;
assign LUT_2[15857] = 32'b11111111111111110011001111101110;
assign LUT_2[15858] = 32'b11111111111111111101010000010001;
assign LUT_2[15859] = 32'b11111111111111111010001000101010;
assign LUT_2[15860] = 32'b11111111111111110010110100111101;
assign LUT_2[15861] = 32'b11111111111111101111101101010110;
assign LUT_2[15862] = 32'b11111111111111111001101101111001;
assign LUT_2[15863] = 32'b11111111111111110110100110010010;
assign LUT_2[15864] = 32'b11111111111111110001001000110010;
assign LUT_2[15865] = 32'b11111111111111101110000001001011;
assign LUT_2[15866] = 32'b11111111111111111000000001101110;
assign LUT_2[15867] = 32'b11111111111111110100111010000111;
assign LUT_2[15868] = 32'b11111111111111101101100110011010;
assign LUT_2[15869] = 32'b11111111111111101010011110110011;
assign LUT_2[15870] = 32'b11111111111111110100011111010110;
assign LUT_2[15871] = 32'b11111111111111110001010111101111;
assign LUT_2[15872] = 32'b11111111111111111111101101111100;
assign LUT_2[15873] = 32'b11111111111111111100100110010101;
assign LUT_2[15874] = 32'b00000000000000000110100110111000;
assign LUT_2[15875] = 32'b00000000000000000011011111010001;
assign LUT_2[15876] = 32'b11111111111111111100001011100100;
assign LUT_2[15877] = 32'b11111111111111111001000011111101;
assign LUT_2[15878] = 32'b00000000000000000011000100100000;
assign LUT_2[15879] = 32'b11111111111111111111111100111001;
assign LUT_2[15880] = 32'b11111111111111111010011111011001;
assign LUT_2[15881] = 32'b11111111111111110111010111110010;
assign LUT_2[15882] = 32'b00000000000000000001011000010101;
assign LUT_2[15883] = 32'b11111111111111111110010000101110;
assign LUT_2[15884] = 32'b11111111111111110110111101000001;
assign LUT_2[15885] = 32'b11111111111111110011110101011010;
assign LUT_2[15886] = 32'b11111111111111111101110101111101;
assign LUT_2[15887] = 32'b11111111111111111010101110010110;
assign LUT_2[15888] = 32'b11111111111111111010010010000110;
assign LUT_2[15889] = 32'b11111111111111110111001010011111;
assign LUT_2[15890] = 32'b00000000000000000001001011000010;
assign LUT_2[15891] = 32'b11111111111111111110000011011011;
assign LUT_2[15892] = 32'b11111111111111110110101111101110;
assign LUT_2[15893] = 32'b11111111111111110011101000000111;
assign LUT_2[15894] = 32'b11111111111111111101101000101010;
assign LUT_2[15895] = 32'b11111111111111111010100001000011;
assign LUT_2[15896] = 32'b11111111111111110101000011100011;
assign LUT_2[15897] = 32'b11111111111111110001111011111100;
assign LUT_2[15898] = 32'b11111111111111111011111100011111;
assign LUT_2[15899] = 32'b11111111111111111000110100111000;
assign LUT_2[15900] = 32'b11111111111111110001100001001011;
assign LUT_2[15901] = 32'b11111111111111101110011001100100;
assign LUT_2[15902] = 32'b11111111111111111000011010000111;
assign LUT_2[15903] = 32'b11111111111111110101010010100000;
assign LUT_2[15904] = 32'b00000000000000000000001001100101;
assign LUT_2[15905] = 32'b11111111111111111101000001111110;
assign LUT_2[15906] = 32'b00000000000000000111000010100001;
assign LUT_2[15907] = 32'b00000000000000000011111010111010;
assign LUT_2[15908] = 32'b11111111111111111100100111001101;
assign LUT_2[15909] = 32'b11111111111111111001011111100110;
assign LUT_2[15910] = 32'b00000000000000000011100000001001;
assign LUT_2[15911] = 32'b00000000000000000000011000100010;
assign LUT_2[15912] = 32'b11111111111111111010111011000010;
assign LUT_2[15913] = 32'b11111111111111110111110011011011;
assign LUT_2[15914] = 32'b00000000000000000001110011111110;
assign LUT_2[15915] = 32'b11111111111111111110101100010111;
assign LUT_2[15916] = 32'b11111111111111110111011000101010;
assign LUT_2[15917] = 32'b11111111111111110100010001000011;
assign LUT_2[15918] = 32'b11111111111111111110010001100110;
assign LUT_2[15919] = 32'b11111111111111111011001001111111;
assign LUT_2[15920] = 32'b11111111111111111010101101101111;
assign LUT_2[15921] = 32'b11111111111111110111100110001000;
assign LUT_2[15922] = 32'b00000000000000000001100110101011;
assign LUT_2[15923] = 32'b11111111111111111110011111000100;
assign LUT_2[15924] = 32'b11111111111111110111001011010111;
assign LUT_2[15925] = 32'b11111111111111110100000011110000;
assign LUT_2[15926] = 32'b11111111111111111110000100010011;
assign LUT_2[15927] = 32'b11111111111111111010111100101100;
assign LUT_2[15928] = 32'b11111111111111110101011111001100;
assign LUT_2[15929] = 32'b11111111111111110010010111100101;
assign LUT_2[15930] = 32'b11111111111111111100011000001000;
assign LUT_2[15931] = 32'b11111111111111111001010000100001;
assign LUT_2[15932] = 32'b11111111111111110001111100110100;
assign LUT_2[15933] = 32'b11111111111111101110110101001101;
assign LUT_2[15934] = 32'b11111111111111111000110101110000;
assign LUT_2[15935] = 32'b11111111111111110101101110001001;
assign LUT_2[15936] = 32'b11111111111111110111110110011111;
assign LUT_2[15937] = 32'b11111111111111110100101110111000;
assign LUT_2[15938] = 32'b11111111111111111110101111011011;
assign LUT_2[15939] = 32'b11111111111111111011100111110100;
assign LUT_2[15940] = 32'b11111111111111110100010100000111;
assign LUT_2[15941] = 32'b11111111111111110001001100100000;
assign LUT_2[15942] = 32'b11111111111111111011001101000011;
assign LUT_2[15943] = 32'b11111111111111111000000101011100;
assign LUT_2[15944] = 32'b11111111111111110010100111111100;
assign LUT_2[15945] = 32'b11111111111111101111100000010101;
assign LUT_2[15946] = 32'b11111111111111111001100000111000;
assign LUT_2[15947] = 32'b11111111111111110110011001010001;
assign LUT_2[15948] = 32'b11111111111111101111000101100100;
assign LUT_2[15949] = 32'b11111111111111101011111101111101;
assign LUT_2[15950] = 32'b11111111111111110101111110100000;
assign LUT_2[15951] = 32'b11111111111111110010110110111001;
assign LUT_2[15952] = 32'b11111111111111110010011010101001;
assign LUT_2[15953] = 32'b11111111111111101111010011000010;
assign LUT_2[15954] = 32'b11111111111111111001010011100101;
assign LUT_2[15955] = 32'b11111111111111110110001011111110;
assign LUT_2[15956] = 32'b11111111111111101110111000010001;
assign LUT_2[15957] = 32'b11111111111111101011110000101010;
assign LUT_2[15958] = 32'b11111111111111110101110001001101;
assign LUT_2[15959] = 32'b11111111111111110010101001100110;
assign LUT_2[15960] = 32'b11111111111111101101001100000110;
assign LUT_2[15961] = 32'b11111111111111101010000100011111;
assign LUT_2[15962] = 32'b11111111111111110100000101000010;
assign LUT_2[15963] = 32'b11111111111111110000111101011011;
assign LUT_2[15964] = 32'b11111111111111101001101001101110;
assign LUT_2[15965] = 32'b11111111111111100110100010000111;
assign LUT_2[15966] = 32'b11111111111111110000100010101010;
assign LUT_2[15967] = 32'b11111111111111101101011011000011;
assign LUT_2[15968] = 32'b11111111111111111000010010001000;
assign LUT_2[15969] = 32'b11111111111111110101001010100001;
assign LUT_2[15970] = 32'b11111111111111111111001011000100;
assign LUT_2[15971] = 32'b11111111111111111100000011011101;
assign LUT_2[15972] = 32'b11111111111111110100101111110000;
assign LUT_2[15973] = 32'b11111111111111110001101000001001;
assign LUT_2[15974] = 32'b11111111111111111011101000101100;
assign LUT_2[15975] = 32'b11111111111111111000100001000101;
assign LUT_2[15976] = 32'b11111111111111110011000011100101;
assign LUT_2[15977] = 32'b11111111111111101111111011111110;
assign LUT_2[15978] = 32'b11111111111111111001111100100001;
assign LUT_2[15979] = 32'b11111111111111110110110100111010;
assign LUT_2[15980] = 32'b11111111111111101111100001001101;
assign LUT_2[15981] = 32'b11111111111111101100011001100110;
assign LUT_2[15982] = 32'b11111111111111110110011010001001;
assign LUT_2[15983] = 32'b11111111111111110011010010100010;
assign LUT_2[15984] = 32'b11111111111111110010110110010010;
assign LUT_2[15985] = 32'b11111111111111101111101110101011;
assign LUT_2[15986] = 32'b11111111111111111001101111001110;
assign LUT_2[15987] = 32'b11111111111111110110100111100111;
assign LUT_2[15988] = 32'b11111111111111101111010011111010;
assign LUT_2[15989] = 32'b11111111111111101100001100010011;
assign LUT_2[15990] = 32'b11111111111111110110001100110110;
assign LUT_2[15991] = 32'b11111111111111110011000101001111;
assign LUT_2[15992] = 32'b11111111111111101101100111101111;
assign LUT_2[15993] = 32'b11111111111111101010100000001000;
assign LUT_2[15994] = 32'b11111111111111110100100000101011;
assign LUT_2[15995] = 32'b11111111111111110001011001000100;
assign LUT_2[15996] = 32'b11111111111111101010000101010111;
assign LUT_2[15997] = 32'b11111111111111100110111101110000;
assign LUT_2[15998] = 32'b11111111111111110000111110010011;
assign LUT_2[15999] = 32'b11111111111111101101110110101100;
assign LUT_2[16000] = 32'b00000000000000000100000010001011;
assign LUT_2[16001] = 32'b00000000000000000000111010100100;
assign LUT_2[16002] = 32'b00000000000000001010111011000111;
assign LUT_2[16003] = 32'b00000000000000000111110011100000;
assign LUT_2[16004] = 32'b00000000000000000000011111110011;
assign LUT_2[16005] = 32'b11111111111111111101011000001100;
assign LUT_2[16006] = 32'b00000000000000000111011000101111;
assign LUT_2[16007] = 32'b00000000000000000100010001001000;
assign LUT_2[16008] = 32'b11111111111111111110110011101000;
assign LUT_2[16009] = 32'b11111111111111111011101100000001;
assign LUT_2[16010] = 32'b00000000000000000101101100100100;
assign LUT_2[16011] = 32'b00000000000000000010100100111101;
assign LUT_2[16012] = 32'b11111111111111111011010001010000;
assign LUT_2[16013] = 32'b11111111111111111000001001101001;
assign LUT_2[16014] = 32'b00000000000000000010001010001100;
assign LUT_2[16015] = 32'b11111111111111111111000010100101;
assign LUT_2[16016] = 32'b11111111111111111110100110010101;
assign LUT_2[16017] = 32'b11111111111111111011011110101110;
assign LUT_2[16018] = 32'b00000000000000000101011111010001;
assign LUT_2[16019] = 32'b00000000000000000010010111101010;
assign LUT_2[16020] = 32'b11111111111111111011000011111101;
assign LUT_2[16021] = 32'b11111111111111110111111100010110;
assign LUT_2[16022] = 32'b00000000000000000001111100111001;
assign LUT_2[16023] = 32'b11111111111111111110110101010010;
assign LUT_2[16024] = 32'b11111111111111111001010111110010;
assign LUT_2[16025] = 32'b11111111111111110110010000001011;
assign LUT_2[16026] = 32'b00000000000000000000010000101110;
assign LUT_2[16027] = 32'b11111111111111111101001001000111;
assign LUT_2[16028] = 32'b11111111111111110101110101011010;
assign LUT_2[16029] = 32'b11111111111111110010101101110011;
assign LUT_2[16030] = 32'b11111111111111111100101110010110;
assign LUT_2[16031] = 32'b11111111111111111001100110101111;
assign LUT_2[16032] = 32'b00000000000000000100011101110100;
assign LUT_2[16033] = 32'b00000000000000000001010110001101;
assign LUT_2[16034] = 32'b00000000000000001011010110110000;
assign LUT_2[16035] = 32'b00000000000000001000001111001001;
assign LUT_2[16036] = 32'b00000000000000000000111011011100;
assign LUT_2[16037] = 32'b11111111111111111101110011110101;
assign LUT_2[16038] = 32'b00000000000000000111110100011000;
assign LUT_2[16039] = 32'b00000000000000000100101100110001;
assign LUT_2[16040] = 32'b11111111111111111111001111010001;
assign LUT_2[16041] = 32'b11111111111111111100000111101010;
assign LUT_2[16042] = 32'b00000000000000000110001000001101;
assign LUT_2[16043] = 32'b00000000000000000011000000100110;
assign LUT_2[16044] = 32'b11111111111111111011101100111001;
assign LUT_2[16045] = 32'b11111111111111111000100101010010;
assign LUT_2[16046] = 32'b00000000000000000010100101110101;
assign LUT_2[16047] = 32'b11111111111111111111011110001110;
assign LUT_2[16048] = 32'b11111111111111111111000001111110;
assign LUT_2[16049] = 32'b11111111111111111011111010010111;
assign LUT_2[16050] = 32'b00000000000000000101111010111010;
assign LUT_2[16051] = 32'b00000000000000000010110011010011;
assign LUT_2[16052] = 32'b11111111111111111011011111100110;
assign LUT_2[16053] = 32'b11111111111111111000010111111111;
assign LUT_2[16054] = 32'b00000000000000000010011000100010;
assign LUT_2[16055] = 32'b11111111111111111111010000111011;
assign LUT_2[16056] = 32'b11111111111111111001110011011011;
assign LUT_2[16057] = 32'b11111111111111110110101011110100;
assign LUT_2[16058] = 32'b00000000000000000000101100010111;
assign LUT_2[16059] = 32'b11111111111111111101100100110000;
assign LUT_2[16060] = 32'b11111111111111110110010001000011;
assign LUT_2[16061] = 32'b11111111111111110011001001011100;
assign LUT_2[16062] = 32'b11111111111111111101001001111111;
assign LUT_2[16063] = 32'b11111111111111111010000010011000;
assign LUT_2[16064] = 32'b11111111111111111100001010101110;
assign LUT_2[16065] = 32'b11111111111111111001000011000111;
assign LUT_2[16066] = 32'b00000000000000000011000011101010;
assign LUT_2[16067] = 32'b11111111111111111111111100000011;
assign LUT_2[16068] = 32'b11111111111111111000101000010110;
assign LUT_2[16069] = 32'b11111111111111110101100000101111;
assign LUT_2[16070] = 32'b11111111111111111111100001010010;
assign LUT_2[16071] = 32'b11111111111111111100011001101011;
assign LUT_2[16072] = 32'b11111111111111110110111100001011;
assign LUT_2[16073] = 32'b11111111111111110011110100100100;
assign LUT_2[16074] = 32'b11111111111111111101110101000111;
assign LUT_2[16075] = 32'b11111111111111111010101101100000;
assign LUT_2[16076] = 32'b11111111111111110011011001110011;
assign LUT_2[16077] = 32'b11111111111111110000010010001100;
assign LUT_2[16078] = 32'b11111111111111111010010010101111;
assign LUT_2[16079] = 32'b11111111111111110111001011001000;
assign LUT_2[16080] = 32'b11111111111111110110101110111000;
assign LUT_2[16081] = 32'b11111111111111110011100111010001;
assign LUT_2[16082] = 32'b11111111111111111101100111110100;
assign LUT_2[16083] = 32'b11111111111111111010100000001101;
assign LUT_2[16084] = 32'b11111111111111110011001100100000;
assign LUT_2[16085] = 32'b11111111111111110000000100111001;
assign LUT_2[16086] = 32'b11111111111111111010000101011100;
assign LUT_2[16087] = 32'b11111111111111110110111101110101;
assign LUT_2[16088] = 32'b11111111111111110001100000010101;
assign LUT_2[16089] = 32'b11111111111111101110011000101110;
assign LUT_2[16090] = 32'b11111111111111111000011001010001;
assign LUT_2[16091] = 32'b11111111111111110101010001101010;
assign LUT_2[16092] = 32'b11111111111111101101111101111101;
assign LUT_2[16093] = 32'b11111111111111101010110110010110;
assign LUT_2[16094] = 32'b11111111111111110100110110111001;
assign LUT_2[16095] = 32'b11111111111111110001101111010010;
assign LUT_2[16096] = 32'b11111111111111111100100110010111;
assign LUT_2[16097] = 32'b11111111111111111001011110110000;
assign LUT_2[16098] = 32'b00000000000000000011011111010011;
assign LUT_2[16099] = 32'b00000000000000000000010111101100;
assign LUT_2[16100] = 32'b11111111111111111001000011111111;
assign LUT_2[16101] = 32'b11111111111111110101111100011000;
assign LUT_2[16102] = 32'b11111111111111111111111100111011;
assign LUT_2[16103] = 32'b11111111111111111100110101010100;
assign LUT_2[16104] = 32'b11111111111111110111010111110100;
assign LUT_2[16105] = 32'b11111111111111110100010000001101;
assign LUT_2[16106] = 32'b11111111111111111110010000110000;
assign LUT_2[16107] = 32'b11111111111111111011001001001001;
assign LUT_2[16108] = 32'b11111111111111110011110101011100;
assign LUT_2[16109] = 32'b11111111111111110000101101110101;
assign LUT_2[16110] = 32'b11111111111111111010101110011000;
assign LUT_2[16111] = 32'b11111111111111110111100110110001;
assign LUT_2[16112] = 32'b11111111111111110111001010100001;
assign LUT_2[16113] = 32'b11111111111111110100000010111010;
assign LUT_2[16114] = 32'b11111111111111111110000011011101;
assign LUT_2[16115] = 32'b11111111111111111010111011110110;
assign LUT_2[16116] = 32'b11111111111111110011101000001001;
assign LUT_2[16117] = 32'b11111111111111110000100000100010;
assign LUT_2[16118] = 32'b11111111111111111010100001000101;
assign LUT_2[16119] = 32'b11111111111111110111011001011110;
assign LUT_2[16120] = 32'b11111111111111110001111011111110;
assign LUT_2[16121] = 32'b11111111111111101110110100010111;
assign LUT_2[16122] = 32'b11111111111111111000110100111010;
assign LUT_2[16123] = 32'b11111111111111110101101101010011;
assign LUT_2[16124] = 32'b11111111111111101110011001100110;
assign LUT_2[16125] = 32'b11111111111111101011010001111111;
assign LUT_2[16126] = 32'b11111111111111110101010010100010;
assign LUT_2[16127] = 32'b11111111111111110010001010111011;
assign LUT_2[16128] = 32'b00000000000000000011101100100010;
assign LUT_2[16129] = 32'b00000000000000000000100100111011;
assign LUT_2[16130] = 32'b00000000000000001010100101011110;
assign LUT_2[16131] = 32'b00000000000000000111011101110111;
assign LUT_2[16132] = 32'b00000000000000000000001010001010;
assign LUT_2[16133] = 32'b11111111111111111101000010100011;
assign LUT_2[16134] = 32'b00000000000000000111000011000110;
assign LUT_2[16135] = 32'b00000000000000000011111011011111;
assign LUT_2[16136] = 32'b11111111111111111110011101111111;
assign LUT_2[16137] = 32'b11111111111111111011010110011000;
assign LUT_2[16138] = 32'b00000000000000000101010110111011;
assign LUT_2[16139] = 32'b00000000000000000010001111010100;
assign LUT_2[16140] = 32'b11111111111111111010111011100111;
assign LUT_2[16141] = 32'b11111111111111110111110100000000;
assign LUT_2[16142] = 32'b00000000000000000001110100100011;
assign LUT_2[16143] = 32'b11111111111111111110101100111100;
assign LUT_2[16144] = 32'b11111111111111111110010000101100;
assign LUT_2[16145] = 32'b11111111111111111011001001000101;
assign LUT_2[16146] = 32'b00000000000000000101001001101000;
assign LUT_2[16147] = 32'b00000000000000000010000010000001;
assign LUT_2[16148] = 32'b11111111111111111010101110010100;
assign LUT_2[16149] = 32'b11111111111111110111100110101101;
assign LUT_2[16150] = 32'b00000000000000000001100111010000;
assign LUT_2[16151] = 32'b11111111111111111110011111101001;
assign LUT_2[16152] = 32'b11111111111111111001000010001001;
assign LUT_2[16153] = 32'b11111111111111110101111010100010;
assign LUT_2[16154] = 32'b11111111111111111111111011000101;
assign LUT_2[16155] = 32'b11111111111111111100110011011110;
assign LUT_2[16156] = 32'b11111111111111110101011111110001;
assign LUT_2[16157] = 32'b11111111111111110010011000001010;
assign LUT_2[16158] = 32'b11111111111111111100011000101101;
assign LUT_2[16159] = 32'b11111111111111111001010001000110;
assign LUT_2[16160] = 32'b00000000000000000100001000001011;
assign LUT_2[16161] = 32'b00000000000000000001000000100100;
assign LUT_2[16162] = 32'b00000000000000001011000001000111;
assign LUT_2[16163] = 32'b00000000000000000111111001100000;
assign LUT_2[16164] = 32'b00000000000000000000100101110011;
assign LUT_2[16165] = 32'b11111111111111111101011110001100;
assign LUT_2[16166] = 32'b00000000000000000111011110101111;
assign LUT_2[16167] = 32'b00000000000000000100010111001000;
assign LUT_2[16168] = 32'b11111111111111111110111001101000;
assign LUT_2[16169] = 32'b11111111111111111011110010000001;
assign LUT_2[16170] = 32'b00000000000000000101110010100100;
assign LUT_2[16171] = 32'b00000000000000000010101010111101;
assign LUT_2[16172] = 32'b11111111111111111011010111010000;
assign LUT_2[16173] = 32'b11111111111111111000001111101001;
assign LUT_2[16174] = 32'b00000000000000000010010000001100;
assign LUT_2[16175] = 32'b11111111111111111111001000100101;
assign LUT_2[16176] = 32'b11111111111111111110101100010101;
assign LUT_2[16177] = 32'b11111111111111111011100100101110;
assign LUT_2[16178] = 32'b00000000000000000101100101010001;
assign LUT_2[16179] = 32'b00000000000000000010011101101010;
assign LUT_2[16180] = 32'b11111111111111111011001001111101;
assign LUT_2[16181] = 32'b11111111111111111000000010010110;
assign LUT_2[16182] = 32'b00000000000000000010000010111001;
assign LUT_2[16183] = 32'b11111111111111111110111011010010;
assign LUT_2[16184] = 32'b11111111111111111001011101110010;
assign LUT_2[16185] = 32'b11111111111111110110010110001011;
assign LUT_2[16186] = 32'b00000000000000000000010110101110;
assign LUT_2[16187] = 32'b11111111111111111101001111000111;
assign LUT_2[16188] = 32'b11111111111111110101111011011010;
assign LUT_2[16189] = 32'b11111111111111110010110011110011;
assign LUT_2[16190] = 32'b11111111111111111100110100010110;
assign LUT_2[16191] = 32'b11111111111111111001101100101111;
assign LUT_2[16192] = 32'b11111111111111111011110101000101;
assign LUT_2[16193] = 32'b11111111111111111000101101011110;
assign LUT_2[16194] = 32'b00000000000000000010101110000001;
assign LUT_2[16195] = 32'b11111111111111111111100110011010;
assign LUT_2[16196] = 32'b11111111111111111000010010101101;
assign LUT_2[16197] = 32'b11111111111111110101001011000110;
assign LUT_2[16198] = 32'b11111111111111111111001011101001;
assign LUT_2[16199] = 32'b11111111111111111100000100000010;
assign LUT_2[16200] = 32'b11111111111111110110100110100010;
assign LUT_2[16201] = 32'b11111111111111110011011110111011;
assign LUT_2[16202] = 32'b11111111111111111101011111011110;
assign LUT_2[16203] = 32'b11111111111111111010010111110111;
assign LUT_2[16204] = 32'b11111111111111110011000100001010;
assign LUT_2[16205] = 32'b11111111111111101111111100100011;
assign LUT_2[16206] = 32'b11111111111111111001111101000110;
assign LUT_2[16207] = 32'b11111111111111110110110101011111;
assign LUT_2[16208] = 32'b11111111111111110110011001001111;
assign LUT_2[16209] = 32'b11111111111111110011010001101000;
assign LUT_2[16210] = 32'b11111111111111111101010010001011;
assign LUT_2[16211] = 32'b11111111111111111010001010100100;
assign LUT_2[16212] = 32'b11111111111111110010110110110111;
assign LUT_2[16213] = 32'b11111111111111101111101111010000;
assign LUT_2[16214] = 32'b11111111111111111001101111110011;
assign LUT_2[16215] = 32'b11111111111111110110101000001100;
assign LUT_2[16216] = 32'b11111111111111110001001010101100;
assign LUT_2[16217] = 32'b11111111111111101110000011000101;
assign LUT_2[16218] = 32'b11111111111111111000000011101000;
assign LUT_2[16219] = 32'b11111111111111110100111100000001;
assign LUT_2[16220] = 32'b11111111111111101101101000010100;
assign LUT_2[16221] = 32'b11111111111111101010100000101101;
assign LUT_2[16222] = 32'b11111111111111110100100001010000;
assign LUT_2[16223] = 32'b11111111111111110001011001101001;
assign LUT_2[16224] = 32'b11111111111111111100010000101110;
assign LUT_2[16225] = 32'b11111111111111111001001001000111;
assign LUT_2[16226] = 32'b00000000000000000011001001101010;
assign LUT_2[16227] = 32'b00000000000000000000000010000011;
assign LUT_2[16228] = 32'b11111111111111111000101110010110;
assign LUT_2[16229] = 32'b11111111111111110101100110101111;
assign LUT_2[16230] = 32'b11111111111111111111100111010010;
assign LUT_2[16231] = 32'b11111111111111111100011111101011;
assign LUT_2[16232] = 32'b11111111111111110111000010001011;
assign LUT_2[16233] = 32'b11111111111111110011111010100100;
assign LUT_2[16234] = 32'b11111111111111111101111011000111;
assign LUT_2[16235] = 32'b11111111111111111010110011100000;
assign LUT_2[16236] = 32'b11111111111111110011011111110011;
assign LUT_2[16237] = 32'b11111111111111110000011000001100;
assign LUT_2[16238] = 32'b11111111111111111010011000101111;
assign LUT_2[16239] = 32'b11111111111111110111010001001000;
assign LUT_2[16240] = 32'b11111111111111110110110100111000;
assign LUT_2[16241] = 32'b11111111111111110011101101010001;
assign LUT_2[16242] = 32'b11111111111111111101101101110100;
assign LUT_2[16243] = 32'b11111111111111111010100110001101;
assign LUT_2[16244] = 32'b11111111111111110011010010100000;
assign LUT_2[16245] = 32'b11111111111111110000001010111001;
assign LUT_2[16246] = 32'b11111111111111111010001011011100;
assign LUT_2[16247] = 32'b11111111111111110111000011110101;
assign LUT_2[16248] = 32'b11111111111111110001100110010101;
assign LUT_2[16249] = 32'b11111111111111101110011110101110;
assign LUT_2[16250] = 32'b11111111111111111000011111010001;
assign LUT_2[16251] = 32'b11111111111111110101010111101010;
assign LUT_2[16252] = 32'b11111111111111101110000011111101;
assign LUT_2[16253] = 32'b11111111111111101010111100010110;
assign LUT_2[16254] = 32'b11111111111111110100111100111001;
assign LUT_2[16255] = 32'b11111111111111110001110101010010;
assign LUT_2[16256] = 32'b00000000000000001000000000110001;
assign LUT_2[16257] = 32'b00000000000000000100111001001010;
assign LUT_2[16258] = 32'b00000000000000001110111001101101;
assign LUT_2[16259] = 32'b00000000000000001011110010000110;
assign LUT_2[16260] = 32'b00000000000000000100011110011001;
assign LUT_2[16261] = 32'b00000000000000000001010110110010;
assign LUT_2[16262] = 32'b00000000000000001011010111010101;
assign LUT_2[16263] = 32'b00000000000000001000001111101110;
assign LUT_2[16264] = 32'b00000000000000000010110010001110;
assign LUT_2[16265] = 32'b11111111111111111111101010100111;
assign LUT_2[16266] = 32'b00000000000000001001101011001010;
assign LUT_2[16267] = 32'b00000000000000000110100011100011;
assign LUT_2[16268] = 32'b11111111111111111111001111110110;
assign LUT_2[16269] = 32'b11111111111111111100001000001111;
assign LUT_2[16270] = 32'b00000000000000000110001000110010;
assign LUT_2[16271] = 32'b00000000000000000011000001001011;
assign LUT_2[16272] = 32'b00000000000000000010100100111011;
assign LUT_2[16273] = 32'b11111111111111111111011101010100;
assign LUT_2[16274] = 32'b00000000000000001001011101110111;
assign LUT_2[16275] = 32'b00000000000000000110010110010000;
assign LUT_2[16276] = 32'b11111111111111111111000010100011;
assign LUT_2[16277] = 32'b11111111111111111011111010111100;
assign LUT_2[16278] = 32'b00000000000000000101111011011111;
assign LUT_2[16279] = 32'b00000000000000000010110011111000;
assign LUT_2[16280] = 32'b11111111111111111101010110011000;
assign LUT_2[16281] = 32'b11111111111111111010001110110001;
assign LUT_2[16282] = 32'b00000000000000000100001111010100;
assign LUT_2[16283] = 32'b00000000000000000001000111101101;
assign LUT_2[16284] = 32'b11111111111111111001110100000000;
assign LUT_2[16285] = 32'b11111111111111110110101100011001;
assign LUT_2[16286] = 32'b00000000000000000000101100111100;
assign LUT_2[16287] = 32'b11111111111111111101100101010101;
assign LUT_2[16288] = 32'b00000000000000001000011100011010;
assign LUT_2[16289] = 32'b00000000000000000101010100110011;
assign LUT_2[16290] = 32'b00000000000000001111010101010110;
assign LUT_2[16291] = 32'b00000000000000001100001101101111;
assign LUT_2[16292] = 32'b00000000000000000100111010000010;
assign LUT_2[16293] = 32'b00000000000000000001110010011011;
assign LUT_2[16294] = 32'b00000000000000001011110010111110;
assign LUT_2[16295] = 32'b00000000000000001000101011010111;
assign LUT_2[16296] = 32'b00000000000000000011001101110111;
assign LUT_2[16297] = 32'b00000000000000000000000110010000;
assign LUT_2[16298] = 32'b00000000000000001010000110110011;
assign LUT_2[16299] = 32'b00000000000000000110111111001100;
assign LUT_2[16300] = 32'b11111111111111111111101011011111;
assign LUT_2[16301] = 32'b11111111111111111100100011111000;
assign LUT_2[16302] = 32'b00000000000000000110100100011011;
assign LUT_2[16303] = 32'b00000000000000000011011100110100;
assign LUT_2[16304] = 32'b00000000000000000011000000100100;
assign LUT_2[16305] = 32'b11111111111111111111111000111101;
assign LUT_2[16306] = 32'b00000000000000001001111001100000;
assign LUT_2[16307] = 32'b00000000000000000110110001111001;
assign LUT_2[16308] = 32'b11111111111111111111011110001100;
assign LUT_2[16309] = 32'b11111111111111111100010110100101;
assign LUT_2[16310] = 32'b00000000000000000110010111001000;
assign LUT_2[16311] = 32'b00000000000000000011001111100001;
assign LUT_2[16312] = 32'b11111111111111111101110010000001;
assign LUT_2[16313] = 32'b11111111111111111010101010011010;
assign LUT_2[16314] = 32'b00000000000000000100101010111101;
assign LUT_2[16315] = 32'b00000000000000000001100011010110;
assign LUT_2[16316] = 32'b11111111111111111010001111101001;
assign LUT_2[16317] = 32'b11111111111111110111001000000010;
assign LUT_2[16318] = 32'b00000000000000000001001000100101;
assign LUT_2[16319] = 32'b11111111111111111110000000111110;
assign LUT_2[16320] = 32'b00000000000000000000001001010100;
assign LUT_2[16321] = 32'b11111111111111111101000001101101;
assign LUT_2[16322] = 32'b00000000000000000111000010010000;
assign LUT_2[16323] = 32'b00000000000000000011111010101001;
assign LUT_2[16324] = 32'b11111111111111111100100110111100;
assign LUT_2[16325] = 32'b11111111111111111001011111010101;
assign LUT_2[16326] = 32'b00000000000000000011011111111000;
assign LUT_2[16327] = 32'b00000000000000000000011000010001;
assign LUT_2[16328] = 32'b11111111111111111010111010110001;
assign LUT_2[16329] = 32'b11111111111111110111110011001010;
assign LUT_2[16330] = 32'b00000000000000000001110011101101;
assign LUT_2[16331] = 32'b11111111111111111110101100000110;
assign LUT_2[16332] = 32'b11111111111111110111011000011001;
assign LUT_2[16333] = 32'b11111111111111110100010000110010;
assign LUT_2[16334] = 32'b11111111111111111110010001010101;
assign LUT_2[16335] = 32'b11111111111111111011001001101110;
assign LUT_2[16336] = 32'b11111111111111111010101101011110;
assign LUT_2[16337] = 32'b11111111111111110111100101110111;
assign LUT_2[16338] = 32'b00000000000000000001100110011010;
assign LUT_2[16339] = 32'b11111111111111111110011110110011;
assign LUT_2[16340] = 32'b11111111111111110111001011000110;
assign LUT_2[16341] = 32'b11111111111111110100000011011111;
assign LUT_2[16342] = 32'b11111111111111111110000100000010;
assign LUT_2[16343] = 32'b11111111111111111010111100011011;
assign LUT_2[16344] = 32'b11111111111111110101011110111011;
assign LUT_2[16345] = 32'b11111111111111110010010111010100;
assign LUT_2[16346] = 32'b11111111111111111100010111110111;
assign LUT_2[16347] = 32'b11111111111111111001010000010000;
assign LUT_2[16348] = 32'b11111111111111110001111100100011;
assign LUT_2[16349] = 32'b11111111111111101110110100111100;
assign LUT_2[16350] = 32'b11111111111111111000110101011111;
assign LUT_2[16351] = 32'b11111111111111110101101101111000;
assign LUT_2[16352] = 32'b00000000000000000000100100111101;
assign LUT_2[16353] = 32'b11111111111111111101011101010110;
assign LUT_2[16354] = 32'b00000000000000000111011101111001;
assign LUT_2[16355] = 32'b00000000000000000100010110010010;
assign LUT_2[16356] = 32'b11111111111111111101000010100101;
assign LUT_2[16357] = 32'b11111111111111111001111010111110;
assign LUT_2[16358] = 32'b00000000000000000011111011100001;
assign LUT_2[16359] = 32'b00000000000000000000110011111010;
assign LUT_2[16360] = 32'b11111111111111111011010110011010;
assign LUT_2[16361] = 32'b11111111111111111000001110110011;
assign LUT_2[16362] = 32'b00000000000000000010001111010110;
assign LUT_2[16363] = 32'b11111111111111111111000111101111;
assign LUT_2[16364] = 32'b11111111111111110111110100000010;
assign LUT_2[16365] = 32'b11111111111111110100101100011011;
assign LUT_2[16366] = 32'b11111111111111111110101100111110;
assign LUT_2[16367] = 32'b11111111111111111011100101010111;
assign LUT_2[16368] = 32'b11111111111111111011001001000111;
assign LUT_2[16369] = 32'b11111111111111111000000001100000;
assign LUT_2[16370] = 32'b00000000000000000010000010000011;
assign LUT_2[16371] = 32'b11111111111111111110111010011100;
assign LUT_2[16372] = 32'b11111111111111110111100110101111;
assign LUT_2[16373] = 32'b11111111111111110100011111001000;
assign LUT_2[16374] = 32'b11111111111111111110011111101011;
assign LUT_2[16375] = 32'b11111111111111111011011000000100;
assign LUT_2[16376] = 32'b11111111111111110101111010100100;
assign LUT_2[16377] = 32'b11111111111111110010110010111101;
assign LUT_2[16378] = 32'b11111111111111111100110011100000;
assign LUT_2[16379] = 32'b11111111111111111001101011111001;
assign LUT_2[16380] = 32'b11111111111111110010011000001100;
assign LUT_2[16381] = 32'b11111111111111101111010000100101;
assign LUT_2[16382] = 32'b11111111111111111001010001001000;
assign LUT_2[16383] = 32'b11111111111111110110001001100001;
assign LUT_2[16384] = 32'b11111111111111111011101001110011;
assign LUT_2[16385] = 32'b11111111111111111000100010001100;
assign LUT_2[16386] = 32'b00000000000000000010100010101111;
assign LUT_2[16387] = 32'b11111111111111111111011011001000;
assign LUT_2[16388] = 32'b11111111111111111000000111011011;
assign LUT_2[16389] = 32'b11111111111111110100111111110100;
assign LUT_2[16390] = 32'b11111111111111111111000000010111;
assign LUT_2[16391] = 32'b11111111111111111011111000110000;
assign LUT_2[16392] = 32'b11111111111111110110011011010000;
assign LUT_2[16393] = 32'b11111111111111110011010011101001;
assign LUT_2[16394] = 32'b11111111111111111101010100001100;
assign LUT_2[16395] = 32'b11111111111111111010001100100101;
assign LUT_2[16396] = 32'b11111111111111110010111000111000;
assign LUT_2[16397] = 32'b11111111111111101111110001010001;
assign LUT_2[16398] = 32'b11111111111111111001110001110100;
assign LUT_2[16399] = 32'b11111111111111110110101010001101;
assign LUT_2[16400] = 32'b11111111111111110110001101111101;
assign LUT_2[16401] = 32'b11111111111111110011000110010110;
assign LUT_2[16402] = 32'b11111111111111111101000110111001;
assign LUT_2[16403] = 32'b11111111111111111001111111010010;
assign LUT_2[16404] = 32'b11111111111111110010101011100101;
assign LUT_2[16405] = 32'b11111111111111101111100011111110;
assign LUT_2[16406] = 32'b11111111111111111001100100100001;
assign LUT_2[16407] = 32'b11111111111111110110011100111010;
assign LUT_2[16408] = 32'b11111111111111110000111111011010;
assign LUT_2[16409] = 32'b11111111111111101101110111110011;
assign LUT_2[16410] = 32'b11111111111111110111111000010110;
assign LUT_2[16411] = 32'b11111111111111110100110000101111;
assign LUT_2[16412] = 32'b11111111111111101101011101000010;
assign LUT_2[16413] = 32'b11111111111111101010010101011011;
assign LUT_2[16414] = 32'b11111111111111110100010101111110;
assign LUT_2[16415] = 32'b11111111111111110001001110010111;
assign LUT_2[16416] = 32'b11111111111111111100000101011100;
assign LUT_2[16417] = 32'b11111111111111111000111101110101;
assign LUT_2[16418] = 32'b00000000000000000010111110011000;
assign LUT_2[16419] = 32'b11111111111111111111110110110001;
assign LUT_2[16420] = 32'b11111111111111111000100011000100;
assign LUT_2[16421] = 32'b11111111111111110101011011011101;
assign LUT_2[16422] = 32'b11111111111111111111011100000000;
assign LUT_2[16423] = 32'b11111111111111111100010100011001;
assign LUT_2[16424] = 32'b11111111111111110110110110111001;
assign LUT_2[16425] = 32'b11111111111111110011101111010010;
assign LUT_2[16426] = 32'b11111111111111111101101111110101;
assign LUT_2[16427] = 32'b11111111111111111010101000001110;
assign LUT_2[16428] = 32'b11111111111111110011010100100001;
assign LUT_2[16429] = 32'b11111111111111110000001100111010;
assign LUT_2[16430] = 32'b11111111111111111010001101011101;
assign LUT_2[16431] = 32'b11111111111111110111000101110110;
assign LUT_2[16432] = 32'b11111111111111110110101001100110;
assign LUT_2[16433] = 32'b11111111111111110011100001111111;
assign LUT_2[16434] = 32'b11111111111111111101100010100010;
assign LUT_2[16435] = 32'b11111111111111111010011010111011;
assign LUT_2[16436] = 32'b11111111111111110011000111001110;
assign LUT_2[16437] = 32'b11111111111111101111111111100111;
assign LUT_2[16438] = 32'b11111111111111111010000000001010;
assign LUT_2[16439] = 32'b11111111111111110110111000100011;
assign LUT_2[16440] = 32'b11111111111111110001011011000011;
assign LUT_2[16441] = 32'b11111111111111101110010011011100;
assign LUT_2[16442] = 32'b11111111111111111000010011111111;
assign LUT_2[16443] = 32'b11111111111111110101001100011000;
assign LUT_2[16444] = 32'b11111111111111101101111000101011;
assign LUT_2[16445] = 32'b11111111111111101010110001000100;
assign LUT_2[16446] = 32'b11111111111111110100110001100111;
assign LUT_2[16447] = 32'b11111111111111110001101010000000;
assign LUT_2[16448] = 32'b11111111111111110011110010010110;
assign LUT_2[16449] = 32'b11111111111111110000101010101111;
assign LUT_2[16450] = 32'b11111111111111111010101011010010;
assign LUT_2[16451] = 32'b11111111111111110111100011101011;
assign LUT_2[16452] = 32'b11111111111111110000001111111110;
assign LUT_2[16453] = 32'b11111111111111101101001000010111;
assign LUT_2[16454] = 32'b11111111111111110111001000111010;
assign LUT_2[16455] = 32'b11111111111111110100000001010011;
assign LUT_2[16456] = 32'b11111111111111101110100011110011;
assign LUT_2[16457] = 32'b11111111111111101011011100001100;
assign LUT_2[16458] = 32'b11111111111111110101011100101111;
assign LUT_2[16459] = 32'b11111111111111110010010101001000;
assign LUT_2[16460] = 32'b11111111111111101011000001011011;
assign LUT_2[16461] = 32'b11111111111111100111111001110100;
assign LUT_2[16462] = 32'b11111111111111110001111010010111;
assign LUT_2[16463] = 32'b11111111111111101110110010110000;
assign LUT_2[16464] = 32'b11111111111111101110010110100000;
assign LUT_2[16465] = 32'b11111111111111101011001110111001;
assign LUT_2[16466] = 32'b11111111111111110101001111011100;
assign LUT_2[16467] = 32'b11111111111111110010000111110101;
assign LUT_2[16468] = 32'b11111111111111101010110100001000;
assign LUT_2[16469] = 32'b11111111111111100111101100100001;
assign LUT_2[16470] = 32'b11111111111111110001101101000100;
assign LUT_2[16471] = 32'b11111111111111101110100101011101;
assign LUT_2[16472] = 32'b11111111111111101001000111111101;
assign LUT_2[16473] = 32'b11111111111111100110000000010110;
assign LUT_2[16474] = 32'b11111111111111110000000000111001;
assign LUT_2[16475] = 32'b11111111111111101100111001010010;
assign LUT_2[16476] = 32'b11111111111111100101100101100101;
assign LUT_2[16477] = 32'b11111111111111100010011101111110;
assign LUT_2[16478] = 32'b11111111111111101100011110100001;
assign LUT_2[16479] = 32'b11111111111111101001010110111010;
assign LUT_2[16480] = 32'b11111111111111110100001101111111;
assign LUT_2[16481] = 32'b11111111111111110001000110011000;
assign LUT_2[16482] = 32'b11111111111111111011000110111011;
assign LUT_2[16483] = 32'b11111111111111110111111111010100;
assign LUT_2[16484] = 32'b11111111111111110000101011100111;
assign LUT_2[16485] = 32'b11111111111111101101100100000000;
assign LUT_2[16486] = 32'b11111111111111110111100100100011;
assign LUT_2[16487] = 32'b11111111111111110100011100111100;
assign LUT_2[16488] = 32'b11111111111111101110111111011100;
assign LUT_2[16489] = 32'b11111111111111101011110111110101;
assign LUT_2[16490] = 32'b11111111111111110101111000011000;
assign LUT_2[16491] = 32'b11111111111111110010110000110001;
assign LUT_2[16492] = 32'b11111111111111101011011101000100;
assign LUT_2[16493] = 32'b11111111111111101000010101011101;
assign LUT_2[16494] = 32'b11111111111111110010010110000000;
assign LUT_2[16495] = 32'b11111111111111101111001110011001;
assign LUT_2[16496] = 32'b11111111111111101110110010001001;
assign LUT_2[16497] = 32'b11111111111111101011101010100010;
assign LUT_2[16498] = 32'b11111111111111110101101011000101;
assign LUT_2[16499] = 32'b11111111111111110010100011011110;
assign LUT_2[16500] = 32'b11111111111111101011001111110001;
assign LUT_2[16501] = 32'b11111111111111101000001000001010;
assign LUT_2[16502] = 32'b11111111111111110010001000101101;
assign LUT_2[16503] = 32'b11111111111111101111000001000110;
assign LUT_2[16504] = 32'b11111111111111101001100011100110;
assign LUT_2[16505] = 32'b11111111111111100110011011111111;
assign LUT_2[16506] = 32'b11111111111111110000011100100010;
assign LUT_2[16507] = 32'b11111111111111101101010100111011;
assign LUT_2[16508] = 32'b11111111111111100110000001001110;
assign LUT_2[16509] = 32'b11111111111111100010111001100111;
assign LUT_2[16510] = 32'b11111111111111101100111010001010;
assign LUT_2[16511] = 32'b11111111111111101001110010100011;
assign LUT_2[16512] = 32'b11111111111111111111111110000010;
assign LUT_2[16513] = 32'b11111111111111111100110110011011;
assign LUT_2[16514] = 32'b00000000000000000110110110111110;
assign LUT_2[16515] = 32'b00000000000000000011101111010111;
assign LUT_2[16516] = 32'b11111111111111111100011011101010;
assign LUT_2[16517] = 32'b11111111111111111001010100000011;
assign LUT_2[16518] = 32'b00000000000000000011010100100110;
assign LUT_2[16519] = 32'b00000000000000000000001100111111;
assign LUT_2[16520] = 32'b11111111111111111010101111011111;
assign LUT_2[16521] = 32'b11111111111111110111100111111000;
assign LUT_2[16522] = 32'b00000000000000000001101000011011;
assign LUT_2[16523] = 32'b11111111111111111110100000110100;
assign LUT_2[16524] = 32'b11111111111111110111001101000111;
assign LUT_2[16525] = 32'b11111111111111110100000101100000;
assign LUT_2[16526] = 32'b11111111111111111110000110000011;
assign LUT_2[16527] = 32'b11111111111111111010111110011100;
assign LUT_2[16528] = 32'b11111111111111111010100010001100;
assign LUT_2[16529] = 32'b11111111111111110111011010100101;
assign LUT_2[16530] = 32'b00000000000000000001011011001000;
assign LUT_2[16531] = 32'b11111111111111111110010011100001;
assign LUT_2[16532] = 32'b11111111111111110110111111110100;
assign LUT_2[16533] = 32'b11111111111111110011111000001101;
assign LUT_2[16534] = 32'b11111111111111111101111000110000;
assign LUT_2[16535] = 32'b11111111111111111010110001001001;
assign LUT_2[16536] = 32'b11111111111111110101010011101001;
assign LUT_2[16537] = 32'b11111111111111110010001100000010;
assign LUT_2[16538] = 32'b11111111111111111100001100100101;
assign LUT_2[16539] = 32'b11111111111111111001000100111110;
assign LUT_2[16540] = 32'b11111111111111110001110001010001;
assign LUT_2[16541] = 32'b11111111111111101110101001101010;
assign LUT_2[16542] = 32'b11111111111111111000101010001101;
assign LUT_2[16543] = 32'b11111111111111110101100010100110;
assign LUT_2[16544] = 32'b00000000000000000000011001101011;
assign LUT_2[16545] = 32'b11111111111111111101010010000100;
assign LUT_2[16546] = 32'b00000000000000000111010010100111;
assign LUT_2[16547] = 32'b00000000000000000100001011000000;
assign LUT_2[16548] = 32'b11111111111111111100110111010011;
assign LUT_2[16549] = 32'b11111111111111111001101111101100;
assign LUT_2[16550] = 32'b00000000000000000011110000001111;
assign LUT_2[16551] = 32'b00000000000000000000101000101000;
assign LUT_2[16552] = 32'b11111111111111111011001011001000;
assign LUT_2[16553] = 32'b11111111111111111000000011100001;
assign LUT_2[16554] = 32'b00000000000000000010000100000100;
assign LUT_2[16555] = 32'b11111111111111111110111100011101;
assign LUT_2[16556] = 32'b11111111111111110111101000110000;
assign LUT_2[16557] = 32'b11111111111111110100100001001001;
assign LUT_2[16558] = 32'b11111111111111111110100001101100;
assign LUT_2[16559] = 32'b11111111111111111011011010000101;
assign LUT_2[16560] = 32'b11111111111111111010111101110101;
assign LUT_2[16561] = 32'b11111111111111110111110110001110;
assign LUT_2[16562] = 32'b00000000000000000001110110110001;
assign LUT_2[16563] = 32'b11111111111111111110101111001010;
assign LUT_2[16564] = 32'b11111111111111110111011011011101;
assign LUT_2[16565] = 32'b11111111111111110100010011110110;
assign LUT_2[16566] = 32'b11111111111111111110010100011001;
assign LUT_2[16567] = 32'b11111111111111111011001100110010;
assign LUT_2[16568] = 32'b11111111111111110101101111010010;
assign LUT_2[16569] = 32'b11111111111111110010100111101011;
assign LUT_2[16570] = 32'b11111111111111111100101000001110;
assign LUT_2[16571] = 32'b11111111111111111001100000100111;
assign LUT_2[16572] = 32'b11111111111111110010001100111010;
assign LUT_2[16573] = 32'b11111111111111101111000101010011;
assign LUT_2[16574] = 32'b11111111111111111001000101110110;
assign LUT_2[16575] = 32'b11111111111111110101111110001111;
assign LUT_2[16576] = 32'b11111111111111111000000110100101;
assign LUT_2[16577] = 32'b11111111111111110100111110111110;
assign LUT_2[16578] = 32'b11111111111111111110111111100001;
assign LUT_2[16579] = 32'b11111111111111111011110111111010;
assign LUT_2[16580] = 32'b11111111111111110100100100001101;
assign LUT_2[16581] = 32'b11111111111111110001011100100110;
assign LUT_2[16582] = 32'b11111111111111111011011101001001;
assign LUT_2[16583] = 32'b11111111111111111000010101100010;
assign LUT_2[16584] = 32'b11111111111111110010111000000010;
assign LUT_2[16585] = 32'b11111111111111101111110000011011;
assign LUT_2[16586] = 32'b11111111111111111001110000111110;
assign LUT_2[16587] = 32'b11111111111111110110101001010111;
assign LUT_2[16588] = 32'b11111111111111101111010101101010;
assign LUT_2[16589] = 32'b11111111111111101100001110000011;
assign LUT_2[16590] = 32'b11111111111111110110001110100110;
assign LUT_2[16591] = 32'b11111111111111110011000110111111;
assign LUT_2[16592] = 32'b11111111111111110010101010101111;
assign LUT_2[16593] = 32'b11111111111111101111100011001000;
assign LUT_2[16594] = 32'b11111111111111111001100011101011;
assign LUT_2[16595] = 32'b11111111111111110110011100000100;
assign LUT_2[16596] = 32'b11111111111111101111001000010111;
assign LUT_2[16597] = 32'b11111111111111101100000000110000;
assign LUT_2[16598] = 32'b11111111111111110110000001010011;
assign LUT_2[16599] = 32'b11111111111111110010111001101100;
assign LUT_2[16600] = 32'b11111111111111101101011100001100;
assign LUT_2[16601] = 32'b11111111111111101010010100100101;
assign LUT_2[16602] = 32'b11111111111111110100010101001000;
assign LUT_2[16603] = 32'b11111111111111110001001101100001;
assign LUT_2[16604] = 32'b11111111111111101001111001110100;
assign LUT_2[16605] = 32'b11111111111111100110110010001101;
assign LUT_2[16606] = 32'b11111111111111110000110010110000;
assign LUT_2[16607] = 32'b11111111111111101101101011001001;
assign LUT_2[16608] = 32'b11111111111111111000100010001110;
assign LUT_2[16609] = 32'b11111111111111110101011010100111;
assign LUT_2[16610] = 32'b11111111111111111111011011001010;
assign LUT_2[16611] = 32'b11111111111111111100010011100011;
assign LUT_2[16612] = 32'b11111111111111110100111111110110;
assign LUT_2[16613] = 32'b11111111111111110001111000001111;
assign LUT_2[16614] = 32'b11111111111111111011111000110010;
assign LUT_2[16615] = 32'b11111111111111111000110001001011;
assign LUT_2[16616] = 32'b11111111111111110011010011101011;
assign LUT_2[16617] = 32'b11111111111111110000001100000100;
assign LUT_2[16618] = 32'b11111111111111111010001100100111;
assign LUT_2[16619] = 32'b11111111111111110111000101000000;
assign LUT_2[16620] = 32'b11111111111111101111110001010011;
assign LUT_2[16621] = 32'b11111111111111101100101001101100;
assign LUT_2[16622] = 32'b11111111111111110110101010001111;
assign LUT_2[16623] = 32'b11111111111111110011100010101000;
assign LUT_2[16624] = 32'b11111111111111110011000110011000;
assign LUT_2[16625] = 32'b11111111111111101111111110110001;
assign LUT_2[16626] = 32'b11111111111111111001111111010100;
assign LUT_2[16627] = 32'b11111111111111110110110111101101;
assign LUT_2[16628] = 32'b11111111111111101111100100000000;
assign LUT_2[16629] = 32'b11111111111111101100011100011001;
assign LUT_2[16630] = 32'b11111111111111110110011100111100;
assign LUT_2[16631] = 32'b11111111111111110011010101010101;
assign LUT_2[16632] = 32'b11111111111111101101110111110101;
assign LUT_2[16633] = 32'b11111111111111101010110000001110;
assign LUT_2[16634] = 32'b11111111111111110100110000110001;
assign LUT_2[16635] = 32'b11111111111111110001101001001010;
assign LUT_2[16636] = 32'b11111111111111101010010101011101;
assign LUT_2[16637] = 32'b11111111111111100111001101110110;
assign LUT_2[16638] = 32'b11111111111111110001001110011001;
assign LUT_2[16639] = 32'b11111111111111101110000110110010;
assign LUT_2[16640] = 32'b11111111111111111111101000011001;
assign LUT_2[16641] = 32'b11111111111111111100100000110010;
assign LUT_2[16642] = 32'b00000000000000000110100001010101;
assign LUT_2[16643] = 32'b00000000000000000011011001101110;
assign LUT_2[16644] = 32'b11111111111111111100000110000001;
assign LUT_2[16645] = 32'b11111111111111111000111110011010;
assign LUT_2[16646] = 32'b00000000000000000010111110111101;
assign LUT_2[16647] = 32'b11111111111111111111110111010110;
assign LUT_2[16648] = 32'b11111111111111111010011001110110;
assign LUT_2[16649] = 32'b11111111111111110111010010001111;
assign LUT_2[16650] = 32'b00000000000000000001010010110010;
assign LUT_2[16651] = 32'b11111111111111111110001011001011;
assign LUT_2[16652] = 32'b11111111111111110110110111011110;
assign LUT_2[16653] = 32'b11111111111111110011101111110111;
assign LUT_2[16654] = 32'b11111111111111111101110000011010;
assign LUT_2[16655] = 32'b11111111111111111010101000110011;
assign LUT_2[16656] = 32'b11111111111111111010001100100011;
assign LUT_2[16657] = 32'b11111111111111110111000100111100;
assign LUT_2[16658] = 32'b00000000000000000001000101011111;
assign LUT_2[16659] = 32'b11111111111111111101111101111000;
assign LUT_2[16660] = 32'b11111111111111110110101010001011;
assign LUT_2[16661] = 32'b11111111111111110011100010100100;
assign LUT_2[16662] = 32'b11111111111111111101100011000111;
assign LUT_2[16663] = 32'b11111111111111111010011011100000;
assign LUT_2[16664] = 32'b11111111111111110100111110000000;
assign LUT_2[16665] = 32'b11111111111111110001110110011001;
assign LUT_2[16666] = 32'b11111111111111111011110110111100;
assign LUT_2[16667] = 32'b11111111111111111000101111010101;
assign LUT_2[16668] = 32'b11111111111111110001011011101000;
assign LUT_2[16669] = 32'b11111111111111101110010100000001;
assign LUT_2[16670] = 32'b11111111111111111000010100100100;
assign LUT_2[16671] = 32'b11111111111111110101001100111101;
assign LUT_2[16672] = 32'b00000000000000000000000100000010;
assign LUT_2[16673] = 32'b11111111111111111100111100011011;
assign LUT_2[16674] = 32'b00000000000000000110111100111110;
assign LUT_2[16675] = 32'b00000000000000000011110101010111;
assign LUT_2[16676] = 32'b11111111111111111100100001101010;
assign LUT_2[16677] = 32'b11111111111111111001011010000011;
assign LUT_2[16678] = 32'b00000000000000000011011010100110;
assign LUT_2[16679] = 32'b00000000000000000000010010111111;
assign LUT_2[16680] = 32'b11111111111111111010110101011111;
assign LUT_2[16681] = 32'b11111111111111110111101101111000;
assign LUT_2[16682] = 32'b00000000000000000001101110011011;
assign LUT_2[16683] = 32'b11111111111111111110100110110100;
assign LUT_2[16684] = 32'b11111111111111110111010011000111;
assign LUT_2[16685] = 32'b11111111111111110100001011100000;
assign LUT_2[16686] = 32'b11111111111111111110001100000011;
assign LUT_2[16687] = 32'b11111111111111111011000100011100;
assign LUT_2[16688] = 32'b11111111111111111010101000001100;
assign LUT_2[16689] = 32'b11111111111111110111100000100101;
assign LUT_2[16690] = 32'b00000000000000000001100001001000;
assign LUT_2[16691] = 32'b11111111111111111110011001100001;
assign LUT_2[16692] = 32'b11111111111111110111000101110100;
assign LUT_2[16693] = 32'b11111111111111110011111110001101;
assign LUT_2[16694] = 32'b11111111111111111101111110110000;
assign LUT_2[16695] = 32'b11111111111111111010110111001001;
assign LUT_2[16696] = 32'b11111111111111110101011001101001;
assign LUT_2[16697] = 32'b11111111111111110010010010000010;
assign LUT_2[16698] = 32'b11111111111111111100010010100101;
assign LUT_2[16699] = 32'b11111111111111111001001010111110;
assign LUT_2[16700] = 32'b11111111111111110001110111010001;
assign LUT_2[16701] = 32'b11111111111111101110101111101010;
assign LUT_2[16702] = 32'b11111111111111111000110000001101;
assign LUT_2[16703] = 32'b11111111111111110101101000100110;
assign LUT_2[16704] = 32'b11111111111111110111110000111100;
assign LUT_2[16705] = 32'b11111111111111110100101001010101;
assign LUT_2[16706] = 32'b11111111111111111110101001111000;
assign LUT_2[16707] = 32'b11111111111111111011100010010001;
assign LUT_2[16708] = 32'b11111111111111110100001110100100;
assign LUT_2[16709] = 32'b11111111111111110001000110111101;
assign LUT_2[16710] = 32'b11111111111111111011000111100000;
assign LUT_2[16711] = 32'b11111111111111110111111111111001;
assign LUT_2[16712] = 32'b11111111111111110010100010011001;
assign LUT_2[16713] = 32'b11111111111111101111011010110010;
assign LUT_2[16714] = 32'b11111111111111111001011011010101;
assign LUT_2[16715] = 32'b11111111111111110110010011101110;
assign LUT_2[16716] = 32'b11111111111111101111000000000001;
assign LUT_2[16717] = 32'b11111111111111101011111000011010;
assign LUT_2[16718] = 32'b11111111111111110101111000111101;
assign LUT_2[16719] = 32'b11111111111111110010110001010110;
assign LUT_2[16720] = 32'b11111111111111110010010101000110;
assign LUT_2[16721] = 32'b11111111111111101111001101011111;
assign LUT_2[16722] = 32'b11111111111111111001001110000010;
assign LUT_2[16723] = 32'b11111111111111110110000110011011;
assign LUT_2[16724] = 32'b11111111111111101110110010101110;
assign LUT_2[16725] = 32'b11111111111111101011101011000111;
assign LUT_2[16726] = 32'b11111111111111110101101011101010;
assign LUT_2[16727] = 32'b11111111111111110010100100000011;
assign LUT_2[16728] = 32'b11111111111111101101000110100011;
assign LUT_2[16729] = 32'b11111111111111101001111110111100;
assign LUT_2[16730] = 32'b11111111111111110011111111011111;
assign LUT_2[16731] = 32'b11111111111111110000110111111000;
assign LUT_2[16732] = 32'b11111111111111101001100100001011;
assign LUT_2[16733] = 32'b11111111111111100110011100100100;
assign LUT_2[16734] = 32'b11111111111111110000011101000111;
assign LUT_2[16735] = 32'b11111111111111101101010101100000;
assign LUT_2[16736] = 32'b11111111111111111000001100100101;
assign LUT_2[16737] = 32'b11111111111111110101000100111110;
assign LUT_2[16738] = 32'b11111111111111111111000101100001;
assign LUT_2[16739] = 32'b11111111111111111011111101111010;
assign LUT_2[16740] = 32'b11111111111111110100101010001101;
assign LUT_2[16741] = 32'b11111111111111110001100010100110;
assign LUT_2[16742] = 32'b11111111111111111011100011001001;
assign LUT_2[16743] = 32'b11111111111111111000011011100010;
assign LUT_2[16744] = 32'b11111111111111110010111110000010;
assign LUT_2[16745] = 32'b11111111111111101111110110011011;
assign LUT_2[16746] = 32'b11111111111111111001110110111110;
assign LUT_2[16747] = 32'b11111111111111110110101111010111;
assign LUT_2[16748] = 32'b11111111111111101111011011101010;
assign LUT_2[16749] = 32'b11111111111111101100010100000011;
assign LUT_2[16750] = 32'b11111111111111110110010100100110;
assign LUT_2[16751] = 32'b11111111111111110011001100111111;
assign LUT_2[16752] = 32'b11111111111111110010110000101111;
assign LUT_2[16753] = 32'b11111111111111101111101001001000;
assign LUT_2[16754] = 32'b11111111111111111001101001101011;
assign LUT_2[16755] = 32'b11111111111111110110100010000100;
assign LUT_2[16756] = 32'b11111111111111101111001110010111;
assign LUT_2[16757] = 32'b11111111111111101100000110110000;
assign LUT_2[16758] = 32'b11111111111111110110000111010011;
assign LUT_2[16759] = 32'b11111111111111110010111111101100;
assign LUT_2[16760] = 32'b11111111111111101101100010001100;
assign LUT_2[16761] = 32'b11111111111111101010011010100101;
assign LUT_2[16762] = 32'b11111111111111110100011011001000;
assign LUT_2[16763] = 32'b11111111111111110001010011100001;
assign LUT_2[16764] = 32'b11111111111111101001111111110100;
assign LUT_2[16765] = 32'b11111111111111100110111000001101;
assign LUT_2[16766] = 32'b11111111111111110000111000110000;
assign LUT_2[16767] = 32'b11111111111111101101110001001001;
assign LUT_2[16768] = 32'b00000000000000000011111100101000;
assign LUT_2[16769] = 32'b00000000000000000000110101000001;
assign LUT_2[16770] = 32'b00000000000000001010110101100100;
assign LUT_2[16771] = 32'b00000000000000000111101101111101;
assign LUT_2[16772] = 32'b00000000000000000000011010010000;
assign LUT_2[16773] = 32'b11111111111111111101010010101001;
assign LUT_2[16774] = 32'b00000000000000000111010011001100;
assign LUT_2[16775] = 32'b00000000000000000100001011100101;
assign LUT_2[16776] = 32'b11111111111111111110101110000101;
assign LUT_2[16777] = 32'b11111111111111111011100110011110;
assign LUT_2[16778] = 32'b00000000000000000101100111000001;
assign LUT_2[16779] = 32'b00000000000000000010011111011010;
assign LUT_2[16780] = 32'b11111111111111111011001011101101;
assign LUT_2[16781] = 32'b11111111111111111000000100000110;
assign LUT_2[16782] = 32'b00000000000000000010000100101001;
assign LUT_2[16783] = 32'b11111111111111111110111101000010;
assign LUT_2[16784] = 32'b11111111111111111110100000110010;
assign LUT_2[16785] = 32'b11111111111111111011011001001011;
assign LUT_2[16786] = 32'b00000000000000000101011001101110;
assign LUT_2[16787] = 32'b00000000000000000010010010000111;
assign LUT_2[16788] = 32'b11111111111111111010111110011010;
assign LUT_2[16789] = 32'b11111111111111110111110110110011;
assign LUT_2[16790] = 32'b00000000000000000001110111010110;
assign LUT_2[16791] = 32'b11111111111111111110101111101111;
assign LUT_2[16792] = 32'b11111111111111111001010010001111;
assign LUT_2[16793] = 32'b11111111111111110110001010101000;
assign LUT_2[16794] = 32'b00000000000000000000001011001011;
assign LUT_2[16795] = 32'b11111111111111111101000011100100;
assign LUT_2[16796] = 32'b11111111111111110101101111110111;
assign LUT_2[16797] = 32'b11111111111111110010101000010000;
assign LUT_2[16798] = 32'b11111111111111111100101000110011;
assign LUT_2[16799] = 32'b11111111111111111001100001001100;
assign LUT_2[16800] = 32'b00000000000000000100011000010001;
assign LUT_2[16801] = 32'b00000000000000000001010000101010;
assign LUT_2[16802] = 32'b00000000000000001011010001001101;
assign LUT_2[16803] = 32'b00000000000000001000001001100110;
assign LUT_2[16804] = 32'b00000000000000000000110101111001;
assign LUT_2[16805] = 32'b11111111111111111101101110010010;
assign LUT_2[16806] = 32'b00000000000000000111101110110101;
assign LUT_2[16807] = 32'b00000000000000000100100111001110;
assign LUT_2[16808] = 32'b11111111111111111111001001101110;
assign LUT_2[16809] = 32'b11111111111111111100000010000111;
assign LUT_2[16810] = 32'b00000000000000000110000010101010;
assign LUT_2[16811] = 32'b00000000000000000010111011000011;
assign LUT_2[16812] = 32'b11111111111111111011100111010110;
assign LUT_2[16813] = 32'b11111111111111111000011111101111;
assign LUT_2[16814] = 32'b00000000000000000010100000010010;
assign LUT_2[16815] = 32'b11111111111111111111011000101011;
assign LUT_2[16816] = 32'b11111111111111111110111100011011;
assign LUT_2[16817] = 32'b11111111111111111011110100110100;
assign LUT_2[16818] = 32'b00000000000000000101110101010111;
assign LUT_2[16819] = 32'b00000000000000000010101101110000;
assign LUT_2[16820] = 32'b11111111111111111011011010000011;
assign LUT_2[16821] = 32'b11111111111111111000010010011100;
assign LUT_2[16822] = 32'b00000000000000000010010010111111;
assign LUT_2[16823] = 32'b11111111111111111111001011011000;
assign LUT_2[16824] = 32'b11111111111111111001101101111000;
assign LUT_2[16825] = 32'b11111111111111110110100110010001;
assign LUT_2[16826] = 32'b00000000000000000000100110110100;
assign LUT_2[16827] = 32'b11111111111111111101011111001101;
assign LUT_2[16828] = 32'b11111111111111110110001011100000;
assign LUT_2[16829] = 32'b11111111111111110011000011111001;
assign LUT_2[16830] = 32'b11111111111111111101000100011100;
assign LUT_2[16831] = 32'b11111111111111111001111100110101;
assign LUT_2[16832] = 32'b11111111111111111100000101001011;
assign LUT_2[16833] = 32'b11111111111111111000111101100100;
assign LUT_2[16834] = 32'b00000000000000000010111110000111;
assign LUT_2[16835] = 32'b11111111111111111111110110100000;
assign LUT_2[16836] = 32'b11111111111111111000100010110011;
assign LUT_2[16837] = 32'b11111111111111110101011011001100;
assign LUT_2[16838] = 32'b11111111111111111111011011101111;
assign LUT_2[16839] = 32'b11111111111111111100010100001000;
assign LUT_2[16840] = 32'b11111111111111110110110110101000;
assign LUT_2[16841] = 32'b11111111111111110011101111000001;
assign LUT_2[16842] = 32'b11111111111111111101101111100100;
assign LUT_2[16843] = 32'b11111111111111111010100111111101;
assign LUT_2[16844] = 32'b11111111111111110011010100010000;
assign LUT_2[16845] = 32'b11111111111111110000001100101001;
assign LUT_2[16846] = 32'b11111111111111111010001101001100;
assign LUT_2[16847] = 32'b11111111111111110111000101100101;
assign LUT_2[16848] = 32'b11111111111111110110101001010101;
assign LUT_2[16849] = 32'b11111111111111110011100001101110;
assign LUT_2[16850] = 32'b11111111111111111101100010010001;
assign LUT_2[16851] = 32'b11111111111111111010011010101010;
assign LUT_2[16852] = 32'b11111111111111110011000110111101;
assign LUT_2[16853] = 32'b11111111111111101111111111010110;
assign LUT_2[16854] = 32'b11111111111111111001111111111001;
assign LUT_2[16855] = 32'b11111111111111110110111000010010;
assign LUT_2[16856] = 32'b11111111111111110001011010110010;
assign LUT_2[16857] = 32'b11111111111111101110010011001011;
assign LUT_2[16858] = 32'b11111111111111111000010011101110;
assign LUT_2[16859] = 32'b11111111111111110101001100000111;
assign LUT_2[16860] = 32'b11111111111111101101111000011010;
assign LUT_2[16861] = 32'b11111111111111101010110000110011;
assign LUT_2[16862] = 32'b11111111111111110100110001010110;
assign LUT_2[16863] = 32'b11111111111111110001101001101111;
assign LUT_2[16864] = 32'b11111111111111111100100000110100;
assign LUT_2[16865] = 32'b11111111111111111001011001001101;
assign LUT_2[16866] = 32'b00000000000000000011011001110000;
assign LUT_2[16867] = 32'b00000000000000000000010010001001;
assign LUT_2[16868] = 32'b11111111111111111000111110011100;
assign LUT_2[16869] = 32'b11111111111111110101110110110101;
assign LUT_2[16870] = 32'b11111111111111111111110111011000;
assign LUT_2[16871] = 32'b11111111111111111100101111110001;
assign LUT_2[16872] = 32'b11111111111111110111010010010001;
assign LUT_2[16873] = 32'b11111111111111110100001010101010;
assign LUT_2[16874] = 32'b11111111111111111110001011001101;
assign LUT_2[16875] = 32'b11111111111111111011000011100110;
assign LUT_2[16876] = 32'b11111111111111110011101111111001;
assign LUT_2[16877] = 32'b11111111111111110000101000010010;
assign LUT_2[16878] = 32'b11111111111111111010101000110101;
assign LUT_2[16879] = 32'b11111111111111110111100001001110;
assign LUT_2[16880] = 32'b11111111111111110111000100111110;
assign LUT_2[16881] = 32'b11111111111111110011111101010111;
assign LUT_2[16882] = 32'b11111111111111111101111101111010;
assign LUT_2[16883] = 32'b11111111111111111010110110010011;
assign LUT_2[16884] = 32'b11111111111111110011100010100110;
assign LUT_2[16885] = 32'b11111111111111110000011010111111;
assign LUT_2[16886] = 32'b11111111111111111010011011100010;
assign LUT_2[16887] = 32'b11111111111111110111010011111011;
assign LUT_2[16888] = 32'b11111111111111110001110110011011;
assign LUT_2[16889] = 32'b11111111111111101110101110110100;
assign LUT_2[16890] = 32'b11111111111111111000101111010111;
assign LUT_2[16891] = 32'b11111111111111110101100111110000;
assign LUT_2[16892] = 32'b11111111111111101110010100000011;
assign LUT_2[16893] = 32'b11111111111111101011001100011100;
assign LUT_2[16894] = 32'b11111111111111110101001100111111;
assign LUT_2[16895] = 32'b11111111111111110010000101011000;
assign LUT_2[16896] = 32'b00000000000000000000011011100101;
assign LUT_2[16897] = 32'b11111111111111111101010011111110;
assign LUT_2[16898] = 32'b00000000000000000111010100100001;
assign LUT_2[16899] = 32'b00000000000000000100001100111010;
assign LUT_2[16900] = 32'b11111111111111111100111001001101;
assign LUT_2[16901] = 32'b11111111111111111001110001100110;
assign LUT_2[16902] = 32'b00000000000000000011110010001001;
assign LUT_2[16903] = 32'b00000000000000000000101010100010;
assign LUT_2[16904] = 32'b11111111111111111011001101000010;
assign LUT_2[16905] = 32'b11111111111111111000000101011011;
assign LUT_2[16906] = 32'b00000000000000000010000101111110;
assign LUT_2[16907] = 32'b11111111111111111110111110010111;
assign LUT_2[16908] = 32'b11111111111111110111101010101010;
assign LUT_2[16909] = 32'b11111111111111110100100011000011;
assign LUT_2[16910] = 32'b11111111111111111110100011100110;
assign LUT_2[16911] = 32'b11111111111111111011011011111111;
assign LUT_2[16912] = 32'b11111111111111111010111111101111;
assign LUT_2[16913] = 32'b11111111111111110111111000001000;
assign LUT_2[16914] = 32'b00000000000000000001111000101011;
assign LUT_2[16915] = 32'b11111111111111111110110001000100;
assign LUT_2[16916] = 32'b11111111111111110111011101010111;
assign LUT_2[16917] = 32'b11111111111111110100010101110000;
assign LUT_2[16918] = 32'b11111111111111111110010110010011;
assign LUT_2[16919] = 32'b11111111111111111011001110101100;
assign LUT_2[16920] = 32'b11111111111111110101110001001100;
assign LUT_2[16921] = 32'b11111111111111110010101001100101;
assign LUT_2[16922] = 32'b11111111111111111100101010001000;
assign LUT_2[16923] = 32'b11111111111111111001100010100001;
assign LUT_2[16924] = 32'b11111111111111110010001110110100;
assign LUT_2[16925] = 32'b11111111111111101111000111001101;
assign LUT_2[16926] = 32'b11111111111111111001000111110000;
assign LUT_2[16927] = 32'b11111111111111110110000000001001;
assign LUT_2[16928] = 32'b00000000000000000000110111001110;
assign LUT_2[16929] = 32'b11111111111111111101101111100111;
assign LUT_2[16930] = 32'b00000000000000000111110000001010;
assign LUT_2[16931] = 32'b00000000000000000100101000100011;
assign LUT_2[16932] = 32'b11111111111111111101010100110110;
assign LUT_2[16933] = 32'b11111111111111111010001101001111;
assign LUT_2[16934] = 32'b00000000000000000100001101110010;
assign LUT_2[16935] = 32'b00000000000000000001000110001011;
assign LUT_2[16936] = 32'b11111111111111111011101000101011;
assign LUT_2[16937] = 32'b11111111111111111000100001000100;
assign LUT_2[16938] = 32'b00000000000000000010100001100111;
assign LUT_2[16939] = 32'b11111111111111111111011010000000;
assign LUT_2[16940] = 32'b11111111111111111000000110010011;
assign LUT_2[16941] = 32'b11111111111111110100111110101100;
assign LUT_2[16942] = 32'b11111111111111111110111111001111;
assign LUT_2[16943] = 32'b11111111111111111011110111101000;
assign LUT_2[16944] = 32'b11111111111111111011011011011000;
assign LUT_2[16945] = 32'b11111111111111111000010011110001;
assign LUT_2[16946] = 32'b00000000000000000010010100010100;
assign LUT_2[16947] = 32'b11111111111111111111001100101101;
assign LUT_2[16948] = 32'b11111111111111110111111001000000;
assign LUT_2[16949] = 32'b11111111111111110100110001011001;
assign LUT_2[16950] = 32'b11111111111111111110110001111100;
assign LUT_2[16951] = 32'b11111111111111111011101010010101;
assign LUT_2[16952] = 32'b11111111111111110110001100110101;
assign LUT_2[16953] = 32'b11111111111111110011000101001110;
assign LUT_2[16954] = 32'b11111111111111111101000101110001;
assign LUT_2[16955] = 32'b11111111111111111001111110001010;
assign LUT_2[16956] = 32'b11111111111111110010101010011101;
assign LUT_2[16957] = 32'b11111111111111101111100010110110;
assign LUT_2[16958] = 32'b11111111111111111001100011011001;
assign LUT_2[16959] = 32'b11111111111111110110011011110010;
assign LUT_2[16960] = 32'b11111111111111111000100100001000;
assign LUT_2[16961] = 32'b11111111111111110101011100100001;
assign LUT_2[16962] = 32'b11111111111111111111011101000100;
assign LUT_2[16963] = 32'b11111111111111111100010101011101;
assign LUT_2[16964] = 32'b11111111111111110101000001110000;
assign LUT_2[16965] = 32'b11111111111111110001111010001001;
assign LUT_2[16966] = 32'b11111111111111111011111010101100;
assign LUT_2[16967] = 32'b11111111111111111000110011000101;
assign LUT_2[16968] = 32'b11111111111111110011010101100101;
assign LUT_2[16969] = 32'b11111111111111110000001101111110;
assign LUT_2[16970] = 32'b11111111111111111010001110100001;
assign LUT_2[16971] = 32'b11111111111111110111000110111010;
assign LUT_2[16972] = 32'b11111111111111101111110011001101;
assign LUT_2[16973] = 32'b11111111111111101100101011100110;
assign LUT_2[16974] = 32'b11111111111111110110101100001001;
assign LUT_2[16975] = 32'b11111111111111110011100100100010;
assign LUT_2[16976] = 32'b11111111111111110011001000010010;
assign LUT_2[16977] = 32'b11111111111111110000000000101011;
assign LUT_2[16978] = 32'b11111111111111111010000001001110;
assign LUT_2[16979] = 32'b11111111111111110110111001100111;
assign LUT_2[16980] = 32'b11111111111111101111100101111010;
assign LUT_2[16981] = 32'b11111111111111101100011110010011;
assign LUT_2[16982] = 32'b11111111111111110110011110110110;
assign LUT_2[16983] = 32'b11111111111111110011010111001111;
assign LUT_2[16984] = 32'b11111111111111101101111001101111;
assign LUT_2[16985] = 32'b11111111111111101010110010001000;
assign LUT_2[16986] = 32'b11111111111111110100110010101011;
assign LUT_2[16987] = 32'b11111111111111110001101011000100;
assign LUT_2[16988] = 32'b11111111111111101010010111010111;
assign LUT_2[16989] = 32'b11111111111111100111001111110000;
assign LUT_2[16990] = 32'b11111111111111110001010000010011;
assign LUT_2[16991] = 32'b11111111111111101110001000101100;
assign LUT_2[16992] = 32'b11111111111111111000111111110001;
assign LUT_2[16993] = 32'b11111111111111110101111000001010;
assign LUT_2[16994] = 32'b11111111111111111111111000101101;
assign LUT_2[16995] = 32'b11111111111111111100110001000110;
assign LUT_2[16996] = 32'b11111111111111110101011101011001;
assign LUT_2[16997] = 32'b11111111111111110010010101110010;
assign LUT_2[16998] = 32'b11111111111111111100010110010101;
assign LUT_2[16999] = 32'b11111111111111111001001110101110;
assign LUT_2[17000] = 32'b11111111111111110011110001001110;
assign LUT_2[17001] = 32'b11111111111111110000101001100111;
assign LUT_2[17002] = 32'b11111111111111111010101010001010;
assign LUT_2[17003] = 32'b11111111111111110111100010100011;
assign LUT_2[17004] = 32'b11111111111111110000001110110110;
assign LUT_2[17005] = 32'b11111111111111101101000111001111;
assign LUT_2[17006] = 32'b11111111111111110111000111110010;
assign LUT_2[17007] = 32'b11111111111111110100000000001011;
assign LUT_2[17008] = 32'b11111111111111110011100011111011;
assign LUT_2[17009] = 32'b11111111111111110000011100010100;
assign LUT_2[17010] = 32'b11111111111111111010011100110111;
assign LUT_2[17011] = 32'b11111111111111110111010101010000;
assign LUT_2[17012] = 32'b11111111111111110000000001100011;
assign LUT_2[17013] = 32'b11111111111111101100111001111100;
assign LUT_2[17014] = 32'b11111111111111110110111010011111;
assign LUT_2[17015] = 32'b11111111111111110011110010111000;
assign LUT_2[17016] = 32'b11111111111111101110010101011000;
assign LUT_2[17017] = 32'b11111111111111101011001101110001;
assign LUT_2[17018] = 32'b11111111111111110101001110010100;
assign LUT_2[17019] = 32'b11111111111111110010000110101101;
assign LUT_2[17020] = 32'b11111111111111101010110011000000;
assign LUT_2[17021] = 32'b11111111111111100111101011011001;
assign LUT_2[17022] = 32'b11111111111111110001101011111100;
assign LUT_2[17023] = 32'b11111111111111101110100100010101;
assign LUT_2[17024] = 32'b00000000000000000100101111110100;
assign LUT_2[17025] = 32'b00000000000000000001101000001101;
assign LUT_2[17026] = 32'b00000000000000001011101000110000;
assign LUT_2[17027] = 32'b00000000000000001000100001001001;
assign LUT_2[17028] = 32'b00000000000000000001001101011100;
assign LUT_2[17029] = 32'b11111111111111111110000101110101;
assign LUT_2[17030] = 32'b00000000000000001000000110011000;
assign LUT_2[17031] = 32'b00000000000000000100111110110001;
assign LUT_2[17032] = 32'b11111111111111111111100001010001;
assign LUT_2[17033] = 32'b11111111111111111100011001101010;
assign LUT_2[17034] = 32'b00000000000000000110011010001101;
assign LUT_2[17035] = 32'b00000000000000000011010010100110;
assign LUT_2[17036] = 32'b11111111111111111011111110111001;
assign LUT_2[17037] = 32'b11111111111111111000110111010010;
assign LUT_2[17038] = 32'b00000000000000000010110111110101;
assign LUT_2[17039] = 32'b11111111111111111111110000001110;
assign LUT_2[17040] = 32'b11111111111111111111010011111110;
assign LUT_2[17041] = 32'b11111111111111111100001100010111;
assign LUT_2[17042] = 32'b00000000000000000110001100111010;
assign LUT_2[17043] = 32'b00000000000000000011000101010011;
assign LUT_2[17044] = 32'b11111111111111111011110001100110;
assign LUT_2[17045] = 32'b11111111111111111000101001111111;
assign LUT_2[17046] = 32'b00000000000000000010101010100010;
assign LUT_2[17047] = 32'b11111111111111111111100010111011;
assign LUT_2[17048] = 32'b11111111111111111010000101011011;
assign LUT_2[17049] = 32'b11111111111111110110111101110100;
assign LUT_2[17050] = 32'b00000000000000000000111110010111;
assign LUT_2[17051] = 32'b11111111111111111101110110110000;
assign LUT_2[17052] = 32'b11111111111111110110100011000011;
assign LUT_2[17053] = 32'b11111111111111110011011011011100;
assign LUT_2[17054] = 32'b11111111111111111101011011111111;
assign LUT_2[17055] = 32'b11111111111111111010010100011000;
assign LUT_2[17056] = 32'b00000000000000000101001011011101;
assign LUT_2[17057] = 32'b00000000000000000010000011110110;
assign LUT_2[17058] = 32'b00000000000000001100000100011001;
assign LUT_2[17059] = 32'b00000000000000001000111100110010;
assign LUT_2[17060] = 32'b00000000000000000001101001000101;
assign LUT_2[17061] = 32'b11111111111111111110100001011110;
assign LUT_2[17062] = 32'b00000000000000001000100010000001;
assign LUT_2[17063] = 32'b00000000000000000101011010011010;
assign LUT_2[17064] = 32'b11111111111111111111111100111010;
assign LUT_2[17065] = 32'b11111111111111111100110101010011;
assign LUT_2[17066] = 32'b00000000000000000110110101110110;
assign LUT_2[17067] = 32'b00000000000000000011101110001111;
assign LUT_2[17068] = 32'b11111111111111111100011010100010;
assign LUT_2[17069] = 32'b11111111111111111001010010111011;
assign LUT_2[17070] = 32'b00000000000000000011010011011110;
assign LUT_2[17071] = 32'b00000000000000000000001011110111;
assign LUT_2[17072] = 32'b11111111111111111111101111100111;
assign LUT_2[17073] = 32'b11111111111111111100101000000000;
assign LUT_2[17074] = 32'b00000000000000000110101000100011;
assign LUT_2[17075] = 32'b00000000000000000011100000111100;
assign LUT_2[17076] = 32'b11111111111111111100001101001111;
assign LUT_2[17077] = 32'b11111111111111111001000101101000;
assign LUT_2[17078] = 32'b00000000000000000011000110001011;
assign LUT_2[17079] = 32'b11111111111111111111111110100100;
assign LUT_2[17080] = 32'b11111111111111111010100001000100;
assign LUT_2[17081] = 32'b11111111111111110111011001011101;
assign LUT_2[17082] = 32'b00000000000000000001011010000000;
assign LUT_2[17083] = 32'b11111111111111111110010010011001;
assign LUT_2[17084] = 32'b11111111111111110110111110101100;
assign LUT_2[17085] = 32'b11111111111111110011110111000101;
assign LUT_2[17086] = 32'b11111111111111111101110111101000;
assign LUT_2[17087] = 32'b11111111111111111010110000000001;
assign LUT_2[17088] = 32'b11111111111111111100111000010111;
assign LUT_2[17089] = 32'b11111111111111111001110000110000;
assign LUT_2[17090] = 32'b00000000000000000011110001010011;
assign LUT_2[17091] = 32'b00000000000000000000101001101100;
assign LUT_2[17092] = 32'b11111111111111111001010101111111;
assign LUT_2[17093] = 32'b11111111111111110110001110011000;
assign LUT_2[17094] = 32'b00000000000000000000001110111011;
assign LUT_2[17095] = 32'b11111111111111111101000111010100;
assign LUT_2[17096] = 32'b11111111111111110111101001110100;
assign LUT_2[17097] = 32'b11111111111111110100100010001101;
assign LUT_2[17098] = 32'b11111111111111111110100010110000;
assign LUT_2[17099] = 32'b11111111111111111011011011001001;
assign LUT_2[17100] = 32'b11111111111111110100000111011100;
assign LUT_2[17101] = 32'b11111111111111110000111111110101;
assign LUT_2[17102] = 32'b11111111111111111011000000011000;
assign LUT_2[17103] = 32'b11111111111111110111111000110001;
assign LUT_2[17104] = 32'b11111111111111110111011100100001;
assign LUT_2[17105] = 32'b11111111111111110100010100111010;
assign LUT_2[17106] = 32'b11111111111111111110010101011101;
assign LUT_2[17107] = 32'b11111111111111111011001101110110;
assign LUT_2[17108] = 32'b11111111111111110011111010001001;
assign LUT_2[17109] = 32'b11111111111111110000110010100010;
assign LUT_2[17110] = 32'b11111111111111111010110011000101;
assign LUT_2[17111] = 32'b11111111111111110111101011011110;
assign LUT_2[17112] = 32'b11111111111111110010001101111110;
assign LUT_2[17113] = 32'b11111111111111101111000110010111;
assign LUT_2[17114] = 32'b11111111111111111001000110111010;
assign LUT_2[17115] = 32'b11111111111111110101111111010011;
assign LUT_2[17116] = 32'b11111111111111101110101011100110;
assign LUT_2[17117] = 32'b11111111111111101011100011111111;
assign LUT_2[17118] = 32'b11111111111111110101100100100010;
assign LUT_2[17119] = 32'b11111111111111110010011100111011;
assign LUT_2[17120] = 32'b11111111111111111101010100000000;
assign LUT_2[17121] = 32'b11111111111111111010001100011001;
assign LUT_2[17122] = 32'b00000000000000000100001100111100;
assign LUT_2[17123] = 32'b00000000000000000001000101010101;
assign LUT_2[17124] = 32'b11111111111111111001110001101000;
assign LUT_2[17125] = 32'b11111111111111110110101010000001;
assign LUT_2[17126] = 32'b00000000000000000000101010100100;
assign LUT_2[17127] = 32'b11111111111111111101100010111101;
assign LUT_2[17128] = 32'b11111111111111111000000101011101;
assign LUT_2[17129] = 32'b11111111111111110100111101110110;
assign LUT_2[17130] = 32'b11111111111111111110111110011001;
assign LUT_2[17131] = 32'b11111111111111111011110110110010;
assign LUT_2[17132] = 32'b11111111111111110100100011000101;
assign LUT_2[17133] = 32'b11111111111111110001011011011110;
assign LUT_2[17134] = 32'b11111111111111111011011100000001;
assign LUT_2[17135] = 32'b11111111111111111000010100011010;
assign LUT_2[17136] = 32'b11111111111111110111111000001010;
assign LUT_2[17137] = 32'b11111111111111110100110000100011;
assign LUT_2[17138] = 32'b11111111111111111110110001000110;
assign LUT_2[17139] = 32'b11111111111111111011101001011111;
assign LUT_2[17140] = 32'b11111111111111110100010101110010;
assign LUT_2[17141] = 32'b11111111111111110001001110001011;
assign LUT_2[17142] = 32'b11111111111111111011001110101110;
assign LUT_2[17143] = 32'b11111111111111111000000111000111;
assign LUT_2[17144] = 32'b11111111111111110010101001100111;
assign LUT_2[17145] = 32'b11111111111111101111100010000000;
assign LUT_2[17146] = 32'b11111111111111111001100010100011;
assign LUT_2[17147] = 32'b11111111111111110110011010111100;
assign LUT_2[17148] = 32'b11111111111111101111000111001111;
assign LUT_2[17149] = 32'b11111111111111101011111111101000;
assign LUT_2[17150] = 32'b11111111111111110110000000001011;
assign LUT_2[17151] = 32'b11111111111111110010111000100100;
assign LUT_2[17152] = 32'b00000000000000000100011010001011;
assign LUT_2[17153] = 32'b00000000000000000001010010100100;
assign LUT_2[17154] = 32'b00000000000000001011010011000111;
assign LUT_2[17155] = 32'b00000000000000001000001011100000;
assign LUT_2[17156] = 32'b00000000000000000000110111110011;
assign LUT_2[17157] = 32'b11111111111111111101110000001100;
assign LUT_2[17158] = 32'b00000000000000000111110000101111;
assign LUT_2[17159] = 32'b00000000000000000100101001001000;
assign LUT_2[17160] = 32'b11111111111111111111001011101000;
assign LUT_2[17161] = 32'b11111111111111111100000100000001;
assign LUT_2[17162] = 32'b00000000000000000110000100100100;
assign LUT_2[17163] = 32'b00000000000000000010111100111101;
assign LUT_2[17164] = 32'b11111111111111111011101001010000;
assign LUT_2[17165] = 32'b11111111111111111000100001101001;
assign LUT_2[17166] = 32'b00000000000000000010100010001100;
assign LUT_2[17167] = 32'b11111111111111111111011010100101;
assign LUT_2[17168] = 32'b11111111111111111110111110010101;
assign LUT_2[17169] = 32'b11111111111111111011110110101110;
assign LUT_2[17170] = 32'b00000000000000000101110111010001;
assign LUT_2[17171] = 32'b00000000000000000010101111101010;
assign LUT_2[17172] = 32'b11111111111111111011011011111101;
assign LUT_2[17173] = 32'b11111111111111111000010100010110;
assign LUT_2[17174] = 32'b00000000000000000010010100111001;
assign LUT_2[17175] = 32'b11111111111111111111001101010010;
assign LUT_2[17176] = 32'b11111111111111111001101111110010;
assign LUT_2[17177] = 32'b11111111111111110110101000001011;
assign LUT_2[17178] = 32'b00000000000000000000101000101110;
assign LUT_2[17179] = 32'b11111111111111111101100001000111;
assign LUT_2[17180] = 32'b11111111111111110110001101011010;
assign LUT_2[17181] = 32'b11111111111111110011000101110011;
assign LUT_2[17182] = 32'b11111111111111111101000110010110;
assign LUT_2[17183] = 32'b11111111111111111001111110101111;
assign LUT_2[17184] = 32'b00000000000000000100110101110100;
assign LUT_2[17185] = 32'b00000000000000000001101110001101;
assign LUT_2[17186] = 32'b00000000000000001011101110110000;
assign LUT_2[17187] = 32'b00000000000000001000100111001001;
assign LUT_2[17188] = 32'b00000000000000000001010011011100;
assign LUT_2[17189] = 32'b11111111111111111110001011110101;
assign LUT_2[17190] = 32'b00000000000000001000001100011000;
assign LUT_2[17191] = 32'b00000000000000000101000100110001;
assign LUT_2[17192] = 32'b11111111111111111111100111010001;
assign LUT_2[17193] = 32'b11111111111111111100011111101010;
assign LUT_2[17194] = 32'b00000000000000000110100000001101;
assign LUT_2[17195] = 32'b00000000000000000011011000100110;
assign LUT_2[17196] = 32'b11111111111111111100000100111001;
assign LUT_2[17197] = 32'b11111111111111111000111101010010;
assign LUT_2[17198] = 32'b00000000000000000010111101110101;
assign LUT_2[17199] = 32'b11111111111111111111110110001110;
assign LUT_2[17200] = 32'b11111111111111111111011001111110;
assign LUT_2[17201] = 32'b11111111111111111100010010010111;
assign LUT_2[17202] = 32'b00000000000000000110010010111010;
assign LUT_2[17203] = 32'b00000000000000000011001011010011;
assign LUT_2[17204] = 32'b11111111111111111011110111100110;
assign LUT_2[17205] = 32'b11111111111111111000101111111111;
assign LUT_2[17206] = 32'b00000000000000000010110000100010;
assign LUT_2[17207] = 32'b11111111111111111111101000111011;
assign LUT_2[17208] = 32'b11111111111111111010001011011011;
assign LUT_2[17209] = 32'b11111111111111110111000011110100;
assign LUT_2[17210] = 32'b00000000000000000001000100010111;
assign LUT_2[17211] = 32'b11111111111111111101111100110000;
assign LUT_2[17212] = 32'b11111111111111110110101001000011;
assign LUT_2[17213] = 32'b11111111111111110011100001011100;
assign LUT_2[17214] = 32'b11111111111111111101100001111111;
assign LUT_2[17215] = 32'b11111111111111111010011010011000;
assign LUT_2[17216] = 32'b11111111111111111100100010101110;
assign LUT_2[17217] = 32'b11111111111111111001011011000111;
assign LUT_2[17218] = 32'b00000000000000000011011011101010;
assign LUT_2[17219] = 32'b00000000000000000000010100000011;
assign LUT_2[17220] = 32'b11111111111111111001000000010110;
assign LUT_2[17221] = 32'b11111111111111110101111000101111;
assign LUT_2[17222] = 32'b11111111111111111111111001010010;
assign LUT_2[17223] = 32'b11111111111111111100110001101011;
assign LUT_2[17224] = 32'b11111111111111110111010100001011;
assign LUT_2[17225] = 32'b11111111111111110100001100100100;
assign LUT_2[17226] = 32'b11111111111111111110001101000111;
assign LUT_2[17227] = 32'b11111111111111111011000101100000;
assign LUT_2[17228] = 32'b11111111111111110011110001110011;
assign LUT_2[17229] = 32'b11111111111111110000101010001100;
assign LUT_2[17230] = 32'b11111111111111111010101010101111;
assign LUT_2[17231] = 32'b11111111111111110111100011001000;
assign LUT_2[17232] = 32'b11111111111111110111000110111000;
assign LUT_2[17233] = 32'b11111111111111110011111111010001;
assign LUT_2[17234] = 32'b11111111111111111101111111110100;
assign LUT_2[17235] = 32'b11111111111111111010111000001101;
assign LUT_2[17236] = 32'b11111111111111110011100100100000;
assign LUT_2[17237] = 32'b11111111111111110000011100111001;
assign LUT_2[17238] = 32'b11111111111111111010011101011100;
assign LUT_2[17239] = 32'b11111111111111110111010101110101;
assign LUT_2[17240] = 32'b11111111111111110001111000010101;
assign LUT_2[17241] = 32'b11111111111111101110110000101110;
assign LUT_2[17242] = 32'b11111111111111111000110001010001;
assign LUT_2[17243] = 32'b11111111111111110101101001101010;
assign LUT_2[17244] = 32'b11111111111111101110010101111101;
assign LUT_2[17245] = 32'b11111111111111101011001110010110;
assign LUT_2[17246] = 32'b11111111111111110101001110111001;
assign LUT_2[17247] = 32'b11111111111111110010000111010010;
assign LUT_2[17248] = 32'b11111111111111111100111110010111;
assign LUT_2[17249] = 32'b11111111111111111001110110110000;
assign LUT_2[17250] = 32'b00000000000000000011110111010011;
assign LUT_2[17251] = 32'b00000000000000000000101111101100;
assign LUT_2[17252] = 32'b11111111111111111001011011111111;
assign LUT_2[17253] = 32'b11111111111111110110010100011000;
assign LUT_2[17254] = 32'b00000000000000000000010100111011;
assign LUT_2[17255] = 32'b11111111111111111101001101010100;
assign LUT_2[17256] = 32'b11111111111111110111101111110100;
assign LUT_2[17257] = 32'b11111111111111110100101000001101;
assign LUT_2[17258] = 32'b11111111111111111110101000110000;
assign LUT_2[17259] = 32'b11111111111111111011100001001001;
assign LUT_2[17260] = 32'b11111111111111110100001101011100;
assign LUT_2[17261] = 32'b11111111111111110001000101110101;
assign LUT_2[17262] = 32'b11111111111111111011000110011000;
assign LUT_2[17263] = 32'b11111111111111110111111110110001;
assign LUT_2[17264] = 32'b11111111111111110111100010100001;
assign LUT_2[17265] = 32'b11111111111111110100011010111010;
assign LUT_2[17266] = 32'b11111111111111111110011011011101;
assign LUT_2[17267] = 32'b11111111111111111011010011110110;
assign LUT_2[17268] = 32'b11111111111111110100000000001001;
assign LUT_2[17269] = 32'b11111111111111110000111000100010;
assign LUT_2[17270] = 32'b11111111111111111010111001000101;
assign LUT_2[17271] = 32'b11111111111111110111110001011110;
assign LUT_2[17272] = 32'b11111111111111110010010011111110;
assign LUT_2[17273] = 32'b11111111111111101111001100010111;
assign LUT_2[17274] = 32'b11111111111111111001001100111010;
assign LUT_2[17275] = 32'b11111111111111110110000101010011;
assign LUT_2[17276] = 32'b11111111111111101110110001100110;
assign LUT_2[17277] = 32'b11111111111111101011101001111111;
assign LUT_2[17278] = 32'b11111111111111110101101010100010;
assign LUT_2[17279] = 32'b11111111111111110010100010111011;
assign LUT_2[17280] = 32'b00000000000000001000101110011010;
assign LUT_2[17281] = 32'b00000000000000000101100110110011;
assign LUT_2[17282] = 32'b00000000000000001111100111010110;
assign LUT_2[17283] = 32'b00000000000000001100011111101111;
assign LUT_2[17284] = 32'b00000000000000000101001100000010;
assign LUT_2[17285] = 32'b00000000000000000010000100011011;
assign LUT_2[17286] = 32'b00000000000000001100000100111110;
assign LUT_2[17287] = 32'b00000000000000001000111101010111;
assign LUT_2[17288] = 32'b00000000000000000011011111110111;
assign LUT_2[17289] = 32'b00000000000000000000011000010000;
assign LUT_2[17290] = 32'b00000000000000001010011000110011;
assign LUT_2[17291] = 32'b00000000000000000111010001001100;
assign LUT_2[17292] = 32'b11111111111111111111111101011111;
assign LUT_2[17293] = 32'b11111111111111111100110101111000;
assign LUT_2[17294] = 32'b00000000000000000110110110011011;
assign LUT_2[17295] = 32'b00000000000000000011101110110100;
assign LUT_2[17296] = 32'b00000000000000000011010010100100;
assign LUT_2[17297] = 32'b00000000000000000000001010111101;
assign LUT_2[17298] = 32'b00000000000000001010001011100000;
assign LUT_2[17299] = 32'b00000000000000000111000011111001;
assign LUT_2[17300] = 32'b11111111111111111111110000001100;
assign LUT_2[17301] = 32'b11111111111111111100101000100101;
assign LUT_2[17302] = 32'b00000000000000000110101001001000;
assign LUT_2[17303] = 32'b00000000000000000011100001100001;
assign LUT_2[17304] = 32'b11111111111111111110000100000001;
assign LUT_2[17305] = 32'b11111111111111111010111100011010;
assign LUT_2[17306] = 32'b00000000000000000100111100111101;
assign LUT_2[17307] = 32'b00000000000000000001110101010110;
assign LUT_2[17308] = 32'b11111111111111111010100001101001;
assign LUT_2[17309] = 32'b11111111111111110111011010000010;
assign LUT_2[17310] = 32'b00000000000000000001011010100101;
assign LUT_2[17311] = 32'b11111111111111111110010010111110;
assign LUT_2[17312] = 32'b00000000000000001001001010000011;
assign LUT_2[17313] = 32'b00000000000000000110000010011100;
assign LUT_2[17314] = 32'b00000000000000010000000010111111;
assign LUT_2[17315] = 32'b00000000000000001100111011011000;
assign LUT_2[17316] = 32'b00000000000000000101100111101011;
assign LUT_2[17317] = 32'b00000000000000000010100000000100;
assign LUT_2[17318] = 32'b00000000000000001100100000100111;
assign LUT_2[17319] = 32'b00000000000000001001011001000000;
assign LUT_2[17320] = 32'b00000000000000000011111011100000;
assign LUT_2[17321] = 32'b00000000000000000000110011111001;
assign LUT_2[17322] = 32'b00000000000000001010110100011100;
assign LUT_2[17323] = 32'b00000000000000000111101100110101;
assign LUT_2[17324] = 32'b00000000000000000000011001001000;
assign LUT_2[17325] = 32'b11111111111111111101010001100001;
assign LUT_2[17326] = 32'b00000000000000000111010010000100;
assign LUT_2[17327] = 32'b00000000000000000100001010011101;
assign LUT_2[17328] = 32'b00000000000000000011101110001101;
assign LUT_2[17329] = 32'b00000000000000000000100110100110;
assign LUT_2[17330] = 32'b00000000000000001010100111001001;
assign LUT_2[17331] = 32'b00000000000000000111011111100010;
assign LUT_2[17332] = 32'b00000000000000000000001011110101;
assign LUT_2[17333] = 32'b11111111111111111101000100001110;
assign LUT_2[17334] = 32'b00000000000000000111000100110001;
assign LUT_2[17335] = 32'b00000000000000000011111101001010;
assign LUT_2[17336] = 32'b11111111111111111110011111101010;
assign LUT_2[17337] = 32'b11111111111111111011011000000011;
assign LUT_2[17338] = 32'b00000000000000000101011000100110;
assign LUT_2[17339] = 32'b00000000000000000010010000111111;
assign LUT_2[17340] = 32'b11111111111111111010111101010010;
assign LUT_2[17341] = 32'b11111111111111110111110101101011;
assign LUT_2[17342] = 32'b00000000000000000001110110001110;
assign LUT_2[17343] = 32'b11111111111111111110101110100111;
assign LUT_2[17344] = 32'b00000000000000000000110110111101;
assign LUT_2[17345] = 32'b11111111111111111101101111010110;
assign LUT_2[17346] = 32'b00000000000000000111101111111001;
assign LUT_2[17347] = 32'b00000000000000000100101000010010;
assign LUT_2[17348] = 32'b11111111111111111101010100100101;
assign LUT_2[17349] = 32'b11111111111111111010001100111110;
assign LUT_2[17350] = 32'b00000000000000000100001101100001;
assign LUT_2[17351] = 32'b00000000000000000001000101111010;
assign LUT_2[17352] = 32'b11111111111111111011101000011010;
assign LUT_2[17353] = 32'b11111111111111111000100000110011;
assign LUT_2[17354] = 32'b00000000000000000010100001010110;
assign LUT_2[17355] = 32'b11111111111111111111011001101111;
assign LUT_2[17356] = 32'b11111111111111111000000110000010;
assign LUT_2[17357] = 32'b11111111111111110100111110011011;
assign LUT_2[17358] = 32'b11111111111111111110111110111110;
assign LUT_2[17359] = 32'b11111111111111111011110111010111;
assign LUT_2[17360] = 32'b11111111111111111011011011000111;
assign LUT_2[17361] = 32'b11111111111111111000010011100000;
assign LUT_2[17362] = 32'b00000000000000000010010100000011;
assign LUT_2[17363] = 32'b11111111111111111111001100011100;
assign LUT_2[17364] = 32'b11111111111111110111111000101111;
assign LUT_2[17365] = 32'b11111111111111110100110001001000;
assign LUT_2[17366] = 32'b11111111111111111110110001101011;
assign LUT_2[17367] = 32'b11111111111111111011101010000100;
assign LUT_2[17368] = 32'b11111111111111110110001100100100;
assign LUT_2[17369] = 32'b11111111111111110011000100111101;
assign LUT_2[17370] = 32'b11111111111111111101000101100000;
assign LUT_2[17371] = 32'b11111111111111111001111101111001;
assign LUT_2[17372] = 32'b11111111111111110010101010001100;
assign LUT_2[17373] = 32'b11111111111111101111100010100101;
assign LUT_2[17374] = 32'b11111111111111111001100011001000;
assign LUT_2[17375] = 32'b11111111111111110110011011100001;
assign LUT_2[17376] = 32'b00000000000000000001010010100110;
assign LUT_2[17377] = 32'b11111111111111111110001010111111;
assign LUT_2[17378] = 32'b00000000000000001000001011100010;
assign LUT_2[17379] = 32'b00000000000000000101000011111011;
assign LUT_2[17380] = 32'b11111111111111111101110000001110;
assign LUT_2[17381] = 32'b11111111111111111010101000100111;
assign LUT_2[17382] = 32'b00000000000000000100101001001010;
assign LUT_2[17383] = 32'b00000000000000000001100001100011;
assign LUT_2[17384] = 32'b11111111111111111100000100000011;
assign LUT_2[17385] = 32'b11111111111111111000111100011100;
assign LUT_2[17386] = 32'b00000000000000000010111100111111;
assign LUT_2[17387] = 32'b11111111111111111111110101011000;
assign LUT_2[17388] = 32'b11111111111111111000100001101011;
assign LUT_2[17389] = 32'b11111111111111110101011010000100;
assign LUT_2[17390] = 32'b11111111111111111111011010100111;
assign LUT_2[17391] = 32'b11111111111111111100010011000000;
assign LUT_2[17392] = 32'b11111111111111111011110110110000;
assign LUT_2[17393] = 32'b11111111111111111000101111001001;
assign LUT_2[17394] = 32'b00000000000000000010101111101100;
assign LUT_2[17395] = 32'b11111111111111111111101000000101;
assign LUT_2[17396] = 32'b11111111111111111000010100011000;
assign LUT_2[17397] = 32'b11111111111111110101001100110001;
assign LUT_2[17398] = 32'b11111111111111111111001101010100;
assign LUT_2[17399] = 32'b11111111111111111100000101101101;
assign LUT_2[17400] = 32'b11111111111111110110101000001101;
assign LUT_2[17401] = 32'b11111111111111110011100000100110;
assign LUT_2[17402] = 32'b11111111111111111101100001001001;
assign LUT_2[17403] = 32'b11111111111111111010011001100010;
assign LUT_2[17404] = 32'b11111111111111110011000101110101;
assign LUT_2[17405] = 32'b11111111111111101111111110001110;
assign LUT_2[17406] = 32'b11111111111111111001111110110001;
assign LUT_2[17407] = 32'b11111111111111110110110111001010;
assign LUT_2[17408] = 32'b00000000000000000010010101111000;
assign LUT_2[17409] = 32'b11111111111111111111001110010001;
assign LUT_2[17410] = 32'b00000000000000001001001110110100;
assign LUT_2[17411] = 32'b00000000000000000110000111001101;
assign LUT_2[17412] = 32'b11111111111111111110110011100000;
assign LUT_2[17413] = 32'b11111111111111111011101011111001;
assign LUT_2[17414] = 32'b00000000000000000101101100011100;
assign LUT_2[17415] = 32'b00000000000000000010100100110101;
assign LUT_2[17416] = 32'b11111111111111111101000111010101;
assign LUT_2[17417] = 32'b11111111111111111001111111101110;
assign LUT_2[17418] = 32'b00000000000000000100000000010001;
assign LUT_2[17419] = 32'b00000000000000000000111000101010;
assign LUT_2[17420] = 32'b11111111111111111001100100111101;
assign LUT_2[17421] = 32'b11111111111111110110011101010110;
assign LUT_2[17422] = 32'b00000000000000000000011101111001;
assign LUT_2[17423] = 32'b11111111111111111101010110010010;
assign LUT_2[17424] = 32'b11111111111111111100111010000010;
assign LUT_2[17425] = 32'b11111111111111111001110010011011;
assign LUT_2[17426] = 32'b00000000000000000011110010111110;
assign LUT_2[17427] = 32'b00000000000000000000101011010111;
assign LUT_2[17428] = 32'b11111111111111111001010111101010;
assign LUT_2[17429] = 32'b11111111111111110110010000000011;
assign LUT_2[17430] = 32'b00000000000000000000010000100110;
assign LUT_2[17431] = 32'b11111111111111111101001000111111;
assign LUT_2[17432] = 32'b11111111111111110111101011011111;
assign LUT_2[17433] = 32'b11111111111111110100100011111000;
assign LUT_2[17434] = 32'b11111111111111111110100100011011;
assign LUT_2[17435] = 32'b11111111111111111011011100110100;
assign LUT_2[17436] = 32'b11111111111111110100001001000111;
assign LUT_2[17437] = 32'b11111111111111110001000001100000;
assign LUT_2[17438] = 32'b11111111111111111011000010000011;
assign LUT_2[17439] = 32'b11111111111111110111111010011100;
assign LUT_2[17440] = 32'b00000000000000000010110001100001;
assign LUT_2[17441] = 32'b11111111111111111111101001111010;
assign LUT_2[17442] = 32'b00000000000000001001101010011101;
assign LUT_2[17443] = 32'b00000000000000000110100010110110;
assign LUT_2[17444] = 32'b11111111111111111111001111001001;
assign LUT_2[17445] = 32'b11111111111111111100000111100010;
assign LUT_2[17446] = 32'b00000000000000000110001000000101;
assign LUT_2[17447] = 32'b00000000000000000011000000011110;
assign LUT_2[17448] = 32'b11111111111111111101100010111110;
assign LUT_2[17449] = 32'b11111111111111111010011011010111;
assign LUT_2[17450] = 32'b00000000000000000100011011111010;
assign LUT_2[17451] = 32'b00000000000000000001010100010011;
assign LUT_2[17452] = 32'b11111111111111111010000000100110;
assign LUT_2[17453] = 32'b11111111111111110110111000111111;
assign LUT_2[17454] = 32'b00000000000000000000111001100010;
assign LUT_2[17455] = 32'b11111111111111111101110001111011;
assign LUT_2[17456] = 32'b11111111111111111101010101101011;
assign LUT_2[17457] = 32'b11111111111111111010001110000100;
assign LUT_2[17458] = 32'b00000000000000000100001110100111;
assign LUT_2[17459] = 32'b00000000000000000001000111000000;
assign LUT_2[17460] = 32'b11111111111111111001110011010011;
assign LUT_2[17461] = 32'b11111111111111110110101011101100;
assign LUT_2[17462] = 32'b00000000000000000000101100001111;
assign LUT_2[17463] = 32'b11111111111111111101100100101000;
assign LUT_2[17464] = 32'b11111111111111111000000111001000;
assign LUT_2[17465] = 32'b11111111111111110100111111100001;
assign LUT_2[17466] = 32'b11111111111111111111000000000100;
assign LUT_2[17467] = 32'b11111111111111111011111000011101;
assign LUT_2[17468] = 32'b11111111111111110100100100110000;
assign LUT_2[17469] = 32'b11111111111111110001011101001001;
assign LUT_2[17470] = 32'b11111111111111111011011101101100;
assign LUT_2[17471] = 32'b11111111111111111000010110000101;
assign LUT_2[17472] = 32'b11111111111111111010011110011011;
assign LUT_2[17473] = 32'b11111111111111110111010110110100;
assign LUT_2[17474] = 32'b00000000000000000001010111010111;
assign LUT_2[17475] = 32'b11111111111111111110001111110000;
assign LUT_2[17476] = 32'b11111111111111110110111100000011;
assign LUT_2[17477] = 32'b11111111111111110011110100011100;
assign LUT_2[17478] = 32'b11111111111111111101110100111111;
assign LUT_2[17479] = 32'b11111111111111111010101101011000;
assign LUT_2[17480] = 32'b11111111111111110101001111111000;
assign LUT_2[17481] = 32'b11111111111111110010001000010001;
assign LUT_2[17482] = 32'b11111111111111111100001000110100;
assign LUT_2[17483] = 32'b11111111111111111001000001001101;
assign LUT_2[17484] = 32'b11111111111111110001101101100000;
assign LUT_2[17485] = 32'b11111111111111101110100101111001;
assign LUT_2[17486] = 32'b11111111111111111000100110011100;
assign LUT_2[17487] = 32'b11111111111111110101011110110101;
assign LUT_2[17488] = 32'b11111111111111110101000010100101;
assign LUT_2[17489] = 32'b11111111111111110001111010111110;
assign LUT_2[17490] = 32'b11111111111111111011111011100001;
assign LUT_2[17491] = 32'b11111111111111111000110011111010;
assign LUT_2[17492] = 32'b11111111111111110001100000001101;
assign LUT_2[17493] = 32'b11111111111111101110011000100110;
assign LUT_2[17494] = 32'b11111111111111111000011001001001;
assign LUT_2[17495] = 32'b11111111111111110101010001100010;
assign LUT_2[17496] = 32'b11111111111111101111110100000010;
assign LUT_2[17497] = 32'b11111111111111101100101100011011;
assign LUT_2[17498] = 32'b11111111111111110110101100111110;
assign LUT_2[17499] = 32'b11111111111111110011100101010111;
assign LUT_2[17500] = 32'b11111111111111101100010001101010;
assign LUT_2[17501] = 32'b11111111111111101001001010000011;
assign LUT_2[17502] = 32'b11111111111111110011001010100110;
assign LUT_2[17503] = 32'b11111111111111110000000010111111;
assign LUT_2[17504] = 32'b11111111111111111010111010000100;
assign LUT_2[17505] = 32'b11111111111111110111110010011101;
assign LUT_2[17506] = 32'b00000000000000000001110011000000;
assign LUT_2[17507] = 32'b11111111111111111110101011011001;
assign LUT_2[17508] = 32'b11111111111111110111010111101100;
assign LUT_2[17509] = 32'b11111111111111110100010000000101;
assign LUT_2[17510] = 32'b11111111111111111110010000101000;
assign LUT_2[17511] = 32'b11111111111111111011001001000001;
assign LUT_2[17512] = 32'b11111111111111110101101011100001;
assign LUT_2[17513] = 32'b11111111111111110010100011111010;
assign LUT_2[17514] = 32'b11111111111111111100100100011101;
assign LUT_2[17515] = 32'b11111111111111111001011100110110;
assign LUT_2[17516] = 32'b11111111111111110010001001001001;
assign LUT_2[17517] = 32'b11111111111111101111000001100010;
assign LUT_2[17518] = 32'b11111111111111111001000010000101;
assign LUT_2[17519] = 32'b11111111111111110101111010011110;
assign LUT_2[17520] = 32'b11111111111111110101011110001110;
assign LUT_2[17521] = 32'b11111111111111110010010110100111;
assign LUT_2[17522] = 32'b11111111111111111100010111001010;
assign LUT_2[17523] = 32'b11111111111111111001001111100011;
assign LUT_2[17524] = 32'b11111111111111110001111011110110;
assign LUT_2[17525] = 32'b11111111111111101110110100001111;
assign LUT_2[17526] = 32'b11111111111111111000110100110010;
assign LUT_2[17527] = 32'b11111111111111110101101101001011;
assign LUT_2[17528] = 32'b11111111111111110000001111101011;
assign LUT_2[17529] = 32'b11111111111111101101001000000100;
assign LUT_2[17530] = 32'b11111111111111110111001000100111;
assign LUT_2[17531] = 32'b11111111111111110100000001000000;
assign LUT_2[17532] = 32'b11111111111111101100101101010011;
assign LUT_2[17533] = 32'b11111111111111101001100101101100;
assign LUT_2[17534] = 32'b11111111111111110011100110001111;
assign LUT_2[17535] = 32'b11111111111111110000011110101000;
assign LUT_2[17536] = 32'b00000000000000000110101010000111;
assign LUT_2[17537] = 32'b00000000000000000011100010100000;
assign LUT_2[17538] = 32'b00000000000000001101100011000011;
assign LUT_2[17539] = 32'b00000000000000001010011011011100;
assign LUT_2[17540] = 32'b00000000000000000011000111101111;
assign LUT_2[17541] = 32'b00000000000000000000000000001000;
assign LUT_2[17542] = 32'b00000000000000001010000000101011;
assign LUT_2[17543] = 32'b00000000000000000110111001000100;
assign LUT_2[17544] = 32'b00000000000000000001011011100100;
assign LUT_2[17545] = 32'b11111111111111111110010011111101;
assign LUT_2[17546] = 32'b00000000000000001000010100100000;
assign LUT_2[17547] = 32'b00000000000000000101001100111001;
assign LUT_2[17548] = 32'b11111111111111111101111001001100;
assign LUT_2[17549] = 32'b11111111111111111010110001100101;
assign LUT_2[17550] = 32'b00000000000000000100110010001000;
assign LUT_2[17551] = 32'b00000000000000000001101010100001;
assign LUT_2[17552] = 32'b00000000000000000001001110010001;
assign LUT_2[17553] = 32'b11111111111111111110000110101010;
assign LUT_2[17554] = 32'b00000000000000001000000111001101;
assign LUT_2[17555] = 32'b00000000000000000100111111100110;
assign LUT_2[17556] = 32'b11111111111111111101101011111001;
assign LUT_2[17557] = 32'b11111111111111111010100100010010;
assign LUT_2[17558] = 32'b00000000000000000100100100110101;
assign LUT_2[17559] = 32'b00000000000000000001011101001110;
assign LUT_2[17560] = 32'b11111111111111111011111111101110;
assign LUT_2[17561] = 32'b11111111111111111000111000000111;
assign LUT_2[17562] = 32'b00000000000000000010111000101010;
assign LUT_2[17563] = 32'b11111111111111111111110001000011;
assign LUT_2[17564] = 32'b11111111111111111000011101010110;
assign LUT_2[17565] = 32'b11111111111111110101010101101111;
assign LUT_2[17566] = 32'b11111111111111111111010110010010;
assign LUT_2[17567] = 32'b11111111111111111100001110101011;
assign LUT_2[17568] = 32'b00000000000000000111000101110000;
assign LUT_2[17569] = 32'b00000000000000000011111110001001;
assign LUT_2[17570] = 32'b00000000000000001101111110101100;
assign LUT_2[17571] = 32'b00000000000000001010110111000101;
assign LUT_2[17572] = 32'b00000000000000000011100011011000;
assign LUT_2[17573] = 32'b00000000000000000000011011110001;
assign LUT_2[17574] = 32'b00000000000000001010011100010100;
assign LUT_2[17575] = 32'b00000000000000000111010100101101;
assign LUT_2[17576] = 32'b00000000000000000001110111001101;
assign LUT_2[17577] = 32'b11111111111111111110101111100110;
assign LUT_2[17578] = 32'b00000000000000001000110000001001;
assign LUT_2[17579] = 32'b00000000000000000101101000100010;
assign LUT_2[17580] = 32'b11111111111111111110010100110101;
assign LUT_2[17581] = 32'b11111111111111111011001101001110;
assign LUT_2[17582] = 32'b00000000000000000101001101110001;
assign LUT_2[17583] = 32'b00000000000000000010000110001010;
assign LUT_2[17584] = 32'b00000000000000000001101001111010;
assign LUT_2[17585] = 32'b11111111111111111110100010010011;
assign LUT_2[17586] = 32'b00000000000000001000100010110110;
assign LUT_2[17587] = 32'b00000000000000000101011011001111;
assign LUT_2[17588] = 32'b11111111111111111110000111100010;
assign LUT_2[17589] = 32'b11111111111111111010111111111011;
assign LUT_2[17590] = 32'b00000000000000000101000000011110;
assign LUT_2[17591] = 32'b00000000000000000001111000110111;
assign LUT_2[17592] = 32'b11111111111111111100011011010111;
assign LUT_2[17593] = 32'b11111111111111111001010011110000;
assign LUT_2[17594] = 32'b00000000000000000011010100010011;
assign LUT_2[17595] = 32'b00000000000000000000001100101100;
assign LUT_2[17596] = 32'b11111111111111111000111000111111;
assign LUT_2[17597] = 32'b11111111111111110101110001011000;
assign LUT_2[17598] = 32'b11111111111111111111110001111011;
assign LUT_2[17599] = 32'b11111111111111111100101010010100;
assign LUT_2[17600] = 32'b11111111111111111110110010101010;
assign LUT_2[17601] = 32'b11111111111111111011101011000011;
assign LUT_2[17602] = 32'b00000000000000000101101011100110;
assign LUT_2[17603] = 32'b00000000000000000010100011111111;
assign LUT_2[17604] = 32'b11111111111111111011010000010010;
assign LUT_2[17605] = 32'b11111111111111111000001000101011;
assign LUT_2[17606] = 32'b00000000000000000010001001001110;
assign LUT_2[17607] = 32'b11111111111111111111000001100111;
assign LUT_2[17608] = 32'b11111111111111111001100100000111;
assign LUT_2[17609] = 32'b11111111111111110110011100100000;
assign LUT_2[17610] = 32'b00000000000000000000011101000011;
assign LUT_2[17611] = 32'b11111111111111111101010101011100;
assign LUT_2[17612] = 32'b11111111111111110110000001101111;
assign LUT_2[17613] = 32'b11111111111111110010111010001000;
assign LUT_2[17614] = 32'b11111111111111111100111010101011;
assign LUT_2[17615] = 32'b11111111111111111001110011000100;
assign LUT_2[17616] = 32'b11111111111111111001010110110100;
assign LUT_2[17617] = 32'b11111111111111110110001111001101;
assign LUT_2[17618] = 32'b00000000000000000000001111110000;
assign LUT_2[17619] = 32'b11111111111111111101001000001001;
assign LUT_2[17620] = 32'b11111111111111110101110100011100;
assign LUT_2[17621] = 32'b11111111111111110010101100110101;
assign LUT_2[17622] = 32'b11111111111111111100101101011000;
assign LUT_2[17623] = 32'b11111111111111111001100101110001;
assign LUT_2[17624] = 32'b11111111111111110100001000010001;
assign LUT_2[17625] = 32'b11111111111111110001000000101010;
assign LUT_2[17626] = 32'b11111111111111111011000001001101;
assign LUT_2[17627] = 32'b11111111111111110111111001100110;
assign LUT_2[17628] = 32'b11111111111111110000100101111001;
assign LUT_2[17629] = 32'b11111111111111101101011110010010;
assign LUT_2[17630] = 32'b11111111111111110111011110110101;
assign LUT_2[17631] = 32'b11111111111111110100010111001110;
assign LUT_2[17632] = 32'b11111111111111111111001110010011;
assign LUT_2[17633] = 32'b11111111111111111100000110101100;
assign LUT_2[17634] = 32'b00000000000000000110000111001111;
assign LUT_2[17635] = 32'b00000000000000000010111111101000;
assign LUT_2[17636] = 32'b11111111111111111011101011111011;
assign LUT_2[17637] = 32'b11111111111111111000100100010100;
assign LUT_2[17638] = 32'b00000000000000000010100100110111;
assign LUT_2[17639] = 32'b11111111111111111111011101010000;
assign LUT_2[17640] = 32'b11111111111111111001111111110000;
assign LUT_2[17641] = 32'b11111111111111110110111000001001;
assign LUT_2[17642] = 32'b00000000000000000000111000101100;
assign LUT_2[17643] = 32'b11111111111111111101110001000101;
assign LUT_2[17644] = 32'b11111111111111110110011101011000;
assign LUT_2[17645] = 32'b11111111111111110011010101110001;
assign LUT_2[17646] = 32'b11111111111111111101010110010100;
assign LUT_2[17647] = 32'b11111111111111111010001110101101;
assign LUT_2[17648] = 32'b11111111111111111001110010011101;
assign LUT_2[17649] = 32'b11111111111111110110101010110110;
assign LUT_2[17650] = 32'b00000000000000000000101011011001;
assign LUT_2[17651] = 32'b11111111111111111101100011110010;
assign LUT_2[17652] = 32'b11111111111111110110010000000101;
assign LUT_2[17653] = 32'b11111111111111110011001000011110;
assign LUT_2[17654] = 32'b11111111111111111101001001000001;
assign LUT_2[17655] = 32'b11111111111111111010000001011010;
assign LUT_2[17656] = 32'b11111111111111110100100011111010;
assign LUT_2[17657] = 32'b11111111111111110001011100010011;
assign LUT_2[17658] = 32'b11111111111111111011011100110110;
assign LUT_2[17659] = 32'b11111111111111111000010101001111;
assign LUT_2[17660] = 32'b11111111111111110001000001100010;
assign LUT_2[17661] = 32'b11111111111111101101111001111011;
assign LUT_2[17662] = 32'b11111111111111110111111010011110;
assign LUT_2[17663] = 32'b11111111111111110100110010110111;
assign LUT_2[17664] = 32'b00000000000000000110010100011110;
assign LUT_2[17665] = 32'b00000000000000000011001100110111;
assign LUT_2[17666] = 32'b00000000000000001101001101011010;
assign LUT_2[17667] = 32'b00000000000000001010000101110011;
assign LUT_2[17668] = 32'b00000000000000000010110010000110;
assign LUT_2[17669] = 32'b11111111111111111111101010011111;
assign LUT_2[17670] = 32'b00000000000000001001101011000010;
assign LUT_2[17671] = 32'b00000000000000000110100011011011;
assign LUT_2[17672] = 32'b00000000000000000001000101111011;
assign LUT_2[17673] = 32'b11111111111111111101111110010100;
assign LUT_2[17674] = 32'b00000000000000000111111110110111;
assign LUT_2[17675] = 32'b00000000000000000100110111010000;
assign LUT_2[17676] = 32'b11111111111111111101100011100011;
assign LUT_2[17677] = 32'b11111111111111111010011011111100;
assign LUT_2[17678] = 32'b00000000000000000100011100011111;
assign LUT_2[17679] = 32'b00000000000000000001010100111000;
assign LUT_2[17680] = 32'b00000000000000000000111000101000;
assign LUT_2[17681] = 32'b11111111111111111101110001000001;
assign LUT_2[17682] = 32'b00000000000000000111110001100100;
assign LUT_2[17683] = 32'b00000000000000000100101001111101;
assign LUT_2[17684] = 32'b11111111111111111101010110010000;
assign LUT_2[17685] = 32'b11111111111111111010001110101001;
assign LUT_2[17686] = 32'b00000000000000000100001111001100;
assign LUT_2[17687] = 32'b00000000000000000001000111100101;
assign LUT_2[17688] = 32'b11111111111111111011101010000101;
assign LUT_2[17689] = 32'b11111111111111111000100010011110;
assign LUT_2[17690] = 32'b00000000000000000010100011000001;
assign LUT_2[17691] = 32'b11111111111111111111011011011010;
assign LUT_2[17692] = 32'b11111111111111111000000111101101;
assign LUT_2[17693] = 32'b11111111111111110101000000000110;
assign LUT_2[17694] = 32'b11111111111111111111000000101001;
assign LUT_2[17695] = 32'b11111111111111111011111001000010;
assign LUT_2[17696] = 32'b00000000000000000110110000000111;
assign LUT_2[17697] = 32'b00000000000000000011101000100000;
assign LUT_2[17698] = 32'b00000000000000001101101001000011;
assign LUT_2[17699] = 32'b00000000000000001010100001011100;
assign LUT_2[17700] = 32'b00000000000000000011001101101111;
assign LUT_2[17701] = 32'b00000000000000000000000110001000;
assign LUT_2[17702] = 32'b00000000000000001010000110101011;
assign LUT_2[17703] = 32'b00000000000000000110111111000100;
assign LUT_2[17704] = 32'b00000000000000000001100001100100;
assign LUT_2[17705] = 32'b11111111111111111110011001111101;
assign LUT_2[17706] = 32'b00000000000000001000011010100000;
assign LUT_2[17707] = 32'b00000000000000000101010010111001;
assign LUT_2[17708] = 32'b11111111111111111101111111001100;
assign LUT_2[17709] = 32'b11111111111111111010110111100101;
assign LUT_2[17710] = 32'b00000000000000000100111000001000;
assign LUT_2[17711] = 32'b00000000000000000001110000100001;
assign LUT_2[17712] = 32'b00000000000000000001010100010001;
assign LUT_2[17713] = 32'b11111111111111111110001100101010;
assign LUT_2[17714] = 32'b00000000000000001000001101001101;
assign LUT_2[17715] = 32'b00000000000000000101000101100110;
assign LUT_2[17716] = 32'b11111111111111111101110001111001;
assign LUT_2[17717] = 32'b11111111111111111010101010010010;
assign LUT_2[17718] = 32'b00000000000000000100101010110101;
assign LUT_2[17719] = 32'b00000000000000000001100011001110;
assign LUT_2[17720] = 32'b11111111111111111100000101101110;
assign LUT_2[17721] = 32'b11111111111111111000111110000111;
assign LUT_2[17722] = 32'b00000000000000000010111110101010;
assign LUT_2[17723] = 32'b11111111111111111111110111000011;
assign LUT_2[17724] = 32'b11111111111111111000100011010110;
assign LUT_2[17725] = 32'b11111111111111110101011011101111;
assign LUT_2[17726] = 32'b11111111111111111111011100010010;
assign LUT_2[17727] = 32'b11111111111111111100010100101011;
assign LUT_2[17728] = 32'b11111111111111111110011101000001;
assign LUT_2[17729] = 32'b11111111111111111011010101011010;
assign LUT_2[17730] = 32'b00000000000000000101010101111101;
assign LUT_2[17731] = 32'b00000000000000000010001110010110;
assign LUT_2[17732] = 32'b11111111111111111010111010101001;
assign LUT_2[17733] = 32'b11111111111111110111110011000010;
assign LUT_2[17734] = 32'b00000000000000000001110011100101;
assign LUT_2[17735] = 32'b11111111111111111110101011111110;
assign LUT_2[17736] = 32'b11111111111111111001001110011110;
assign LUT_2[17737] = 32'b11111111111111110110000110110111;
assign LUT_2[17738] = 32'b00000000000000000000000111011010;
assign LUT_2[17739] = 32'b11111111111111111100111111110011;
assign LUT_2[17740] = 32'b11111111111111110101101100000110;
assign LUT_2[17741] = 32'b11111111111111110010100100011111;
assign LUT_2[17742] = 32'b11111111111111111100100101000010;
assign LUT_2[17743] = 32'b11111111111111111001011101011011;
assign LUT_2[17744] = 32'b11111111111111111001000001001011;
assign LUT_2[17745] = 32'b11111111111111110101111001100100;
assign LUT_2[17746] = 32'b11111111111111111111111010000111;
assign LUT_2[17747] = 32'b11111111111111111100110010100000;
assign LUT_2[17748] = 32'b11111111111111110101011110110011;
assign LUT_2[17749] = 32'b11111111111111110010010111001100;
assign LUT_2[17750] = 32'b11111111111111111100010111101111;
assign LUT_2[17751] = 32'b11111111111111111001010000001000;
assign LUT_2[17752] = 32'b11111111111111110011110010101000;
assign LUT_2[17753] = 32'b11111111111111110000101011000001;
assign LUT_2[17754] = 32'b11111111111111111010101011100100;
assign LUT_2[17755] = 32'b11111111111111110111100011111101;
assign LUT_2[17756] = 32'b11111111111111110000010000010000;
assign LUT_2[17757] = 32'b11111111111111101101001000101001;
assign LUT_2[17758] = 32'b11111111111111110111001001001100;
assign LUT_2[17759] = 32'b11111111111111110100000001100101;
assign LUT_2[17760] = 32'b11111111111111111110111000101010;
assign LUT_2[17761] = 32'b11111111111111111011110001000011;
assign LUT_2[17762] = 32'b00000000000000000101110001100110;
assign LUT_2[17763] = 32'b00000000000000000010101001111111;
assign LUT_2[17764] = 32'b11111111111111111011010110010010;
assign LUT_2[17765] = 32'b11111111111111111000001110101011;
assign LUT_2[17766] = 32'b00000000000000000010001111001110;
assign LUT_2[17767] = 32'b11111111111111111111000111100111;
assign LUT_2[17768] = 32'b11111111111111111001101010000111;
assign LUT_2[17769] = 32'b11111111111111110110100010100000;
assign LUT_2[17770] = 32'b00000000000000000000100011000011;
assign LUT_2[17771] = 32'b11111111111111111101011011011100;
assign LUT_2[17772] = 32'b11111111111111110110000111101111;
assign LUT_2[17773] = 32'b11111111111111110011000000001000;
assign LUT_2[17774] = 32'b11111111111111111101000000101011;
assign LUT_2[17775] = 32'b11111111111111111001111001000100;
assign LUT_2[17776] = 32'b11111111111111111001011100110100;
assign LUT_2[17777] = 32'b11111111111111110110010101001101;
assign LUT_2[17778] = 32'b00000000000000000000010101110000;
assign LUT_2[17779] = 32'b11111111111111111101001110001001;
assign LUT_2[17780] = 32'b11111111111111110101111010011100;
assign LUT_2[17781] = 32'b11111111111111110010110010110101;
assign LUT_2[17782] = 32'b11111111111111111100110011011000;
assign LUT_2[17783] = 32'b11111111111111111001101011110001;
assign LUT_2[17784] = 32'b11111111111111110100001110010001;
assign LUT_2[17785] = 32'b11111111111111110001000110101010;
assign LUT_2[17786] = 32'b11111111111111111011000111001101;
assign LUT_2[17787] = 32'b11111111111111110111111111100110;
assign LUT_2[17788] = 32'b11111111111111110000101011111001;
assign LUT_2[17789] = 32'b11111111111111101101100100010010;
assign LUT_2[17790] = 32'b11111111111111110111100100110101;
assign LUT_2[17791] = 32'b11111111111111110100011101001110;
assign LUT_2[17792] = 32'b00000000000000001010101000101101;
assign LUT_2[17793] = 32'b00000000000000000111100001000110;
assign LUT_2[17794] = 32'b00000000000000010001100001101001;
assign LUT_2[17795] = 32'b00000000000000001110011010000010;
assign LUT_2[17796] = 32'b00000000000000000111000110010101;
assign LUT_2[17797] = 32'b00000000000000000011111110101110;
assign LUT_2[17798] = 32'b00000000000000001101111111010001;
assign LUT_2[17799] = 32'b00000000000000001010110111101010;
assign LUT_2[17800] = 32'b00000000000000000101011010001010;
assign LUT_2[17801] = 32'b00000000000000000010010010100011;
assign LUT_2[17802] = 32'b00000000000000001100010011000110;
assign LUT_2[17803] = 32'b00000000000000001001001011011111;
assign LUT_2[17804] = 32'b00000000000000000001110111110010;
assign LUT_2[17805] = 32'b11111111111111111110110000001011;
assign LUT_2[17806] = 32'b00000000000000001000110000101110;
assign LUT_2[17807] = 32'b00000000000000000101101001000111;
assign LUT_2[17808] = 32'b00000000000000000101001100110111;
assign LUT_2[17809] = 32'b00000000000000000010000101010000;
assign LUT_2[17810] = 32'b00000000000000001100000101110011;
assign LUT_2[17811] = 32'b00000000000000001000111110001100;
assign LUT_2[17812] = 32'b00000000000000000001101010011111;
assign LUT_2[17813] = 32'b11111111111111111110100010111000;
assign LUT_2[17814] = 32'b00000000000000001000100011011011;
assign LUT_2[17815] = 32'b00000000000000000101011011110100;
assign LUT_2[17816] = 32'b11111111111111111111111110010100;
assign LUT_2[17817] = 32'b11111111111111111100110110101101;
assign LUT_2[17818] = 32'b00000000000000000110110111010000;
assign LUT_2[17819] = 32'b00000000000000000011101111101001;
assign LUT_2[17820] = 32'b11111111111111111100011011111100;
assign LUT_2[17821] = 32'b11111111111111111001010100010101;
assign LUT_2[17822] = 32'b00000000000000000011010100111000;
assign LUT_2[17823] = 32'b00000000000000000000001101010001;
assign LUT_2[17824] = 32'b00000000000000001011000100010110;
assign LUT_2[17825] = 32'b00000000000000000111111100101111;
assign LUT_2[17826] = 32'b00000000000000010001111101010010;
assign LUT_2[17827] = 32'b00000000000000001110110101101011;
assign LUT_2[17828] = 32'b00000000000000000111100001111110;
assign LUT_2[17829] = 32'b00000000000000000100011010010111;
assign LUT_2[17830] = 32'b00000000000000001110011010111010;
assign LUT_2[17831] = 32'b00000000000000001011010011010011;
assign LUT_2[17832] = 32'b00000000000000000101110101110011;
assign LUT_2[17833] = 32'b00000000000000000010101110001100;
assign LUT_2[17834] = 32'b00000000000000001100101110101111;
assign LUT_2[17835] = 32'b00000000000000001001100111001000;
assign LUT_2[17836] = 32'b00000000000000000010010011011011;
assign LUT_2[17837] = 32'b11111111111111111111001011110100;
assign LUT_2[17838] = 32'b00000000000000001001001100010111;
assign LUT_2[17839] = 32'b00000000000000000110000100110000;
assign LUT_2[17840] = 32'b00000000000000000101101000100000;
assign LUT_2[17841] = 32'b00000000000000000010100000111001;
assign LUT_2[17842] = 32'b00000000000000001100100001011100;
assign LUT_2[17843] = 32'b00000000000000001001011001110101;
assign LUT_2[17844] = 32'b00000000000000000010000110001000;
assign LUT_2[17845] = 32'b11111111111111111110111110100001;
assign LUT_2[17846] = 32'b00000000000000001000111111000100;
assign LUT_2[17847] = 32'b00000000000000000101110111011101;
assign LUT_2[17848] = 32'b00000000000000000000011001111101;
assign LUT_2[17849] = 32'b11111111111111111101010010010110;
assign LUT_2[17850] = 32'b00000000000000000111010010111001;
assign LUT_2[17851] = 32'b00000000000000000100001011010010;
assign LUT_2[17852] = 32'b11111111111111111100110111100101;
assign LUT_2[17853] = 32'b11111111111111111001101111111110;
assign LUT_2[17854] = 32'b00000000000000000011110000100001;
assign LUT_2[17855] = 32'b00000000000000000000101000111010;
assign LUT_2[17856] = 32'b00000000000000000010110001010000;
assign LUT_2[17857] = 32'b11111111111111111111101001101001;
assign LUT_2[17858] = 32'b00000000000000001001101010001100;
assign LUT_2[17859] = 32'b00000000000000000110100010100101;
assign LUT_2[17860] = 32'b11111111111111111111001110111000;
assign LUT_2[17861] = 32'b11111111111111111100000111010001;
assign LUT_2[17862] = 32'b00000000000000000110000111110100;
assign LUT_2[17863] = 32'b00000000000000000011000000001101;
assign LUT_2[17864] = 32'b11111111111111111101100010101101;
assign LUT_2[17865] = 32'b11111111111111111010011011000110;
assign LUT_2[17866] = 32'b00000000000000000100011011101001;
assign LUT_2[17867] = 32'b00000000000000000001010100000010;
assign LUT_2[17868] = 32'b11111111111111111010000000010101;
assign LUT_2[17869] = 32'b11111111111111110110111000101110;
assign LUT_2[17870] = 32'b00000000000000000000111001010001;
assign LUT_2[17871] = 32'b11111111111111111101110001101010;
assign LUT_2[17872] = 32'b11111111111111111101010101011010;
assign LUT_2[17873] = 32'b11111111111111111010001101110011;
assign LUT_2[17874] = 32'b00000000000000000100001110010110;
assign LUT_2[17875] = 32'b00000000000000000001000110101111;
assign LUT_2[17876] = 32'b11111111111111111001110011000010;
assign LUT_2[17877] = 32'b11111111111111110110101011011011;
assign LUT_2[17878] = 32'b00000000000000000000101011111110;
assign LUT_2[17879] = 32'b11111111111111111101100100010111;
assign LUT_2[17880] = 32'b11111111111111111000000110110111;
assign LUT_2[17881] = 32'b11111111111111110100111111010000;
assign LUT_2[17882] = 32'b11111111111111111110111111110011;
assign LUT_2[17883] = 32'b11111111111111111011111000001100;
assign LUT_2[17884] = 32'b11111111111111110100100100011111;
assign LUT_2[17885] = 32'b11111111111111110001011100111000;
assign LUT_2[17886] = 32'b11111111111111111011011101011011;
assign LUT_2[17887] = 32'b11111111111111111000010101110100;
assign LUT_2[17888] = 32'b00000000000000000011001100111001;
assign LUT_2[17889] = 32'b00000000000000000000000101010010;
assign LUT_2[17890] = 32'b00000000000000001010000101110101;
assign LUT_2[17891] = 32'b00000000000000000110111110001110;
assign LUT_2[17892] = 32'b11111111111111111111101010100001;
assign LUT_2[17893] = 32'b11111111111111111100100010111010;
assign LUT_2[17894] = 32'b00000000000000000110100011011101;
assign LUT_2[17895] = 32'b00000000000000000011011011110110;
assign LUT_2[17896] = 32'b11111111111111111101111110010110;
assign LUT_2[17897] = 32'b11111111111111111010110110101111;
assign LUT_2[17898] = 32'b00000000000000000100110111010010;
assign LUT_2[17899] = 32'b00000000000000000001101111101011;
assign LUT_2[17900] = 32'b11111111111111111010011011111110;
assign LUT_2[17901] = 32'b11111111111111110111010100010111;
assign LUT_2[17902] = 32'b00000000000000000001010100111010;
assign LUT_2[17903] = 32'b11111111111111111110001101010011;
assign LUT_2[17904] = 32'b11111111111111111101110001000011;
assign LUT_2[17905] = 32'b11111111111111111010101001011100;
assign LUT_2[17906] = 32'b00000000000000000100101001111111;
assign LUT_2[17907] = 32'b00000000000000000001100010011000;
assign LUT_2[17908] = 32'b11111111111111111010001110101011;
assign LUT_2[17909] = 32'b11111111111111110111000111000100;
assign LUT_2[17910] = 32'b00000000000000000001000111100111;
assign LUT_2[17911] = 32'b11111111111111111110000000000000;
assign LUT_2[17912] = 32'b11111111111111111000100010100000;
assign LUT_2[17913] = 32'b11111111111111110101011010111001;
assign LUT_2[17914] = 32'b11111111111111111111011011011100;
assign LUT_2[17915] = 32'b11111111111111111100010011110101;
assign LUT_2[17916] = 32'b11111111111111110101000000001000;
assign LUT_2[17917] = 32'b11111111111111110001111000100001;
assign LUT_2[17918] = 32'b11111111111111111011111001000100;
assign LUT_2[17919] = 32'b11111111111111111000110001011101;
assign LUT_2[17920] = 32'b00000000000000000111000111101010;
assign LUT_2[17921] = 32'b00000000000000000100000000000011;
assign LUT_2[17922] = 32'b00000000000000001110000000100110;
assign LUT_2[17923] = 32'b00000000000000001010111000111111;
assign LUT_2[17924] = 32'b00000000000000000011100101010010;
assign LUT_2[17925] = 32'b00000000000000000000011101101011;
assign LUT_2[17926] = 32'b00000000000000001010011110001110;
assign LUT_2[17927] = 32'b00000000000000000111010110100111;
assign LUT_2[17928] = 32'b00000000000000000001111001000111;
assign LUT_2[17929] = 32'b11111111111111111110110001100000;
assign LUT_2[17930] = 32'b00000000000000001000110010000011;
assign LUT_2[17931] = 32'b00000000000000000101101010011100;
assign LUT_2[17932] = 32'b11111111111111111110010110101111;
assign LUT_2[17933] = 32'b11111111111111111011001111001000;
assign LUT_2[17934] = 32'b00000000000000000101001111101011;
assign LUT_2[17935] = 32'b00000000000000000010001000000100;
assign LUT_2[17936] = 32'b00000000000000000001101011110100;
assign LUT_2[17937] = 32'b11111111111111111110100100001101;
assign LUT_2[17938] = 32'b00000000000000001000100100110000;
assign LUT_2[17939] = 32'b00000000000000000101011101001001;
assign LUT_2[17940] = 32'b11111111111111111110001001011100;
assign LUT_2[17941] = 32'b11111111111111111011000001110101;
assign LUT_2[17942] = 32'b00000000000000000101000010011000;
assign LUT_2[17943] = 32'b00000000000000000001111010110001;
assign LUT_2[17944] = 32'b11111111111111111100011101010001;
assign LUT_2[17945] = 32'b11111111111111111001010101101010;
assign LUT_2[17946] = 32'b00000000000000000011010110001101;
assign LUT_2[17947] = 32'b00000000000000000000001110100110;
assign LUT_2[17948] = 32'b11111111111111111000111010111001;
assign LUT_2[17949] = 32'b11111111111111110101110011010010;
assign LUT_2[17950] = 32'b11111111111111111111110011110101;
assign LUT_2[17951] = 32'b11111111111111111100101100001110;
assign LUT_2[17952] = 32'b00000000000000000111100011010011;
assign LUT_2[17953] = 32'b00000000000000000100011011101100;
assign LUT_2[17954] = 32'b00000000000000001110011100001111;
assign LUT_2[17955] = 32'b00000000000000001011010100101000;
assign LUT_2[17956] = 32'b00000000000000000100000000111011;
assign LUT_2[17957] = 32'b00000000000000000000111001010100;
assign LUT_2[17958] = 32'b00000000000000001010111001110111;
assign LUT_2[17959] = 32'b00000000000000000111110010010000;
assign LUT_2[17960] = 32'b00000000000000000010010100110000;
assign LUT_2[17961] = 32'b11111111111111111111001101001001;
assign LUT_2[17962] = 32'b00000000000000001001001101101100;
assign LUT_2[17963] = 32'b00000000000000000110000110000101;
assign LUT_2[17964] = 32'b11111111111111111110110010011000;
assign LUT_2[17965] = 32'b11111111111111111011101010110001;
assign LUT_2[17966] = 32'b00000000000000000101101011010100;
assign LUT_2[17967] = 32'b00000000000000000010100011101101;
assign LUT_2[17968] = 32'b00000000000000000010000111011101;
assign LUT_2[17969] = 32'b11111111111111111110111111110110;
assign LUT_2[17970] = 32'b00000000000000001001000000011001;
assign LUT_2[17971] = 32'b00000000000000000101111000110010;
assign LUT_2[17972] = 32'b11111111111111111110100101000101;
assign LUT_2[17973] = 32'b11111111111111111011011101011110;
assign LUT_2[17974] = 32'b00000000000000000101011110000001;
assign LUT_2[17975] = 32'b00000000000000000010010110011010;
assign LUT_2[17976] = 32'b11111111111111111100111000111010;
assign LUT_2[17977] = 32'b11111111111111111001110001010011;
assign LUT_2[17978] = 32'b00000000000000000011110001110110;
assign LUT_2[17979] = 32'b00000000000000000000101010001111;
assign LUT_2[17980] = 32'b11111111111111111001010110100010;
assign LUT_2[17981] = 32'b11111111111111110110001110111011;
assign LUT_2[17982] = 32'b00000000000000000000001111011110;
assign LUT_2[17983] = 32'b11111111111111111101000111110111;
assign LUT_2[17984] = 32'b11111111111111111111010000001101;
assign LUT_2[17985] = 32'b11111111111111111100001000100110;
assign LUT_2[17986] = 32'b00000000000000000110001001001001;
assign LUT_2[17987] = 32'b00000000000000000011000001100010;
assign LUT_2[17988] = 32'b11111111111111111011101101110101;
assign LUT_2[17989] = 32'b11111111111111111000100110001110;
assign LUT_2[17990] = 32'b00000000000000000010100110110001;
assign LUT_2[17991] = 32'b11111111111111111111011111001010;
assign LUT_2[17992] = 32'b11111111111111111010000001101010;
assign LUT_2[17993] = 32'b11111111111111110110111010000011;
assign LUT_2[17994] = 32'b00000000000000000000111010100110;
assign LUT_2[17995] = 32'b11111111111111111101110010111111;
assign LUT_2[17996] = 32'b11111111111111110110011111010010;
assign LUT_2[17997] = 32'b11111111111111110011010111101011;
assign LUT_2[17998] = 32'b11111111111111111101011000001110;
assign LUT_2[17999] = 32'b11111111111111111010010000100111;
assign LUT_2[18000] = 32'b11111111111111111001110100010111;
assign LUT_2[18001] = 32'b11111111111111110110101100110000;
assign LUT_2[18002] = 32'b00000000000000000000101101010011;
assign LUT_2[18003] = 32'b11111111111111111101100101101100;
assign LUT_2[18004] = 32'b11111111111111110110010001111111;
assign LUT_2[18005] = 32'b11111111111111110011001010011000;
assign LUT_2[18006] = 32'b11111111111111111101001010111011;
assign LUT_2[18007] = 32'b11111111111111111010000011010100;
assign LUT_2[18008] = 32'b11111111111111110100100101110100;
assign LUT_2[18009] = 32'b11111111111111110001011110001101;
assign LUT_2[18010] = 32'b11111111111111111011011110110000;
assign LUT_2[18011] = 32'b11111111111111111000010111001001;
assign LUT_2[18012] = 32'b11111111111111110001000011011100;
assign LUT_2[18013] = 32'b11111111111111101101111011110101;
assign LUT_2[18014] = 32'b11111111111111110111111100011000;
assign LUT_2[18015] = 32'b11111111111111110100110100110001;
assign LUT_2[18016] = 32'b11111111111111111111101011110110;
assign LUT_2[18017] = 32'b11111111111111111100100100001111;
assign LUT_2[18018] = 32'b00000000000000000110100100110010;
assign LUT_2[18019] = 32'b00000000000000000011011101001011;
assign LUT_2[18020] = 32'b11111111111111111100001001011110;
assign LUT_2[18021] = 32'b11111111111111111001000001110111;
assign LUT_2[18022] = 32'b00000000000000000011000010011010;
assign LUT_2[18023] = 32'b11111111111111111111111010110011;
assign LUT_2[18024] = 32'b11111111111111111010011101010011;
assign LUT_2[18025] = 32'b11111111111111110111010101101100;
assign LUT_2[18026] = 32'b00000000000000000001010110001111;
assign LUT_2[18027] = 32'b11111111111111111110001110101000;
assign LUT_2[18028] = 32'b11111111111111110110111010111011;
assign LUT_2[18029] = 32'b11111111111111110011110011010100;
assign LUT_2[18030] = 32'b11111111111111111101110011110111;
assign LUT_2[18031] = 32'b11111111111111111010101100010000;
assign LUT_2[18032] = 32'b11111111111111111010010000000000;
assign LUT_2[18033] = 32'b11111111111111110111001000011001;
assign LUT_2[18034] = 32'b00000000000000000001001000111100;
assign LUT_2[18035] = 32'b11111111111111111110000001010101;
assign LUT_2[18036] = 32'b11111111111111110110101101101000;
assign LUT_2[18037] = 32'b11111111111111110011100110000001;
assign LUT_2[18038] = 32'b11111111111111111101100110100100;
assign LUT_2[18039] = 32'b11111111111111111010011110111101;
assign LUT_2[18040] = 32'b11111111111111110101000001011101;
assign LUT_2[18041] = 32'b11111111111111110001111001110110;
assign LUT_2[18042] = 32'b11111111111111111011111010011001;
assign LUT_2[18043] = 32'b11111111111111111000110010110010;
assign LUT_2[18044] = 32'b11111111111111110001011111000101;
assign LUT_2[18045] = 32'b11111111111111101110010111011110;
assign LUT_2[18046] = 32'b11111111111111111000011000000001;
assign LUT_2[18047] = 32'b11111111111111110101010000011010;
assign LUT_2[18048] = 32'b00000000000000001011011011111001;
assign LUT_2[18049] = 32'b00000000000000001000010100010010;
assign LUT_2[18050] = 32'b00000000000000010010010100110101;
assign LUT_2[18051] = 32'b00000000000000001111001101001110;
assign LUT_2[18052] = 32'b00000000000000000111111001100001;
assign LUT_2[18053] = 32'b00000000000000000100110001111010;
assign LUT_2[18054] = 32'b00000000000000001110110010011101;
assign LUT_2[18055] = 32'b00000000000000001011101010110110;
assign LUT_2[18056] = 32'b00000000000000000110001101010110;
assign LUT_2[18057] = 32'b00000000000000000011000101101111;
assign LUT_2[18058] = 32'b00000000000000001101000110010010;
assign LUT_2[18059] = 32'b00000000000000001001111110101011;
assign LUT_2[18060] = 32'b00000000000000000010101010111110;
assign LUT_2[18061] = 32'b11111111111111111111100011010111;
assign LUT_2[18062] = 32'b00000000000000001001100011111010;
assign LUT_2[18063] = 32'b00000000000000000110011100010011;
assign LUT_2[18064] = 32'b00000000000000000110000000000011;
assign LUT_2[18065] = 32'b00000000000000000010111000011100;
assign LUT_2[18066] = 32'b00000000000000001100111000111111;
assign LUT_2[18067] = 32'b00000000000000001001110001011000;
assign LUT_2[18068] = 32'b00000000000000000010011101101011;
assign LUT_2[18069] = 32'b11111111111111111111010110000100;
assign LUT_2[18070] = 32'b00000000000000001001010110100111;
assign LUT_2[18071] = 32'b00000000000000000110001111000000;
assign LUT_2[18072] = 32'b00000000000000000000110001100000;
assign LUT_2[18073] = 32'b11111111111111111101101001111001;
assign LUT_2[18074] = 32'b00000000000000000111101010011100;
assign LUT_2[18075] = 32'b00000000000000000100100010110101;
assign LUT_2[18076] = 32'b11111111111111111101001111001000;
assign LUT_2[18077] = 32'b11111111111111111010000111100001;
assign LUT_2[18078] = 32'b00000000000000000100001000000100;
assign LUT_2[18079] = 32'b00000000000000000001000000011101;
assign LUT_2[18080] = 32'b00000000000000001011110111100010;
assign LUT_2[18081] = 32'b00000000000000001000101111111011;
assign LUT_2[18082] = 32'b00000000000000010010110000011110;
assign LUT_2[18083] = 32'b00000000000000001111101000110111;
assign LUT_2[18084] = 32'b00000000000000001000010101001010;
assign LUT_2[18085] = 32'b00000000000000000101001101100011;
assign LUT_2[18086] = 32'b00000000000000001111001110000110;
assign LUT_2[18087] = 32'b00000000000000001100000110011111;
assign LUT_2[18088] = 32'b00000000000000000110101000111111;
assign LUT_2[18089] = 32'b00000000000000000011100001011000;
assign LUT_2[18090] = 32'b00000000000000001101100001111011;
assign LUT_2[18091] = 32'b00000000000000001010011010010100;
assign LUT_2[18092] = 32'b00000000000000000011000110100111;
assign LUT_2[18093] = 32'b11111111111111111111111111000000;
assign LUT_2[18094] = 32'b00000000000000001001111111100011;
assign LUT_2[18095] = 32'b00000000000000000110110111111100;
assign LUT_2[18096] = 32'b00000000000000000110011011101100;
assign LUT_2[18097] = 32'b00000000000000000011010100000101;
assign LUT_2[18098] = 32'b00000000000000001101010100101000;
assign LUT_2[18099] = 32'b00000000000000001010001101000001;
assign LUT_2[18100] = 32'b00000000000000000010111001010100;
assign LUT_2[18101] = 32'b11111111111111111111110001101101;
assign LUT_2[18102] = 32'b00000000000000001001110010010000;
assign LUT_2[18103] = 32'b00000000000000000110101010101001;
assign LUT_2[18104] = 32'b00000000000000000001001101001001;
assign LUT_2[18105] = 32'b11111111111111111110000101100010;
assign LUT_2[18106] = 32'b00000000000000001000000110000101;
assign LUT_2[18107] = 32'b00000000000000000100111110011110;
assign LUT_2[18108] = 32'b11111111111111111101101010110001;
assign LUT_2[18109] = 32'b11111111111111111010100011001010;
assign LUT_2[18110] = 32'b00000000000000000100100011101101;
assign LUT_2[18111] = 32'b00000000000000000001011100000110;
assign LUT_2[18112] = 32'b00000000000000000011100100011100;
assign LUT_2[18113] = 32'b00000000000000000000011100110101;
assign LUT_2[18114] = 32'b00000000000000001010011101011000;
assign LUT_2[18115] = 32'b00000000000000000111010101110001;
assign LUT_2[18116] = 32'b00000000000000000000000010000100;
assign LUT_2[18117] = 32'b11111111111111111100111010011101;
assign LUT_2[18118] = 32'b00000000000000000110111011000000;
assign LUT_2[18119] = 32'b00000000000000000011110011011001;
assign LUT_2[18120] = 32'b11111111111111111110010101111001;
assign LUT_2[18121] = 32'b11111111111111111011001110010010;
assign LUT_2[18122] = 32'b00000000000000000101001110110101;
assign LUT_2[18123] = 32'b00000000000000000010000111001110;
assign LUT_2[18124] = 32'b11111111111111111010110011100001;
assign LUT_2[18125] = 32'b11111111111111110111101011111010;
assign LUT_2[18126] = 32'b00000000000000000001101100011101;
assign LUT_2[18127] = 32'b11111111111111111110100100110110;
assign LUT_2[18128] = 32'b11111111111111111110001000100110;
assign LUT_2[18129] = 32'b11111111111111111011000000111111;
assign LUT_2[18130] = 32'b00000000000000000101000001100010;
assign LUT_2[18131] = 32'b00000000000000000001111001111011;
assign LUT_2[18132] = 32'b11111111111111111010100110001110;
assign LUT_2[18133] = 32'b11111111111111110111011110100111;
assign LUT_2[18134] = 32'b00000000000000000001011111001010;
assign LUT_2[18135] = 32'b11111111111111111110010111100011;
assign LUT_2[18136] = 32'b11111111111111111000111010000011;
assign LUT_2[18137] = 32'b11111111111111110101110010011100;
assign LUT_2[18138] = 32'b11111111111111111111110010111111;
assign LUT_2[18139] = 32'b11111111111111111100101011011000;
assign LUT_2[18140] = 32'b11111111111111110101010111101011;
assign LUT_2[18141] = 32'b11111111111111110010010000000100;
assign LUT_2[18142] = 32'b11111111111111111100010000100111;
assign LUT_2[18143] = 32'b11111111111111111001001001000000;
assign LUT_2[18144] = 32'b00000000000000000100000000000101;
assign LUT_2[18145] = 32'b00000000000000000000111000011110;
assign LUT_2[18146] = 32'b00000000000000001010111001000001;
assign LUT_2[18147] = 32'b00000000000000000111110001011010;
assign LUT_2[18148] = 32'b00000000000000000000011101101101;
assign LUT_2[18149] = 32'b11111111111111111101010110000110;
assign LUT_2[18150] = 32'b00000000000000000111010110101001;
assign LUT_2[18151] = 32'b00000000000000000100001111000010;
assign LUT_2[18152] = 32'b11111111111111111110110001100010;
assign LUT_2[18153] = 32'b11111111111111111011101001111011;
assign LUT_2[18154] = 32'b00000000000000000101101010011110;
assign LUT_2[18155] = 32'b00000000000000000010100010110111;
assign LUT_2[18156] = 32'b11111111111111111011001111001010;
assign LUT_2[18157] = 32'b11111111111111111000000111100011;
assign LUT_2[18158] = 32'b00000000000000000010001000000110;
assign LUT_2[18159] = 32'b11111111111111111111000000011111;
assign LUT_2[18160] = 32'b11111111111111111110100100001111;
assign LUT_2[18161] = 32'b11111111111111111011011100101000;
assign LUT_2[18162] = 32'b00000000000000000101011101001011;
assign LUT_2[18163] = 32'b00000000000000000010010101100100;
assign LUT_2[18164] = 32'b11111111111111111011000001110111;
assign LUT_2[18165] = 32'b11111111111111110111111010010000;
assign LUT_2[18166] = 32'b00000000000000000001111010110011;
assign LUT_2[18167] = 32'b11111111111111111110110011001100;
assign LUT_2[18168] = 32'b11111111111111111001010101101100;
assign LUT_2[18169] = 32'b11111111111111110110001110000101;
assign LUT_2[18170] = 32'b00000000000000000000001110101000;
assign LUT_2[18171] = 32'b11111111111111111101000111000001;
assign LUT_2[18172] = 32'b11111111111111110101110011010100;
assign LUT_2[18173] = 32'b11111111111111110010101011101101;
assign LUT_2[18174] = 32'b11111111111111111100101100010000;
assign LUT_2[18175] = 32'b11111111111111111001100100101001;
assign LUT_2[18176] = 32'b00000000000000001011000110010000;
assign LUT_2[18177] = 32'b00000000000000000111111110101001;
assign LUT_2[18178] = 32'b00000000000000010001111111001100;
assign LUT_2[18179] = 32'b00000000000000001110110111100101;
assign LUT_2[18180] = 32'b00000000000000000111100011111000;
assign LUT_2[18181] = 32'b00000000000000000100011100010001;
assign LUT_2[18182] = 32'b00000000000000001110011100110100;
assign LUT_2[18183] = 32'b00000000000000001011010101001101;
assign LUT_2[18184] = 32'b00000000000000000101110111101101;
assign LUT_2[18185] = 32'b00000000000000000010110000000110;
assign LUT_2[18186] = 32'b00000000000000001100110000101001;
assign LUT_2[18187] = 32'b00000000000000001001101001000010;
assign LUT_2[18188] = 32'b00000000000000000010010101010101;
assign LUT_2[18189] = 32'b11111111111111111111001101101110;
assign LUT_2[18190] = 32'b00000000000000001001001110010001;
assign LUT_2[18191] = 32'b00000000000000000110000110101010;
assign LUT_2[18192] = 32'b00000000000000000101101010011010;
assign LUT_2[18193] = 32'b00000000000000000010100010110011;
assign LUT_2[18194] = 32'b00000000000000001100100011010110;
assign LUT_2[18195] = 32'b00000000000000001001011011101111;
assign LUT_2[18196] = 32'b00000000000000000010001000000010;
assign LUT_2[18197] = 32'b11111111111111111111000000011011;
assign LUT_2[18198] = 32'b00000000000000001001000000111110;
assign LUT_2[18199] = 32'b00000000000000000101111001010111;
assign LUT_2[18200] = 32'b00000000000000000000011011110111;
assign LUT_2[18201] = 32'b11111111111111111101010100010000;
assign LUT_2[18202] = 32'b00000000000000000111010100110011;
assign LUT_2[18203] = 32'b00000000000000000100001101001100;
assign LUT_2[18204] = 32'b11111111111111111100111001011111;
assign LUT_2[18205] = 32'b11111111111111111001110001111000;
assign LUT_2[18206] = 32'b00000000000000000011110010011011;
assign LUT_2[18207] = 32'b00000000000000000000101010110100;
assign LUT_2[18208] = 32'b00000000000000001011100001111001;
assign LUT_2[18209] = 32'b00000000000000001000011010010010;
assign LUT_2[18210] = 32'b00000000000000010010011010110101;
assign LUT_2[18211] = 32'b00000000000000001111010011001110;
assign LUT_2[18212] = 32'b00000000000000000111111111100001;
assign LUT_2[18213] = 32'b00000000000000000100110111111010;
assign LUT_2[18214] = 32'b00000000000000001110111000011101;
assign LUT_2[18215] = 32'b00000000000000001011110000110110;
assign LUT_2[18216] = 32'b00000000000000000110010011010110;
assign LUT_2[18217] = 32'b00000000000000000011001011101111;
assign LUT_2[18218] = 32'b00000000000000001101001100010010;
assign LUT_2[18219] = 32'b00000000000000001010000100101011;
assign LUT_2[18220] = 32'b00000000000000000010110000111110;
assign LUT_2[18221] = 32'b11111111111111111111101001010111;
assign LUT_2[18222] = 32'b00000000000000001001101001111010;
assign LUT_2[18223] = 32'b00000000000000000110100010010011;
assign LUT_2[18224] = 32'b00000000000000000110000110000011;
assign LUT_2[18225] = 32'b00000000000000000010111110011100;
assign LUT_2[18226] = 32'b00000000000000001100111110111111;
assign LUT_2[18227] = 32'b00000000000000001001110111011000;
assign LUT_2[18228] = 32'b00000000000000000010100011101011;
assign LUT_2[18229] = 32'b11111111111111111111011100000100;
assign LUT_2[18230] = 32'b00000000000000001001011100100111;
assign LUT_2[18231] = 32'b00000000000000000110010101000000;
assign LUT_2[18232] = 32'b00000000000000000000110111100000;
assign LUT_2[18233] = 32'b11111111111111111101101111111001;
assign LUT_2[18234] = 32'b00000000000000000111110000011100;
assign LUT_2[18235] = 32'b00000000000000000100101000110101;
assign LUT_2[18236] = 32'b11111111111111111101010101001000;
assign LUT_2[18237] = 32'b11111111111111111010001101100001;
assign LUT_2[18238] = 32'b00000000000000000100001110000100;
assign LUT_2[18239] = 32'b00000000000000000001000110011101;
assign LUT_2[18240] = 32'b00000000000000000011001110110011;
assign LUT_2[18241] = 32'b00000000000000000000000111001100;
assign LUT_2[18242] = 32'b00000000000000001010000111101111;
assign LUT_2[18243] = 32'b00000000000000000111000000001000;
assign LUT_2[18244] = 32'b11111111111111111111101100011011;
assign LUT_2[18245] = 32'b11111111111111111100100100110100;
assign LUT_2[18246] = 32'b00000000000000000110100101010111;
assign LUT_2[18247] = 32'b00000000000000000011011101110000;
assign LUT_2[18248] = 32'b11111111111111111110000000010000;
assign LUT_2[18249] = 32'b11111111111111111010111000101001;
assign LUT_2[18250] = 32'b00000000000000000100111001001100;
assign LUT_2[18251] = 32'b00000000000000000001110001100101;
assign LUT_2[18252] = 32'b11111111111111111010011101111000;
assign LUT_2[18253] = 32'b11111111111111110111010110010001;
assign LUT_2[18254] = 32'b00000000000000000001010110110100;
assign LUT_2[18255] = 32'b11111111111111111110001111001101;
assign LUT_2[18256] = 32'b11111111111111111101110010111101;
assign LUT_2[18257] = 32'b11111111111111111010101011010110;
assign LUT_2[18258] = 32'b00000000000000000100101011111001;
assign LUT_2[18259] = 32'b00000000000000000001100100010010;
assign LUT_2[18260] = 32'b11111111111111111010010000100101;
assign LUT_2[18261] = 32'b11111111111111110111001000111110;
assign LUT_2[18262] = 32'b00000000000000000001001001100001;
assign LUT_2[18263] = 32'b11111111111111111110000001111010;
assign LUT_2[18264] = 32'b11111111111111111000100100011010;
assign LUT_2[18265] = 32'b11111111111111110101011100110011;
assign LUT_2[18266] = 32'b11111111111111111111011101010110;
assign LUT_2[18267] = 32'b11111111111111111100010101101111;
assign LUT_2[18268] = 32'b11111111111111110101000010000010;
assign LUT_2[18269] = 32'b11111111111111110001111010011011;
assign LUT_2[18270] = 32'b11111111111111111011111010111110;
assign LUT_2[18271] = 32'b11111111111111111000110011010111;
assign LUT_2[18272] = 32'b00000000000000000011101010011100;
assign LUT_2[18273] = 32'b00000000000000000000100010110101;
assign LUT_2[18274] = 32'b00000000000000001010100011011000;
assign LUT_2[18275] = 32'b00000000000000000111011011110001;
assign LUT_2[18276] = 32'b00000000000000000000001000000100;
assign LUT_2[18277] = 32'b11111111111111111101000000011101;
assign LUT_2[18278] = 32'b00000000000000000111000001000000;
assign LUT_2[18279] = 32'b00000000000000000011111001011001;
assign LUT_2[18280] = 32'b11111111111111111110011011111001;
assign LUT_2[18281] = 32'b11111111111111111011010100010010;
assign LUT_2[18282] = 32'b00000000000000000101010100110101;
assign LUT_2[18283] = 32'b00000000000000000010001101001110;
assign LUT_2[18284] = 32'b11111111111111111010111001100001;
assign LUT_2[18285] = 32'b11111111111111110111110001111010;
assign LUT_2[18286] = 32'b00000000000000000001110010011101;
assign LUT_2[18287] = 32'b11111111111111111110101010110110;
assign LUT_2[18288] = 32'b11111111111111111110001110100110;
assign LUT_2[18289] = 32'b11111111111111111011000110111111;
assign LUT_2[18290] = 32'b00000000000000000101000111100010;
assign LUT_2[18291] = 32'b00000000000000000001111111111011;
assign LUT_2[18292] = 32'b11111111111111111010101100001110;
assign LUT_2[18293] = 32'b11111111111111110111100100100111;
assign LUT_2[18294] = 32'b00000000000000000001100101001010;
assign LUT_2[18295] = 32'b11111111111111111110011101100011;
assign LUT_2[18296] = 32'b11111111111111111001000000000011;
assign LUT_2[18297] = 32'b11111111111111110101111000011100;
assign LUT_2[18298] = 32'b11111111111111111111111000111111;
assign LUT_2[18299] = 32'b11111111111111111100110001011000;
assign LUT_2[18300] = 32'b11111111111111110101011101101011;
assign LUT_2[18301] = 32'b11111111111111110010010110000100;
assign LUT_2[18302] = 32'b11111111111111111100010110100111;
assign LUT_2[18303] = 32'b11111111111111111001001111000000;
assign LUT_2[18304] = 32'b00000000000000001111011010011111;
assign LUT_2[18305] = 32'b00000000000000001100010010111000;
assign LUT_2[18306] = 32'b00000000000000010110010011011011;
assign LUT_2[18307] = 32'b00000000000000010011001011110100;
assign LUT_2[18308] = 32'b00000000000000001011111000000111;
assign LUT_2[18309] = 32'b00000000000000001000110000100000;
assign LUT_2[18310] = 32'b00000000000000010010110001000011;
assign LUT_2[18311] = 32'b00000000000000001111101001011100;
assign LUT_2[18312] = 32'b00000000000000001010001011111100;
assign LUT_2[18313] = 32'b00000000000000000111000100010101;
assign LUT_2[18314] = 32'b00000000000000010001000100111000;
assign LUT_2[18315] = 32'b00000000000000001101111101010001;
assign LUT_2[18316] = 32'b00000000000000000110101001100100;
assign LUT_2[18317] = 32'b00000000000000000011100001111101;
assign LUT_2[18318] = 32'b00000000000000001101100010100000;
assign LUT_2[18319] = 32'b00000000000000001010011010111001;
assign LUT_2[18320] = 32'b00000000000000001001111110101001;
assign LUT_2[18321] = 32'b00000000000000000110110111000010;
assign LUT_2[18322] = 32'b00000000000000010000110111100101;
assign LUT_2[18323] = 32'b00000000000000001101101111111110;
assign LUT_2[18324] = 32'b00000000000000000110011100010001;
assign LUT_2[18325] = 32'b00000000000000000011010100101010;
assign LUT_2[18326] = 32'b00000000000000001101010101001101;
assign LUT_2[18327] = 32'b00000000000000001010001101100110;
assign LUT_2[18328] = 32'b00000000000000000100110000000110;
assign LUT_2[18329] = 32'b00000000000000000001101000011111;
assign LUT_2[18330] = 32'b00000000000000001011101001000010;
assign LUT_2[18331] = 32'b00000000000000001000100001011011;
assign LUT_2[18332] = 32'b00000000000000000001001101101110;
assign LUT_2[18333] = 32'b11111111111111111110000110000111;
assign LUT_2[18334] = 32'b00000000000000001000000110101010;
assign LUT_2[18335] = 32'b00000000000000000100111111000011;
assign LUT_2[18336] = 32'b00000000000000001111110110001000;
assign LUT_2[18337] = 32'b00000000000000001100101110100001;
assign LUT_2[18338] = 32'b00000000000000010110101111000100;
assign LUT_2[18339] = 32'b00000000000000010011100111011101;
assign LUT_2[18340] = 32'b00000000000000001100010011110000;
assign LUT_2[18341] = 32'b00000000000000001001001100001001;
assign LUT_2[18342] = 32'b00000000000000010011001100101100;
assign LUT_2[18343] = 32'b00000000000000010000000101000101;
assign LUT_2[18344] = 32'b00000000000000001010100111100101;
assign LUT_2[18345] = 32'b00000000000000000111011111111110;
assign LUT_2[18346] = 32'b00000000000000010001100000100001;
assign LUT_2[18347] = 32'b00000000000000001110011000111010;
assign LUT_2[18348] = 32'b00000000000000000111000101001101;
assign LUT_2[18349] = 32'b00000000000000000011111101100110;
assign LUT_2[18350] = 32'b00000000000000001101111110001001;
assign LUT_2[18351] = 32'b00000000000000001010110110100010;
assign LUT_2[18352] = 32'b00000000000000001010011010010010;
assign LUT_2[18353] = 32'b00000000000000000111010010101011;
assign LUT_2[18354] = 32'b00000000000000010001010011001110;
assign LUT_2[18355] = 32'b00000000000000001110001011100111;
assign LUT_2[18356] = 32'b00000000000000000110110111111010;
assign LUT_2[18357] = 32'b00000000000000000011110000010011;
assign LUT_2[18358] = 32'b00000000000000001101110000110110;
assign LUT_2[18359] = 32'b00000000000000001010101001001111;
assign LUT_2[18360] = 32'b00000000000000000101001011101111;
assign LUT_2[18361] = 32'b00000000000000000010000100001000;
assign LUT_2[18362] = 32'b00000000000000001100000100101011;
assign LUT_2[18363] = 32'b00000000000000001000111101000100;
assign LUT_2[18364] = 32'b00000000000000000001101001010111;
assign LUT_2[18365] = 32'b11111111111111111110100001110000;
assign LUT_2[18366] = 32'b00000000000000001000100010010011;
assign LUT_2[18367] = 32'b00000000000000000101011010101100;
assign LUT_2[18368] = 32'b00000000000000000111100011000010;
assign LUT_2[18369] = 32'b00000000000000000100011011011011;
assign LUT_2[18370] = 32'b00000000000000001110011011111110;
assign LUT_2[18371] = 32'b00000000000000001011010100010111;
assign LUT_2[18372] = 32'b00000000000000000100000000101010;
assign LUT_2[18373] = 32'b00000000000000000000111001000011;
assign LUT_2[18374] = 32'b00000000000000001010111001100110;
assign LUT_2[18375] = 32'b00000000000000000111110001111111;
assign LUT_2[18376] = 32'b00000000000000000010010100011111;
assign LUT_2[18377] = 32'b11111111111111111111001100111000;
assign LUT_2[18378] = 32'b00000000000000001001001101011011;
assign LUT_2[18379] = 32'b00000000000000000110000101110100;
assign LUT_2[18380] = 32'b11111111111111111110110010000111;
assign LUT_2[18381] = 32'b11111111111111111011101010100000;
assign LUT_2[18382] = 32'b00000000000000000101101011000011;
assign LUT_2[18383] = 32'b00000000000000000010100011011100;
assign LUT_2[18384] = 32'b00000000000000000010000111001100;
assign LUT_2[18385] = 32'b11111111111111111110111111100101;
assign LUT_2[18386] = 32'b00000000000000001001000000001000;
assign LUT_2[18387] = 32'b00000000000000000101111000100001;
assign LUT_2[18388] = 32'b11111111111111111110100100110100;
assign LUT_2[18389] = 32'b11111111111111111011011101001101;
assign LUT_2[18390] = 32'b00000000000000000101011101110000;
assign LUT_2[18391] = 32'b00000000000000000010010110001001;
assign LUT_2[18392] = 32'b11111111111111111100111000101001;
assign LUT_2[18393] = 32'b11111111111111111001110001000010;
assign LUT_2[18394] = 32'b00000000000000000011110001100101;
assign LUT_2[18395] = 32'b00000000000000000000101001111110;
assign LUT_2[18396] = 32'b11111111111111111001010110010001;
assign LUT_2[18397] = 32'b11111111111111110110001110101010;
assign LUT_2[18398] = 32'b00000000000000000000001111001101;
assign LUT_2[18399] = 32'b11111111111111111101000111100110;
assign LUT_2[18400] = 32'b00000000000000000111111110101011;
assign LUT_2[18401] = 32'b00000000000000000100110111000100;
assign LUT_2[18402] = 32'b00000000000000001110110111100111;
assign LUT_2[18403] = 32'b00000000000000001011110000000000;
assign LUT_2[18404] = 32'b00000000000000000100011100010011;
assign LUT_2[18405] = 32'b00000000000000000001010100101100;
assign LUT_2[18406] = 32'b00000000000000001011010101001111;
assign LUT_2[18407] = 32'b00000000000000001000001101101000;
assign LUT_2[18408] = 32'b00000000000000000010110000001000;
assign LUT_2[18409] = 32'b11111111111111111111101000100001;
assign LUT_2[18410] = 32'b00000000000000001001101001000100;
assign LUT_2[18411] = 32'b00000000000000000110100001011101;
assign LUT_2[18412] = 32'b11111111111111111111001101110000;
assign LUT_2[18413] = 32'b11111111111111111100000110001001;
assign LUT_2[18414] = 32'b00000000000000000110000110101100;
assign LUT_2[18415] = 32'b00000000000000000010111111000101;
assign LUT_2[18416] = 32'b00000000000000000010100010110101;
assign LUT_2[18417] = 32'b11111111111111111111011011001110;
assign LUT_2[18418] = 32'b00000000000000001001011011110001;
assign LUT_2[18419] = 32'b00000000000000000110010100001010;
assign LUT_2[18420] = 32'b11111111111111111111000000011101;
assign LUT_2[18421] = 32'b11111111111111111011111000110110;
assign LUT_2[18422] = 32'b00000000000000000101111001011001;
assign LUT_2[18423] = 32'b00000000000000000010110001110010;
assign LUT_2[18424] = 32'b11111111111111111101010100010010;
assign LUT_2[18425] = 32'b11111111111111111010001100101011;
assign LUT_2[18426] = 32'b00000000000000000100001101001110;
assign LUT_2[18427] = 32'b00000000000000000001000101100111;
assign LUT_2[18428] = 32'b11111111111111111001110001111010;
assign LUT_2[18429] = 32'b11111111111111110110101010010011;
assign LUT_2[18430] = 32'b00000000000000000000101010110110;
assign LUT_2[18431] = 32'b11111111111111111101100011001111;
assign LUT_2[18432] = 32'b11111111111111110111011111101111;
assign LUT_2[18433] = 32'b11111111111111110100011000001000;
assign LUT_2[18434] = 32'b11111111111111111110011000101011;
assign LUT_2[18435] = 32'b11111111111111111011010001000100;
assign LUT_2[18436] = 32'b11111111111111110011111101010111;
assign LUT_2[18437] = 32'b11111111111111110000110101110000;
assign LUT_2[18438] = 32'b11111111111111111010110110010011;
assign LUT_2[18439] = 32'b11111111111111110111101110101100;
assign LUT_2[18440] = 32'b11111111111111110010010001001100;
assign LUT_2[18441] = 32'b11111111111111101111001001100101;
assign LUT_2[18442] = 32'b11111111111111111001001010001000;
assign LUT_2[18443] = 32'b11111111111111110110000010100001;
assign LUT_2[18444] = 32'b11111111111111101110101110110100;
assign LUT_2[18445] = 32'b11111111111111101011100111001101;
assign LUT_2[18446] = 32'b11111111111111110101100111110000;
assign LUT_2[18447] = 32'b11111111111111110010100000001001;
assign LUT_2[18448] = 32'b11111111111111110010000011111001;
assign LUT_2[18449] = 32'b11111111111111101110111100010010;
assign LUT_2[18450] = 32'b11111111111111111000111100110101;
assign LUT_2[18451] = 32'b11111111111111110101110101001110;
assign LUT_2[18452] = 32'b11111111111111101110100001100001;
assign LUT_2[18453] = 32'b11111111111111101011011001111010;
assign LUT_2[18454] = 32'b11111111111111110101011010011101;
assign LUT_2[18455] = 32'b11111111111111110010010010110110;
assign LUT_2[18456] = 32'b11111111111111101100110101010110;
assign LUT_2[18457] = 32'b11111111111111101001101101101111;
assign LUT_2[18458] = 32'b11111111111111110011101110010010;
assign LUT_2[18459] = 32'b11111111111111110000100110101011;
assign LUT_2[18460] = 32'b11111111111111101001010010111110;
assign LUT_2[18461] = 32'b11111111111111100110001011010111;
assign LUT_2[18462] = 32'b11111111111111110000001011111010;
assign LUT_2[18463] = 32'b11111111111111101101000100010011;
assign LUT_2[18464] = 32'b11111111111111110111111011011000;
assign LUT_2[18465] = 32'b11111111111111110100110011110001;
assign LUT_2[18466] = 32'b11111111111111111110110100010100;
assign LUT_2[18467] = 32'b11111111111111111011101100101101;
assign LUT_2[18468] = 32'b11111111111111110100011001000000;
assign LUT_2[18469] = 32'b11111111111111110001010001011001;
assign LUT_2[18470] = 32'b11111111111111111011010001111100;
assign LUT_2[18471] = 32'b11111111111111111000001010010101;
assign LUT_2[18472] = 32'b11111111111111110010101100110101;
assign LUT_2[18473] = 32'b11111111111111101111100101001110;
assign LUT_2[18474] = 32'b11111111111111111001100101110001;
assign LUT_2[18475] = 32'b11111111111111110110011110001010;
assign LUT_2[18476] = 32'b11111111111111101111001010011101;
assign LUT_2[18477] = 32'b11111111111111101100000010110110;
assign LUT_2[18478] = 32'b11111111111111110110000011011001;
assign LUT_2[18479] = 32'b11111111111111110010111011110010;
assign LUT_2[18480] = 32'b11111111111111110010011111100010;
assign LUT_2[18481] = 32'b11111111111111101111010111111011;
assign LUT_2[18482] = 32'b11111111111111111001011000011110;
assign LUT_2[18483] = 32'b11111111111111110110010000110111;
assign LUT_2[18484] = 32'b11111111111111101110111101001010;
assign LUT_2[18485] = 32'b11111111111111101011110101100011;
assign LUT_2[18486] = 32'b11111111111111110101110110000110;
assign LUT_2[18487] = 32'b11111111111111110010101110011111;
assign LUT_2[18488] = 32'b11111111111111101101010000111111;
assign LUT_2[18489] = 32'b11111111111111101010001001011000;
assign LUT_2[18490] = 32'b11111111111111110100001001111011;
assign LUT_2[18491] = 32'b11111111111111110001000010010100;
assign LUT_2[18492] = 32'b11111111111111101001101110100111;
assign LUT_2[18493] = 32'b11111111111111100110100111000000;
assign LUT_2[18494] = 32'b11111111111111110000100111100011;
assign LUT_2[18495] = 32'b11111111111111101101011111111100;
assign LUT_2[18496] = 32'b11111111111111101111101000010010;
assign LUT_2[18497] = 32'b11111111111111101100100000101011;
assign LUT_2[18498] = 32'b11111111111111110110100001001110;
assign LUT_2[18499] = 32'b11111111111111110011011001100111;
assign LUT_2[18500] = 32'b11111111111111101100000101111010;
assign LUT_2[18501] = 32'b11111111111111101000111110010011;
assign LUT_2[18502] = 32'b11111111111111110010111110110110;
assign LUT_2[18503] = 32'b11111111111111101111110111001111;
assign LUT_2[18504] = 32'b11111111111111101010011001101111;
assign LUT_2[18505] = 32'b11111111111111100111010010001000;
assign LUT_2[18506] = 32'b11111111111111110001010010101011;
assign LUT_2[18507] = 32'b11111111111111101110001011000100;
assign LUT_2[18508] = 32'b11111111111111100110110111010111;
assign LUT_2[18509] = 32'b11111111111111100011101111110000;
assign LUT_2[18510] = 32'b11111111111111101101110000010011;
assign LUT_2[18511] = 32'b11111111111111101010101000101100;
assign LUT_2[18512] = 32'b11111111111111101010001100011100;
assign LUT_2[18513] = 32'b11111111111111100111000100110101;
assign LUT_2[18514] = 32'b11111111111111110001000101011000;
assign LUT_2[18515] = 32'b11111111111111101101111101110001;
assign LUT_2[18516] = 32'b11111111111111100110101010000100;
assign LUT_2[18517] = 32'b11111111111111100011100010011101;
assign LUT_2[18518] = 32'b11111111111111101101100011000000;
assign LUT_2[18519] = 32'b11111111111111101010011011011001;
assign LUT_2[18520] = 32'b11111111111111100100111101111001;
assign LUT_2[18521] = 32'b11111111111111100001110110010010;
assign LUT_2[18522] = 32'b11111111111111101011110110110101;
assign LUT_2[18523] = 32'b11111111111111101000101111001110;
assign LUT_2[18524] = 32'b11111111111111100001011011100001;
assign LUT_2[18525] = 32'b11111111111111011110010011111010;
assign LUT_2[18526] = 32'b11111111111111101000010100011101;
assign LUT_2[18527] = 32'b11111111111111100101001100110110;
assign LUT_2[18528] = 32'b11111111111111110000000011111011;
assign LUT_2[18529] = 32'b11111111111111101100111100010100;
assign LUT_2[18530] = 32'b11111111111111110110111100110111;
assign LUT_2[18531] = 32'b11111111111111110011110101010000;
assign LUT_2[18532] = 32'b11111111111111101100100001100011;
assign LUT_2[18533] = 32'b11111111111111101001011001111100;
assign LUT_2[18534] = 32'b11111111111111110011011010011111;
assign LUT_2[18535] = 32'b11111111111111110000010010111000;
assign LUT_2[18536] = 32'b11111111111111101010110101011000;
assign LUT_2[18537] = 32'b11111111111111100111101101110001;
assign LUT_2[18538] = 32'b11111111111111110001101110010100;
assign LUT_2[18539] = 32'b11111111111111101110100110101101;
assign LUT_2[18540] = 32'b11111111111111100111010011000000;
assign LUT_2[18541] = 32'b11111111111111100100001011011001;
assign LUT_2[18542] = 32'b11111111111111101110001011111100;
assign LUT_2[18543] = 32'b11111111111111101011000100010101;
assign LUT_2[18544] = 32'b11111111111111101010101000000101;
assign LUT_2[18545] = 32'b11111111111111100111100000011110;
assign LUT_2[18546] = 32'b11111111111111110001100001000001;
assign LUT_2[18547] = 32'b11111111111111101110011001011010;
assign LUT_2[18548] = 32'b11111111111111100111000101101101;
assign LUT_2[18549] = 32'b11111111111111100011111110000110;
assign LUT_2[18550] = 32'b11111111111111101101111110101001;
assign LUT_2[18551] = 32'b11111111111111101010110111000010;
assign LUT_2[18552] = 32'b11111111111111100101011001100010;
assign LUT_2[18553] = 32'b11111111111111100010010001111011;
assign LUT_2[18554] = 32'b11111111111111101100010010011110;
assign LUT_2[18555] = 32'b11111111111111101001001010110111;
assign LUT_2[18556] = 32'b11111111111111100001110111001010;
assign LUT_2[18557] = 32'b11111111111111011110101111100011;
assign LUT_2[18558] = 32'b11111111111111101000110000000110;
assign LUT_2[18559] = 32'b11111111111111100101101000011111;
assign LUT_2[18560] = 32'b11111111111111111011110011111110;
assign LUT_2[18561] = 32'b11111111111111111000101100010111;
assign LUT_2[18562] = 32'b00000000000000000010101100111010;
assign LUT_2[18563] = 32'b11111111111111111111100101010011;
assign LUT_2[18564] = 32'b11111111111111111000010001100110;
assign LUT_2[18565] = 32'b11111111111111110101001001111111;
assign LUT_2[18566] = 32'b11111111111111111111001010100010;
assign LUT_2[18567] = 32'b11111111111111111100000010111011;
assign LUT_2[18568] = 32'b11111111111111110110100101011011;
assign LUT_2[18569] = 32'b11111111111111110011011101110100;
assign LUT_2[18570] = 32'b11111111111111111101011110010111;
assign LUT_2[18571] = 32'b11111111111111111010010110110000;
assign LUT_2[18572] = 32'b11111111111111110011000011000011;
assign LUT_2[18573] = 32'b11111111111111101111111011011100;
assign LUT_2[18574] = 32'b11111111111111111001111011111111;
assign LUT_2[18575] = 32'b11111111111111110110110100011000;
assign LUT_2[18576] = 32'b11111111111111110110011000001000;
assign LUT_2[18577] = 32'b11111111111111110011010000100001;
assign LUT_2[18578] = 32'b11111111111111111101010001000100;
assign LUT_2[18579] = 32'b11111111111111111010001001011101;
assign LUT_2[18580] = 32'b11111111111111110010110101110000;
assign LUT_2[18581] = 32'b11111111111111101111101110001001;
assign LUT_2[18582] = 32'b11111111111111111001101110101100;
assign LUT_2[18583] = 32'b11111111111111110110100111000101;
assign LUT_2[18584] = 32'b11111111111111110001001001100101;
assign LUT_2[18585] = 32'b11111111111111101110000001111110;
assign LUT_2[18586] = 32'b11111111111111111000000010100001;
assign LUT_2[18587] = 32'b11111111111111110100111010111010;
assign LUT_2[18588] = 32'b11111111111111101101100111001101;
assign LUT_2[18589] = 32'b11111111111111101010011111100110;
assign LUT_2[18590] = 32'b11111111111111110100100000001001;
assign LUT_2[18591] = 32'b11111111111111110001011000100010;
assign LUT_2[18592] = 32'b11111111111111111100001111100111;
assign LUT_2[18593] = 32'b11111111111111111001001000000000;
assign LUT_2[18594] = 32'b00000000000000000011001000100011;
assign LUT_2[18595] = 32'b00000000000000000000000000111100;
assign LUT_2[18596] = 32'b11111111111111111000101101001111;
assign LUT_2[18597] = 32'b11111111111111110101100101101000;
assign LUT_2[18598] = 32'b11111111111111111111100110001011;
assign LUT_2[18599] = 32'b11111111111111111100011110100100;
assign LUT_2[18600] = 32'b11111111111111110111000001000100;
assign LUT_2[18601] = 32'b11111111111111110011111001011101;
assign LUT_2[18602] = 32'b11111111111111111101111010000000;
assign LUT_2[18603] = 32'b11111111111111111010110010011001;
assign LUT_2[18604] = 32'b11111111111111110011011110101100;
assign LUT_2[18605] = 32'b11111111111111110000010111000101;
assign LUT_2[18606] = 32'b11111111111111111010010111101000;
assign LUT_2[18607] = 32'b11111111111111110111010000000001;
assign LUT_2[18608] = 32'b11111111111111110110110011110001;
assign LUT_2[18609] = 32'b11111111111111110011101100001010;
assign LUT_2[18610] = 32'b11111111111111111101101100101101;
assign LUT_2[18611] = 32'b11111111111111111010100101000110;
assign LUT_2[18612] = 32'b11111111111111110011010001011001;
assign LUT_2[18613] = 32'b11111111111111110000001001110010;
assign LUT_2[18614] = 32'b11111111111111111010001010010101;
assign LUT_2[18615] = 32'b11111111111111110111000010101110;
assign LUT_2[18616] = 32'b11111111111111110001100101001110;
assign LUT_2[18617] = 32'b11111111111111101110011101100111;
assign LUT_2[18618] = 32'b11111111111111111000011110001010;
assign LUT_2[18619] = 32'b11111111111111110101010110100011;
assign LUT_2[18620] = 32'b11111111111111101110000010110110;
assign LUT_2[18621] = 32'b11111111111111101010111011001111;
assign LUT_2[18622] = 32'b11111111111111110100111011110010;
assign LUT_2[18623] = 32'b11111111111111110001110100001011;
assign LUT_2[18624] = 32'b11111111111111110011111100100001;
assign LUT_2[18625] = 32'b11111111111111110000110100111010;
assign LUT_2[18626] = 32'b11111111111111111010110101011101;
assign LUT_2[18627] = 32'b11111111111111110111101101110110;
assign LUT_2[18628] = 32'b11111111111111110000011010001001;
assign LUT_2[18629] = 32'b11111111111111101101010010100010;
assign LUT_2[18630] = 32'b11111111111111110111010011000101;
assign LUT_2[18631] = 32'b11111111111111110100001011011110;
assign LUT_2[18632] = 32'b11111111111111101110101101111110;
assign LUT_2[18633] = 32'b11111111111111101011100110010111;
assign LUT_2[18634] = 32'b11111111111111110101100110111010;
assign LUT_2[18635] = 32'b11111111111111110010011111010011;
assign LUT_2[18636] = 32'b11111111111111101011001011100110;
assign LUT_2[18637] = 32'b11111111111111101000000011111111;
assign LUT_2[18638] = 32'b11111111111111110010000100100010;
assign LUT_2[18639] = 32'b11111111111111101110111100111011;
assign LUT_2[18640] = 32'b11111111111111101110100000101011;
assign LUT_2[18641] = 32'b11111111111111101011011001000100;
assign LUT_2[18642] = 32'b11111111111111110101011001100111;
assign LUT_2[18643] = 32'b11111111111111110010010010000000;
assign LUT_2[18644] = 32'b11111111111111101010111110010011;
assign LUT_2[18645] = 32'b11111111111111100111110110101100;
assign LUT_2[18646] = 32'b11111111111111110001110111001111;
assign LUT_2[18647] = 32'b11111111111111101110101111101000;
assign LUT_2[18648] = 32'b11111111111111101001010010001000;
assign LUT_2[18649] = 32'b11111111111111100110001010100001;
assign LUT_2[18650] = 32'b11111111111111110000001011000100;
assign LUT_2[18651] = 32'b11111111111111101101000011011101;
assign LUT_2[18652] = 32'b11111111111111100101101111110000;
assign LUT_2[18653] = 32'b11111111111111100010101000001001;
assign LUT_2[18654] = 32'b11111111111111101100101000101100;
assign LUT_2[18655] = 32'b11111111111111101001100001000101;
assign LUT_2[18656] = 32'b11111111111111110100011000001010;
assign LUT_2[18657] = 32'b11111111111111110001010000100011;
assign LUT_2[18658] = 32'b11111111111111111011010001000110;
assign LUT_2[18659] = 32'b11111111111111111000001001011111;
assign LUT_2[18660] = 32'b11111111111111110000110101110010;
assign LUT_2[18661] = 32'b11111111111111101101101110001011;
assign LUT_2[18662] = 32'b11111111111111110111101110101110;
assign LUT_2[18663] = 32'b11111111111111110100100111000111;
assign LUT_2[18664] = 32'b11111111111111101111001001100111;
assign LUT_2[18665] = 32'b11111111111111101100000010000000;
assign LUT_2[18666] = 32'b11111111111111110110000010100011;
assign LUT_2[18667] = 32'b11111111111111110010111010111100;
assign LUT_2[18668] = 32'b11111111111111101011100111001111;
assign LUT_2[18669] = 32'b11111111111111101000011111101000;
assign LUT_2[18670] = 32'b11111111111111110010100000001011;
assign LUT_2[18671] = 32'b11111111111111101111011000100100;
assign LUT_2[18672] = 32'b11111111111111101110111100010100;
assign LUT_2[18673] = 32'b11111111111111101011110100101101;
assign LUT_2[18674] = 32'b11111111111111110101110101010000;
assign LUT_2[18675] = 32'b11111111111111110010101101101001;
assign LUT_2[18676] = 32'b11111111111111101011011001111100;
assign LUT_2[18677] = 32'b11111111111111101000010010010101;
assign LUT_2[18678] = 32'b11111111111111110010010010111000;
assign LUT_2[18679] = 32'b11111111111111101111001011010001;
assign LUT_2[18680] = 32'b11111111111111101001101101110001;
assign LUT_2[18681] = 32'b11111111111111100110100110001010;
assign LUT_2[18682] = 32'b11111111111111110000100110101101;
assign LUT_2[18683] = 32'b11111111111111101101011111000110;
assign LUT_2[18684] = 32'b11111111111111100110001011011001;
assign LUT_2[18685] = 32'b11111111111111100011000011110010;
assign LUT_2[18686] = 32'b11111111111111101101000100010101;
assign LUT_2[18687] = 32'b11111111111111101001111100101110;
assign LUT_2[18688] = 32'b11111111111111111011011110010101;
assign LUT_2[18689] = 32'b11111111111111111000010110101110;
assign LUT_2[18690] = 32'b00000000000000000010010111010001;
assign LUT_2[18691] = 32'b11111111111111111111001111101010;
assign LUT_2[18692] = 32'b11111111111111110111111011111101;
assign LUT_2[18693] = 32'b11111111111111110100110100010110;
assign LUT_2[18694] = 32'b11111111111111111110110100111001;
assign LUT_2[18695] = 32'b11111111111111111011101101010010;
assign LUT_2[18696] = 32'b11111111111111110110001111110010;
assign LUT_2[18697] = 32'b11111111111111110011001000001011;
assign LUT_2[18698] = 32'b11111111111111111101001000101110;
assign LUT_2[18699] = 32'b11111111111111111010000001000111;
assign LUT_2[18700] = 32'b11111111111111110010101101011010;
assign LUT_2[18701] = 32'b11111111111111101111100101110011;
assign LUT_2[18702] = 32'b11111111111111111001100110010110;
assign LUT_2[18703] = 32'b11111111111111110110011110101111;
assign LUT_2[18704] = 32'b11111111111111110110000010011111;
assign LUT_2[18705] = 32'b11111111111111110010111010111000;
assign LUT_2[18706] = 32'b11111111111111111100111011011011;
assign LUT_2[18707] = 32'b11111111111111111001110011110100;
assign LUT_2[18708] = 32'b11111111111111110010100000000111;
assign LUT_2[18709] = 32'b11111111111111101111011000100000;
assign LUT_2[18710] = 32'b11111111111111111001011001000011;
assign LUT_2[18711] = 32'b11111111111111110110010001011100;
assign LUT_2[18712] = 32'b11111111111111110000110011111100;
assign LUT_2[18713] = 32'b11111111111111101101101100010101;
assign LUT_2[18714] = 32'b11111111111111110111101100111000;
assign LUT_2[18715] = 32'b11111111111111110100100101010001;
assign LUT_2[18716] = 32'b11111111111111101101010001100100;
assign LUT_2[18717] = 32'b11111111111111101010001001111101;
assign LUT_2[18718] = 32'b11111111111111110100001010100000;
assign LUT_2[18719] = 32'b11111111111111110001000010111001;
assign LUT_2[18720] = 32'b11111111111111111011111001111110;
assign LUT_2[18721] = 32'b11111111111111111000110010010111;
assign LUT_2[18722] = 32'b00000000000000000010110010111010;
assign LUT_2[18723] = 32'b11111111111111111111101011010011;
assign LUT_2[18724] = 32'b11111111111111111000010111100110;
assign LUT_2[18725] = 32'b11111111111111110101001111111111;
assign LUT_2[18726] = 32'b11111111111111111111010000100010;
assign LUT_2[18727] = 32'b11111111111111111100001000111011;
assign LUT_2[18728] = 32'b11111111111111110110101011011011;
assign LUT_2[18729] = 32'b11111111111111110011100011110100;
assign LUT_2[18730] = 32'b11111111111111111101100100010111;
assign LUT_2[18731] = 32'b11111111111111111010011100110000;
assign LUT_2[18732] = 32'b11111111111111110011001001000011;
assign LUT_2[18733] = 32'b11111111111111110000000001011100;
assign LUT_2[18734] = 32'b11111111111111111010000001111111;
assign LUT_2[18735] = 32'b11111111111111110110111010011000;
assign LUT_2[18736] = 32'b11111111111111110110011110001000;
assign LUT_2[18737] = 32'b11111111111111110011010110100001;
assign LUT_2[18738] = 32'b11111111111111111101010111000100;
assign LUT_2[18739] = 32'b11111111111111111010001111011101;
assign LUT_2[18740] = 32'b11111111111111110010111011110000;
assign LUT_2[18741] = 32'b11111111111111101111110100001001;
assign LUT_2[18742] = 32'b11111111111111111001110100101100;
assign LUT_2[18743] = 32'b11111111111111110110101101000101;
assign LUT_2[18744] = 32'b11111111111111110001001111100101;
assign LUT_2[18745] = 32'b11111111111111101110000111111110;
assign LUT_2[18746] = 32'b11111111111111111000001000100001;
assign LUT_2[18747] = 32'b11111111111111110101000000111010;
assign LUT_2[18748] = 32'b11111111111111101101101101001101;
assign LUT_2[18749] = 32'b11111111111111101010100101100110;
assign LUT_2[18750] = 32'b11111111111111110100100110001001;
assign LUT_2[18751] = 32'b11111111111111110001011110100010;
assign LUT_2[18752] = 32'b11111111111111110011100110111000;
assign LUT_2[18753] = 32'b11111111111111110000011111010001;
assign LUT_2[18754] = 32'b11111111111111111010011111110100;
assign LUT_2[18755] = 32'b11111111111111110111011000001101;
assign LUT_2[18756] = 32'b11111111111111110000000100100000;
assign LUT_2[18757] = 32'b11111111111111101100111100111001;
assign LUT_2[18758] = 32'b11111111111111110110111101011100;
assign LUT_2[18759] = 32'b11111111111111110011110101110101;
assign LUT_2[18760] = 32'b11111111111111101110011000010101;
assign LUT_2[18761] = 32'b11111111111111101011010000101110;
assign LUT_2[18762] = 32'b11111111111111110101010001010001;
assign LUT_2[18763] = 32'b11111111111111110010001001101010;
assign LUT_2[18764] = 32'b11111111111111101010110101111101;
assign LUT_2[18765] = 32'b11111111111111100111101110010110;
assign LUT_2[18766] = 32'b11111111111111110001101110111001;
assign LUT_2[18767] = 32'b11111111111111101110100111010010;
assign LUT_2[18768] = 32'b11111111111111101110001011000010;
assign LUT_2[18769] = 32'b11111111111111101011000011011011;
assign LUT_2[18770] = 32'b11111111111111110101000011111110;
assign LUT_2[18771] = 32'b11111111111111110001111100010111;
assign LUT_2[18772] = 32'b11111111111111101010101000101010;
assign LUT_2[18773] = 32'b11111111111111100111100001000011;
assign LUT_2[18774] = 32'b11111111111111110001100001100110;
assign LUT_2[18775] = 32'b11111111111111101110011001111111;
assign LUT_2[18776] = 32'b11111111111111101000111100011111;
assign LUT_2[18777] = 32'b11111111111111100101110100111000;
assign LUT_2[18778] = 32'b11111111111111101111110101011011;
assign LUT_2[18779] = 32'b11111111111111101100101101110100;
assign LUT_2[18780] = 32'b11111111111111100101011010000111;
assign LUT_2[18781] = 32'b11111111111111100010010010100000;
assign LUT_2[18782] = 32'b11111111111111101100010011000011;
assign LUT_2[18783] = 32'b11111111111111101001001011011100;
assign LUT_2[18784] = 32'b11111111111111110100000010100001;
assign LUT_2[18785] = 32'b11111111111111110000111010111010;
assign LUT_2[18786] = 32'b11111111111111111010111011011101;
assign LUT_2[18787] = 32'b11111111111111110111110011110110;
assign LUT_2[18788] = 32'b11111111111111110000100000001001;
assign LUT_2[18789] = 32'b11111111111111101101011000100010;
assign LUT_2[18790] = 32'b11111111111111110111011001000101;
assign LUT_2[18791] = 32'b11111111111111110100010001011110;
assign LUT_2[18792] = 32'b11111111111111101110110011111110;
assign LUT_2[18793] = 32'b11111111111111101011101100010111;
assign LUT_2[18794] = 32'b11111111111111110101101100111010;
assign LUT_2[18795] = 32'b11111111111111110010100101010011;
assign LUT_2[18796] = 32'b11111111111111101011010001100110;
assign LUT_2[18797] = 32'b11111111111111101000001001111111;
assign LUT_2[18798] = 32'b11111111111111110010001010100010;
assign LUT_2[18799] = 32'b11111111111111101111000010111011;
assign LUT_2[18800] = 32'b11111111111111101110100110101011;
assign LUT_2[18801] = 32'b11111111111111101011011111000100;
assign LUT_2[18802] = 32'b11111111111111110101011111100111;
assign LUT_2[18803] = 32'b11111111111111110010011000000000;
assign LUT_2[18804] = 32'b11111111111111101011000100010011;
assign LUT_2[18805] = 32'b11111111111111100111111100101100;
assign LUT_2[18806] = 32'b11111111111111110001111101001111;
assign LUT_2[18807] = 32'b11111111111111101110110101101000;
assign LUT_2[18808] = 32'b11111111111111101001011000001000;
assign LUT_2[18809] = 32'b11111111111111100110010000100001;
assign LUT_2[18810] = 32'b11111111111111110000010001000100;
assign LUT_2[18811] = 32'b11111111111111101101001001011101;
assign LUT_2[18812] = 32'b11111111111111100101110101110000;
assign LUT_2[18813] = 32'b11111111111111100010101110001001;
assign LUT_2[18814] = 32'b11111111111111101100101110101100;
assign LUT_2[18815] = 32'b11111111111111101001100111000101;
assign LUT_2[18816] = 32'b11111111111111111111110010100100;
assign LUT_2[18817] = 32'b11111111111111111100101010111101;
assign LUT_2[18818] = 32'b00000000000000000110101011100000;
assign LUT_2[18819] = 32'b00000000000000000011100011111001;
assign LUT_2[18820] = 32'b11111111111111111100010000001100;
assign LUT_2[18821] = 32'b11111111111111111001001000100101;
assign LUT_2[18822] = 32'b00000000000000000011001001001000;
assign LUT_2[18823] = 32'b00000000000000000000000001100001;
assign LUT_2[18824] = 32'b11111111111111111010100100000001;
assign LUT_2[18825] = 32'b11111111111111110111011100011010;
assign LUT_2[18826] = 32'b00000000000000000001011100111101;
assign LUT_2[18827] = 32'b11111111111111111110010101010110;
assign LUT_2[18828] = 32'b11111111111111110111000001101001;
assign LUT_2[18829] = 32'b11111111111111110011111010000010;
assign LUT_2[18830] = 32'b11111111111111111101111010100101;
assign LUT_2[18831] = 32'b11111111111111111010110010111110;
assign LUT_2[18832] = 32'b11111111111111111010010110101110;
assign LUT_2[18833] = 32'b11111111111111110111001111000111;
assign LUT_2[18834] = 32'b00000000000000000001001111101010;
assign LUT_2[18835] = 32'b11111111111111111110001000000011;
assign LUT_2[18836] = 32'b11111111111111110110110100010110;
assign LUT_2[18837] = 32'b11111111111111110011101100101111;
assign LUT_2[18838] = 32'b11111111111111111101101101010010;
assign LUT_2[18839] = 32'b11111111111111111010100101101011;
assign LUT_2[18840] = 32'b11111111111111110101001000001011;
assign LUT_2[18841] = 32'b11111111111111110010000000100100;
assign LUT_2[18842] = 32'b11111111111111111100000001000111;
assign LUT_2[18843] = 32'b11111111111111111000111001100000;
assign LUT_2[18844] = 32'b11111111111111110001100101110011;
assign LUT_2[18845] = 32'b11111111111111101110011110001100;
assign LUT_2[18846] = 32'b11111111111111111000011110101111;
assign LUT_2[18847] = 32'b11111111111111110101010111001000;
assign LUT_2[18848] = 32'b00000000000000000000001110001101;
assign LUT_2[18849] = 32'b11111111111111111101000110100110;
assign LUT_2[18850] = 32'b00000000000000000111000111001001;
assign LUT_2[18851] = 32'b00000000000000000011111111100010;
assign LUT_2[18852] = 32'b11111111111111111100101011110101;
assign LUT_2[18853] = 32'b11111111111111111001100100001110;
assign LUT_2[18854] = 32'b00000000000000000011100100110001;
assign LUT_2[18855] = 32'b00000000000000000000011101001010;
assign LUT_2[18856] = 32'b11111111111111111010111111101010;
assign LUT_2[18857] = 32'b11111111111111110111111000000011;
assign LUT_2[18858] = 32'b00000000000000000001111000100110;
assign LUT_2[18859] = 32'b11111111111111111110110000111111;
assign LUT_2[18860] = 32'b11111111111111110111011101010010;
assign LUT_2[18861] = 32'b11111111111111110100010101101011;
assign LUT_2[18862] = 32'b11111111111111111110010110001110;
assign LUT_2[18863] = 32'b11111111111111111011001110100111;
assign LUT_2[18864] = 32'b11111111111111111010110010010111;
assign LUT_2[18865] = 32'b11111111111111110111101010110000;
assign LUT_2[18866] = 32'b00000000000000000001101011010011;
assign LUT_2[18867] = 32'b11111111111111111110100011101100;
assign LUT_2[18868] = 32'b11111111111111110111001111111111;
assign LUT_2[18869] = 32'b11111111111111110100001000011000;
assign LUT_2[18870] = 32'b11111111111111111110001000111011;
assign LUT_2[18871] = 32'b11111111111111111011000001010100;
assign LUT_2[18872] = 32'b11111111111111110101100011110100;
assign LUT_2[18873] = 32'b11111111111111110010011100001101;
assign LUT_2[18874] = 32'b11111111111111111100011100110000;
assign LUT_2[18875] = 32'b11111111111111111001010101001001;
assign LUT_2[18876] = 32'b11111111111111110010000001011100;
assign LUT_2[18877] = 32'b11111111111111101110111001110101;
assign LUT_2[18878] = 32'b11111111111111111000111010011000;
assign LUT_2[18879] = 32'b11111111111111110101110010110001;
assign LUT_2[18880] = 32'b11111111111111110111111011000111;
assign LUT_2[18881] = 32'b11111111111111110100110011100000;
assign LUT_2[18882] = 32'b11111111111111111110110100000011;
assign LUT_2[18883] = 32'b11111111111111111011101100011100;
assign LUT_2[18884] = 32'b11111111111111110100011000101111;
assign LUT_2[18885] = 32'b11111111111111110001010001001000;
assign LUT_2[18886] = 32'b11111111111111111011010001101011;
assign LUT_2[18887] = 32'b11111111111111111000001010000100;
assign LUT_2[18888] = 32'b11111111111111110010101100100100;
assign LUT_2[18889] = 32'b11111111111111101111100100111101;
assign LUT_2[18890] = 32'b11111111111111111001100101100000;
assign LUT_2[18891] = 32'b11111111111111110110011101111001;
assign LUT_2[18892] = 32'b11111111111111101111001010001100;
assign LUT_2[18893] = 32'b11111111111111101100000010100101;
assign LUT_2[18894] = 32'b11111111111111110110000011001000;
assign LUT_2[18895] = 32'b11111111111111110010111011100001;
assign LUT_2[18896] = 32'b11111111111111110010011111010001;
assign LUT_2[18897] = 32'b11111111111111101111010111101010;
assign LUT_2[18898] = 32'b11111111111111111001011000001101;
assign LUT_2[18899] = 32'b11111111111111110110010000100110;
assign LUT_2[18900] = 32'b11111111111111101110111100111001;
assign LUT_2[18901] = 32'b11111111111111101011110101010010;
assign LUT_2[18902] = 32'b11111111111111110101110101110101;
assign LUT_2[18903] = 32'b11111111111111110010101110001110;
assign LUT_2[18904] = 32'b11111111111111101101010000101110;
assign LUT_2[18905] = 32'b11111111111111101010001001000111;
assign LUT_2[18906] = 32'b11111111111111110100001001101010;
assign LUT_2[18907] = 32'b11111111111111110001000010000011;
assign LUT_2[18908] = 32'b11111111111111101001101110010110;
assign LUT_2[18909] = 32'b11111111111111100110100110101111;
assign LUT_2[18910] = 32'b11111111111111110000100111010010;
assign LUT_2[18911] = 32'b11111111111111101101011111101011;
assign LUT_2[18912] = 32'b11111111111111111000010110110000;
assign LUT_2[18913] = 32'b11111111111111110101001111001001;
assign LUT_2[18914] = 32'b11111111111111111111001111101100;
assign LUT_2[18915] = 32'b11111111111111111100001000000101;
assign LUT_2[18916] = 32'b11111111111111110100110100011000;
assign LUT_2[18917] = 32'b11111111111111110001101100110001;
assign LUT_2[18918] = 32'b11111111111111111011101101010100;
assign LUT_2[18919] = 32'b11111111111111111000100101101101;
assign LUT_2[18920] = 32'b11111111111111110011001000001101;
assign LUT_2[18921] = 32'b11111111111111110000000000100110;
assign LUT_2[18922] = 32'b11111111111111111010000001001001;
assign LUT_2[18923] = 32'b11111111111111110110111001100010;
assign LUT_2[18924] = 32'b11111111111111101111100101110101;
assign LUT_2[18925] = 32'b11111111111111101100011110001110;
assign LUT_2[18926] = 32'b11111111111111110110011110110001;
assign LUT_2[18927] = 32'b11111111111111110011010111001010;
assign LUT_2[18928] = 32'b11111111111111110010111010111010;
assign LUT_2[18929] = 32'b11111111111111101111110011010011;
assign LUT_2[18930] = 32'b11111111111111111001110011110110;
assign LUT_2[18931] = 32'b11111111111111110110101100001111;
assign LUT_2[18932] = 32'b11111111111111101111011000100010;
assign LUT_2[18933] = 32'b11111111111111101100010000111011;
assign LUT_2[18934] = 32'b11111111111111110110010001011110;
assign LUT_2[18935] = 32'b11111111111111110011001001110111;
assign LUT_2[18936] = 32'b11111111111111101101101100010111;
assign LUT_2[18937] = 32'b11111111111111101010100100110000;
assign LUT_2[18938] = 32'b11111111111111110100100101010011;
assign LUT_2[18939] = 32'b11111111111111110001011101101100;
assign LUT_2[18940] = 32'b11111111111111101010001001111111;
assign LUT_2[18941] = 32'b11111111111111100111000010011000;
assign LUT_2[18942] = 32'b11111111111111110001000010111011;
assign LUT_2[18943] = 32'b11111111111111101101111011010100;
assign LUT_2[18944] = 32'b11111111111111111100010001100001;
assign LUT_2[18945] = 32'b11111111111111111001001001111010;
assign LUT_2[18946] = 32'b00000000000000000011001010011101;
assign LUT_2[18947] = 32'b00000000000000000000000010110110;
assign LUT_2[18948] = 32'b11111111111111111000101111001001;
assign LUT_2[18949] = 32'b11111111111111110101100111100010;
assign LUT_2[18950] = 32'b11111111111111111111101000000101;
assign LUT_2[18951] = 32'b11111111111111111100100000011110;
assign LUT_2[18952] = 32'b11111111111111110111000010111110;
assign LUT_2[18953] = 32'b11111111111111110011111011010111;
assign LUT_2[18954] = 32'b11111111111111111101111011111010;
assign LUT_2[18955] = 32'b11111111111111111010110100010011;
assign LUT_2[18956] = 32'b11111111111111110011100000100110;
assign LUT_2[18957] = 32'b11111111111111110000011000111111;
assign LUT_2[18958] = 32'b11111111111111111010011001100010;
assign LUT_2[18959] = 32'b11111111111111110111010001111011;
assign LUT_2[18960] = 32'b11111111111111110110110101101011;
assign LUT_2[18961] = 32'b11111111111111110011101110000100;
assign LUT_2[18962] = 32'b11111111111111111101101110100111;
assign LUT_2[18963] = 32'b11111111111111111010100111000000;
assign LUT_2[18964] = 32'b11111111111111110011010011010011;
assign LUT_2[18965] = 32'b11111111111111110000001011101100;
assign LUT_2[18966] = 32'b11111111111111111010001100001111;
assign LUT_2[18967] = 32'b11111111111111110111000100101000;
assign LUT_2[18968] = 32'b11111111111111110001100111001000;
assign LUT_2[18969] = 32'b11111111111111101110011111100001;
assign LUT_2[18970] = 32'b11111111111111111000100000000100;
assign LUT_2[18971] = 32'b11111111111111110101011000011101;
assign LUT_2[18972] = 32'b11111111111111101110000100110000;
assign LUT_2[18973] = 32'b11111111111111101010111101001001;
assign LUT_2[18974] = 32'b11111111111111110100111101101100;
assign LUT_2[18975] = 32'b11111111111111110001110110000101;
assign LUT_2[18976] = 32'b11111111111111111100101101001010;
assign LUT_2[18977] = 32'b11111111111111111001100101100011;
assign LUT_2[18978] = 32'b00000000000000000011100110000110;
assign LUT_2[18979] = 32'b00000000000000000000011110011111;
assign LUT_2[18980] = 32'b11111111111111111001001010110010;
assign LUT_2[18981] = 32'b11111111111111110110000011001011;
assign LUT_2[18982] = 32'b00000000000000000000000011101110;
assign LUT_2[18983] = 32'b11111111111111111100111100000111;
assign LUT_2[18984] = 32'b11111111111111110111011110100111;
assign LUT_2[18985] = 32'b11111111111111110100010111000000;
assign LUT_2[18986] = 32'b11111111111111111110010111100011;
assign LUT_2[18987] = 32'b11111111111111111011001111111100;
assign LUT_2[18988] = 32'b11111111111111110011111100001111;
assign LUT_2[18989] = 32'b11111111111111110000110100101000;
assign LUT_2[18990] = 32'b11111111111111111010110101001011;
assign LUT_2[18991] = 32'b11111111111111110111101101100100;
assign LUT_2[18992] = 32'b11111111111111110111010001010100;
assign LUT_2[18993] = 32'b11111111111111110100001001101101;
assign LUT_2[18994] = 32'b11111111111111111110001010010000;
assign LUT_2[18995] = 32'b11111111111111111011000010101001;
assign LUT_2[18996] = 32'b11111111111111110011101110111100;
assign LUT_2[18997] = 32'b11111111111111110000100111010101;
assign LUT_2[18998] = 32'b11111111111111111010100111111000;
assign LUT_2[18999] = 32'b11111111111111110111100000010001;
assign LUT_2[19000] = 32'b11111111111111110010000010110001;
assign LUT_2[19001] = 32'b11111111111111101110111011001010;
assign LUT_2[19002] = 32'b11111111111111111000111011101101;
assign LUT_2[19003] = 32'b11111111111111110101110100000110;
assign LUT_2[19004] = 32'b11111111111111101110100000011001;
assign LUT_2[19005] = 32'b11111111111111101011011000110010;
assign LUT_2[19006] = 32'b11111111111111110101011001010101;
assign LUT_2[19007] = 32'b11111111111111110010010001101110;
assign LUT_2[19008] = 32'b11111111111111110100011010000100;
assign LUT_2[19009] = 32'b11111111111111110001010010011101;
assign LUT_2[19010] = 32'b11111111111111111011010011000000;
assign LUT_2[19011] = 32'b11111111111111111000001011011001;
assign LUT_2[19012] = 32'b11111111111111110000110111101100;
assign LUT_2[19013] = 32'b11111111111111101101110000000101;
assign LUT_2[19014] = 32'b11111111111111110111110000101000;
assign LUT_2[19015] = 32'b11111111111111110100101001000001;
assign LUT_2[19016] = 32'b11111111111111101111001011100001;
assign LUT_2[19017] = 32'b11111111111111101100000011111010;
assign LUT_2[19018] = 32'b11111111111111110110000100011101;
assign LUT_2[19019] = 32'b11111111111111110010111100110110;
assign LUT_2[19020] = 32'b11111111111111101011101001001001;
assign LUT_2[19021] = 32'b11111111111111101000100001100010;
assign LUT_2[19022] = 32'b11111111111111110010100010000101;
assign LUT_2[19023] = 32'b11111111111111101111011010011110;
assign LUT_2[19024] = 32'b11111111111111101110111110001110;
assign LUT_2[19025] = 32'b11111111111111101011110110100111;
assign LUT_2[19026] = 32'b11111111111111110101110111001010;
assign LUT_2[19027] = 32'b11111111111111110010101111100011;
assign LUT_2[19028] = 32'b11111111111111101011011011110110;
assign LUT_2[19029] = 32'b11111111111111101000010100001111;
assign LUT_2[19030] = 32'b11111111111111110010010100110010;
assign LUT_2[19031] = 32'b11111111111111101111001101001011;
assign LUT_2[19032] = 32'b11111111111111101001101111101011;
assign LUT_2[19033] = 32'b11111111111111100110101000000100;
assign LUT_2[19034] = 32'b11111111111111110000101000100111;
assign LUT_2[19035] = 32'b11111111111111101101100001000000;
assign LUT_2[19036] = 32'b11111111111111100110001101010011;
assign LUT_2[19037] = 32'b11111111111111100011000101101100;
assign LUT_2[19038] = 32'b11111111111111101101000110001111;
assign LUT_2[19039] = 32'b11111111111111101001111110101000;
assign LUT_2[19040] = 32'b11111111111111110100110101101101;
assign LUT_2[19041] = 32'b11111111111111110001101110000110;
assign LUT_2[19042] = 32'b11111111111111111011101110101001;
assign LUT_2[19043] = 32'b11111111111111111000100111000010;
assign LUT_2[19044] = 32'b11111111111111110001010011010101;
assign LUT_2[19045] = 32'b11111111111111101110001011101110;
assign LUT_2[19046] = 32'b11111111111111111000001100010001;
assign LUT_2[19047] = 32'b11111111111111110101000100101010;
assign LUT_2[19048] = 32'b11111111111111101111100111001010;
assign LUT_2[19049] = 32'b11111111111111101100011111100011;
assign LUT_2[19050] = 32'b11111111111111110110100000000110;
assign LUT_2[19051] = 32'b11111111111111110011011000011111;
assign LUT_2[19052] = 32'b11111111111111101100000100110010;
assign LUT_2[19053] = 32'b11111111111111101000111101001011;
assign LUT_2[19054] = 32'b11111111111111110010111101101110;
assign LUT_2[19055] = 32'b11111111111111101111110110000111;
assign LUT_2[19056] = 32'b11111111111111101111011001110111;
assign LUT_2[19057] = 32'b11111111111111101100010010010000;
assign LUT_2[19058] = 32'b11111111111111110110010010110011;
assign LUT_2[19059] = 32'b11111111111111110011001011001100;
assign LUT_2[19060] = 32'b11111111111111101011110111011111;
assign LUT_2[19061] = 32'b11111111111111101000101111111000;
assign LUT_2[19062] = 32'b11111111111111110010110000011011;
assign LUT_2[19063] = 32'b11111111111111101111101000110100;
assign LUT_2[19064] = 32'b11111111111111101010001011010100;
assign LUT_2[19065] = 32'b11111111111111100111000011101101;
assign LUT_2[19066] = 32'b11111111111111110001000100010000;
assign LUT_2[19067] = 32'b11111111111111101101111100101001;
assign LUT_2[19068] = 32'b11111111111111100110101000111100;
assign LUT_2[19069] = 32'b11111111111111100011100001010101;
assign LUT_2[19070] = 32'b11111111111111101101100001111000;
assign LUT_2[19071] = 32'b11111111111111101010011010010001;
assign LUT_2[19072] = 32'b00000000000000000000100101110000;
assign LUT_2[19073] = 32'b11111111111111111101011110001001;
assign LUT_2[19074] = 32'b00000000000000000111011110101100;
assign LUT_2[19075] = 32'b00000000000000000100010111000101;
assign LUT_2[19076] = 32'b11111111111111111101000011011000;
assign LUT_2[19077] = 32'b11111111111111111001111011110001;
assign LUT_2[19078] = 32'b00000000000000000011111100010100;
assign LUT_2[19079] = 32'b00000000000000000000110100101101;
assign LUT_2[19080] = 32'b11111111111111111011010111001101;
assign LUT_2[19081] = 32'b11111111111111111000001111100110;
assign LUT_2[19082] = 32'b00000000000000000010010000001001;
assign LUT_2[19083] = 32'b11111111111111111111001000100010;
assign LUT_2[19084] = 32'b11111111111111110111110100110101;
assign LUT_2[19085] = 32'b11111111111111110100101101001110;
assign LUT_2[19086] = 32'b11111111111111111110101101110001;
assign LUT_2[19087] = 32'b11111111111111111011100110001010;
assign LUT_2[19088] = 32'b11111111111111111011001001111010;
assign LUT_2[19089] = 32'b11111111111111111000000010010011;
assign LUT_2[19090] = 32'b00000000000000000010000010110110;
assign LUT_2[19091] = 32'b11111111111111111110111011001111;
assign LUT_2[19092] = 32'b11111111111111110111100111100010;
assign LUT_2[19093] = 32'b11111111111111110100011111111011;
assign LUT_2[19094] = 32'b11111111111111111110100000011110;
assign LUT_2[19095] = 32'b11111111111111111011011000110111;
assign LUT_2[19096] = 32'b11111111111111110101111011010111;
assign LUT_2[19097] = 32'b11111111111111110010110011110000;
assign LUT_2[19098] = 32'b11111111111111111100110100010011;
assign LUT_2[19099] = 32'b11111111111111111001101100101100;
assign LUT_2[19100] = 32'b11111111111111110010011000111111;
assign LUT_2[19101] = 32'b11111111111111101111010001011000;
assign LUT_2[19102] = 32'b11111111111111111001010001111011;
assign LUT_2[19103] = 32'b11111111111111110110001010010100;
assign LUT_2[19104] = 32'b00000000000000000001000001011001;
assign LUT_2[19105] = 32'b11111111111111111101111001110010;
assign LUT_2[19106] = 32'b00000000000000000111111010010101;
assign LUT_2[19107] = 32'b00000000000000000100110010101110;
assign LUT_2[19108] = 32'b11111111111111111101011111000001;
assign LUT_2[19109] = 32'b11111111111111111010010111011010;
assign LUT_2[19110] = 32'b00000000000000000100010111111101;
assign LUT_2[19111] = 32'b00000000000000000001010000010110;
assign LUT_2[19112] = 32'b11111111111111111011110010110110;
assign LUT_2[19113] = 32'b11111111111111111000101011001111;
assign LUT_2[19114] = 32'b00000000000000000010101011110010;
assign LUT_2[19115] = 32'b11111111111111111111100100001011;
assign LUT_2[19116] = 32'b11111111111111111000010000011110;
assign LUT_2[19117] = 32'b11111111111111110101001000110111;
assign LUT_2[19118] = 32'b11111111111111111111001001011010;
assign LUT_2[19119] = 32'b11111111111111111100000001110011;
assign LUT_2[19120] = 32'b11111111111111111011100101100011;
assign LUT_2[19121] = 32'b11111111111111111000011101111100;
assign LUT_2[19122] = 32'b00000000000000000010011110011111;
assign LUT_2[19123] = 32'b11111111111111111111010110111000;
assign LUT_2[19124] = 32'b11111111111111111000000011001011;
assign LUT_2[19125] = 32'b11111111111111110100111011100100;
assign LUT_2[19126] = 32'b11111111111111111110111100000111;
assign LUT_2[19127] = 32'b11111111111111111011110100100000;
assign LUT_2[19128] = 32'b11111111111111110110010111000000;
assign LUT_2[19129] = 32'b11111111111111110011001111011001;
assign LUT_2[19130] = 32'b11111111111111111101001111111100;
assign LUT_2[19131] = 32'b11111111111111111010001000010101;
assign LUT_2[19132] = 32'b11111111111111110010110100101000;
assign LUT_2[19133] = 32'b11111111111111101111101101000001;
assign LUT_2[19134] = 32'b11111111111111111001101101100100;
assign LUT_2[19135] = 32'b11111111111111110110100101111101;
assign LUT_2[19136] = 32'b11111111111111111000101110010011;
assign LUT_2[19137] = 32'b11111111111111110101100110101100;
assign LUT_2[19138] = 32'b11111111111111111111100111001111;
assign LUT_2[19139] = 32'b11111111111111111100011111101000;
assign LUT_2[19140] = 32'b11111111111111110101001011111011;
assign LUT_2[19141] = 32'b11111111111111110010000100010100;
assign LUT_2[19142] = 32'b11111111111111111100000100110111;
assign LUT_2[19143] = 32'b11111111111111111000111101010000;
assign LUT_2[19144] = 32'b11111111111111110011011111110000;
assign LUT_2[19145] = 32'b11111111111111110000011000001001;
assign LUT_2[19146] = 32'b11111111111111111010011000101100;
assign LUT_2[19147] = 32'b11111111111111110111010001000101;
assign LUT_2[19148] = 32'b11111111111111101111111101011000;
assign LUT_2[19149] = 32'b11111111111111101100110101110001;
assign LUT_2[19150] = 32'b11111111111111110110110110010100;
assign LUT_2[19151] = 32'b11111111111111110011101110101101;
assign LUT_2[19152] = 32'b11111111111111110011010010011101;
assign LUT_2[19153] = 32'b11111111111111110000001010110110;
assign LUT_2[19154] = 32'b11111111111111111010001011011001;
assign LUT_2[19155] = 32'b11111111111111110111000011110010;
assign LUT_2[19156] = 32'b11111111111111101111110000000101;
assign LUT_2[19157] = 32'b11111111111111101100101000011110;
assign LUT_2[19158] = 32'b11111111111111110110101001000001;
assign LUT_2[19159] = 32'b11111111111111110011100001011010;
assign LUT_2[19160] = 32'b11111111111111101110000011111010;
assign LUT_2[19161] = 32'b11111111111111101010111100010011;
assign LUT_2[19162] = 32'b11111111111111110100111100110110;
assign LUT_2[19163] = 32'b11111111111111110001110101001111;
assign LUT_2[19164] = 32'b11111111111111101010100001100010;
assign LUT_2[19165] = 32'b11111111111111100111011001111011;
assign LUT_2[19166] = 32'b11111111111111110001011010011110;
assign LUT_2[19167] = 32'b11111111111111101110010010110111;
assign LUT_2[19168] = 32'b11111111111111111001001001111100;
assign LUT_2[19169] = 32'b11111111111111110110000010010101;
assign LUT_2[19170] = 32'b00000000000000000000000010111000;
assign LUT_2[19171] = 32'b11111111111111111100111011010001;
assign LUT_2[19172] = 32'b11111111111111110101100111100100;
assign LUT_2[19173] = 32'b11111111111111110010011111111101;
assign LUT_2[19174] = 32'b11111111111111111100100000100000;
assign LUT_2[19175] = 32'b11111111111111111001011000111001;
assign LUT_2[19176] = 32'b11111111111111110011111011011001;
assign LUT_2[19177] = 32'b11111111111111110000110011110010;
assign LUT_2[19178] = 32'b11111111111111111010110100010101;
assign LUT_2[19179] = 32'b11111111111111110111101100101110;
assign LUT_2[19180] = 32'b11111111111111110000011001000001;
assign LUT_2[19181] = 32'b11111111111111101101010001011010;
assign LUT_2[19182] = 32'b11111111111111110111010001111101;
assign LUT_2[19183] = 32'b11111111111111110100001010010110;
assign LUT_2[19184] = 32'b11111111111111110011101110000110;
assign LUT_2[19185] = 32'b11111111111111110000100110011111;
assign LUT_2[19186] = 32'b11111111111111111010100111000010;
assign LUT_2[19187] = 32'b11111111111111110111011111011011;
assign LUT_2[19188] = 32'b11111111111111110000001011101110;
assign LUT_2[19189] = 32'b11111111111111101101000100000111;
assign LUT_2[19190] = 32'b11111111111111110111000100101010;
assign LUT_2[19191] = 32'b11111111111111110011111101000011;
assign LUT_2[19192] = 32'b11111111111111101110011111100011;
assign LUT_2[19193] = 32'b11111111111111101011010111111100;
assign LUT_2[19194] = 32'b11111111111111110101011000011111;
assign LUT_2[19195] = 32'b11111111111111110010010000111000;
assign LUT_2[19196] = 32'b11111111111111101010111101001011;
assign LUT_2[19197] = 32'b11111111111111100111110101100100;
assign LUT_2[19198] = 32'b11111111111111110001110110000111;
assign LUT_2[19199] = 32'b11111111111111101110101110100000;
assign LUT_2[19200] = 32'b00000000000000000000010000000111;
assign LUT_2[19201] = 32'b11111111111111111101001000100000;
assign LUT_2[19202] = 32'b00000000000000000111001001000011;
assign LUT_2[19203] = 32'b00000000000000000100000001011100;
assign LUT_2[19204] = 32'b11111111111111111100101101101111;
assign LUT_2[19205] = 32'b11111111111111111001100110001000;
assign LUT_2[19206] = 32'b00000000000000000011100110101011;
assign LUT_2[19207] = 32'b00000000000000000000011111000100;
assign LUT_2[19208] = 32'b11111111111111111011000001100100;
assign LUT_2[19209] = 32'b11111111111111110111111001111101;
assign LUT_2[19210] = 32'b00000000000000000001111010100000;
assign LUT_2[19211] = 32'b11111111111111111110110010111001;
assign LUT_2[19212] = 32'b11111111111111110111011111001100;
assign LUT_2[19213] = 32'b11111111111111110100010111100101;
assign LUT_2[19214] = 32'b11111111111111111110011000001000;
assign LUT_2[19215] = 32'b11111111111111111011010000100001;
assign LUT_2[19216] = 32'b11111111111111111010110100010001;
assign LUT_2[19217] = 32'b11111111111111110111101100101010;
assign LUT_2[19218] = 32'b00000000000000000001101101001101;
assign LUT_2[19219] = 32'b11111111111111111110100101100110;
assign LUT_2[19220] = 32'b11111111111111110111010001111001;
assign LUT_2[19221] = 32'b11111111111111110100001010010010;
assign LUT_2[19222] = 32'b11111111111111111110001010110101;
assign LUT_2[19223] = 32'b11111111111111111011000011001110;
assign LUT_2[19224] = 32'b11111111111111110101100101101110;
assign LUT_2[19225] = 32'b11111111111111110010011110000111;
assign LUT_2[19226] = 32'b11111111111111111100011110101010;
assign LUT_2[19227] = 32'b11111111111111111001010111000011;
assign LUT_2[19228] = 32'b11111111111111110010000011010110;
assign LUT_2[19229] = 32'b11111111111111101110111011101111;
assign LUT_2[19230] = 32'b11111111111111111000111100010010;
assign LUT_2[19231] = 32'b11111111111111110101110100101011;
assign LUT_2[19232] = 32'b00000000000000000000101011110000;
assign LUT_2[19233] = 32'b11111111111111111101100100001001;
assign LUT_2[19234] = 32'b00000000000000000111100100101100;
assign LUT_2[19235] = 32'b00000000000000000100011101000101;
assign LUT_2[19236] = 32'b11111111111111111101001001011000;
assign LUT_2[19237] = 32'b11111111111111111010000001110001;
assign LUT_2[19238] = 32'b00000000000000000100000010010100;
assign LUT_2[19239] = 32'b00000000000000000000111010101101;
assign LUT_2[19240] = 32'b11111111111111111011011101001101;
assign LUT_2[19241] = 32'b11111111111111111000010101100110;
assign LUT_2[19242] = 32'b00000000000000000010010110001001;
assign LUT_2[19243] = 32'b11111111111111111111001110100010;
assign LUT_2[19244] = 32'b11111111111111110111111010110101;
assign LUT_2[19245] = 32'b11111111111111110100110011001110;
assign LUT_2[19246] = 32'b11111111111111111110110011110001;
assign LUT_2[19247] = 32'b11111111111111111011101100001010;
assign LUT_2[19248] = 32'b11111111111111111011001111111010;
assign LUT_2[19249] = 32'b11111111111111111000001000010011;
assign LUT_2[19250] = 32'b00000000000000000010001000110110;
assign LUT_2[19251] = 32'b11111111111111111111000001001111;
assign LUT_2[19252] = 32'b11111111111111110111101101100010;
assign LUT_2[19253] = 32'b11111111111111110100100101111011;
assign LUT_2[19254] = 32'b11111111111111111110100110011110;
assign LUT_2[19255] = 32'b11111111111111111011011110110111;
assign LUT_2[19256] = 32'b11111111111111110110000001010111;
assign LUT_2[19257] = 32'b11111111111111110010111001110000;
assign LUT_2[19258] = 32'b11111111111111111100111010010011;
assign LUT_2[19259] = 32'b11111111111111111001110010101100;
assign LUT_2[19260] = 32'b11111111111111110010011110111111;
assign LUT_2[19261] = 32'b11111111111111101111010111011000;
assign LUT_2[19262] = 32'b11111111111111111001010111111011;
assign LUT_2[19263] = 32'b11111111111111110110010000010100;
assign LUT_2[19264] = 32'b11111111111111111000011000101010;
assign LUT_2[19265] = 32'b11111111111111110101010001000011;
assign LUT_2[19266] = 32'b11111111111111111111010001100110;
assign LUT_2[19267] = 32'b11111111111111111100001001111111;
assign LUT_2[19268] = 32'b11111111111111110100110110010010;
assign LUT_2[19269] = 32'b11111111111111110001101110101011;
assign LUT_2[19270] = 32'b11111111111111111011101111001110;
assign LUT_2[19271] = 32'b11111111111111111000100111100111;
assign LUT_2[19272] = 32'b11111111111111110011001010000111;
assign LUT_2[19273] = 32'b11111111111111110000000010100000;
assign LUT_2[19274] = 32'b11111111111111111010000011000011;
assign LUT_2[19275] = 32'b11111111111111110110111011011100;
assign LUT_2[19276] = 32'b11111111111111101111100111101111;
assign LUT_2[19277] = 32'b11111111111111101100100000001000;
assign LUT_2[19278] = 32'b11111111111111110110100000101011;
assign LUT_2[19279] = 32'b11111111111111110011011001000100;
assign LUT_2[19280] = 32'b11111111111111110010111100110100;
assign LUT_2[19281] = 32'b11111111111111101111110101001101;
assign LUT_2[19282] = 32'b11111111111111111001110101110000;
assign LUT_2[19283] = 32'b11111111111111110110101110001001;
assign LUT_2[19284] = 32'b11111111111111101111011010011100;
assign LUT_2[19285] = 32'b11111111111111101100010010110101;
assign LUT_2[19286] = 32'b11111111111111110110010011011000;
assign LUT_2[19287] = 32'b11111111111111110011001011110001;
assign LUT_2[19288] = 32'b11111111111111101101101110010001;
assign LUT_2[19289] = 32'b11111111111111101010100110101010;
assign LUT_2[19290] = 32'b11111111111111110100100111001101;
assign LUT_2[19291] = 32'b11111111111111110001011111100110;
assign LUT_2[19292] = 32'b11111111111111101010001011111001;
assign LUT_2[19293] = 32'b11111111111111100111000100010010;
assign LUT_2[19294] = 32'b11111111111111110001000100110101;
assign LUT_2[19295] = 32'b11111111111111101101111101001110;
assign LUT_2[19296] = 32'b11111111111111111000110100010011;
assign LUT_2[19297] = 32'b11111111111111110101101100101100;
assign LUT_2[19298] = 32'b11111111111111111111101101001111;
assign LUT_2[19299] = 32'b11111111111111111100100101101000;
assign LUT_2[19300] = 32'b11111111111111110101010001111011;
assign LUT_2[19301] = 32'b11111111111111110010001010010100;
assign LUT_2[19302] = 32'b11111111111111111100001010110111;
assign LUT_2[19303] = 32'b11111111111111111001000011010000;
assign LUT_2[19304] = 32'b11111111111111110011100101110000;
assign LUT_2[19305] = 32'b11111111111111110000011110001001;
assign LUT_2[19306] = 32'b11111111111111111010011110101100;
assign LUT_2[19307] = 32'b11111111111111110111010111000101;
assign LUT_2[19308] = 32'b11111111111111110000000011011000;
assign LUT_2[19309] = 32'b11111111111111101100111011110001;
assign LUT_2[19310] = 32'b11111111111111110110111100010100;
assign LUT_2[19311] = 32'b11111111111111110011110100101101;
assign LUT_2[19312] = 32'b11111111111111110011011000011101;
assign LUT_2[19313] = 32'b11111111111111110000010000110110;
assign LUT_2[19314] = 32'b11111111111111111010010001011001;
assign LUT_2[19315] = 32'b11111111111111110111001001110010;
assign LUT_2[19316] = 32'b11111111111111101111110110000101;
assign LUT_2[19317] = 32'b11111111111111101100101110011110;
assign LUT_2[19318] = 32'b11111111111111110110101111000001;
assign LUT_2[19319] = 32'b11111111111111110011100111011010;
assign LUT_2[19320] = 32'b11111111111111101110001001111010;
assign LUT_2[19321] = 32'b11111111111111101011000010010011;
assign LUT_2[19322] = 32'b11111111111111110101000010110110;
assign LUT_2[19323] = 32'b11111111111111110001111011001111;
assign LUT_2[19324] = 32'b11111111111111101010100111100010;
assign LUT_2[19325] = 32'b11111111111111100111011111111011;
assign LUT_2[19326] = 32'b11111111111111110001100000011110;
assign LUT_2[19327] = 32'b11111111111111101110011000110111;
assign LUT_2[19328] = 32'b00000000000000000100100100010110;
assign LUT_2[19329] = 32'b00000000000000000001011100101111;
assign LUT_2[19330] = 32'b00000000000000001011011101010010;
assign LUT_2[19331] = 32'b00000000000000001000010101101011;
assign LUT_2[19332] = 32'b00000000000000000001000001111110;
assign LUT_2[19333] = 32'b11111111111111111101111010010111;
assign LUT_2[19334] = 32'b00000000000000000111111010111010;
assign LUT_2[19335] = 32'b00000000000000000100110011010011;
assign LUT_2[19336] = 32'b11111111111111111111010101110011;
assign LUT_2[19337] = 32'b11111111111111111100001110001100;
assign LUT_2[19338] = 32'b00000000000000000110001110101111;
assign LUT_2[19339] = 32'b00000000000000000011000111001000;
assign LUT_2[19340] = 32'b11111111111111111011110011011011;
assign LUT_2[19341] = 32'b11111111111111111000101011110100;
assign LUT_2[19342] = 32'b00000000000000000010101100010111;
assign LUT_2[19343] = 32'b11111111111111111111100100110000;
assign LUT_2[19344] = 32'b11111111111111111111001000100000;
assign LUT_2[19345] = 32'b11111111111111111100000000111001;
assign LUT_2[19346] = 32'b00000000000000000110000001011100;
assign LUT_2[19347] = 32'b00000000000000000010111001110101;
assign LUT_2[19348] = 32'b11111111111111111011100110001000;
assign LUT_2[19349] = 32'b11111111111111111000011110100001;
assign LUT_2[19350] = 32'b00000000000000000010011111000100;
assign LUT_2[19351] = 32'b11111111111111111111010111011101;
assign LUT_2[19352] = 32'b11111111111111111001111001111101;
assign LUT_2[19353] = 32'b11111111111111110110110010010110;
assign LUT_2[19354] = 32'b00000000000000000000110010111001;
assign LUT_2[19355] = 32'b11111111111111111101101011010010;
assign LUT_2[19356] = 32'b11111111111111110110010111100101;
assign LUT_2[19357] = 32'b11111111111111110011001111111110;
assign LUT_2[19358] = 32'b11111111111111111101010000100001;
assign LUT_2[19359] = 32'b11111111111111111010001000111010;
assign LUT_2[19360] = 32'b00000000000000000100111111111111;
assign LUT_2[19361] = 32'b00000000000000000001111000011000;
assign LUT_2[19362] = 32'b00000000000000001011111000111011;
assign LUT_2[19363] = 32'b00000000000000001000110001010100;
assign LUT_2[19364] = 32'b00000000000000000001011101100111;
assign LUT_2[19365] = 32'b11111111111111111110010110000000;
assign LUT_2[19366] = 32'b00000000000000001000010110100011;
assign LUT_2[19367] = 32'b00000000000000000101001110111100;
assign LUT_2[19368] = 32'b11111111111111111111110001011100;
assign LUT_2[19369] = 32'b11111111111111111100101001110101;
assign LUT_2[19370] = 32'b00000000000000000110101010011000;
assign LUT_2[19371] = 32'b00000000000000000011100010110001;
assign LUT_2[19372] = 32'b11111111111111111100001111000100;
assign LUT_2[19373] = 32'b11111111111111111001000111011101;
assign LUT_2[19374] = 32'b00000000000000000011001000000000;
assign LUT_2[19375] = 32'b00000000000000000000000000011001;
assign LUT_2[19376] = 32'b11111111111111111111100100001001;
assign LUT_2[19377] = 32'b11111111111111111100011100100010;
assign LUT_2[19378] = 32'b00000000000000000110011101000101;
assign LUT_2[19379] = 32'b00000000000000000011010101011110;
assign LUT_2[19380] = 32'b11111111111111111100000001110001;
assign LUT_2[19381] = 32'b11111111111111111000111010001010;
assign LUT_2[19382] = 32'b00000000000000000010111010101101;
assign LUT_2[19383] = 32'b11111111111111111111110011000110;
assign LUT_2[19384] = 32'b11111111111111111010010101100110;
assign LUT_2[19385] = 32'b11111111111111110111001101111111;
assign LUT_2[19386] = 32'b00000000000000000001001110100010;
assign LUT_2[19387] = 32'b11111111111111111110000110111011;
assign LUT_2[19388] = 32'b11111111111111110110110011001110;
assign LUT_2[19389] = 32'b11111111111111110011101011100111;
assign LUT_2[19390] = 32'b11111111111111111101101100001010;
assign LUT_2[19391] = 32'b11111111111111111010100100100011;
assign LUT_2[19392] = 32'b11111111111111111100101100111001;
assign LUT_2[19393] = 32'b11111111111111111001100101010010;
assign LUT_2[19394] = 32'b00000000000000000011100101110101;
assign LUT_2[19395] = 32'b00000000000000000000011110001110;
assign LUT_2[19396] = 32'b11111111111111111001001010100001;
assign LUT_2[19397] = 32'b11111111111111110110000010111010;
assign LUT_2[19398] = 32'b00000000000000000000000011011101;
assign LUT_2[19399] = 32'b11111111111111111100111011110110;
assign LUT_2[19400] = 32'b11111111111111110111011110010110;
assign LUT_2[19401] = 32'b11111111111111110100010110101111;
assign LUT_2[19402] = 32'b11111111111111111110010111010010;
assign LUT_2[19403] = 32'b11111111111111111011001111101011;
assign LUT_2[19404] = 32'b11111111111111110011111011111110;
assign LUT_2[19405] = 32'b11111111111111110000110100010111;
assign LUT_2[19406] = 32'b11111111111111111010110100111010;
assign LUT_2[19407] = 32'b11111111111111110111101101010011;
assign LUT_2[19408] = 32'b11111111111111110111010001000011;
assign LUT_2[19409] = 32'b11111111111111110100001001011100;
assign LUT_2[19410] = 32'b11111111111111111110001001111111;
assign LUT_2[19411] = 32'b11111111111111111011000010011000;
assign LUT_2[19412] = 32'b11111111111111110011101110101011;
assign LUT_2[19413] = 32'b11111111111111110000100111000100;
assign LUT_2[19414] = 32'b11111111111111111010100111100111;
assign LUT_2[19415] = 32'b11111111111111110111100000000000;
assign LUT_2[19416] = 32'b11111111111111110010000010100000;
assign LUT_2[19417] = 32'b11111111111111101110111010111001;
assign LUT_2[19418] = 32'b11111111111111111000111011011100;
assign LUT_2[19419] = 32'b11111111111111110101110011110101;
assign LUT_2[19420] = 32'b11111111111111101110100000001000;
assign LUT_2[19421] = 32'b11111111111111101011011000100001;
assign LUT_2[19422] = 32'b11111111111111110101011001000100;
assign LUT_2[19423] = 32'b11111111111111110010010001011101;
assign LUT_2[19424] = 32'b11111111111111111101001000100010;
assign LUT_2[19425] = 32'b11111111111111111010000000111011;
assign LUT_2[19426] = 32'b00000000000000000100000001011110;
assign LUT_2[19427] = 32'b00000000000000000000111001110111;
assign LUT_2[19428] = 32'b11111111111111111001100110001010;
assign LUT_2[19429] = 32'b11111111111111110110011110100011;
assign LUT_2[19430] = 32'b00000000000000000000011111000110;
assign LUT_2[19431] = 32'b11111111111111111101010111011111;
assign LUT_2[19432] = 32'b11111111111111110111111001111111;
assign LUT_2[19433] = 32'b11111111111111110100110010011000;
assign LUT_2[19434] = 32'b11111111111111111110110010111011;
assign LUT_2[19435] = 32'b11111111111111111011101011010100;
assign LUT_2[19436] = 32'b11111111111111110100010111100111;
assign LUT_2[19437] = 32'b11111111111111110001010000000000;
assign LUT_2[19438] = 32'b11111111111111111011010000100011;
assign LUT_2[19439] = 32'b11111111111111111000001000111100;
assign LUT_2[19440] = 32'b11111111111111110111101100101100;
assign LUT_2[19441] = 32'b11111111111111110100100101000101;
assign LUT_2[19442] = 32'b11111111111111111110100101101000;
assign LUT_2[19443] = 32'b11111111111111111011011110000001;
assign LUT_2[19444] = 32'b11111111111111110100001010010100;
assign LUT_2[19445] = 32'b11111111111111110001000010101101;
assign LUT_2[19446] = 32'b11111111111111111011000011010000;
assign LUT_2[19447] = 32'b11111111111111110111111011101001;
assign LUT_2[19448] = 32'b11111111111111110010011110001001;
assign LUT_2[19449] = 32'b11111111111111101111010110100010;
assign LUT_2[19450] = 32'b11111111111111111001010111000101;
assign LUT_2[19451] = 32'b11111111111111110110001111011110;
assign LUT_2[19452] = 32'b11111111111111101110111011110001;
assign LUT_2[19453] = 32'b11111111111111101011110100001010;
assign LUT_2[19454] = 32'b11111111111111110101110100101101;
assign LUT_2[19455] = 32'b11111111111111110010101101000110;
assign LUT_2[19456] = 32'b11111111111111111110001011110100;
assign LUT_2[19457] = 32'b11111111111111111011000100001101;
assign LUT_2[19458] = 32'b00000000000000000101000100110000;
assign LUT_2[19459] = 32'b00000000000000000001111101001001;
assign LUT_2[19460] = 32'b11111111111111111010101001011100;
assign LUT_2[19461] = 32'b11111111111111110111100001110101;
assign LUT_2[19462] = 32'b00000000000000000001100010011000;
assign LUT_2[19463] = 32'b11111111111111111110011010110001;
assign LUT_2[19464] = 32'b11111111111111111000111101010001;
assign LUT_2[19465] = 32'b11111111111111110101110101101010;
assign LUT_2[19466] = 32'b11111111111111111111110110001101;
assign LUT_2[19467] = 32'b11111111111111111100101110100110;
assign LUT_2[19468] = 32'b11111111111111110101011010111001;
assign LUT_2[19469] = 32'b11111111111111110010010011010010;
assign LUT_2[19470] = 32'b11111111111111111100010011110101;
assign LUT_2[19471] = 32'b11111111111111111001001100001110;
assign LUT_2[19472] = 32'b11111111111111111000101111111110;
assign LUT_2[19473] = 32'b11111111111111110101101000010111;
assign LUT_2[19474] = 32'b11111111111111111111101000111010;
assign LUT_2[19475] = 32'b11111111111111111100100001010011;
assign LUT_2[19476] = 32'b11111111111111110101001101100110;
assign LUT_2[19477] = 32'b11111111111111110010000101111111;
assign LUT_2[19478] = 32'b11111111111111111100000110100010;
assign LUT_2[19479] = 32'b11111111111111111000111110111011;
assign LUT_2[19480] = 32'b11111111111111110011100001011011;
assign LUT_2[19481] = 32'b11111111111111110000011001110100;
assign LUT_2[19482] = 32'b11111111111111111010011010010111;
assign LUT_2[19483] = 32'b11111111111111110111010010110000;
assign LUT_2[19484] = 32'b11111111111111101111111111000011;
assign LUT_2[19485] = 32'b11111111111111101100110111011100;
assign LUT_2[19486] = 32'b11111111111111110110110111111111;
assign LUT_2[19487] = 32'b11111111111111110011110000011000;
assign LUT_2[19488] = 32'b11111111111111111110100111011101;
assign LUT_2[19489] = 32'b11111111111111111011011111110110;
assign LUT_2[19490] = 32'b00000000000000000101100000011001;
assign LUT_2[19491] = 32'b00000000000000000010011000110010;
assign LUT_2[19492] = 32'b11111111111111111011000101000101;
assign LUT_2[19493] = 32'b11111111111111110111111101011110;
assign LUT_2[19494] = 32'b00000000000000000001111110000001;
assign LUT_2[19495] = 32'b11111111111111111110110110011010;
assign LUT_2[19496] = 32'b11111111111111111001011000111010;
assign LUT_2[19497] = 32'b11111111111111110110010001010011;
assign LUT_2[19498] = 32'b00000000000000000000010001110110;
assign LUT_2[19499] = 32'b11111111111111111101001010001111;
assign LUT_2[19500] = 32'b11111111111111110101110110100010;
assign LUT_2[19501] = 32'b11111111111111110010101110111011;
assign LUT_2[19502] = 32'b11111111111111111100101111011110;
assign LUT_2[19503] = 32'b11111111111111111001100111110111;
assign LUT_2[19504] = 32'b11111111111111111001001011100111;
assign LUT_2[19505] = 32'b11111111111111110110000100000000;
assign LUT_2[19506] = 32'b00000000000000000000000100100011;
assign LUT_2[19507] = 32'b11111111111111111100111100111100;
assign LUT_2[19508] = 32'b11111111111111110101101001001111;
assign LUT_2[19509] = 32'b11111111111111110010100001101000;
assign LUT_2[19510] = 32'b11111111111111111100100010001011;
assign LUT_2[19511] = 32'b11111111111111111001011010100100;
assign LUT_2[19512] = 32'b11111111111111110011111101000100;
assign LUT_2[19513] = 32'b11111111111111110000110101011101;
assign LUT_2[19514] = 32'b11111111111111111010110110000000;
assign LUT_2[19515] = 32'b11111111111111110111101110011001;
assign LUT_2[19516] = 32'b11111111111111110000011010101100;
assign LUT_2[19517] = 32'b11111111111111101101010011000101;
assign LUT_2[19518] = 32'b11111111111111110111010011101000;
assign LUT_2[19519] = 32'b11111111111111110100001100000001;
assign LUT_2[19520] = 32'b11111111111111110110010100010111;
assign LUT_2[19521] = 32'b11111111111111110011001100110000;
assign LUT_2[19522] = 32'b11111111111111111101001101010011;
assign LUT_2[19523] = 32'b11111111111111111010000101101100;
assign LUT_2[19524] = 32'b11111111111111110010110001111111;
assign LUT_2[19525] = 32'b11111111111111101111101010011000;
assign LUT_2[19526] = 32'b11111111111111111001101010111011;
assign LUT_2[19527] = 32'b11111111111111110110100011010100;
assign LUT_2[19528] = 32'b11111111111111110001000101110100;
assign LUT_2[19529] = 32'b11111111111111101101111110001101;
assign LUT_2[19530] = 32'b11111111111111110111111110110000;
assign LUT_2[19531] = 32'b11111111111111110100110111001001;
assign LUT_2[19532] = 32'b11111111111111101101100011011100;
assign LUT_2[19533] = 32'b11111111111111101010011011110101;
assign LUT_2[19534] = 32'b11111111111111110100011100011000;
assign LUT_2[19535] = 32'b11111111111111110001010100110001;
assign LUT_2[19536] = 32'b11111111111111110000111000100001;
assign LUT_2[19537] = 32'b11111111111111101101110000111010;
assign LUT_2[19538] = 32'b11111111111111110111110001011101;
assign LUT_2[19539] = 32'b11111111111111110100101001110110;
assign LUT_2[19540] = 32'b11111111111111101101010110001001;
assign LUT_2[19541] = 32'b11111111111111101010001110100010;
assign LUT_2[19542] = 32'b11111111111111110100001111000101;
assign LUT_2[19543] = 32'b11111111111111110001000111011110;
assign LUT_2[19544] = 32'b11111111111111101011101001111110;
assign LUT_2[19545] = 32'b11111111111111101000100010010111;
assign LUT_2[19546] = 32'b11111111111111110010100010111010;
assign LUT_2[19547] = 32'b11111111111111101111011011010011;
assign LUT_2[19548] = 32'b11111111111111101000000111100110;
assign LUT_2[19549] = 32'b11111111111111100100111111111111;
assign LUT_2[19550] = 32'b11111111111111101111000000100010;
assign LUT_2[19551] = 32'b11111111111111101011111000111011;
assign LUT_2[19552] = 32'b11111111111111110110110000000000;
assign LUT_2[19553] = 32'b11111111111111110011101000011001;
assign LUT_2[19554] = 32'b11111111111111111101101000111100;
assign LUT_2[19555] = 32'b11111111111111111010100001010101;
assign LUT_2[19556] = 32'b11111111111111110011001101101000;
assign LUT_2[19557] = 32'b11111111111111110000000110000001;
assign LUT_2[19558] = 32'b11111111111111111010000110100100;
assign LUT_2[19559] = 32'b11111111111111110110111110111101;
assign LUT_2[19560] = 32'b11111111111111110001100001011101;
assign LUT_2[19561] = 32'b11111111111111101110011001110110;
assign LUT_2[19562] = 32'b11111111111111111000011010011001;
assign LUT_2[19563] = 32'b11111111111111110101010010110010;
assign LUT_2[19564] = 32'b11111111111111101101111111000101;
assign LUT_2[19565] = 32'b11111111111111101010110111011110;
assign LUT_2[19566] = 32'b11111111111111110100111000000001;
assign LUT_2[19567] = 32'b11111111111111110001110000011010;
assign LUT_2[19568] = 32'b11111111111111110001010100001010;
assign LUT_2[19569] = 32'b11111111111111101110001100100011;
assign LUT_2[19570] = 32'b11111111111111111000001101000110;
assign LUT_2[19571] = 32'b11111111111111110101000101011111;
assign LUT_2[19572] = 32'b11111111111111101101110001110010;
assign LUT_2[19573] = 32'b11111111111111101010101010001011;
assign LUT_2[19574] = 32'b11111111111111110100101010101110;
assign LUT_2[19575] = 32'b11111111111111110001100011000111;
assign LUT_2[19576] = 32'b11111111111111101100000101100111;
assign LUT_2[19577] = 32'b11111111111111101000111110000000;
assign LUT_2[19578] = 32'b11111111111111110010111110100011;
assign LUT_2[19579] = 32'b11111111111111101111110110111100;
assign LUT_2[19580] = 32'b11111111111111101000100011001111;
assign LUT_2[19581] = 32'b11111111111111100101011011101000;
assign LUT_2[19582] = 32'b11111111111111101111011100001011;
assign LUT_2[19583] = 32'b11111111111111101100010100100100;
assign LUT_2[19584] = 32'b00000000000000000010100000000011;
assign LUT_2[19585] = 32'b11111111111111111111011000011100;
assign LUT_2[19586] = 32'b00000000000000001001011000111111;
assign LUT_2[19587] = 32'b00000000000000000110010001011000;
assign LUT_2[19588] = 32'b11111111111111111110111101101011;
assign LUT_2[19589] = 32'b11111111111111111011110110000100;
assign LUT_2[19590] = 32'b00000000000000000101110110100111;
assign LUT_2[19591] = 32'b00000000000000000010101111000000;
assign LUT_2[19592] = 32'b11111111111111111101010001100000;
assign LUT_2[19593] = 32'b11111111111111111010001001111001;
assign LUT_2[19594] = 32'b00000000000000000100001010011100;
assign LUT_2[19595] = 32'b00000000000000000001000010110101;
assign LUT_2[19596] = 32'b11111111111111111001101111001000;
assign LUT_2[19597] = 32'b11111111111111110110100111100001;
assign LUT_2[19598] = 32'b00000000000000000000101000000100;
assign LUT_2[19599] = 32'b11111111111111111101100000011101;
assign LUT_2[19600] = 32'b11111111111111111101000100001101;
assign LUT_2[19601] = 32'b11111111111111111001111100100110;
assign LUT_2[19602] = 32'b00000000000000000011111101001001;
assign LUT_2[19603] = 32'b00000000000000000000110101100010;
assign LUT_2[19604] = 32'b11111111111111111001100001110101;
assign LUT_2[19605] = 32'b11111111111111110110011010001110;
assign LUT_2[19606] = 32'b00000000000000000000011010110001;
assign LUT_2[19607] = 32'b11111111111111111101010011001010;
assign LUT_2[19608] = 32'b11111111111111110111110101101010;
assign LUT_2[19609] = 32'b11111111111111110100101110000011;
assign LUT_2[19610] = 32'b11111111111111111110101110100110;
assign LUT_2[19611] = 32'b11111111111111111011100110111111;
assign LUT_2[19612] = 32'b11111111111111110100010011010010;
assign LUT_2[19613] = 32'b11111111111111110001001011101011;
assign LUT_2[19614] = 32'b11111111111111111011001100001110;
assign LUT_2[19615] = 32'b11111111111111111000000100100111;
assign LUT_2[19616] = 32'b00000000000000000010111011101100;
assign LUT_2[19617] = 32'b11111111111111111111110100000101;
assign LUT_2[19618] = 32'b00000000000000001001110100101000;
assign LUT_2[19619] = 32'b00000000000000000110101101000001;
assign LUT_2[19620] = 32'b11111111111111111111011001010100;
assign LUT_2[19621] = 32'b11111111111111111100010001101101;
assign LUT_2[19622] = 32'b00000000000000000110010010010000;
assign LUT_2[19623] = 32'b00000000000000000011001010101001;
assign LUT_2[19624] = 32'b11111111111111111101101101001001;
assign LUT_2[19625] = 32'b11111111111111111010100101100010;
assign LUT_2[19626] = 32'b00000000000000000100100110000101;
assign LUT_2[19627] = 32'b00000000000000000001011110011110;
assign LUT_2[19628] = 32'b11111111111111111010001010110001;
assign LUT_2[19629] = 32'b11111111111111110111000011001010;
assign LUT_2[19630] = 32'b00000000000000000001000011101101;
assign LUT_2[19631] = 32'b11111111111111111101111100000110;
assign LUT_2[19632] = 32'b11111111111111111101011111110110;
assign LUT_2[19633] = 32'b11111111111111111010011000001111;
assign LUT_2[19634] = 32'b00000000000000000100011000110010;
assign LUT_2[19635] = 32'b00000000000000000001010001001011;
assign LUT_2[19636] = 32'b11111111111111111001111101011110;
assign LUT_2[19637] = 32'b11111111111111110110110101110111;
assign LUT_2[19638] = 32'b00000000000000000000110110011010;
assign LUT_2[19639] = 32'b11111111111111111101101110110011;
assign LUT_2[19640] = 32'b11111111111111111000010001010011;
assign LUT_2[19641] = 32'b11111111111111110101001001101100;
assign LUT_2[19642] = 32'b11111111111111111111001010001111;
assign LUT_2[19643] = 32'b11111111111111111100000010101000;
assign LUT_2[19644] = 32'b11111111111111110100101110111011;
assign LUT_2[19645] = 32'b11111111111111110001100111010100;
assign LUT_2[19646] = 32'b11111111111111111011100111110111;
assign LUT_2[19647] = 32'b11111111111111111000100000010000;
assign LUT_2[19648] = 32'b11111111111111111010101000100110;
assign LUT_2[19649] = 32'b11111111111111110111100000111111;
assign LUT_2[19650] = 32'b00000000000000000001100001100010;
assign LUT_2[19651] = 32'b11111111111111111110011001111011;
assign LUT_2[19652] = 32'b11111111111111110111000110001110;
assign LUT_2[19653] = 32'b11111111111111110011111110100111;
assign LUT_2[19654] = 32'b11111111111111111101111111001010;
assign LUT_2[19655] = 32'b11111111111111111010110111100011;
assign LUT_2[19656] = 32'b11111111111111110101011010000011;
assign LUT_2[19657] = 32'b11111111111111110010010010011100;
assign LUT_2[19658] = 32'b11111111111111111100010010111111;
assign LUT_2[19659] = 32'b11111111111111111001001011011000;
assign LUT_2[19660] = 32'b11111111111111110001110111101011;
assign LUT_2[19661] = 32'b11111111111111101110110000000100;
assign LUT_2[19662] = 32'b11111111111111111000110000100111;
assign LUT_2[19663] = 32'b11111111111111110101101001000000;
assign LUT_2[19664] = 32'b11111111111111110101001100110000;
assign LUT_2[19665] = 32'b11111111111111110010000101001001;
assign LUT_2[19666] = 32'b11111111111111111100000101101100;
assign LUT_2[19667] = 32'b11111111111111111000111110000101;
assign LUT_2[19668] = 32'b11111111111111110001101010011000;
assign LUT_2[19669] = 32'b11111111111111101110100010110001;
assign LUT_2[19670] = 32'b11111111111111111000100011010100;
assign LUT_2[19671] = 32'b11111111111111110101011011101101;
assign LUT_2[19672] = 32'b11111111111111101111111110001101;
assign LUT_2[19673] = 32'b11111111111111101100110110100110;
assign LUT_2[19674] = 32'b11111111111111110110110111001001;
assign LUT_2[19675] = 32'b11111111111111110011101111100010;
assign LUT_2[19676] = 32'b11111111111111101100011011110101;
assign LUT_2[19677] = 32'b11111111111111101001010100001110;
assign LUT_2[19678] = 32'b11111111111111110011010100110001;
assign LUT_2[19679] = 32'b11111111111111110000001101001010;
assign LUT_2[19680] = 32'b11111111111111111011000100001111;
assign LUT_2[19681] = 32'b11111111111111110111111100101000;
assign LUT_2[19682] = 32'b00000000000000000001111101001011;
assign LUT_2[19683] = 32'b11111111111111111110110101100100;
assign LUT_2[19684] = 32'b11111111111111110111100001110111;
assign LUT_2[19685] = 32'b11111111111111110100011010010000;
assign LUT_2[19686] = 32'b11111111111111111110011010110011;
assign LUT_2[19687] = 32'b11111111111111111011010011001100;
assign LUT_2[19688] = 32'b11111111111111110101110101101100;
assign LUT_2[19689] = 32'b11111111111111110010101110000101;
assign LUT_2[19690] = 32'b11111111111111111100101110101000;
assign LUT_2[19691] = 32'b11111111111111111001100111000001;
assign LUT_2[19692] = 32'b11111111111111110010010011010100;
assign LUT_2[19693] = 32'b11111111111111101111001011101101;
assign LUT_2[19694] = 32'b11111111111111111001001100010000;
assign LUT_2[19695] = 32'b11111111111111110110000100101001;
assign LUT_2[19696] = 32'b11111111111111110101101000011001;
assign LUT_2[19697] = 32'b11111111111111110010100000110010;
assign LUT_2[19698] = 32'b11111111111111111100100001010101;
assign LUT_2[19699] = 32'b11111111111111111001011001101110;
assign LUT_2[19700] = 32'b11111111111111110010000110000001;
assign LUT_2[19701] = 32'b11111111111111101110111110011010;
assign LUT_2[19702] = 32'b11111111111111111000111110111101;
assign LUT_2[19703] = 32'b11111111111111110101110111010110;
assign LUT_2[19704] = 32'b11111111111111110000011001110110;
assign LUT_2[19705] = 32'b11111111111111101101010010001111;
assign LUT_2[19706] = 32'b11111111111111110111010010110010;
assign LUT_2[19707] = 32'b11111111111111110100001011001011;
assign LUT_2[19708] = 32'b11111111111111101100110111011110;
assign LUT_2[19709] = 32'b11111111111111101001101111110111;
assign LUT_2[19710] = 32'b11111111111111110011110000011010;
assign LUT_2[19711] = 32'b11111111111111110000101000110011;
assign LUT_2[19712] = 32'b00000000000000000010001010011010;
assign LUT_2[19713] = 32'b11111111111111111111000010110011;
assign LUT_2[19714] = 32'b00000000000000001001000011010110;
assign LUT_2[19715] = 32'b00000000000000000101111011101111;
assign LUT_2[19716] = 32'b11111111111111111110101000000010;
assign LUT_2[19717] = 32'b11111111111111111011100000011011;
assign LUT_2[19718] = 32'b00000000000000000101100000111110;
assign LUT_2[19719] = 32'b00000000000000000010011001010111;
assign LUT_2[19720] = 32'b11111111111111111100111011110111;
assign LUT_2[19721] = 32'b11111111111111111001110100010000;
assign LUT_2[19722] = 32'b00000000000000000011110100110011;
assign LUT_2[19723] = 32'b00000000000000000000101101001100;
assign LUT_2[19724] = 32'b11111111111111111001011001011111;
assign LUT_2[19725] = 32'b11111111111111110110010001111000;
assign LUT_2[19726] = 32'b00000000000000000000010010011011;
assign LUT_2[19727] = 32'b11111111111111111101001010110100;
assign LUT_2[19728] = 32'b11111111111111111100101110100100;
assign LUT_2[19729] = 32'b11111111111111111001100110111101;
assign LUT_2[19730] = 32'b00000000000000000011100111100000;
assign LUT_2[19731] = 32'b00000000000000000000011111111001;
assign LUT_2[19732] = 32'b11111111111111111001001100001100;
assign LUT_2[19733] = 32'b11111111111111110110000100100101;
assign LUT_2[19734] = 32'b00000000000000000000000101001000;
assign LUT_2[19735] = 32'b11111111111111111100111101100001;
assign LUT_2[19736] = 32'b11111111111111110111100000000001;
assign LUT_2[19737] = 32'b11111111111111110100011000011010;
assign LUT_2[19738] = 32'b11111111111111111110011000111101;
assign LUT_2[19739] = 32'b11111111111111111011010001010110;
assign LUT_2[19740] = 32'b11111111111111110011111101101001;
assign LUT_2[19741] = 32'b11111111111111110000110110000010;
assign LUT_2[19742] = 32'b11111111111111111010110110100101;
assign LUT_2[19743] = 32'b11111111111111110111101110111110;
assign LUT_2[19744] = 32'b00000000000000000010100110000011;
assign LUT_2[19745] = 32'b11111111111111111111011110011100;
assign LUT_2[19746] = 32'b00000000000000001001011110111111;
assign LUT_2[19747] = 32'b00000000000000000110010111011000;
assign LUT_2[19748] = 32'b11111111111111111111000011101011;
assign LUT_2[19749] = 32'b11111111111111111011111100000100;
assign LUT_2[19750] = 32'b00000000000000000101111100100111;
assign LUT_2[19751] = 32'b00000000000000000010110101000000;
assign LUT_2[19752] = 32'b11111111111111111101010111100000;
assign LUT_2[19753] = 32'b11111111111111111010001111111001;
assign LUT_2[19754] = 32'b00000000000000000100010000011100;
assign LUT_2[19755] = 32'b00000000000000000001001000110101;
assign LUT_2[19756] = 32'b11111111111111111001110101001000;
assign LUT_2[19757] = 32'b11111111111111110110101101100001;
assign LUT_2[19758] = 32'b00000000000000000000101110000100;
assign LUT_2[19759] = 32'b11111111111111111101100110011101;
assign LUT_2[19760] = 32'b11111111111111111101001010001101;
assign LUT_2[19761] = 32'b11111111111111111010000010100110;
assign LUT_2[19762] = 32'b00000000000000000100000011001001;
assign LUT_2[19763] = 32'b00000000000000000000111011100010;
assign LUT_2[19764] = 32'b11111111111111111001100111110101;
assign LUT_2[19765] = 32'b11111111111111110110100000001110;
assign LUT_2[19766] = 32'b00000000000000000000100000110001;
assign LUT_2[19767] = 32'b11111111111111111101011001001010;
assign LUT_2[19768] = 32'b11111111111111110111111011101010;
assign LUT_2[19769] = 32'b11111111111111110100110100000011;
assign LUT_2[19770] = 32'b11111111111111111110110100100110;
assign LUT_2[19771] = 32'b11111111111111111011101100111111;
assign LUT_2[19772] = 32'b11111111111111110100011001010010;
assign LUT_2[19773] = 32'b11111111111111110001010001101011;
assign LUT_2[19774] = 32'b11111111111111111011010010001110;
assign LUT_2[19775] = 32'b11111111111111111000001010100111;
assign LUT_2[19776] = 32'b11111111111111111010010010111101;
assign LUT_2[19777] = 32'b11111111111111110111001011010110;
assign LUT_2[19778] = 32'b00000000000000000001001011111001;
assign LUT_2[19779] = 32'b11111111111111111110000100010010;
assign LUT_2[19780] = 32'b11111111111111110110110000100101;
assign LUT_2[19781] = 32'b11111111111111110011101000111110;
assign LUT_2[19782] = 32'b11111111111111111101101001100001;
assign LUT_2[19783] = 32'b11111111111111111010100001111010;
assign LUT_2[19784] = 32'b11111111111111110101000100011010;
assign LUT_2[19785] = 32'b11111111111111110001111100110011;
assign LUT_2[19786] = 32'b11111111111111111011111101010110;
assign LUT_2[19787] = 32'b11111111111111111000110101101111;
assign LUT_2[19788] = 32'b11111111111111110001100010000010;
assign LUT_2[19789] = 32'b11111111111111101110011010011011;
assign LUT_2[19790] = 32'b11111111111111111000011010111110;
assign LUT_2[19791] = 32'b11111111111111110101010011010111;
assign LUT_2[19792] = 32'b11111111111111110100110111000111;
assign LUT_2[19793] = 32'b11111111111111110001101111100000;
assign LUT_2[19794] = 32'b11111111111111111011110000000011;
assign LUT_2[19795] = 32'b11111111111111111000101000011100;
assign LUT_2[19796] = 32'b11111111111111110001010100101111;
assign LUT_2[19797] = 32'b11111111111111101110001101001000;
assign LUT_2[19798] = 32'b11111111111111111000001101101011;
assign LUT_2[19799] = 32'b11111111111111110101000110000100;
assign LUT_2[19800] = 32'b11111111111111101111101000100100;
assign LUT_2[19801] = 32'b11111111111111101100100000111101;
assign LUT_2[19802] = 32'b11111111111111110110100001100000;
assign LUT_2[19803] = 32'b11111111111111110011011001111001;
assign LUT_2[19804] = 32'b11111111111111101100000110001100;
assign LUT_2[19805] = 32'b11111111111111101000111110100101;
assign LUT_2[19806] = 32'b11111111111111110010111111001000;
assign LUT_2[19807] = 32'b11111111111111101111110111100001;
assign LUT_2[19808] = 32'b11111111111111111010101110100110;
assign LUT_2[19809] = 32'b11111111111111110111100110111111;
assign LUT_2[19810] = 32'b00000000000000000001100111100010;
assign LUT_2[19811] = 32'b11111111111111111110011111111011;
assign LUT_2[19812] = 32'b11111111111111110111001100001110;
assign LUT_2[19813] = 32'b11111111111111110100000100100111;
assign LUT_2[19814] = 32'b11111111111111111110000101001010;
assign LUT_2[19815] = 32'b11111111111111111010111101100011;
assign LUT_2[19816] = 32'b11111111111111110101100000000011;
assign LUT_2[19817] = 32'b11111111111111110010011000011100;
assign LUT_2[19818] = 32'b11111111111111111100011000111111;
assign LUT_2[19819] = 32'b11111111111111111001010001011000;
assign LUT_2[19820] = 32'b11111111111111110001111101101011;
assign LUT_2[19821] = 32'b11111111111111101110110110000100;
assign LUT_2[19822] = 32'b11111111111111111000110110100111;
assign LUT_2[19823] = 32'b11111111111111110101101111000000;
assign LUT_2[19824] = 32'b11111111111111110101010010110000;
assign LUT_2[19825] = 32'b11111111111111110010001011001001;
assign LUT_2[19826] = 32'b11111111111111111100001011101100;
assign LUT_2[19827] = 32'b11111111111111111001000100000101;
assign LUT_2[19828] = 32'b11111111111111110001110000011000;
assign LUT_2[19829] = 32'b11111111111111101110101000110001;
assign LUT_2[19830] = 32'b11111111111111111000101001010100;
assign LUT_2[19831] = 32'b11111111111111110101100001101101;
assign LUT_2[19832] = 32'b11111111111111110000000100001101;
assign LUT_2[19833] = 32'b11111111111111101100111100100110;
assign LUT_2[19834] = 32'b11111111111111110110111101001001;
assign LUT_2[19835] = 32'b11111111111111110011110101100010;
assign LUT_2[19836] = 32'b11111111111111101100100001110101;
assign LUT_2[19837] = 32'b11111111111111101001011010001110;
assign LUT_2[19838] = 32'b11111111111111110011011010110001;
assign LUT_2[19839] = 32'b11111111111111110000010011001010;
assign LUT_2[19840] = 32'b00000000000000000110011110101001;
assign LUT_2[19841] = 32'b00000000000000000011010111000010;
assign LUT_2[19842] = 32'b00000000000000001101010111100101;
assign LUT_2[19843] = 32'b00000000000000001010001111111110;
assign LUT_2[19844] = 32'b00000000000000000010111100010001;
assign LUT_2[19845] = 32'b11111111111111111111110100101010;
assign LUT_2[19846] = 32'b00000000000000001001110101001101;
assign LUT_2[19847] = 32'b00000000000000000110101101100110;
assign LUT_2[19848] = 32'b00000000000000000001010000000110;
assign LUT_2[19849] = 32'b11111111111111111110001000011111;
assign LUT_2[19850] = 32'b00000000000000001000001001000010;
assign LUT_2[19851] = 32'b00000000000000000101000001011011;
assign LUT_2[19852] = 32'b11111111111111111101101101101110;
assign LUT_2[19853] = 32'b11111111111111111010100110000111;
assign LUT_2[19854] = 32'b00000000000000000100100110101010;
assign LUT_2[19855] = 32'b00000000000000000001011111000011;
assign LUT_2[19856] = 32'b00000000000000000001000010110011;
assign LUT_2[19857] = 32'b11111111111111111101111011001100;
assign LUT_2[19858] = 32'b00000000000000000111111011101111;
assign LUT_2[19859] = 32'b00000000000000000100110100001000;
assign LUT_2[19860] = 32'b11111111111111111101100000011011;
assign LUT_2[19861] = 32'b11111111111111111010011000110100;
assign LUT_2[19862] = 32'b00000000000000000100011001010111;
assign LUT_2[19863] = 32'b00000000000000000001010001110000;
assign LUT_2[19864] = 32'b11111111111111111011110100010000;
assign LUT_2[19865] = 32'b11111111111111111000101100101001;
assign LUT_2[19866] = 32'b00000000000000000010101101001100;
assign LUT_2[19867] = 32'b11111111111111111111100101100101;
assign LUT_2[19868] = 32'b11111111111111111000010001111000;
assign LUT_2[19869] = 32'b11111111111111110101001010010001;
assign LUT_2[19870] = 32'b11111111111111111111001010110100;
assign LUT_2[19871] = 32'b11111111111111111100000011001101;
assign LUT_2[19872] = 32'b00000000000000000110111010010010;
assign LUT_2[19873] = 32'b00000000000000000011110010101011;
assign LUT_2[19874] = 32'b00000000000000001101110011001110;
assign LUT_2[19875] = 32'b00000000000000001010101011100111;
assign LUT_2[19876] = 32'b00000000000000000011010111111010;
assign LUT_2[19877] = 32'b00000000000000000000010000010011;
assign LUT_2[19878] = 32'b00000000000000001010010000110110;
assign LUT_2[19879] = 32'b00000000000000000111001001001111;
assign LUT_2[19880] = 32'b00000000000000000001101011101111;
assign LUT_2[19881] = 32'b11111111111111111110100100001000;
assign LUT_2[19882] = 32'b00000000000000001000100100101011;
assign LUT_2[19883] = 32'b00000000000000000101011101000100;
assign LUT_2[19884] = 32'b11111111111111111110001001010111;
assign LUT_2[19885] = 32'b11111111111111111011000001110000;
assign LUT_2[19886] = 32'b00000000000000000101000010010011;
assign LUT_2[19887] = 32'b00000000000000000001111010101100;
assign LUT_2[19888] = 32'b00000000000000000001011110011100;
assign LUT_2[19889] = 32'b11111111111111111110010110110101;
assign LUT_2[19890] = 32'b00000000000000001000010111011000;
assign LUT_2[19891] = 32'b00000000000000000101001111110001;
assign LUT_2[19892] = 32'b11111111111111111101111100000100;
assign LUT_2[19893] = 32'b11111111111111111010110100011101;
assign LUT_2[19894] = 32'b00000000000000000100110101000000;
assign LUT_2[19895] = 32'b00000000000000000001101101011001;
assign LUT_2[19896] = 32'b11111111111111111100001111111001;
assign LUT_2[19897] = 32'b11111111111111111001001000010010;
assign LUT_2[19898] = 32'b00000000000000000011001000110101;
assign LUT_2[19899] = 32'b00000000000000000000000001001110;
assign LUT_2[19900] = 32'b11111111111111111000101101100001;
assign LUT_2[19901] = 32'b11111111111111110101100101111010;
assign LUT_2[19902] = 32'b11111111111111111111100110011101;
assign LUT_2[19903] = 32'b11111111111111111100011110110110;
assign LUT_2[19904] = 32'b11111111111111111110100111001100;
assign LUT_2[19905] = 32'b11111111111111111011011111100101;
assign LUT_2[19906] = 32'b00000000000000000101100000001000;
assign LUT_2[19907] = 32'b00000000000000000010011000100001;
assign LUT_2[19908] = 32'b11111111111111111011000100110100;
assign LUT_2[19909] = 32'b11111111111111110111111101001101;
assign LUT_2[19910] = 32'b00000000000000000001111101110000;
assign LUT_2[19911] = 32'b11111111111111111110110110001001;
assign LUT_2[19912] = 32'b11111111111111111001011000101001;
assign LUT_2[19913] = 32'b11111111111111110110010001000010;
assign LUT_2[19914] = 32'b00000000000000000000010001100101;
assign LUT_2[19915] = 32'b11111111111111111101001001111110;
assign LUT_2[19916] = 32'b11111111111111110101110110010001;
assign LUT_2[19917] = 32'b11111111111111110010101110101010;
assign LUT_2[19918] = 32'b11111111111111111100101111001101;
assign LUT_2[19919] = 32'b11111111111111111001100111100110;
assign LUT_2[19920] = 32'b11111111111111111001001011010110;
assign LUT_2[19921] = 32'b11111111111111110110000011101111;
assign LUT_2[19922] = 32'b00000000000000000000000100010010;
assign LUT_2[19923] = 32'b11111111111111111100111100101011;
assign LUT_2[19924] = 32'b11111111111111110101101000111110;
assign LUT_2[19925] = 32'b11111111111111110010100001010111;
assign LUT_2[19926] = 32'b11111111111111111100100001111010;
assign LUT_2[19927] = 32'b11111111111111111001011010010011;
assign LUT_2[19928] = 32'b11111111111111110011111100110011;
assign LUT_2[19929] = 32'b11111111111111110000110101001100;
assign LUT_2[19930] = 32'b11111111111111111010110101101111;
assign LUT_2[19931] = 32'b11111111111111110111101110001000;
assign LUT_2[19932] = 32'b11111111111111110000011010011011;
assign LUT_2[19933] = 32'b11111111111111101101010010110100;
assign LUT_2[19934] = 32'b11111111111111110111010011010111;
assign LUT_2[19935] = 32'b11111111111111110100001011110000;
assign LUT_2[19936] = 32'b11111111111111111111000010110101;
assign LUT_2[19937] = 32'b11111111111111111011111011001110;
assign LUT_2[19938] = 32'b00000000000000000101111011110001;
assign LUT_2[19939] = 32'b00000000000000000010110100001010;
assign LUT_2[19940] = 32'b11111111111111111011100000011101;
assign LUT_2[19941] = 32'b11111111111111111000011000110110;
assign LUT_2[19942] = 32'b00000000000000000010011001011001;
assign LUT_2[19943] = 32'b11111111111111111111010001110010;
assign LUT_2[19944] = 32'b11111111111111111001110100010010;
assign LUT_2[19945] = 32'b11111111111111110110101100101011;
assign LUT_2[19946] = 32'b00000000000000000000101101001110;
assign LUT_2[19947] = 32'b11111111111111111101100101100111;
assign LUT_2[19948] = 32'b11111111111111110110010001111010;
assign LUT_2[19949] = 32'b11111111111111110011001010010011;
assign LUT_2[19950] = 32'b11111111111111111101001010110110;
assign LUT_2[19951] = 32'b11111111111111111010000011001111;
assign LUT_2[19952] = 32'b11111111111111111001100110111111;
assign LUT_2[19953] = 32'b11111111111111110110011111011000;
assign LUT_2[19954] = 32'b00000000000000000000011111111011;
assign LUT_2[19955] = 32'b11111111111111111101011000010100;
assign LUT_2[19956] = 32'b11111111111111110110000100100111;
assign LUT_2[19957] = 32'b11111111111111110010111101000000;
assign LUT_2[19958] = 32'b11111111111111111100111101100011;
assign LUT_2[19959] = 32'b11111111111111111001110101111100;
assign LUT_2[19960] = 32'b11111111111111110100011000011100;
assign LUT_2[19961] = 32'b11111111111111110001010000110101;
assign LUT_2[19962] = 32'b11111111111111111011010001011000;
assign LUT_2[19963] = 32'b11111111111111111000001001110001;
assign LUT_2[19964] = 32'b11111111111111110000110110000100;
assign LUT_2[19965] = 32'b11111111111111101101101110011101;
assign LUT_2[19966] = 32'b11111111111111110111101111000000;
assign LUT_2[19967] = 32'b11111111111111110100100111011001;
assign LUT_2[19968] = 32'b00000000000000000010111101100110;
assign LUT_2[19969] = 32'b11111111111111111111110101111111;
assign LUT_2[19970] = 32'b00000000000000001001110110100010;
assign LUT_2[19971] = 32'b00000000000000000110101110111011;
assign LUT_2[19972] = 32'b11111111111111111111011011001110;
assign LUT_2[19973] = 32'b11111111111111111100010011100111;
assign LUT_2[19974] = 32'b00000000000000000110010100001010;
assign LUT_2[19975] = 32'b00000000000000000011001100100011;
assign LUT_2[19976] = 32'b11111111111111111101101111000011;
assign LUT_2[19977] = 32'b11111111111111111010100111011100;
assign LUT_2[19978] = 32'b00000000000000000100100111111111;
assign LUT_2[19979] = 32'b00000000000000000001100000011000;
assign LUT_2[19980] = 32'b11111111111111111010001100101011;
assign LUT_2[19981] = 32'b11111111111111110111000101000100;
assign LUT_2[19982] = 32'b00000000000000000001000101100111;
assign LUT_2[19983] = 32'b11111111111111111101111110000000;
assign LUT_2[19984] = 32'b11111111111111111101100001110000;
assign LUT_2[19985] = 32'b11111111111111111010011010001001;
assign LUT_2[19986] = 32'b00000000000000000100011010101100;
assign LUT_2[19987] = 32'b00000000000000000001010011000101;
assign LUT_2[19988] = 32'b11111111111111111001111111011000;
assign LUT_2[19989] = 32'b11111111111111110110110111110001;
assign LUT_2[19990] = 32'b00000000000000000000111000010100;
assign LUT_2[19991] = 32'b11111111111111111101110000101101;
assign LUT_2[19992] = 32'b11111111111111111000010011001101;
assign LUT_2[19993] = 32'b11111111111111110101001011100110;
assign LUT_2[19994] = 32'b11111111111111111111001100001001;
assign LUT_2[19995] = 32'b11111111111111111100000100100010;
assign LUT_2[19996] = 32'b11111111111111110100110000110101;
assign LUT_2[19997] = 32'b11111111111111110001101001001110;
assign LUT_2[19998] = 32'b11111111111111111011101001110001;
assign LUT_2[19999] = 32'b11111111111111111000100010001010;
assign LUT_2[20000] = 32'b00000000000000000011011001001111;
assign LUT_2[20001] = 32'b00000000000000000000010001101000;
assign LUT_2[20002] = 32'b00000000000000001010010010001011;
assign LUT_2[20003] = 32'b00000000000000000111001010100100;
assign LUT_2[20004] = 32'b11111111111111111111110110110111;
assign LUT_2[20005] = 32'b11111111111111111100101111010000;
assign LUT_2[20006] = 32'b00000000000000000110101111110011;
assign LUT_2[20007] = 32'b00000000000000000011101000001100;
assign LUT_2[20008] = 32'b11111111111111111110001010101100;
assign LUT_2[20009] = 32'b11111111111111111011000011000101;
assign LUT_2[20010] = 32'b00000000000000000101000011101000;
assign LUT_2[20011] = 32'b00000000000000000001111100000001;
assign LUT_2[20012] = 32'b11111111111111111010101000010100;
assign LUT_2[20013] = 32'b11111111111111110111100000101101;
assign LUT_2[20014] = 32'b00000000000000000001100001010000;
assign LUT_2[20015] = 32'b11111111111111111110011001101001;
assign LUT_2[20016] = 32'b11111111111111111101111101011001;
assign LUT_2[20017] = 32'b11111111111111111010110101110010;
assign LUT_2[20018] = 32'b00000000000000000100110110010101;
assign LUT_2[20019] = 32'b00000000000000000001101110101110;
assign LUT_2[20020] = 32'b11111111111111111010011011000001;
assign LUT_2[20021] = 32'b11111111111111110111010011011010;
assign LUT_2[20022] = 32'b00000000000000000001010011111101;
assign LUT_2[20023] = 32'b11111111111111111110001100010110;
assign LUT_2[20024] = 32'b11111111111111111000101110110110;
assign LUT_2[20025] = 32'b11111111111111110101100111001111;
assign LUT_2[20026] = 32'b11111111111111111111100111110010;
assign LUT_2[20027] = 32'b11111111111111111100100000001011;
assign LUT_2[20028] = 32'b11111111111111110101001100011110;
assign LUT_2[20029] = 32'b11111111111111110010000100110111;
assign LUT_2[20030] = 32'b11111111111111111100000101011010;
assign LUT_2[20031] = 32'b11111111111111111000111101110011;
assign LUT_2[20032] = 32'b11111111111111111011000110001001;
assign LUT_2[20033] = 32'b11111111111111110111111110100010;
assign LUT_2[20034] = 32'b00000000000000000001111111000101;
assign LUT_2[20035] = 32'b11111111111111111110110111011110;
assign LUT_2[20036] = 32'b11111111111111110111100011110001;
assign LUT_2[20037] = 32'b11111111111111110100011100001010;
assign LUT_2[20038] = 32'b11111111111111111110011100101101;
assign LUT_2[20039] = 32'b11111111111111111011010101000110;
assign LUT_2[20040] = 32'b11111111111111110101110111100110;
assign LUT_2[20041] = 32'b11111111111111110010101111111111;
assign LUT_2[20042] = 32'b11111111111111111100110000100010;
assign LUT_2[20043] = 32'b11111111111111111001101000111011;
assign LUT_2[20044] = 32'b11111111111111110010010101001110;
assign LUT_2[20045] = 32'b11111111111111101111001101100111;
assign LUT_2[20046] = 32'b11111111111111111001001110001010;
assign LUT_2[20047] = 32'b11111111111111110110000110100011;
assign LUT_2[20048] = 32'b11111111111111110101101010010011;
assign LUT_2[20049] = 32'b11111111111111110010100010101100;
assign LUT_2[20050] = 32'b11111111111111111100100011001111;
assign LUT_2[20051] = 32'b11111111111111111001011011101000;
assign LUT_2[20052] = 32'b11111111111111110010000111111011;
assign LUT_2[20053] = 32'b11111111111111101111000000010100;
assign LUT_2[20054] = 32'b11111111111111111001000000110111;
assign LUT_2[20055] = 32'b11111111111111110101111001010000;
assign LUT_2[20056] = 32'b11111111111111110000011011110000;
assign LUT_2[20057] = 32'b11111111111111101101010100001001;
assign LUT_2[20058] = 32'b11111111111111110111010100101100;
assign LUT_2[20059] = 32'b11111111111111110100001101000101;
assign LUT_2[20060] = 32'b11111111111111101100111001011000;
assign LUT_2[20061] = 32'b11111111111111101001110001110001;
assign LUT_2[20062] = 32'b11111111111111110011110010010100;
assign LUT_2[20063] = 32'b11111111111111110000101010101101;
assign LUT_2[20064] = 32'b11111111111111111011100001110010;
assign LUT_2[20065] = 32'b11111111111111111000011010001011;
assign LUT_2[20066] = 32'b00000000000000000010011010101110;
assign LUT_2[20067] = 32'b11111111111111111111010011000111;
assign LUT_2[20068] = 32'b11111111111111110111111111011010;
assign LUT_2[20069] = 32'b11111111111111110100110111110011;
assign LUT_2[20070] = 32'b11111111111111111110111000010110;
assign LUT_2[20071] = 32'b11111111111111111011110000101111;
assign LUT_2[20072] = 32'b11111111111111110110010011001111;
assign LUT_2[20073] = 32'b11111111111111110011001011101000;
assign LUT_2[20074] = 32'b11111111111111111101001100001011;
assign LUT_2[20075] = 32'b11111111111111111010000100100100;
assign LUT_2[20076] = 32'b11111111111111110010110000110111;
assign LUT_2[20077] = 32'b11111111111111101111101001010000;
assign LUT_2[20078] = 32'b11111111111111111001101001110011;
assign LUT_2[20079] = 32'b11111111111111110110100010001100;
assign LUT_2[20080] = 32'b11111111111111110110000101111100;
assign LUT_2[20081] = 32'b11111111111111110010111110010101;
assign LUT_2[20082] = 32'b11111111111111111100111110111000;
assign LUT_2[20083] = 32'b11111111111111111001110111010001;
assign LUT_2[20084] = 32'b11111111111111110010100011100100;
assign LUT_2[20085] = 32'b11111111111111101111011011111101;
assign LUT_2[20086] = 32'b11111111111111111001011100100000;
assign LUT_2[20087] = 32'b11111111111111110110010100111001;
assign LUT_2[20088] = 32'b11111111111111110000110111011001;
assign LUT_2[20089] = 32'b11111111111111101101101111110010;
assign LUT_2[20090] = 32'b11111111111111110111110000010101;
assign LUT_2[20091] = 32'b11111111111111110100101000101110;
assign LUT_2[20092] = 32'b11111111111111101101010101000001;
assign LUT_2[20093] = 32'b11111111111111101010001101011010;
assign LUT_2[20094] = 32'b11111111111111110100001101111101;
assign LUT_2[20095] = 32'b11111111111111110001000110010110;
assign LUT_2[20096] = 32'b00000000000000000111010001110101;
assign LUT_2[20097] = 32'b00000000000000000100001010001110;
assign LUT_2[20098] = 32'b00000000000000001110001010110001;
assign LUT_2[20099] = 32'b00000000000000001011000011001010;
assign LUT_2[20100] = 32'b00000000000000000011101111011101;
assign LUT_2[20101] = 32'b00000000000000000000100111110110;
assign LUT_2[20102] = 32'b00000000000000001010101000011001;
assign LUT_2[20103] = 32'b00000000000000000111100000110010;
assign LUT_2[20104] = 32'b00000000000000000010000011010010;
assign LUT_2[20105] = 32'b11111111111111111110111011101011;
assign LUT_2[20106] = 32'b00000000000000001000111100001110;
assign LUT_2[20107] = 32'b00000000000000000101110100100111;
assign LUT_2[20108] = 32'b11111111111111111110100000111010;
assign LUT_2[20109] = 32'b11111111111111111011011001010011;
assign LUT_2[20110] = 32'b00000000000000000101011001110110;
assign LUT_2[20111] = 32'b00000000000000000010010010001111;
assign LUT_2[20112] = 32'b00000000000000000001110101111111;
assign LUT_2[20113] = 32'b11111111111111111110101110011000;
assign LUT_2[20114] = 32'b00000000000000001000101110111011;
assign LUT_2[20115] = 32'b00000000000000000101100111010100;
assign LUT_2[20116] = 32'b11111111111111111110010011100111;
assign LUT_2[20117] = 32'b11111111111111111011001100000000;
assign LUT_2[20118] = 32'b00000000000000000101001100100011;
assign LUT_2[20119] = 32'b00000000000000000010000100111100;
assign LUT_2[20120] = 32'b11111111111111111100100111011100;
assign LUT_2[20121] = 32'b11111111111111111001011111110101;
assign LUT_2[20122] = 32'b00000000000000000011100000011000;
assign LUT_2[20123] = 32'b00000000000000000000011000110001;
assign LUT_2[20124] = 32'b11111111111111111001000101000100;
assign LUT_2[20125] = 32'b11111111111111110101111101011101;
assign LUT_2[20126] = 32'b11111111111111111111111110000000;
assign LUT_2[20127] = 32'b11111111111111111100110110011001;
assign LUT_2[20128] = 32'b00000000000000000111101101011110;
assign LUT_2[20129] = 32'b00000000000000000100100101110111;
assign LUT_2[20130] = 32'b00000000000000001110100110011010;
assign LUT_2[20131] = 32'b00000000000000001011011110110011;
assign LUT_2[20132] = 32'b00000000000000000100001011000110;
assign LUT_2[20133] = 32'b00000000000000000001000011011111;
assign LUT_2[20134] = 32'b00000000000000001011000100000010;
assign LUT_2[20135] = 32'b00000000000000000111111100011011;
assign LUT_2[20136] = 32'b00000000000000000010011110111011;
assign LUT_2[20137] = 32'b11111111111111111111010111010100;
assign LUT_2[20138] = 32'b00000000000000001001010111110111;
assign LUT_2[20139] = 32'b00000000000000000110010000010000;
assign LUT_2[20140] = 32'b11111111111111111110111100100011;
assign LUT_2[20141] = 32'b11111111111111111011110100111100;
assign LUT_2[20142] = 32'b00000000000000000101110101011111;
assign LUT_2[20143] = 32'b00000000000000000010101101111000;
assign LUT_2[20144] = 32'b00000000000000000010010001101000;
assign LUT_2[20145] = 32'b11111111111111111111001010000001;
assign LUT_2[20146] = 32'b00000000000000001001001010100100;
assign LUT_2[20147] = 32'b00000000000000000110000010111101;
assign LUT_2[20148] = 32'b11111111111111111110101111010000;
assign LUT_2[20149] = 32'b11111111111111111011100111101001;
assign LUT_2[20150] = 32'b00000000000000000101101000001100;
assign LUT_2[20151] = 32'b00000000000000000010100000100101;
assign LUT_2[20152] = 32'b11111111111111111101000011000101;
assign LUT_2[20153] = 32'b11111111111111111001111011011110;
assign LUT_2[20154] = 32'b00000000000000000011111100000001;
assign LUT_2[20155] = 32'b00000000000000000000110100011010;
assign LUT_2[20156] = 32'b11111111111111111001100000101101;
assign LUT_2[20157] = 32'b11111111111111110110011001000110;
assign LUT_2[20158] = 32'b00000000000000000000011001101001;
assign LUT_2[20159] = 32'b11111111111111111101010010000010;
assign LUT_2[20160] = 32'b11111111111111111111011010011000;
assign LUT_2[20161] = 32'b11111111111111111100010010110001;
assign LUT_2[20162] = 32'b00000000000000000110010011010100;
assign LUT_2[20163] = 32'b00000000000000000011001011101101;
assign LUT_2[20164] = 32'b11111111111111111011111000000000;
assign LUT_2[20165] = 32'b11111111111111111000110000011001;
assign LUT_2[20166] = 32'b00000000000000000010110000111100;
assign LUT_2[20167] = 32'b11111111111111111111101001010101;
assign LUT_2[20168] = 32'b11111111111111111010001011110101;
assign LUT_2[20169] = 32'b11111111111111110111000100001110;
assign LUT_2[20170] = 32'b00000000000000000001000100110001;
assign LUT_2[20171] = 32'b11111111111111111101111101001010;
assign LUT_2[20172] = 32'b11111111111111110110101001011101;
assign LUT_2[20173] = 32'b11111111111111110011100001110110;
assign LUT_2[20174] = 32'b11111111111111111101100010011001;
assign LUT_2[20175] = 32'b11111111111111111010011010110010;
assign LUT_2[20176] = 32'b11111111111111111001111110100010;
assign LUT_2[20177] = 32'b11111111111111110110110110111011;
assign LUT_2[20178] = 32'b00000000000000000000110111011110;
assign LUT_2[20179] = 32'b11111111111111111101101111110111;
assign LUT_2[20180] = 32'b11111111111111110110011100001010;
assign LUT_2[20181] = 32'b11111111111111110011010100100011;
assign LUT_2[20182] = 32'b11111111111111111101010101000110;
assign LUT_2[20183] = 32'b11111111111111111010001101011111;
assign LUT_2[20184] = 32'b11111111111111110100101111111111;
assign LUT_2[20185] = 32'b11111111111111110001101000011000;
assign LUT_2[20186] = 32'b11111111111111111011101000111011;
assign LUT_2[20187] = 32'b11111111111111111000100001010100;
assign LUT_2[20188] = 32'b11111111111111110001001101100111;
assign LUT_2[20189] = 32'b11111111111111101110000110000000;
assign LUT_2[20190] = 32'b11111111111111111000000110100011;
assign LUT_2[20191] = 32'b11111111111111110100111110111100;
assign LUT_2[20192] = 32'b11111111111111111111110110000001;
assign LUT_2[20193] = 32'b11111111111111111100101110011010;
assign LUT_2[20194] = 32'b00000000000000000110101110111101;
assign LUT_2[20195] = 32'b00000000000000000011100111010110;
assign LUT_2[20196] = 32'b11111111111111111100010011101001;
assign LUT_2[20197] = 32'b11111111111111111001001100000010;
assign LUT_2[20198] = 32'b00000000000000000011001100100101;
assign LUT_2[20199] = 32'b00000000000000000000000100111110;
assign LUT_2[20200] = 32'b11111111111111111010100111011110;
assign LUT_2[20201] = 32'b11111111111111110111011111110111;
assign LUT_2[20202] = 32'b00000000000000000001100000011010;
assign LUT_2[20203] = 32'b11111111111111111110011000110011;
assign LUT_2[20204] = 32'b11111111111111110111000101000110;
assign LUT_2[20205] = 32'b11111111111111110011111101011111;
assign LUT_2[20206] = 32'b11111111111111111101111110000010;
assign LUT_2[20207] = 32'b11111111111111111010110110011011;
assign LUT_2[20208] = 32'b11111111111111111010011010001011;
assign LUT_2[20209] = 32'b11111111111111110111010010100100;
assign LUT_2[20210] = 32'b00000000000000000001010011000111;
assign LUT_2[20211] = 32'b11111111111111111110001011100000;
assign LUT_2[20212] = 32'b11111111111111110110110111110011;
assign LUT_2[20213] = 32'b11111111111111110011110000001100;
assign LUT_2[20214] = 32'b11111111111111111101110000101111;
assign LUT_2[20215] = 32'b11111111111111111010101001001000;
assign LUT_2[20216] = 32'b11111111111111110101001011101000;
assign LUT_2[20217] = 32'b11111111111111110010000100000001;
assign LUT_2[20218] = 32'b11111111111111111100000100100100;
assign LUT_2[20219] = 32'b11111111111111111000111100111101;
assign LUT_2[20220] = 32'b11111111111111110001101001010000;
assign LUT_2[20221] = 32'b11111111111111101110100001101001;
assign LUT_2[20222] = 32'b11111111111111111000100010001100;
assign LUT_2[20223] = 32'b11111111111111110101011010100101;
assign LUT_2[20224] = 32'b00000000000000000110111100001100;
assign LUT_2[20225] = 32'b00000000000000000011110100100101;
assign LUT_2[20226] = 32'b00000000000000001101110101001000;
assign LUT_2[20227] = 32'b00000000000000001010101101100001;
assign LUT_2[20228] = 32'b00000000000000000011011001110100;
assign LUT_2[20229] = 32'b00000000000000000000010010001101;
assign LUT_2[20230] = 32'b00000000000000001010010010110000;
assign LUT_2[20231] = 32'b00000000000000000111001011001001;
assign LUT_2[20232] = 32'b00000000000000000001101101101001;
assign LUT_2[20233] = 32'b11111111111111111110100110000010;
assign LUT_2[20234] = 32'b00000000000000001000100110100101;
assign LUT_2[20235] = 32'b00000000000000000101011110111110;
assign LUT_2[20236] = 32'b11111111111111111110001011010001;
assign LUT_2[20237] = 32'b11111111111111111011000011101010;
assign LUT_2[20238] = 32'b00000000000000000101000100001101;
assign LUT_2[20239] = 32'b00000000000000000001111100100110;
assign LUT_2[20240] = 32'b00000000000000000001100000010110;
assign LUT_2[20241] = 32'b11111111111111111110011000101111;
assign LUT_2[20242] = 32'b00000000000000001000011001010010;
assign LUT_2[20243] = 32'b00000000000000000101010001101011;
assign LUT_2[20244] = 32'b11111111111111111101111101111110;
assign LUT_2[20245] = 32'b11111111111111111010110110010111;
assign LUT_2[20246] = 32'b00000000000000000100110110111010;
assign LUT_2[20247] = 32'b00000000000000000001101111010011;
assign LUT_2[20248] = 32'b11111111111111111100010001110011;
assign LUT_2[20249] = 32'b11111111111111111001001010001100;
assign LUT_2[20250] = 32'b00000000000000000011001010101111;
assign LUT_2[20251] = 32'b00000000000000000000000011001000;
assign LUT_2[20252] = 32'b11111111111111111000101111011011;
assign LUT_2[20253] = 32'b11111111111111110101100111110100;
assign LUT_2[20254] = 32'b11111111111111111111101000010111;
assign LUT_2[20255] = 32'b11111111111111111100100000110000;
assign LUT_2[20256] = 32'b00000000000000000111010111110101;
assign LUT_2[20257] = 32'b00000000000000000100010000001110;
assign LUT_2[20258] = 32'b00000000000000001110010000110001;
assign LUT_2[20259] = 32'b00000000000000001011001001001010;
assign LUT_2[20260] = 32'b00000000000000000011110101011101;
assign LUT_2[20261] = 32'b00000000000000000000101101110110;
assign LUT_2[20262] = 32'b00000000000000001010101110011001;
assign LUT_2[20263] = 32'b00000000000000000111100110110010;
assign LUT_2[20264] = 32'b00000000000000000010001001010010;
assign LUT_2[20265] = 32'b11111111111111111111000001101011;
assign LUT_2[20266] = 32'b00000000000000001001000010001110;
assign LUT_2[20267] = 32'b00000000000000000101111010100111;
assign LUT_2[20268] = 32'b11111111111111111110100110111010;
assign LUT_2[20269] = 32'b11111111111111111011011111010011;
assign LUT_2[20270] = 32'b00000000000000000101011111110110;
assign LUT_2[20271] = 32'b00000000000000000010011000001111;
assign LUT_2[20272] = 32'b00000000000000000001111011111111;
assign LUT_2[20273] = 32'b11111111111111111110110100011000;
assign LUT_2[20274] = 32'b00000000000000001000110100111011;
assign LUT_2[20275] = 32'b00000000000000000101101101010100;
assign LUT_2[20276] = 32'b11111111111111111110011001100111;
assign LUT_2[20277] = 32'b11111111111111111011010010000000;
assign LUT_2[20278] = 32'b00000000000000000101010010100011;
assign LUT_2[20279] = 32'b00000000000000000010001010111100;
assign LUT_2[20280] = 32'b11111111111111111100101101011100;
assign LUT_2[20281] = 32'b11111111111111111001100101110101;
assign LUT_2[20282] = 32'b00000000000000000011100110011000;
assign LUT_2[20283] = 32'b00000000000000000000011110110001;
assign LUT_2[20284] = 32'b11111111111111111001001011000100;
assign LUT_2[20285] = 32'b11111111111111110110000011011101;
assign LUT_2[20286] = 32'b00000000000000000000000100000000;
assign LUT_2[20287] = 32'b11111111111111111100111100011001;
assign LUT_2[20288] = 32'b11111111111111111111000100101111;
assign LUT_2[20289] = 32'b11111111111111111011111101001000;
assign LUT_2[20290] = 32'b00000000000000000101111101101011;
assign LUT_2[20291] = 32'b00000000000000000010110110000100;
assign LUT_2[20292] = 32'b11111111111111111011100010010111;
assign LUT_2[20293] = 32'b11111111111111111000011010110000;
assign LUT_2[20294] = 32'b00000000000000000010011011010011;
assign LUT_2[20295] = 32'b11111111111111111111010011101100;
assign LUT_2[20296] = 32'b11111111111111111001110110001100;
assign LUT_2[20297] = 32'b11111111111111110110101110100101;
assign LUT_2[20298] = 32'b00000000000000000000101111001000;
assign LUT_2[20299] = 32'b11111111111111111101100111100001;
assign LUT_2[20300] = 32'b11111111111111110110010011110100;
assign LUT_2[20301] = 32'b11111111111111110011001100001101;
assign LUT_2[20302] = 32'b11111111111111111101001100110000;
assign LUT_2[20303] = 32'b11111111111111111010000101001001;
assign LUT_2[20304] = 32'b11111111111111111001101000111001;
assign LUT_2[20305] = 32'b11111111111111110110100001010010;
assign LUT_2[20306] = 32'b00000000000000000000100001110101;
assign LUT_2[20307] = 32'b11111111111111111101011010001110;
assign LUT_2[20308] = 32'b11111111111111110110000110100001;
assign LUT_2[20309] = 32'b11111111111111110010111110111010;
assign LUT_2[20310] = 32'b11111111111111111100111111011101;
assign LUT_2[20311] = 32'b11111111111111111001110111110110;
assign LUT_2[20312] = 32'b11111111111111110100011010010110;
assign LUT_2[20313] = 32'b11111111111111110001010010101111;
assign LUT_2[20314] = 32'b11111111111111111011010011010010;
assign LUT_2[20315] = 32'b11111111111111111000001011101011;
assign LUT_2[20316] = 32'b11111111111111110000110111111110;
assign LUT_2[20317] = 32'b11111111111111101101110000010111;
assign LUT_2[20318] = 32'b11111111111111110111110000111010;
assign LUT_2[20319] = 32'b11111111111111110100101001010011;
assign LUT_2[20320] = 32'b11111111111111111111100000011000;
assign LUT_2[20321] = 32'b11111111111111111100011000110001;
assign LUT_2[20322] = 32'b00000000000000000110011001010100;
assign LUT_2[20323] = 32'b00000000000000000011010001101101;
assign LUT_2[20324] = 32'b11111111111111111011111110000000;
assign LUT_2[20325] = 32'b11111111111111111000110110011001;
assign LUT_2[20326] = 32'b00000000000000000010110110111100;
assign LUT_2[20327] = 32'b11111111111111111111101111010101;
assign LUT_2[20328] = 32'b11111111111111111010010001110101;
assign LUT_2[20329] = 32'b11111111111111110111001010001110;
assign LUT_2[20330] = 32'b00000000000000000001001010110001;
assign LUT_2[20331] = 32'b11111111111111111110000011001010;
assign LUT_2[20332] = 32'b11111111111111110110101111011101;
assign LUT_2[20333] = 32'b11111111111111110011100111110110;
assign LUT_2[20334] = 32'b11111111111111111101101000011001;
assign LUT_2[20335] = 32'b11111111111111111010100000110010;
assign LUT_2[20336] = 32'b11111111111111111010000100100010;
assign LUT_2[20337] = 32'b11111111111111110110111100111011;
assign LUT_2[20338] = 32'b00000000000000000000111101011110;
assign LUT_2[20339] = 32'b11111111111111111101110101110111;
assign LUT_2[20340] = 32'b11111111111111110110100010001010;
assign LUT_2[20341] = 32'b11111111111111110011011010100011;
assign LUT_2[20342] = 32'b11111111111111111101011011000110;
assign LUT_2[20343] = 32'b11111111111111111010010011011111;
assign LUT_2[20344] = 32'b11111111111111110100110101111111;
assign LUT_2[20345] = 32'b11111111111111110001101110011000;
assign LUT_2[20346] = 32'b11111111111111111011101110111011;
assign LUT_2[20347] = 32'b11111111111111111000100111010100;
assign LUT_2[20348] = 32'b11111111111111110001010011100111;
assign LUT_2[20349] = 32'b11111111111111101110001100000000;
assign LUT_2[20350] = 32'b11111111111111111000001100100011;
assign LUT_2[20351] = 32'b11111111111111110101000100111100;
assign LUT_2[20352] = 32'b00000000000000001011010000011011;
assign LUT_2[20353] = 32'b00000000000000001000001000110100;
assign LUT_2[20354] = 32'b00000000000000010010001001010111;
assign LUT_2[20355] = 32'b00000000000000001111000001110000;
assign LUT_2[20356] = 32'b00000000000000000111101110000011;
assign LUT_2[20357] = 32'b00000000000000000100100110011100;
assign LUT_2[20358] = 32'b00000000000000001110100110111111;
assign LUT_2[20359] = 32'b00000000000000001011011111011000;
assign LUT_2[20360] = 32'b00000000000000000110000001111000;
assign LUT_2[20361] = 32'b00000000000000000010111010010001;
assign LUT_2[20362] = 32'b00000000000000001100111010110100;
assign LUT_2[20363] = 32'b00000000000000001001110011001101;
assign LUT_2[20364] = 32'b00000000000000000010011111100000;
assign LUT_2[20365] = 32'b11111111111111111111010111111001;
assign LUT_2[20366] = 32'b00000000000000001001011000011100;
assign LUT_2[20367] = 32'b00000000000000000110010000110101;
assign LUT_2[20368] = 32'b00000000000000000101110100100101;
assign LUT_2[20369] = 32'b00000000000000000010101100111110;
assign LUT_2[20370] = 32'b00000000000000001100101101100001;
assign LUT_2[20371] = 32'b00000000000000001001100101111010;
assign LUT_2[20372] = 32'b00000000000000000010010010001101;
assign LUT_2[20373] = 32'b11111111111111111111001010100110;
assign LUT_2[20374] = 32'b00000000000000001001001011001001;
assign LUT_2[20375] = 32'b00000000000000000110000011100010;
assign LUT_2[20376] = 32'b00000000000000000000100110000010;
assign LUT_2[20377] = 32'b11111111111111111101011110011011;
assign LUT_2[20378] = 32'b00000000000000000111011110111110;
assign LUT_2[20379] = 32'b00000000000000000100010111010111;
assign LUT_2[20380] = 32'b11111111111111111101000011101010;
assign LUT_2[20381] = 32'b11111111111111111001111100000011;
assign LUT_2[20382] = 32'b00000000000000000011111100100110;
assign LUT_2[20383] = 32'b00000000000000000000110100111111;
assign LUT_2[20384] = 32'b00000000000000001011101100000100;
assign LUT_2[20385] = 32'b00000000000000001000100100011101;
assign LUT_2[20386] = 32'b00000000000000010010100101000000;
assign LUT_2[20387] = 32'b00000000000000001111011101011001;
assign LUT_2[20388] = 32'b00000000000000001000001001101100;
assign LUT_2[20389] = 32'b00000000000000000101000010000101;
assign LUT_2[20390] = 32'b00000000000000001111000010101000;
assign LUT_2[20391] = 32'b00000000000000001011111011000001;
assign LUT_2[20392] = 32'b00000000000000000110011101100001;
assign LUT_2[20393] = 32'b00000000000000000011010101111010;
assign LUT_2[20394] = 32'b00000000000000001101010110011101;
assign LUT_2[20395] = 32'b00000000000000001010001110110110;
assign LUT_2[20396] = 32'b00000000000000000010111011001001;
assign LUT_2[20397] = 32'b11111111111111111111110011100010;
assign LUT_2[20398] = 32'b00000000000000001001110100000101;
assign LUT_2[20399] = 32'b00000000000000000110101100011110;
assign LUT_2[20400] = 32'b00000000000000000110010000001110;
assign LUT_2[20401] = 32'b00000000000000000011001000100111;
assign LUT_2[20402] = 32'b00000000000000001101001001001010;
assign LUT_2[20403] = 32'b00000000000000001010000001100011;
assign LUT_2[20404] = 32'b00000000000000000010101101110110;
assign LUT_2[20405] = 32'b11111111111111111111100110001111;
assign LUT_2[20406] = 32'b00000000000000001001100110110010;
assign LUT_2[20407] = 32'b00000000000000000110011111001011;
assign LUT_2[20408] = 32'b00000000000000000001000001101011;
assign LUT_2[20409] = 32'b11111111111111111101111010000100;
assign LUT_2[20410] = 32'b00000000000000000111111010100111;
assign LUT_2[20411] = 32'b00000000000000000100110011000000;
assign LUT_2[20412] = 32'b11111111111111111101011111010011;
assign LUT_2[20413] = 32'b11111111111111111010010111101100;
assign LUT_2[20414] = 32'b00000000000000000100011000001111;
assign LUT_2[20415] = 32'b00000000000000000001010000101000;
assign LUT_2[20416] = 32'b00000000000000000011011000111110;
assign LUT_2[20417] = 32'b00000000000000000000010001010111;
assign LUT_2[20418] = 32'b00000000000000001010010001111010;
assign LUT_2[20419] = 32'b00000000000000000111001010010011;
assign LUT_2[20420] = 32'b11111111111111111111110110100110;
assign LUT_2[20421] = 32'b11111111111111111100101110111111;
assign LUT_2[20422] = 32'b00000000000000000110101111100010;
assign LUT_2[20423] = 32'b00000000000000000011100111111011;
assign LUT_2[20424] = 32'b11111111111111111110001010011011;
assign LUT_2[20425] = 32'b11111111111111111011000010110100;
assign LUT_2[20426] = 32'b00000000000000000101000011010111;
assign LUT_2[20427] = 32'b00000000000000000001111011110000;
assign LUT_2[20428] = 32'b11111111111111111010101000000011;
assign LUT_2[20429] = 32'b11111111111111110111100000011100;
assign LUT_2[20430] = 32'b00000000000000000001100000111111;
assign LUT_2[20431] = 32'b11111111111111111110011001011000;
assign LUT_2[20432] = 32'b11111111111111111101111101001000;
assign LUT_2[20433] = 32'b11111111111111111010110101100001;
assign LUT_2[20434] = 32'b00000000000000000100110110000100;
assign LUT_2[20435] = 32'b00000000000000000001101110011101;
assign LUT_2[20436] = 32'b11111111111111111010011010110000;
assign LUT_2[20437] = 32'b11111111111111110111010011001001;
assign LUT_2[20438] = 32'b00000000000000000001010011101100;
assign LUT_2[20439] = 32'b11111111111111111110001100000101;
assign LUT_2[20440] = 32'b11111111111111111000101110100101;
assign LUT_2[20441] = 32'b11111111111111110101100110111110;
assign LUT_2[20442] = 32'b11111111111111111111100111100001;
assign LUT_2[20443] = 32'b11111111111111111100011111111010;
assign LUT_2[20444] = 32'b11111111111111110101001100001101;
assign LUT_2[20445] = 32'b11111111111111110010000100100110;
assign LUT_2[20446] = 32'b11111111111111111100000101001001;
assign LUT_2[20447] = 32'b11111111111111111000111101100010;
assign LUT_2[20448] = 32'b00000000000000000011110100100111;
assign LUT_2[20449] = 32'b00000000000000000000101101000000;
assign LUT_2[20450] = 32'b00000000000000001010101101100011;
assign LUT_2[20451] = 32'b00000000000000000111100101111100;
assign LUT_2[20452] = 32'b00000000000000000000010010001111;
assign LUT_2[20453] = 32'b11111111111111111101001010101000;
assign LUT_2[20454] = 32'b00000000000000000111001011001011;
assign LUT_2[20455] = 32'b00000000000000000100000011100100;
assign LUT_2[20456] = 32'b11111111111111111110100110000100;
assign LUT_2[20457] = 32'b11111111111111111011011110011101;
assign LUT_2[20458] = 32'b00000000000000000101011111000000;
assign LUT_2[20459] = 32'b00000000000000000010010111011001;
assign LUT_2[20460] = 32'b11111111111111111011000011101100;
assign LUT_2[20461] = 32'b11111111111111110111111100000101;
assign LUT_2[20462] = 32'b00000000000000000001111100101000;
assign LUT_2[20463] = 32'b11111111111111111110110101000001;
assign LUT_2[20464] = 32'b11111111111111111110011000110001;
assign LUT_2[20465] = 32'b11111111111111111011010001001010;
assign LUT_2[20466] = 32'b00000000000000000101010001101101;
assign LUT_2[20467] = 32'b00000000000000000010001010000110;
assign LUT_2[20468] = 32'b11111111111111111010110110011001;
assign LUT_2[20469] = 32'b11111111111111110111101110110010;
assign LUT_2[20470] = 32'b00000000000000000001101111010101;
assign LUT_2[20471] = 32'b11111111111111111110100111101110;
assign LUT_2[20472] = 32'b11111111111111111001001010001110;
assign LUT_2[20473] = 32'b11111111111111110110000010100111;
assign LUT_2[20474] = 32'b00000000000000000000000011001010;
assign LUT_2[20475] = 32'b11111111111111111100111011100011;
assign LUT_2[20476] = 32'b11111111111111110101100111110110;
assign LUT_2[20477] = 32'b11111111111111110010100000001111;
assign LUT_2[20478] = 32'b11111111111111111100100000110010;
assign LUT_2[20479] = 32'b11111111111111111001011001001011;
assign LUT_2[20480] = 32'b11111111111111111010101101111110;
assign LUT_2[20481] = 32'b11111111111111110111100110010111;
assign LUT_2[20482] = 32'b00000000000000000001100110111010;
assign LUT_2[20483] = 32'b11111111111111111110011111010011;
assign LUT_2[20484] = 32'b11111111111111110111001011100110;
assign LUT_2[20485] = 32'b11111111111111110100000011111111;
assign LUT_2[20486] = 32'b11111111111111111110000100100010;
assign LUT_2[20487] = 32'b11111111111111111010111100111011;
assign LUT_2[20488] = 32'b11111111111111110101011111011011;
assign LUT_2[20489] = 32'b11111111111111110010010111110100;
assign LUT_2[20490] = 32'b11111111111111111100011000010111;
assign LUT_2[20491] = 32'b11111111111111111001010000110000;
assign LUT_2[20492] = 32'b11111111111111110001111101000011;
assign LUT_2[20493] = 32'b11111111111111101110110101011100;
assign LUT_2[20494] = 32'b11111111111111111000110101111111;
assign LUT_2[20495] = 32'b11111111111111110101101110011000;
assign LUT_2[20496] = 32'b11111111111111110101010010001000;
assign LUT_2[20497] = 32'b11111111111111110010001010100001;
assign LUT_2[20498] = 32'b11111111111111111100001011000100;
assign LUT_2[20499] = 32'b11111111111111111001000011011101;
assign LUT_2[20500] = 32'b11111111111111110001101111110000;
assign LUT_2[20501] = 32'b11111111111111101110101000001001;
assign LUT_2[20502] = 32'b11111111111111111000101000101100;
assign LUT_2[20503] = 32'b11111111111111110101100001000101;
assign LUT_2[20504] = 32'b11111111111111110000000011100101;
assign LUT_2[20505] = 32'b11111111111111101100111011111110;
assign LUT_2[20506] = 32'b11111111111111110110111100100001;
assign LUT_2[20507] = 32'b11111111111111110011110100111010;
assign LUT_2[20508] = 32'b11111111111111101100100001001101;
assign LUT_2[20509] = 32'b11111111111111101001011001100110;
assign LUT_2[20510] = 32'b11111111111111110011011010001001;
assign LUT_2[20511] = 32'b11111111111111110000010010100010;
assign LUT_2[20512] = 32'b11111111111111111011001001100111;
assign LUT_2[20513] = 32'b11111111111111111000000010000000;
assign LUT_2[20514] = 32'b00000000000000000010000010100011;
assign LUT_2[20515] = 32'b11111111111111111110111010111100;
assign LUT_2[20516] = 32'b11111111111111110111100111001111;
assign LUT_2[20517] = 32'b11111111111111110100011111101000;
assign LUT_2[20518] = 32'b11111111111111111110100000001011;
assign LUT_2[20519] = 32'b11111111111111111011011000100100;
assign LUT_2[20520] = 32'b11111111111111110101111011000100;
assign LUT_2[20521] = 32'b11111111111111110010110011011101;
assign LUT_2[20522] = 32'b11111111111111111100110100000000;
assign LUT_2[20523] = 32'b11111111111111111001101100011001;
assign LUT_2[20524] = 32'b11111111111111110010011000101100;
assign LUT_2[20525] = 32'b11111111111111101111010001000101;
assign LUT_2[20526] = 32'b11111111111111111001010001101000;
assign LUT_2[20527] = 32'b11111111111111110110001010000001;
assign LUT_2[20528] = 32'b11111111111111110101101101110001;
assign LUT_2[20529] = 32'b11111111111111110010100110001010;
assign LUT_2[20530] = 32'b11111111111111111100100110101101;
assign LUT_2[20531] = 32'b11111111111111111001011111000110;
assign LUT_2[20532] = 32'b11111111111111110010001011011001;
assign LUT_2[20533] = 32'b11111111111111101111000011110010;
assign LUT_2[20534] = 32'b11111111111111111001000100010101;
assign LUT_2[20535] = 32'b11111111111111110101111100101110;
assign LUT_2[20536] = 32'b11111111111111110000011111001110;
assign LUT_2[20537] = 32'b11111111111111101101010111100111;
assign LUT_2[20538] = 32'b11111111111111110111011000001010;
assign LUT_2[20539] = 32'b11111111111111110100010000100011;
assign LUT_2[20540] = 32'b11111111111111101100111100110110;
assign LUT_2[20541] = 32'b11111111111111101001110101001111;
assign LUT_2[20542] = 32'b11111111111111110011110101110010;
assign LUT_2[20543] = 32'b11111111111111110000101110001011;
assign LUT_2[20544] = 32'b11111111111111110010110110100001;
assign LUT_2[20545] = 32'b11111111111111101111101110111010;
assign LUT_2[20546] = 32'b11111111111111111001101111011101;
assign LUT_2[20547] = 32'b11111111111111110110100111110110;
assign LUT_2[20548] = 32'b11111111111111101111010100001001;
assign LUT_2[20549] = 32'b11111111111111101100001100100010;
assign LUT_2[20550] = 32'b11111111111111110110001101000101;
assign LUT_2[20551] = 32'b11111111111111110011000101011110;
assign LUT_2[20552] = 32'b11111111111111101101100111111110;
assign LUT_2[20553] = 32'b11111111111111101010100000010111;
assign LUT_2[20554] = 32'b11111111111111110100100000111010;
assign LUT_2[20555] = 32'b11111111111111110001011001010011;
assign LUT_2[20556] = 32'b11111111111111101010000101100110;
assign LUT_2[20557] = 32'b11111111111111100110111101111111;
assign LUT_2[20558] = 32'b11111111111111110000111110100010;
assign LUT_2[20559] = 32'b11111111111111101101110110111011;
assign LUT_2[20560] = 32'b11111111111111101101011010101011;
assign LUT_2[20561] = 32'b11111111111111101010010011000100;
assign LUT_2[20562] = 32'b11111111111111110100010011100111;
assign LUT_2[20563] = 32'b11111111111111110001001100000000;
assign LUT_2[20564] = 32'b11111111111111101001111000010011;
assign LUT_2[20565] = 32'b11111111111111100110110000101100;
assign LUT_2[20566] = 32'b11111111111111110000110001001111;
assign LUT_2[20567] = 32'b11111111111111101101101001101000;
assign LUT_2[20568] = 32'b11111111111111101000001100001000;
assign LUT_2[20569] = 32'b11111111111111100101000100100001;
assign LUT_2[20570] = 32'b11111111111111101111000101000100;
assign LUT_2[20571] = 32'b11111111111111101011111101011101;
assign LUT_2[20572] = 32'b11111111111111100100101001110000;
assign LUT_2[20573] = 32'b11111111111111100001100010001001;
assign LUT_2[20574] = 32'b11111111111111101011100010101100;
assign LUT_2[20575] = 32'b11111111111111101000011011000101;
assign LUT_2[20576] = 32'b11111111111111110011010010001010;
assign LUT_2[20577] = 32'b11111111111111110000001010100011;
assign LUT_2[20578] = 32'b11111111111111111010001011000110;
assign LUT_2[20579] = 32'b11111111111111110111000011011111;
assign LUT_2[20580] = 32'b11111111111111101111101111110010;
assign LUT_2[20581] = 32'b11111111111111101100101000001011;
assign LUT_2[20582] = 32'b11111111111111110110101000101110;
assign LUT_2[20583] = 32'b11111111111111110011100001000111;
assign LUT_2[20584] = 32'b11111111111111101110000011100111;
assign LUT_2[20585] = 32'b11111111111111101010111100000000;
assign LUT_2[20586] = 32'b11111111111111110100111100100011;
assign LUT_2[20587] = 32'b11111111111111110001110100111100;
assign LUT_2[20588] = 32'b11111111111111101010100001001111;
assign LUT_2[20589] = 32'b11111111111111100111011001101000;
assign LUT_2[20590] = 32'b11111111111111110001011010001011;
assign LUT_2[20591] = 32'b11111111111111101110010010100100;
assign LUT_2[20592] = 32'b11111111111111101101110110010100;
assign LUT_2[20593] = 32'b11111111111111101010101110101101;
assign LUT_2[20594] = 32'b11111111111111110100101111010000;
assign LUT_2[20595] = 32'b11111111111111110001100111101001;
assign LUT_2[20596] = 32'b11111111111111101010010011111100;
assign LUT_2[20597] = 32'b11111111111111100111001100010101;
assign LUT_2[20598] = 32'b11111111111111110001001100111000;
assign LUT_2[20599] = 32'b11111111111111101110000101010001;
assign LUT_2[20600] = 32'b11111111111111101000100111110001;
assign LUT_2[20601] = 32'b11111111111111100101100000001010;
assign LUT_2[20602] = 32'b11111111111111101111100000101101;
assign LUT_2[20603] = 32'b11111111111111101100011001000110;
assign LUT_2[20604] = 32'b11111111111111100101000101011001;
assign LUT_2[20605] = 32'b11111111111111100001111101110010;
assign LUT_2[20606] = 32'b11111111111111101011111110010101;
assign LUT_2[20607] = 32'b11111111111111101000110110101110;
assign LUT_2[20608] = 32'b11111111111111111111000010001101;
assign LUT_2[20609] = 32'b11111111111111111011111010100110;
assign LUT_2[20610] = 32'b00000000000000000101111011001001;
assign LUT_2[20611] = 32'b00000000000000000010110011100010;
assign LUT_2[20612] = 32'b11111111111111111011011111110101;
assign LUT_2[20613] = 32'b11111111111111111000011000001110;
assign LUT_2[20614] = 32'b00000000000000000010011000110001;
assign LUT_2[20615] = 32'b11111111111111111111010001001010;
assign LUT_2[20616] = 32'b11111111111111111001110011101010;
assign LUT_2[20617] = 32'b11111111111111110110101100000011;
assign LUT_2[20618] = 32'b00000000000000000000101100100110;
assign LUT_2[20619] = 32'b11111111111111111101100100111111;
assign LUT_2[20620] = 32'b11111111111111110110010001010010;
assign LUT_2[20621] = 32'b11111111111111110011001001101011;
assign LUT_2[20622] = 32'b11111111111111111101001010001110;
assign LUT_2[20623] = 32'b11111111111111111010000010100111;
assign LUT_2[20624] = 32'b11111111111111111001100110010111;
assign LUT_2[20625] = 32'b11111111111111110110011110110000;
assign LUT_2[20626] = 32'b00000000000000000000011111010011;
assign LUT_2[20627] = 32'b11111111111111111101010111101100;
assign LUT_2[20628] = 32'b11111111111111110110000011111111;
assign LUT_2[20629] = 32'b11111111111111110010111100011000;
assign LUT_2[20630] = 32'b11111111111111111100111100111011;
assign LUT_2[20631] = 32'b11111111111111111001110101010100;
assign LUT_2[20632] = 32'b11111111111111110100010111110100;
assign LUT_2[20633] = 32'b11111111111111110001010000001101;
assign LUT_2[20634] = 32'b11111111111111111011010000110000;
assign LUT_2[20635] = 32'b11111111111111111000001001001001;
assign LUT_2[20636] = 32'b11111111111111110000110101011100;
assign LUT_2[20637] = 32'b11111111111111101101101101110101;
assign LUT_2[20638] = 32'b11111111111111110111101110011000;
assign LUT_2[20639] = 32'b11111111111111110100100110110001;
assign LUT_2[20640] = 32'b11111111111111111111011101110110;
assign LUT_2[20641] = 32'b11111111111111111100010110001111;
assign LUT_2[20642] = 32'b00000000000000000110010110110010;
assign LUT_2[20643] = 32'b00000000000000000011001111001011;
assign LUT_2[20644] = 32'b11111111111111111011111011011110;
assign LUT_2[20645] = 32'b11111111111111111000110011110111;
assign LUT_2[20646] = 32'b00000000000000000010110100011010;
assign LUT_2[20647] = 32'b11111111111111111111101100110011;
assign LUT_2[20648] = 32'b11111111111111111010001111010011;
assign LUT_2[20649] = 32'b11111111111111110111000111101100;
assign LUT_2[20650] = 32'b00000000000000000001001000001111;
assign LUT_2[20651] = 32'b11111111111111111110000000101000;
assign LUT_2[20652] = 32'b11111111111111110110101100111011;
assign LUT_2[20653] = 32'b11111111111111110011100101010100;
assign LUT_2[20654] = 32'b11111111111111111101100101110111;
assign LUT_2[20655] = 32'b11111111111111111010011110010000;
assign LUT_2[20656] = 32'b11111111111111111010000010000000;
assign LUT_2[20657] = 32'b11111111111111110110111010011001;
assign LUT_2[20658] = 32'b00000000000000000000111010111100;
assign LUT_2[20659] = 32'b11111111111111111101110011010101;
assign LUT_2[20660] = 32'b11111111111111110110011111101000;
assign LUT_2[20661] = 32'b11111111111111110011011000000001;
assign LUT_2[20662] = 32'b11111111111111111101011000100100;
assign LUT_2[20663] = 32'b11111111111111111010010000111101;
assign LUT_2[20664] = 32'b11111111111111110100110011011101;
assign LUT_2[20665] = 32'b11111111111111110001101011110110;
assign LUT_2[20666] = 32'b11111111111111111011101100011001;
assign LUT_2[20667] = 32'b11111111111111111000100100110010;
assign LUT_2[20668] = 32'b11111111111111110001010001000101;
assign LUT_2[20669] = 32'b11111111111111101110001001011110;
assign LUT_2[20670] = 32'b11111111111111111000001010000001;
assign LUT_2[20671] = 32'b11111111111111110101000010011010;
assign LUT_2[20672] = 32'b11111111111111110111001010110000;
assign LUT_2[20673] = 32'b11111111111111110100000011001001;
assign LUT_2[20674] = 32'b11111111111111111110000011101100;
assign LUT_2[20675] = 32'b11111111111111111010111100000101;
assign LUT_2[20676] = 32'b11111111111111110011101000011000;
assign LUT_2[20677] = 32'b11111111111111110000100000110001;
assign LUT_2[20678] = 32'b11111111111111111010100001010100;
assign LUT_2[20679] = 32'b11111111111111110111011001101101;
assign LUT_2[20680] = 32'b11111111111111110001111100001101;
assign LUT_2[20681] = 32'b11111111111111101110110100100110;
assign LUT_2[20682] = 32'b11111111111111111000110101001001;
assign LUT_2[20683] = 32'b11111111111111110101101101100010;
assign LUT_2[20684] = 32'b11111111111111101110011001110101;
assign LUT_2[20685] = 32'b11111111111111101011010010001110;
assign LUT_2[20686] = 32'b11111111111111110101010010110001;
assign LUT_2[20687] = 32'b11111111111111110010001011001010;
assign LUT_2[20688] = 32'b11111111111111110001101110111010;
assign LUT_2[20689] = 32'b11111111111111101110100111010011;
assign LUT_2[20690] = 32'b11111111111111111000100111110110;
assign LUT_2[20691] = 32'b11111111111111110101100000001111;
assign LUT_2[20692] = 32'b11111111111111101110001100100010;
assign LUT_2[20693] = 32'b11111111111111101011000100111011;
assign LUT_2[20694] = 32'b11111111111111110101000101011110;
assign LUT_2[20695] = 32'b11111111111111110001111101110111;
assign LUT_2[20696] = 32'b11111111111111101100100000010111;
assign LUT_2[20697] = 32'b11111111111111101001011000110000;
assign LUT_2[20698] = 32'b11111111111111110011011001010011;
assign LUT_2[20699] = 32'b11111111111111110000010001101100;
assign LUT_2[20700] = 32'b11111111111111101000111101111111;
assign LUT_2[20701] = 32'b11111111111111100101110110011000;
assign LUT_2[20702] = 32'b11111111111111101111110110111011;
assign LUT_2[20703] = 32'b11111111111111101100101111010100;
assign LUT_2[20704] = 32'b11111111111111110111100110011001;
assign LUT_2[20705] = 32'b11111111111111110100011110110010;
assign LUT_2[20706] = 32'b11111111111111111110011111010101;
assign LUT_2[20707] = 32'b11111111111111111011010111101110;
assign LUT_2[20708] = 32'b11111111111111110100000100000001;
assign LUT_2[20709] = 32'b11111111111111110000111100011010;
assign LUT_2[20710] = 32'b11111111111111111010111100111101;
assign LUT_2[20711] = 32'b11111111111111110111110101010110;
assign LUT_2[20712] = 32'b11111111111111110010010111110110;
assign LUT_2[20713] = 32'b11111111111111101111010000001111;
assign LUT_2[20714] = 32'b11111111111111111001010000110010;
assign LUT_2[20715] = 32'b11111111111111110110001001001011;
assign LUT_2[20716] = 32'b11111111111111101110110101011110;
assign LUT_2[20717] = 32'b11111111111111101011101101110111;
assign LUT_2[20718] = 32'b11111111111111110101101110011010;
assign LUT_2[20719] = 32'b11111111111111110010100110110011;
assign LUT_2[20720] = 32'b11111111111111110010001010100011;
assign LUT_2[20721] = 32'b11111111111111101111000010111100;
assign LUT_2[20722] = 32'b11111111111111111001000011011111;
assign LUT_2[20723] = 32'b11111111111111110101111011111000;
assign LUT_2[20724] = 32'b11111111111111101110101000001011;
assign LUT_2[20725] = 32'b11111111111111101011100000100100;
assign LUT_2[20726] = 32'b11111111111111110101100001000111;
assign LUT_2[20727] = 32'b11111111111111110010011001100000;
assign LUT_2[20728] = 32'b11111111111111101100111100000000;
assign LUT_2[20729] = 32'b11111111111111101001110100011001;
assign LUT_2[20730] = 32'b11111111111111110011110100111100;
assign LUT_2[20731] = 32'b11111111111111110000101101010101;
assign LUT_2[20732] = 32'b11111111111111101001011001101000;
assign LUT_2[20733] = 32'b11111111111111100110010010000001;
assign LUT_2[20734] = 32'b11111111111111110000010010100100;
assign LUT_2[20735] = 32'b11111111111111101101001010111101;
assign LUT_2[20736] = 32'b11111111111111111110101100100100;
assign LUT_2[20737] = 32'b11111111111111111011100100111101;
assign LUT_2[20738] = 32'b00000000000000000101100101100000;
assign LUT_2[20739] = 32'b00000000000000000010011101111001;
assign LUT_2[20740] = 32'b11111111111111111011001010001100;
assign LUT_2[20741] = 32'b11111111111111111000000010100101;
assign LUT_2[20742] = 32'b00000000000000000010000011001000;
assign LUT_2[20743] = 32'b11111111111111111110111011100001;
assign LUT_2[20744] = 32'b11111111111111111001011110000001;
assign LUT_2[20745] = 32'b11111111111111110110010110011010;
assign LUT_2[20746] = 32'b00000000000000000000010110111101;
assign LUT_2[20747] = 32'b11111111111111111101001111010110;
assign LUT_2[20748] = 32'b11111111111111110101111011101001;
assign LUT_2[20749] = 32'b11111111111111110010110100000010;
assign LUT_2[20750] = 32'b11111111111111111100110100100101;
assign LUT_2[20751] = 32'b11111111111111111001101100111110;
assign LUT_2[20752] = 32'b11111111111111111001010000101110;
assign LUT_2[20753] = 32'b11111111111111110110001001000111;
assign LUT_2[20754] = 32'b00000000000000000000001001101010;
assign LUT_2[20755] = 32'b11111111111111111101000010000011;
assign LUT_2[20756] = 32'b11111111111111110101101110010110;
assign LUT_2[20757] = 32'b11111111111111110010100110101111;
assign LUT_2[20758] = 32'b11111111111111111100100111010010;
assign LUT_2[20759] = 32'b11111111111111111001011111101011;
assign LUT_2[20760] = 32'b11111111111111110100000010001011;
assign LUT_2[20761] = 32'b11111111111111110000111010100100;
assign LUT_2[20762] = 32'b11111111111111111010111011000111;
assign LUT_2[20763] = 32'b11111111111111110111110011100000;
assign LUT_2[20764] = 32'b11111111111111110000011111110011;
assign LUT_2[20765] = 32'b11111111111111101101011000001100;
assign LUT_2[20766] = 32'b11111111111111110111011000101111;
assign LUT_2[20767] = 32'b11111111111111110100010001001000;
assign LUT_2[20768] = 32'b11111111111111111111001000001101;
assign LUT_2[20769] = 32'b11111111111111111100000000100110;
assign LUT_2[20770] = 32'b00000000000000000110000001001001;
assign LUT_2[20771] = 32'b00000000000000000010111001100010;
assign LUT_2[20772] = 32'b11111111111111111011100101110101;
assign LUT_2[20773] = 32'b11111111111111111000011110001110;
assign LUT_2[20774] = 32'b00000000000000000010011110110001;
assign LUT_2[20775] = 32'b11111111111111111111010111001010;
assign LUT_2[20776] = 32'b11111111111111111001111001101010;
assign LUT_2[20777] = 32'b11111111111111110110110010000011;
assign LUT_2[20778] = 32'b00000000000000000000110010100110;
assign LUT_2[20779] = 32'b11111111111111111101101010111111;
assign LUT_2[20780] = 32'b11111111111111110110010111010010;
assign LUT_2[20781] = 32'b11111111111111110011001111101011;
assign LUT_2[20782] = 32'b11111111111111111101010000001110;
assign LUT_2[20783] = 32'b11111111111111111010001000100111;
assign LUT_2[20784] = 32'b11111111111111111001101100010111;
assign LUT_2[20785] = 32'b11111111111111110110100100110000;
assign LUT_2[20786] = 32'b00000000000000000000100101010011;
assign LUT_2[20787] = 32'b11111111111111111101011101101100;
assign LUT_2[20788] = 32'b11111111111111110110001001111111;
assign LUT_2[20789] = 32'b11111111111111110011000010011000;
assign LUT_2[20790] = 32'b11111111111111111101000010111011;
assign LUT_2[20791] = 32'b11111111111111111001111011010100;
assign LUT_2[20792] = 32'b11111111111111110100011101110100;
assign LUT_2[20793] = 32'b11111111111111110001010110001101;
assign LUT_2[20794] = 32'b11111111111111111011010110110000;
assign LUT_2[20795] = 32'b11111111111111111000001111001001;
assign LUT_2[20796] = 32'b11111111111111110000111011011100;
assign LUT_2[20797] = 32'b11111111111111101101110011110101;
assign LUT_2[20798] = 32'b11111111111111110111110100011000;
assign LUT_2[20799] = 32'b11111111111111110100101100110001;
assign LUT_2[20800] = 32'b11111111111111110110110101000111;
assign LUT_2[20801] = 32'b11111111111111110011101101100000;
assign LUT_2[20802] = 32'b11111111111111111101101110000011;
assign LUT_2[20803] = 32'b11111111111111111010100110011100;
assign LUT_2[20804] = 32'b11111111111111110011010010101111;
assign LUT_2[20805] = 32'b11111111111111110000001011001000;
assign LUT_2[20806] = 32'b11111111111111111010001011101011;
assign LUT_2[20807] = 32'b11111111111111110111000100000100;
assign LUT_2[20808] = 32'b11111111111111110001100110100100;
assign LUT_2[20809] = 32'b11111111111111101110011110111101;
assign LUT_2[20810] = 32'b11111111111111111000011111100000;
assign LUT_2[20811] = 32'b11111111111111110101010111111001;
assign LUT_2[20812] = 32'b11111111111111101110000100001100;
assign LUT_2[20813] = 32'b11111111111111101010111100100101;
assign LUT_2[20814] = 32'b11111111111111110100111101001000;
assign LUT_2[20815] = 32'b11111111111111110001110101100001;
assign LUT_2[20816] = 32'b11111111111111110001011001010001;
assign LUT_2[20817] = 32'b11111111111111101110010001101010;
assign LUT_2[20818] = 32'b11111111111111111000010010001101;
assign LUT_2[20819] = 32'b11111111111111110101001010100110;
assign LUT_2[20820] = 32'b11111111111111101101110110111001;
assign LUT_2[20821] = 32'b11111111111111101010101111010010;
assign LUT_2[20822] = 32'b11111111111111110100101111110101;
assign LUT_2[20823] = 32'b11111111111111110001101000001110;
assign LUT_2[20824] = 32'b11111111111111101100001010101110;
assign LUT_2[20825] = 32'b11111111111111101001000011000111;
assign LUT_2[20826] = 32'b11111111111111110011000011101010;
assign LUT_2[20827] = 32'b11111111111111101111111100000011;
assign LUT_2[20828] = 32'b11111111111111101000101000010110;
assign LUT_2[20829] = 32'b11111111111111100101100000101111;
assign LUT_2[20830] = 32'b11111111111111101111100001010010;
assign LUT_2[20831] = 32'b11111111111111101100011001101011;
assign LUT_2[20832] = 32'b11111111111111110111010000110000;
assign LUT_2[20833] = 32'b11111111111111110100001001001001;
assign LUT_2[20834] = 32'b11111111111111111110001001101100;
assign LUT_2[20835] = 32'b11111111111111111011000010000101;
assign LUT_2[20836] = 32'b11111111111111110011101110011000;
assign LUT_2[20837] = 32'b11111111111111110000100110110001;
assign LUT_2[20838] = 32'b11111111111111111010100111010100;
assign LUT_2[20839] = 32'b11111111111111110111011111101101;
assign LUT_2[20840] = 32'b11111111111111110010000010001101;
assign LUT_2[20841] = 32'b11111111111111101110111010100110;
assign LUT_2[20842] = 32'b11111111111111111000111011001001;
assign LUT_2[20843] = 32'b11111111111111110101110011100010;
assign LUT_2[20844] = 32'b11111111111111101110011111110101;
assign LUT_2[20845] = 32'b11111111111111101011011000001110;
assign LUT_2[20846] = 32'b11111111111111110101011000110001;
assign LUT_2[20847] = 32'b11111111111111110010010001001010;
assign LUT_2[20848] = 32'b11111111111111110001110100111010;
assign LUT_2[20849] = 32'b11111111111111101110101101010011;
assign LUT_2[20850] = 32'b11111111111111111000101101110110;
assign LUT_2[20851] = 32'b11111111111111110101100110001111;
assign LUT_2[20852] = 32'b11111111111111101110010010100010;
assign LUT_2[20853] = 32'b11111111111111101011001010111011;
assign LUT_2[20854] = 32'b11111111111111110101001011011110;
assign LUT_2[20855] = 32'b11111111111111110010000011110111;
assign LUT_2[20856] = 32'b11111111111111101100100110010111;
assign LUT_2[20857] = 32'b11111111111111101001011110110000;
assign LUT_2[20858] = 32'b11111111111111110011011111010011;
assign LUT_2[20859] = 32'b11111111111111110000010111101100;
assign LUT_2[20860] = 32'b11111111111111101001000011111111;
assign LUT_2[20861] = 32'b11111111111111100101111100011000;
assign LUT_2[20862] = 32'b11111111111111101111111100111011;
assign LUT_2[20863] = 32'b11111111111111101100110101010100;
assign LUT_2[20864] = 32'b00000000000000000011000000110011;
assign LUT_2[20865] = 32'b11111111111111111111111001001100;
assign LUT_2[20866] = 32'b00000000000000001001111001101111;
assign LUT_2[20867] = 32'b00000000000000000110110010001000;
assign LUT_2[20868] = 32'b11111111111111111111011110011011;
assign LUT_2[20869] = 32'b11111111111111111100010110110100;
assign LUT_2[20870] = 32'b00000000000000000110010111010111;
assign LUT_2[20871] = 32'b00000000000000000011001111110000;
assign LUT_2[20872] = 32'b11111111111111111101110010010000;
assign LUT_2[20873] = 32'b11111111111111111010101010101001;
assign LUT_2[20874] = 32'b00000000000000000100101011001100;
assign LUT_2[20875] = 32'b00000000000000000001100011100101;
assign LUT_2[20876] = 32'b11111111111111111010001111111000;
assign LUT_2[20877] = 32'b11111111111111110111001000010001;
assign LUT_2[20878] = 32'b00000000000000000001001000110100;
assign LUT_2[20879] = 32'b11111111111111111110000001001101;
assign LUT_2[20880] = 32'b11111111111111111101100100111101;
assign LUT_2[20881] = 32'b11111111111111111010011101010110;
assign LUT_2[20882] = 32'b00000000000000000100011101111001;
assign LUT_2[20883] = 32'b00000000000000000001010110010010;
assign LUT_2[20884] = 32'b11111111111111111010000010100101;
assign LUT_2[20885] = 32'b11111111111111110110111010111110;
assign LUT_2[20886] = 32'b00000000000000000000111011100001;
assign LUT_2[20887] = 32'b11111111111111111101110011111010;
assign LUT_2[20888] = 32'b11111111111111111000010110011010;
assign LUT_2[20889] = 32'b11111111111111110101001110110011;
assign LUT_2[20890] = 32'b11111111111111111111001111010110;
assign LUT_2[20891] = 32'b11111111111111111100000111101111;
assign LUT_2[20892] = 32'b11111111111111110100110100000010;
assign LUT_2[20893] = 32'b11111111111111110001101100011011;
assign LUT_2[20894] = 32'b11111111111111111011101100111110;
assign LUT_2[20895] = 32'b11111111111111111000100101010111;
assign LUT_2[20896] = 32'b00000000000000000011011100011100;
assign LUT_2[20897] = 32'b00000000000000000000010100110101;
assign LUT_2[20898] = 32'b00000000000000001010010101011000;
assign LUT_2[20899] = 32'b00000000000000000111001101110001;
assign LUT_2[20900] = 32'b11111111111111111111111010000100;
assign LUT_2[20901] = 32'b11111111111111111100110010011101;
assign LUT_2[20902] = 32'b00000000000000000110110011000000;
assign LUT_2[20903] = 32'b00000000000000000011101011011001;
assign LUT_2[20904] = 32'b11111111111111111110001101111001;
assign LUT_2[20905] = 32'b11111111111111111011000110010010;
assign LUT_2[20906] = 32'b00000000000000000101000110110101;
assign LUT_2[20907] = 32'b00000000000000000001111111001110;
assign LUT_2[20908] = 32'b11111111111111111010101011100001;
assign LUT_2[20909] = 32'b11111111111111110111100011111010;
assign LUT_2[20910] = 32'b00000000000000000001100100011101;
assign LUT_2[20911] = 32'b11111111111111111110011100110110;
assign LUT_2[20912] = 32'b11111111111111111110000000100110;
assign LUT_2[20913] = 32'b11111111111111111010111000111111;
assign LUT_2[20914] = 32'b00000000000000000100111001100010;
assign LUT_2[20915] = 32'b00000000000000000001110001111011;
assign LUT_2[20916] = 32'b11111111111111111010011110001110;
assign LUT_2[20917] = 32'b11111111111111110111010110100111;
assign LUT_2[20918] = 32'b00000000000000000001010111001010;
assign LUT_2[20919] = 32'b11111111111111111110001111100011;
assign LUT_2[20920] = 32'b11111111111111111000110010000011;
assign LUT_2[20921] = 32'b11111111111111110101101010011100;
assign LUT_2[20922] = 32'b11111111111111111111101010111111;
assign LUT_2[20923] = 32'b11111111111111111100100011011000;
assign LUT_2[20924] = 32'b11111111111111110101001111101011;
assign LUT_2[20925] = 32'b11111111111111110010001000000100;
assign LUT_2[20926] = 32'b11111111111111111100001000100111;
assign LUT_2[20927] = 32'b11111111111111111001000001000000;
assign LUT_2[20928] = 32'b11111111111111111011001001010110;
assign LUT_2[20929] = 32'b11111111111111111000000001101111;
assign LUT_2[20930] = 32'b00000000000000000010000010010010;
assign LUT_2[20931] = 32'b11111111111111111110111010101011;
assign LUT_2[20932] = 32'b11111111111111110111100110111110;
assign LUT_2[20933] = 32'b11111111111111110100011111010111;
assign LUT_2[20934] = 32'b11111111111111111110011111111010;
assign LUT_2[20935] = 32'b11111111111111111011011000010011;
assign LUT_2[20936] = 32'b11111111111111110101111010110011;
assign LUT_2[20937] = 32'b11111111111111110010110011001100;
assign LUT_2[20938] = 32'b11111111111111111100110011101111;
assign LUT_2[20939] = 32'b11111111111111111001101100001000;
assign LUT_2[20940] = 32'b11111111111111110010011000011011;
assign LUT_2[20941] = 32'b11111111111111101111010000110100;
assign LUT_2[20942] = 32'b11111111111111111001010001010111;
assign LUT_2[20943] = 32'b11111111111111110110001001110000;
assign LUT_2[20944] = 32'b11111111111111110101101101100000;
assign LUT_2[20945] = 32'b11111111111111110010100101111001;
assign LUT_2[20946] = 32'b11111111111111111100100110011100;
assign LUT_2[20947] = 32'b11111111111111111001011110110101;
assign LUT_2[20948] = 32'b11111111111111110010001011001000;
assign LUT_2[20949] = 32'b11111111111111101111000011100001;
assign LUT_2[20950] = 32'b11111111111111111001000100000100;
assign LUT_2[20951] = 32'b11111111111111110101111100011101;
assign LUT_2[20952] = 32'b11111111111111110000011110111101;
assign LUT_2[20953] = 32'b11111111111111101101010111010110;
assign LUT_2[20954] = 32'b11111111111111110111010111111001;
assign LUT_2[20955] = 32'b11111111111111110100010000010010;
assign LUT_2[20956] = 32'b11111111111111101100111100100101;
assign LUT_2[20957] = 32'b11111111111111101001110100111110;
assign LUT_2[20958] = 32'b11111111111111110011110101100001;
assign LUT_2[20959] = 32'b11111111111111110000101101111010;
assign LUT_2[20960] = 32'b11111111111111111011100100111111;
assign LUT_2[20961] = 32'b11111111111111111000011101011000;
assign LUT_2[20962] = 32'b00000000000000000010011101111011;
assign LUT_2[20963] = 32'b11111111111111111111010110010100;
assign LUT_2[20964] = 32'b11111111111111111000000010100111;
assign LUT_2[20965] = 32'b11111111111111110100111011000000;
assign LUT_2[20966] = 32'b11111111111111111110111011100011;
assign LUT_2[20967] = 32'b11111111111111111011110011111100;
assign LUT_2[20968] = 32'b11111111111111110110010110011100;
assign LUT_2[20969] = 32'b11111111111111110011001110110101;
assign LUT_2[20970] = 32'b11111111111111111101001111011000;
assign LUT_2[20971] = 32'b11111111111111111010000111110001;
assign LUT_2[20972] = 32'b11111111111111110010110100000100;
assign LUT_2[20973] = 32'b11111111111111101111101100011101;
assign LUT_2[20974] = 32'b11111111111111111001101101000000;
assign LUT_2[20975] = 32'b11111111111111110110100101011001;
assign LUT_2[20976] = 32'b11111111111111110110001001001001;
assign LUT_2[20977] = 32'b11111111111111110011000001100010;
assign LUT_2[20978] = 32'b11111111111111111101000010000101;
assign LUT_2[20979] = 32'b11111111111111111001111010011110;
assign LUT_2[20980] = 32'b11111111111111110010100110110001;
assign LUT_2[20981] = 32'b11111111111111101111011111001010;
assign LUT_2[20982] = 32'b11111111111111111001011111101101;
assign LUT_2[20983] = 32'b11111111111111110110011000000110;
assign LUT_2[20984] = 32'b11111111111111110000111010100110;
assign LUT_2[20985] = 32'b11111111111111101101110010111111;
assign LUT_2[20986] = 32'b11111111111111110111110011100010;
assign LUT_2[20987] = 32'b11111111111111110100101011111011;
assign LUT_2[20988] = 32'b11111111111111101101011000001110;
assign LUT_2[20989] = 32'b11111111111111101010010000100111;
assign LUT_2[20990] = 32'b11111111111111110100010001001010;
assign LUT_2[20991] = 32'b11111111111111110001001001100011;
assign LUT_2[20992] = 32'b11111111111111111111011111110000;
assign LUT_2[20993] = 32'b11111111111111111100011000001001;
assign LUT_2[20994] = 32'b00000000000000000110011000101100;
assign LUT_2[20995] = 32'b00000000000000000011010001000101;
assign LUT_2[20996] = 32'b11111111111111111011111101011000;
assign LUT_2[20997] = 32'b11111111111111111000110101110001;
assign LUT_2[20998] = 32'b00000000000000000010110110010100;
assign LUT_2[20999] = 32'b11111111111111111111101110101101;
assign LUT_2[21000] = 32'b11111111111111111010010001001101;
assign LUT_2[21001] = 32'b11111111111111110111001001100110;
assign LUT_2[21002] = 32'b00000000000000000001001010001001;
assign LUT_2[21003] = 32'b11111111111111111110000010100010;
assign LUT_2[21004] = 32'b11111111111111110110101110110101;
assign LUT_2[21005] = 32'b11111111111111110011100111001110;
assign LUT_2[21006] = 32'b11111111111111111101100111110001;
assign LUT_2[21007] = 32'b11111111111111111010100000001010;
assign LUT_2[21008] = 32'b11111111111111111010000011111010;
assign LUT_2[21009] = 32'b11111111111111110110111100010011;
assign LUT_2[21010] = 32'b00000000000000000000111100110110;
assign LUT_2[21011] = 32'b11111111111111111101110101001111;
assign LUT_2[21012] = 32'b11111111111111110110100001100010;
assign LUT_2[21013] = 32'b11111111111111110011011001111011;
assign LUT_2[21014] = 32'b11111111111111111101011010011110;
assign LUT_2[21015] = 32'b11111111111111111010010010110111;
assign LUT_2[21016] = 32'b11111111111111110100110101010111;
assign LUT_2[21017] = 32'b11111111111111110001101101110000;
assign LUT_2[21018] = 32'b11111111111111111011101110010011;
assign LUT_2[21019] = 32'b11111111111111111000100110101100;
assign LUT_2[21020] = 32'b11111111111111110001010010111111;
assign LUT_2[21021] = 32'b11111111111111101110001011011000;
assign LUT_2[21022] = 32'b11111111111111111000001011111011;
assign LUT_2[21023] = 32'b11111111111111110101000100010100;
assign LUT_2[21024] = 32'b11111111111111111111111011011001;
assign LUT_2[21025] = 32'b11111111111111111100110011110010;
assign LUT_2[21026] = 32'b00000000000000000110110100010101;
assign LUT_2[21027] = 32'b00000000000000000011101100101110;
assign LUT_2[21028] = 32'b11111111111111111100011001000001;
assign LUT_2[21029] = 32'b11111111111111111001010001011010;
assign LUT_2[21030] = 32'b00000000000000000011010001111101;
assign LUT_2[21031] = 32'b00000000000000000000001010010110;
assign LUT_2[21032] = 32'b11111111111111111010101100110110;
assign LUT_2[21033] = 32'b11111111111111110111100101001111;
assign LUT_2[21034] = 32'b00000000000000000001100101110010;
assign LUT_2[21035] = 32'b11111111111111111110011110001011;
assign LUT_2[21036] = 32'b11111111111111110111001010011110;
assign LUT_2[21037] = 32'b11111111111111110100000010110111;
assign LUT_2[21038] = 32'b11111111111111111110000011011010;
assign LUT_2[21039] = 32'b11111111111111111010111011110011;
assign LUT_2[21040] = 32'b11111111111111111010011111100011;
assign LUT_2[21041] = 32'b11111111111111110111010111111100;
assign LUT_2[21042] = 32'b00000000000000000001011000011111;
assign LUT_2[21043] = 32'b11111111111111111110010000111000;
assign LUT_2[21044] = 32'b11111111111111110110111101001011;
assign LUT_2[21045] = 32'b11111111111111110011110101100100;
assign LUT_2[21046] = 32'b11111111111111111101110110000111;
assign LUT_2[21047] = 32'b11111111111111111010101110100000;
assign LUT_2[21048] = 32'b11111111111111110101010001000000;
assign LUT_2[21049] = 32'b11111111111111110010001001011001;
assign LUT_2[21050] = 32'b11111111111111111100001001111100;
assign LUT_2[21051] = 32'b11111111111111111001000010010101;
assign LUT_2[21052] = 32'b11111111111111110001101110101000;
assign LUT_2[21053] = 32'b11111111111111101110100111000001;
assign LUT_2[21054] = 32'b11111111111111111000100111100100;
assign LUT_2[21055] = 32'b11111111111111110101011111111101;
assign LUT_2[21056] = 32'b11111111111111110111101000010011;
assign LUT_2[21057] = 32'b11111111111111110100100000101100;
assign LUT_2[21058] = 32'b11111111111111111110100001001111;
assign LUT_2[21059] = 32'b11111111111111111011011001101000;
assign LUT_2[21060] = 32'b11111111111111110100000101111011;
assign LUT_2[21061] = 32'b11111111111111110000111110010100;
assign LUT_2[21062] = 32'b11111111111111111010111110110111;
assign LUT_2[21063] = 32'b11111111111111110111110111010000;
assign LUT_2[21064] = 32'b11111111111111110010011001110000;
assign LUT_2[21065] = 32'b11111111111111101111010010001001;
assign LUT_2[21066] = 32'b11111111111111111001010010101100;
assign LUT_2[21067] = 32'b11111111111111110110001011000101;
assign LUT_2[21068] = 32'b11111111111111101110110111011000;
assign LUT_2[21069] = 32'b11111111111111101011101111110001;
assign LUT_2[21070] = 32'b11111111111111110101110000010100;
assign LUT_2[21071] = 32'b11111111111111110010101000101101;
assign LUT_2[21072] = 32'b11111111111111110010001100011101;
assign LUT_2[21073] = 32'b11111111111111101111000100110110;
assign LUT_2[21074] = 32'b11111111111111111001000101011001;
assign LUT_2[21075] = 32'b11111111111111110101111101110010;
assign LUT_2[21076] = 32'b11111111111111101110101010000101;
assign LUT_2[21077] = 32'b11111111111111101011100010011110;
assign LUT_2[21078] = 32'b11111111111111110101100011000001;
assign LUT_2[21079] = 32'b11111111111111110010011011011010;
assign LUT_2[21080] = 32'b11111111111111101100111101111010;
assign LUT_2[21081] = 32'b11111111111111101001110110010011;
assign LUT_2[21082] = 32'b11111111111111110011110110110110;
assign LUT_2[21083] = 32'b11111111111111110000101111001111;
assign LUT_2[21084] = 32'b11111111111111101001011011100010;
assign LUT_2[21085] = 32'b11111111111111100110010011111011;
assign LUT_2[21086] = 32'b11111111111111110000010100011110;
assign LUT_2[21087] = 32'b11111111111111101101001100110111;
assign LUT_2[21088] = 32'b11111111111111111000000011111100;
assign LUT_2[21089] = 32'b11111111111111110100111100010101;
assign LUT_2[21090] = 32'b11111111111111111110111100111000;
assign LUT_2[21091] = 32'b11111111111111111011110101010001;
assign LUT_2[21092] = 32'b11111111111111110100100001100100;
assign LUT_2[21093] = 32'b11111111111111110001011001111101;
assign LUT_2[21094] = 32'b11111111111111111011011010100000;
assign LUT_2[21095] = 32'b11111111111111111000010010111001;
assign LUT_2[21096] = 32'b11111111111111110010110101011001;
assign LUT_2[21097] = 32'b11111111111111101111101101110010;
assign LUT_2[21098] = 32'b11111111111111111001101110010101;
assign LUT_2[21099] = 32'b11111111111111110110100110101110;
assign LUT_2[21100] = 32'b11111111111111101111010011000001;
assign LUT_2[21101] = 32'b11111111111111101100001011011010;
assign LUT_2[21102] = 32'b11111111111111110110001011111101;
assign LUT_2[21103] = 32'b11111111111111110011000100010110;
assign LUT_2[21104] = 32'b11111111111111110010101000000110;
assign LUT_2[21105] = 32'b11111111111111101111100000011111;
assign LUT_2[21106] = 32'b11111111111111111001100001000010;
assign LUT_2[21107] = 32'b11111111111111110110011001011011;
assign LUT_2[21108] = 32'b11111111111111101111000101101110;
assign LUT_2[21109] = 32'b11111111111111101011111110000111;
assign LUT_2[21110] = 32'b11111111111111110101111110101010;
assign LUT_2[21111] = 32'b11111111111111110010110111000011;
assign LUT_2[21112] = 32'b11111111111111101101011001100011;
assign LUT_2[21113] = 32'b11111111111111101010010001111100;
assign LUT_2[21114] = 32'b11111111111111110100010010011111;
assign LUT_2[21115] = 32'b11111111111111110001001010111000;
assign LUT_2[21116] = 32'b11111111111111101001110111001011;
assign LUT_2[21117] = 32'b11111111111111100110101111100100;
assign LUT_2[21118] = 32'b11111111111111110000110000000111;
assign LUT_2[21119] = 32'b11111111111111101101101000100000;
assign LUT_2[21120] = 32'b00000000000000000011110011111111;
assign LUT_2[21121] = 32'b00000000000000000000101100011000;
assign LUT_2[21122] = 32'b00000000000000001010101100111011;
assign LUT_2[21123] = 32'b00000000000000000111100101010100;
assign LUT_2[21124] = 32'b00000000000000000000010001100111;
assign LUT_2[21125] = 32'b11111111111111111101001010000000;
assign LUT_2[21126] = 32'b00000000000000000111001010100011;
assign LUT_2[21127] = 32'b00000000000000000100000010111100;
assign LUT_2[21128] = 32'b11111111111111111110100101011100;
assign LUT_2[21129] = 32'b11111111111111111011011101110101;
assign LUT_2[21130] = 32'b00000000000000000101011110011000;
assign LUT_2[21131] = 32'b00000000000000000010010110110001;
assign LUT_2[21132] = 32'b11111111111111111011000011000100;
assign LUT_2[21133] = 32'b11111111111111110111111011011101;
assign LUT_2[21134] = 32'b00000000000000000001111100000000;
assign LUT_2[21135] = 32'b11111111111111111110110100011001;
assign LUT_2[21136] = 32'b11111111111111111110011000001001;
assign LUT_2[21137] = 32'b11111111111111111011010000100010;
assign LUT_2[21138] = 32'b00000000000000000101010001000101;
assign LUT_2[21139] = 32'b00000000000000000010001001011110;
assign LUT_2[21140] = 32'b11111111111111111010110101110001;
assign LUT_2[21141] = 32'b11111111111111110111101110001010;
assign LUT_2[21142] = 32'b00000000000000000001101110101101;
assign LUT_2[21143] = 32'b11111111111111111110100111000110;
assign LUT_2[21144] = 32'b11111111111111111001001001100110;
assign LUT_2[21145] = 32'b11111111111111110110000001111111;
assign LUT_2[21146] = 32'b00000000000000000000000010100010;
assign LUT_2[21147] = 32'b11111111111111111100111010111011;
assign LUT_2[21148] = 32'b11111111111111110101100111001110;
assign LUT_2[21149] = 32'b11111111111111110010011111100111;
assign LUT_2[21150] = 32'b11111111111111111100100000001010;
assign LUT_2[21151] = 32'b11111111111111111001011000100011;
assign LUT_2[21152] = 32'b00000000000000000100001111101000;
assign LUT_2[21153] = 32'b00000000000000000001001000000001;
assign LUT_2[21154] = 32'b00000000000000001011001000100100;
assign LUT_2[21155] = 32'b00000000000000001000000000111101;
assign LUT_2[21156] = 32'b00000000000000000000101101010000;
assign LUT_2[21157] = 32'b11111111111111111101100101101001;
assign LUT_2[21158] = 32'b00000000000000000111100110001100;
assign LUT_2[21159] = 32'b00000000000000000100011110100101;
assign LUT_2[21160] = 32'b11111111111111111111000001000101;
assign LUT_2[21161] = 32'b11111111111111111011111001011110;
assign LUT_2[21162] = 32'b00000000000000000101111010000001;
assign LUT_2[21163] = 32'b00000000000000000010110010011010;
assign LUT_2[21164] = 32'b11111111111111111011011110101101;
assign LUT_2[21165] = 32'b11111111111111111000010111000110;
assign LUT_2[21166] = 32'b00000000000000000010010111101001;
assign LUT_2[21167] = 32'b11111111111111111111010000000010;
assign LUT_2[21168] = 32'b11111111111111111110110011110010;
assign LUT_2[21169] = 32'b11111111111111111011101100001011;
assign LUT_2[21170] = 32'b00000000000000000101101100101110;
assign LUT_2[21171] = 32'b00000000000000000010100101000111;
assign LUT_2[21172] = 32'b11111111111111111011010001011010;
assign LUT_2[21173] = 32'b11111111111111111000001001110011;
assign LUT_2[21174] = 32'b00000000000000000010001010010110;
assign LUT_2[21175] = 32'b11111111111111111111000010101111;
assign LUT_2[21176] = 32'b11111111111111111001100101001111;
assign LUT_2[21177] = 32'b11111111111111110110011101101000;
assign LUT_2[21178] = 32'b00000000000000000000011110001011;
assign LUT_2[21179] = 32'b11111111111111111101010110100100;
assign LUT_2[21180] = 32'b11111111111111110110000010110111;
assign LUT_2[21181] = 32'b11111111111111110010111011010000;
assign LUT_2[21182] = 32'b11111111111111111100111011110011;
assign LUT_2[21183] = 32'b11111111111111111001110100001100;
assign LUT_2[21184] = 32'b11111111111111111011111100100010;
assign LUT_2[21185] = 32'b11111111111111111000110100111011;
assign LUT_2[21186] = 32'b00000000000000000010110101011110;
assign LUT_2[21187] = 32'b11111111111111111111101101110111;
assign LUT_2[21188] = 32'b11111111111111111000011010001010;
assign LUT_2[21189] = 32'b11111111111111110101010010100011;
assign LUT_2[21190] = 32'b11111111111111111111010011000110;
assign LUT_2[21191] = 32'b11111111111111111100001011011111;
assign LUT_2[21192] = 32'b11111111111111110110101101111111;
assign LUT_2[21193] = 32'b11111111111111110011100110011000;
assign LUT_2[21194] = 32'b11111111111111111101100110111011;
assign LUT_2[21195] = 32'b11111111111111111010011111010100;
assign LUT_2[21196] = 32'b11111111111111110011001011100111;
assign LUT_2[21197] = 32'b11111111111111110000000100000000;
assign LUT_2[21198] = 32'b11111111111111111010000100100011;
assign LUT_2[21199] = 32'b11111111111111110110111100111100;
assign LUT_2[21200] = 32'b11111111111111110110100000101100;
assign LUT_2[21201] = 32'b11111111111111110011011001000101;
assign LUT_2[21202] = 32'b11111111111111111101011001101000;
assign LUT_2[21203] = 32'b11111111111111111010010010000001;
assign LUT_2[21204] = 32'b11111111111111110010111110010100;
assign LUT_2[21205] = 32'b11111111111111101111110110101101;
assign LUT_2[21206] = 32'b11111111111111111001110111010000;
assign LUT_2[21207] = 32'b11111111111111110110101111101001;
assign LUT_2[21208] = 32'b11111111111111110001010010001001;
assign LUT_2[21209] = 32'b11111111111111101110001010100010;
assign LUT_2[21210] = 32'b11111111111111111000001011000101;
assign LUT_2[21211] = 32'b11111111111111110101000011011110;
assign LUT_2[21212] = 32'b11111111111111101101101111110001;
assign LUT_2[21213] = 32'b11111111111111101010101000001010;
assign LUT_2[21214] = 32'b11111111111111110100101000101101;
assign LUT_2[21215] = 32'b11111111111111110001100001000110;
assign LUT_2[21216] = 32'b11111111111111111100011000001011;
assign LUT_2[21217] = 32'b11111111111111111001010000100100;
assign LUT_2[21218] = 32'b00000000000000000011010001000111;
assign LUT_2[21219] = 32'b00000000000000000000001001100000;
assign LUT_2[21220] = 32'b11111111111111111000110101110011;
assign LUT_2[21221] = 32'b11111111111111110101101110001100;
assign LUT_2[21222] = 32'b11111111111111111111101110101111;
assign LUT_2[21223] = 32'b11111111111111111100100111001000;
assign LUT_2[21224] = 32'b11111111111111110111001001101000;
assign LUT_2[21225] = 32'b11111111111111110100000010000001;
assign LUT_2[21226] = 32'b11111111111111111110000010100100;
assign LUT_2[21227] = 32'b11111111111111111010111010111101;
assign LUT_2[21228] = 32'b11111111111111110011100111010000;
assign LUT_2[21229] = 32'b11111111111111110000011111101001;
assign LUT_2[21230] = 32'b11111111111111111010100000001100;
assign LUT_2[21231] = 32'b11111111111111110111011000100101;
assign LUT_2[21232] = 32'b11111111111111110110111100010101;
assign LUT_2[21233] = 32'b11111111111111110011110100101110;
assign LUT_2[21234] = 32'b11111111111111111101110101010001;
assign LUT_2[21235] = 32'b11111111111111111010101101101010;
assign LUT_2[21236] = 32'b11111111111111110011011001111101;
assign LUT_2[21237] = 32'b11111111111111110000010010010110;
assign LUT_2[21238] = 32'b11111111111111111010010010111001;
assign LUT_2[21239] = 32'b11111111111111110111001011010010;
assign LUT_2[21240] = 32'b11111111111111110001101101110010;
assign LUT_2[21241] = 32'b11111111111111101110100110001011;
assign LUT_2[21242] = 32'b11111111111111111000100110101110;
assign LUT_2[21243] = 32'b11111111111111110101011111000111;
assign LUT_2[21244] = 32'b11111111111111101110001011011010;
assign LUT_2[21245] = 32'b11111111111111101011000011110011;
assign LUT_2[21246] = 32'b11111111111111110101000100010110;
assign LUT_2[21247] = 32'b11111111111111110001111100101111;
assign LUT_2[21248] = 32'b00000000000000000011011110010110;
assign LUT_2[21249] = 32'b00000000000000000000010110101111;
assign LUT_2[21250] = 32'b00000000000000001010010111010010;
assign LUT_2[21251] = 32'b00000000000000000111001111101011;
assign LUT_2[21252] = 32'b11111111111111111111111011111110;
assign LUT_2[21253] = 32'b11111111111111111100110100010111;
assign LUT_2[21254] = 32'b00000000000000000110110100111010;
assign LUT_2[21255] = 32'b00000000000000000011101101010011;
assign LUT_2[21256] = 32'b11111111111111111110001111110011;
assign LUT_2[21257] = 32'b11111111111111111011001000001100;
assign LUT_2[21258] = 32'b00000000000000000101001000101111;
assign LUT_2[21259] = 32'b00000000000000000010000001001000;
assign LUT_2[21260] = 32'b11111111111111111010101101011011;
assign LUT_2[21261] = 32'b11111111111111110111100101110100;
assign LUT_2[21262] = 32'b00000000000000000001100110010111;
assign LUT_2[21263] = 32'b11111111111111111110011110110000;
assign LUT_2[21264] = 32'b11111111111111111110000010100000;
assign LUT_2[21265] = 32'b11111111111111111010111010111001;
assign LUT_2[21266] = 32'b00000000000000000100111011011100;
assign LUT_2[21267] = 32'b00000000000000000001110011110101;
assign LUT_2[21268] = 32'b11111111111111111010100000001000;
assign LUT_2[21269] = 32'b11111111111111110111011000100001;
assign LUT_2[21270] = 32'b00000000000000000001011001000100;
assign LUT_2[21271] = 32'b11111111111111111110010001011101;
assign LUT_2[21272] = 32'b11111111111111111000110011111101;
assign LUT_2[21273] = 32'b11111111111111110101101100010110;
assign LUT_2[21274] = 32'b11111111111111111111101100111001;
assign LUT_2[21275] = 32'b11111111111111111100100101010010;
assign LUT_2[21276] = 32'b11111111111111110101010001100101;
assign LUT_2[21277] = 32'b11111111111111110010001001111110;
assign LUT_2[21278] = 32'b11111111111111111100001010100001;
assign LUT_2[21279] = 32'b11111111111111111001000010111010;
assign LUT_2[21280] = 32'b00000000000000000011111001111111;
assign LUT_2[21281] = 32'b00000000000000000000110010011000;
assign LUT_2[21282] = 32'b00000000000000001010110010111011;
assign LUT_2[21283] = 32'b00000000000000000111101011010100;
assign LUT_2[21284] = 32'b00000000000000000000010111100111;
assign LUT_2[21285] = 32'b11111111111111111101010000000000;
assign LUT_2[21286] = 32'b00000000000000000111010000100011;
assign LUT_2[21287] = 32'b00000000000000000100001000111100;
assign LUT_2[21288] = 32'b11111111111111111110101011011100;
assign LUT_2[21289] = 32'b11111111111111111011100011110101;
assign LUT_2[21290] = 32'b00000000000000000101100100011000;
assign LUT_2[21291] = 32'b00000000000000000010011100110001;
assign LUT_2[21292] = 32'b11111111111111111011001001000100;
assign LUT_2[21293] = 32'b11111111111111111000000001011101;
assign LUT_2[21294] = 32'b00000000000000000010000010000000;
assign LUT_2[21295] = 32'b11111111111111111110111010011001;
assign LUT_2[21296] = 32'b11111111111111111110011110001001;
assign LUT_2[21297] = 32'b11111111111111111011010110100010;
assign LUT_2[21298] = 32'b00000000000000000101010111000101;
assign LUT_2[21299] = 32'b00000000000000000010001111011110;
assign LUT_2[21300] = 32'b11111111111111111010111011110001;
assign LUT_2[21301] = 32'b11111111111111110111110100001010;
assign LUT_2[21302] = 32'b00000000000000000001110100101101;
assign LUT_2[21303] = 32'b11111111111111111110101101000110;
assign LUT_2[21304] = 32'b11111111111111111001001111100110;
assign LUT_2[21305] = 32'b11111111111111110110000111111111;
assign LUT_2[21306] = 32'b00000000000000000000001000100010;
assign LUT_2[21307] = 32'b11111111111111111101000000111011;
assign LUT_2[21308] = 32'b11111111111111110101101101001110;
assign LUT_2[21309] = 32'b11111111111111110010100101100111;
assign LUT_2[21310] = 32'b11111111111111111100100110001010;
assign LUT_2[21311] = 32'b11111111111111111001011110100011;
assign LUT_2[21312] = 32'b11111111111111111011100110111001;
assign LUT_2[21313] = 32'b11111111111111111000011111010010;
assign LUT_2[21314] = 32'b00000000000000000010011111110101;
assign LUT_2[21315] = 32'b11111111111111111111011000001110;
assign LUT_2[21316] = 32'b11111111111111111000000100100001;
assign LUT_2[21317] = 32'b11111111111111110100111100111010;
assign LUT_2[21318] = 32'b11111111111111111110111101011101;
assign LUT_2[21319] = 32'b11111111111111111011110101110110;
assign LUT_2[21320] = 32'b11111111111111110110011000010110;
assign LUT_2[21321] = 32'b11111111111111110011010000101111;
assign LUT_2[21322] = 32'b11111111111111111101010001010010;
assign LUT_2[21323] = 32'b11111111111111111010001001101011;
assign LUT_2[21324] = 32'b11111111111111110010110101111110;
assign LUT_2[21325] = 32'b11111111111111101111101110010111;
assign LUT_2[21326] = 32'b11111111111111111001101110111010;
assign LUT_2[21327] = 32'b11111111111111110110100111010011;
assign LUT_2[21328] = 32'b11111111111111110110001011000011;
assign LUT_2[21329] = 32'b11111111111111110011000011011100;
assign LUT_2[21330] = 32'b11111111111111111101000011111111;
assign LUT_2[21331] = 32'b11111111111111111001111100011000;
assign LUT_2[21332] = 32'b11111111111111110010101000101011;
assign LUT_2[21333] = 32'b11111111111111101111100001000100;
assign LUT_2[21334] = 32'b11111111111111111001100001100111;
assign LUT_2[21335] = 32'b11111111111111110110011010000000;
assign LUT_2[21336] = 32'b11111111111111110000111100100000;
assign LUT_2[21337] = 32'b11111111111111101101110100111001;
assign LUT_2[21338] = 32'b11111111111111110111110101011100;
assign LUT_2[21339] = 32'b11111111111111110100101101110101;
assign LUT_2[21340] = 32'b11111111111111101101011010001000;
assign LUT_2[21341] = 32'b11111111111111101010010010100001;
assign LUT_2[21342] = 32'b11111111111111110100010011000100;
assign LUT_2[21343] = 32'b11111111111111110001001011011101;
assign LUT_2[21344] = 32'b11111111111111111100000010100010;
assign LUT_2[21345] = 32'b11111111111111111000111010111011;
assign LUT_2[21346] = 32'b00000000000000000010111011011110;
assign LUT_2[21347] = 32'b11111111111111111111110011110111;
assign LUT_2[21348] = 32'b11111111111111111000100000001010;
assign LUT_2[21349] = 32'b11111111111111110101011000100011;
assign LUT_2[21350] = 32'b11111111111111111111011001000110;
assign LUT_2[21351] = 32'b11111111111111111100010001011111;
assign LUT_2[21352] = 32'b11111111111111110110110011111111;
assign LUT_2[21353] = 32'b11111111111111110011101100011000;
assign LUT_2[21354] = 32'b11111111111111111101101100111011;
assign LUT_2[21355] = 32'b11111111111111111010100101010100;
assign LUT_2[21356] = 32'b11111111111111110011010001100111;
assign LUT_2[21357] = 32'b11111111111111110000001010000000;
assign LUT_2[21358] = 32'b11111111111111111010001010100011;
assign LUT_2[21359] = 32'b11111111111111110111000010111100;
assign LUT_2[21360] = 32'b11111111111111110110100110101100;
assign LUT_2[21361] = 32'b11111111111111110011011111000101;
assign LUT_2[21362] = 32'b11111111111111111101011111101000;
assign LUT_2[21363] = 32'b11111111111111111010011000000001;
assign LUT_2[21364] = 32'b11111111111111110011000100010100;
assign LUT_2[21365] = 32'b11111111111111101111111100101101;
assign LUT_2[21366] = 32'b11111111111111111001111101010000;
assign LUT_2[21367] = 32'b11111111111111110110110101101001;
assign LUT_2[21368] = 32'b11111111111111110001011000001001;
assign LUT_2[21369] = 32'b11111111111111101110010000100010;
assign LUT_2[21370] = 32'b11111111111111111000010001000101;
assign LUT_2[21371] = 32'b11111111111111110101001001011110;
assign LUT_2[21372] = 32'b11111111111111101101110101110001;
assign LUT_2[21373] = 32'b11111111111111101010101110001010;
assign LUT_2[21374] = 32'b11111111111111110100101110101101;
assign LUT_2[21375] = 32'b11111111111111110001100111000110;
assign LUT_2[21376] = 32'b00000000000000000111110010100101;
assign LUT_2[21377] = 32'b00000000000000000100101010111110;
assign LUT_2[21378] = 32'b00000000000000001110101011100001;
assign LUT_2[21379] = 32'b00000000000000001011100011111010;
assign LUT_2[21380] = 32'b00000000000000000100010000001101;
assign LUT_2[21381] = 32'b00000000000000000001001000100110;
assign LUT_2[21382] = 32'b00000000000000001011001001001001;
assign LUT_2[21383] = 32'b00000000000000001000000001100010;
assign LUT_2[21384] = 32'b00000000000000000010100100000010;
assign LUT_2[21385] = 32'b11111111111111111111011100011011;
assign LUT_2[21386] = 32'b00000000000000001001011100111110;
assign LUT_2[21387] = 32'b00000000000000000110010101010111;
assign LUT_2[21388] = 32'b11111111111111111111000001101010;
assign LUT_2[21389] = 32'b11111111111111111011111010000011;
assign LUT_2[21390] = 32'b00000000000000000101111010100110;
assign LUT_2[21391] = 32'b00000000000000000010110010111111;
assign LUT_2[21392] = 32'b00000000000000000010010110101111;
assign LUT_2[21393] = 32'b11111111111111111111001111001000;
assign LUT_2[21394] = 32'b00000000000000001001001111101011;
assign LUT_2[21395] = 32'b00000000000000000110001000000100;
assign LUT_2[21396] = 32'b11111111111111111110110100010111;
assign LUT_2[21397] = 32'b11111111111111111011101100110000;
assign LUT_2[21398] = 32'b00000000000000000101101101010011;
assign LUT_2[21399] = 32'b00000000000000000010100101101100;
assign LUT_2[21400] = 32'b11111111111111111101001000001100;
assign LUT_2[21401] = 32'b11111111111111111010000000100101;
assign LUT_2[21402] = 32'b00000000000000000100000001001000;
assign LUT_2[21403] = 32'b00000000000000000000111001100001;
assign LUT_2[21404] = 32'b11111111111111111001100101110100;
assign LUT_2[21405] = 32'b11111111111111110110011110001101;
assign LUT_2[21406] = 32'b00000000000000000000011110110000;
assign LUT_2[21407] = 32'b11111111111111111101010111001001;
assign LUT_2[21408] = 32'b00000000000000001000001110001110;
assign LUT_2[21409] = 32'b00000000000000000101000110100111;
assign LUT_2[21410] = 32'b00000000000000001111000111001010;
assign LUT_2[21411] = 32'b00000000000000001011111111100011;
assign LUT_2[21412] = 32'b00000000000000000100101011110110;
assign LUT_2[21413] = 32'b00000000000000000001100100001111;
assign LUT_2[21414] = 32'b00000000000000001011100100110010;
assign LUT_2[21415] = 32'b00000000000000001000011101001011;
assign LUT_2[21416] = 32'b00000000000000000010111111101011;
assign LUT_2[21417] = 32'b11111111111111111111111000000100;
assign LUT_2[21418] = 32'b00000000000000001001111000100111;
assign LUT_2[21419] = 32'b00000000000000000110110001000000;
assign LUT_2[21420] = 32'b11111111111111111111011101010011;
assign LUT_2[21421] = 32'b11111111111111111100010101101100;
assign LUT_2[21422] = 32'b00000000000000000110010110001111;
assign LUT_2[21423] = 32'b00000000000000000011001110101000;
assign LUT_2[21424] = 32'b00000000000000000010110010011000;
assign LUT_2[21425] = 32'b11111111111111111111101010110001;
assign LUT_2[21426] = 32'b00000000000000001001101011010100;
assign LUT_2[21427] = 32'b00000000000000000110100011101101;
assign LUT_2[21428] = 32'b11111111111111111111010000000000;
assign LUT_2[21429] = 32'b11111111111111111100001000011001;
assign LUT_2[21430] = 32'b00000000000000000110001000111100;
assign LUT_2[21431] = 32'b00000000000000000011000001010101;
assign LUT_2[21432] = 32'b11111111111111111101100011110101;
assign LUT_2[21433] = 32'b11111111111111111010011100001110;
assign LUT_2[21434] = 32'b00000000000000000100011100110001;
assign LUT_2[21435] = 32'b00000000000000000001010101001010;
assign LUT_2[21436] = 32'b11111111111111111010000001011101;
assign LUT_2[21437] = 32'b11111111111111110110111001110110;
assign LUT_2[21438] = 32'b00000000000000000000111010011001;
assign LUT_2[21439] = 32'b11111111111111111101110010110010;
assign LUT_2[21440] = 32'b11111111111111111111111011001000;
assign LUT_2[21441] = 32'b11111111111111111100110011100001;
assign LUT_2[21442] = 32'b00000000000000000110110100000100;
assign LUT_2[21443] = 32'b00000000000000000011101100011101;
assign LUT_2[21444] = 32'b11111111111111111100011000110000;
assign LUT_2[21445] = 32'b11111111111111111001010001001001;
assign LUT_2[21446] = 32'b00000000000000000011010001101100;
assign LUT_2[21447] = 32'b00000000000000000000001010000101;
assign LUT_2[21448] = 32'b11111111111111111010101100100101;
assign LUT_2[21449] = 32'b11111111111111110111100100111110;
assign LUT_2[21450] = 32'b00000000000000000001100101100001;
assign LUT_2[21451] = 32'b11111111111111111110011101111010;
assign LUT_2[21452] = 32'b11111111111111110111001010001101;
assign LUT_2[21453] = 32'b11111111111111110100000010100110;
assign LUT_2[21454] = 32'b11111111111111111110000011001001;
assign LUT_2[21455] = 32'b11111111111111111010111011100010;
assign LUT_2[21456] = 32'b11111111111111111010011111010010;
assign LUT_2[21457] = 32'b11111111111111110111010111101011;
assign LUT_2[21458] = 32'b00000000000000000001011000001110;
assign LUT_2[21459] = 32'b11111111111111111110010000100111;
assign LUT_2[21460] = 32'b11111111111111110110111100111010;
assign LUT_2[21461] = 32'b11111111111111110011110101010011;
assign LUT_2[21462] = 32'b11111111111111111101110101110110;
assign LUT_2[21463] = 32'b11111111111111111010101110001111;
assign LUT_2[21464] = 32'b11111111111111110101010000101111;
assign LUT_2[21465] = 32'b11111111111111110010001001001000;
assign LUT_2[21466] = 32'b11111111111111111100001001101011;
assign LUT_2[21467] = 32'b11111111111111111001000010000100;
assign LUT_2[21468] = 32'b11111111111111110001101110010111;
assign LUT_2[21469] = 32'b11111111111111101110100110110000;
assign LUT_2[21470] = 32'b11111111111111111000100111010011;
assign LUT_2[21471] = 32'b11111111111111110101011111101100;
assign LUT_2[21472] = 32'b00000000000000000000010110110001;
assign LUT_2[21473] = 32'b11111111111111111101001111001010;
assign LUT_2[21474] = 32'b00000000000000000111001111101101;
assign LUT_2[21475] = 32'b00000000000000000100001000000110;
assign LUT_2[21476] = 32'b11111111111111111100110100011001;
assign LUT_2[21477] = 32'b11111111111111111001101100110010;
assign LUT_2[21478] = 32'b00000000000000000011101101010101;
assign LUT_2[21479] = 32'b00000000000000000000100101101110;
assign LUT_2[21480] = 32'b11111111111111111011001000001110;
assign LUT_2[21481] = 32'b11111111111111111000000000100111;
assign LUT_2[21482] = 32'b00000000000000000010000001001010;
assign LUT_2[21483] = 32'b11111111111111111110111001100011;
assign LUT_2[21484] = 32'b11111111111111110111100101110110;
assign LUT_2[21485] = 32'b11111111111111110100011110001111;
assign LUT_2[21486] = 32'b11111111111111111110011110110010;
assign LUT_2[21487] = 32'b11111111111111111011010111001011;
assign LUT_2[21488] = 32'b11111111111111111010111010111011;
assign LUT_2[21489] = 32'b11111111111111110111110011010100;
assign LUT_2[21490] = 32'b00000000000000000001110011110111;
assign LUT_2[21491] = 32'b11111111111111111110101100010000;
assign LUT_2[21492] = 32'b11111111111111110111011000100011;
assign LUT_2[21493] = 32'b11111111111111110100010000111100;
assign LUT_2[21494] = 32'b11111111111111111110010001011111;
assign LUT_2[21495] = 32'b11111111111111111011001001111000;
assign LUT_2[21496] = 32'b11111111111111110101101100011000;
assign LUT_2[21497] = 32'b11111111111111110010100100110001;
assign LUT_2[21498] = 32'b11111111111111111100100101010100;
assign LUT_2[21499] = 32'b11111111111111111001011101101101;
assign LUT_2[21500] = 32'b11111111111111110010001010000000;
assign LUT_2[21501] = 32'b11111111111111101111000010011001;
assign LUT_2[21502] = 32'b11111111111111111001000010111100;
assign LUT_2[21503] = 32'b11111111111111110101111011010101;
assign LUT_2[21504] = 32'b00000000000000000001011010000011;
assign LUT_2[21505] = 32'b11111111111111111110010010011100;
assign LUT_2[21506] = 32'b00000000000000001000010010111111;
assign LUT_2[21507] = 32'b00000000000000000101001011011000;
assign LUT_2[21508] = 32'b11111111111111111101110111101011;
assign LUT_2[21509] = 32'b11111111111111111010110000000100;
assign LUT_2[21510] = 32'b00000000000000000100110000100111;
assign LUT_2[21511] = 32'b00000000000000000001101001000000;
assign LUT_2[21512] = 32'b11111111111111111100001011100000;
assign LUT_2[21513] = 32'b11111111111111111001000011111001;
assign LUT_2[21514] = 32'b00000000000000000011000100011100;
assign LUT_2[21515] = 32'b11111111111111111111111100110101;
assign LUT_2[21516] = 32'b11111111111111111000101001001000;
assign LUT_2[21517] = 32'b11111111111111110101100001100001;
assign LUT_2[21518] = 32'b11111111111111111111100010000100;
assign LUT_2[21519] = 32'b11111111111111111100011010011101;
assign LUT_2[21520] = 32'b11111111111111111011111110001101;
assign LUT_2[21521] = 32'b11111111111111111000110110100110;
assign LUT_2[21522] = 32'b00000000000000000010110111001001;
assign LUT_2[21523] = 32'b11111111111111111111101111100010;
assign LUT_2[21524] = 32'b11111111111111111000011011110101;
assign LUT_2[21525] = 32'b11111111111111110101010100001110;
assign LUT_2[21526] = 32'b11111111111111111111010100110001;
assign LUT_2[21527] = 32'b11111111111111111100001101001010;
assign LUT_2[21528] = 32'b11111111111111110110101111101010;
assign LUT_2[21529] = 32'b11111111111111110011101000000011;
assign LUT_2[21530] = 32'b11111111111111111101101000100110;
assign LUT_2[21531] = 32'b11111111111111111010100000111111;
assign LUT_2[21532] = 32'b11111111111111110011001101010010;
assign LUT_2[21533] = 32'b11111111111111110000000101101011;
assign LUT_2[21534] = 32'b11111111111111111010000110001110;
assign LUT_2[21535] = 32'b11111111111111110110111110100111;
assign LUT_2[21536] = 32'b00000000000000000001110101101100;
assign LUT_2[21537] = 32'b11111111111111111110101110000101;
assign LUT_2[21538] = 32'b00000000000000001000101110101000;
assign LUT_2[21539] = 32'b00000000000000000101100111000001;
assign LUT_2[21540] = 32'b11111111111111111110010011010100;
assign LUT_2[21541] = 32'b11111111111111111011001011101101;
assign LUT_2[21542] = 32'b00000000000000000101001100010000;
assign LUT_2[21543] = 32'b00000000000000000010000100101001;
assign LUT_2[21544] = 32'b11111111111111111100100111001001;
assign LUT_2[21545] = 32'b11111111111111111001011111100010;
assign LUT_2[21546] = 32'b00000000000000000011100000000101;
assign LUT_2[21547] = 32'b00000000000000000000011000011110;
assign LUT_2[21548] = 32'b11111111111111111001000100110001;
assign LUT_2[21549] = 32'b11111111111111110101111101001010;
assign LUT_2[21550] = 32'b11111111111111111111111101101101;
assign LUT_2[21551] = 32'b11111111111111111100110110000110;
assign LUT_2[21552] = 32'b11111111111111111100011001110110;
assign LUT_2[21553] = 32'b11111111111111111001010010001111;
assign LUT_2[21554] = 32'b00000000000000000011010010110010;
assign LUT_2[21555] = 32'b00000000000000000000001011001011;
assign LUT_2[21556] = 32'b11111111111111111000110111011110;
assign LUT_2[21557] = 32'b11111111111111110101101111110111;
assign LUT_2[21558] = 32'b11111111111111111111110000011010;
assign LUT_2[21559] = 32'b11111111111111111100101000110011;
assign LUT_2[21560] = 32'b11111111111111110111001011010011;
assign LUT_2[21561] = 32'b11111111111111110100000011101100;
assign LUT_2[21562] = 32'b11111111111111111110000100001111;
assign LUT_2[21563] = 32'b11111111111111111010111100101000;
assign LUT_2[21564] = 32'b11111111111111110011101000111011;
assign LUT_2[21565] = 32'b11111111111111110000100001010100;
assign LUT_2[21566] = 32'b11111111111111111010100001110111;
assign LUT_2[21567] = 32'b11111111111111110111011010010000;
assign LUT_2[21568] = 32'b11111111111111111001100010100110;
assign LUT_2[21569] = 32'b11111111111111110110011010111111;
assign LUT_2[21570] = 32'b00000000000000000000011011100010;
assign LUT_2[21571] = 32'b11111111111111111101010011111011;
assign LUT_2[21572] = 32'b11111111111111110110000000001110;
assign LUT_2[21573] = 32'b11111111111111110010111000100111;
assign LUT_2[21574] = 32'b11111111111111111100111001001010;
assign LUT_2[21575] = 32'b11111111111111111001110001100011;
assign LUT_2[21576] = 32'b11111111111111110100010100000011;
assign LUT_2[21577] = 32'b11111111111111110001001100011100;
assign LUT_2[21578] = 32'b11111111111111111011001100111111;
assign LUT_2[21579] = 32'b11111111111111111000000101011000;
assign LUT_2[21580] = 32'b11111111111111110000110001101011;
assign LUT_2[21581] = 32'b11111111111111101101101010000100;
assign LUT_2[21582] = 32'b11111111111111110111101010100111;
assign LUT_2[21583] = 32'b11111111111111110100100011000000;
assign LUT_2[21584] = 32'b11111111111111110100000110110000;
assign LUT_2[21585] = 32'b11111111111111110000111111001001;
assign LUT_2[21586] = 32'b11111111111111111010111111101100;
assign LUT_2[21587] = 32'b11111111111111110111111000000101;
assign LUT_2[21588] = 32'b11111111111111110000100100011000;
assign LUT_2[21589] = 32'b11111111111111101101011100110001;
assign LUT_2[21590] = 32'b11111111111111110111011101010100;
assign LUT_2[21591] = 32'b11111111111111110100010101101101;
assign LUT_2[21592] = 32'b11111111111111101110111000001101;
assign LUT_2[21593] = 32'b11111111111111101011110000100110;
assign LUT_2[21594] = 32'b11111111111111110101110001001001;
assign LUT_2[21595] = 32'b11111111111111110010101001100010;
assign LUT_2[21596] = 32'b11111111111111101011010101110101;
assign LUT_2[21597] = 32'b11111111111111101000001110001110;
assign LUT_2[21598] = 32'b11111111111111110010001110110001;
assign LUT_2[21599] = 32'b11111111111111101111000111001010;
assign LUT_2[21600] = 32'b11111111111111111001111110001111;
assign LUT_2[21601] = 32'b11111111111111110110110110101000;
assign LUT_2[21602] = 32'b00000000000000000000110111001011;
assign LUT_2[21603] = 32'b11111111111111111101101111100100;
assign LUT_2[21604] = 32'b11111111111111110110011011110111;
assign LUT_2[21605] = 32'b11111111111111110011010100010000;
assign LUT_2[21606] = 32'b11111111111111111101010100110011;
assign LUT_2[21607] = 32'b11111111111111111010001101001100;
assign LUT_2[21608] = 32'b11111111111111110100101111101100;
assign LUT_2[21609] = 32'b11111111111111110001101000000101;
assign LUT_2[21610] = 32'b11111111111111111011101000101000;
assign LUT_2[21611] = 32'b11111111111111111000100001000001;
assign LUT_2[21612] = 32'b11111111111111110001001101010100;
assign LUT_2[21613] = 32'b11111111111111101110000101101101;
assign LUT_2[21614] = 32'b11111111111111111000000110010000;
assign LUT_2[21615] = 32'b11111111111111110100111110101001;
assign LUT_2[21616] = 32'b11111111111111110100100010011001;
assign LUT_2[21617] = 32'b11111111111111110001011010110010;
assign LUT_2[21618] = 32'b11111111111111111011011011010101;
assign LUT_2[21619] = 32'b11111111111111111000010011101110;
assign LUT_2[21620] = 32'b11111111111111110001000000000001;
assign LUT_2[21621] = 32'b11111111111111101101111000011010;
assign LUT_2[21622] = 32'b11111111111111110111111000111101;
assign LUT_2[21623] = 32'b11111111111111110100110001010110;
assign LUT_2[21624] = 32'b11111111111111101111010011110110;
assign LUT_2[21625] = 32'b11111111111111101100001100001111;
assign LUT_2[21626] = 32'b11111111111111110110001100110010;
assign LUT_2[21627] = 32'b11111111111111110011000101001011;
assign LUT_2[21628] = 32'b11111111111111101011110001011110;
assign LUT_2[21629] = 32'b11111111111111101000101001110111;
assign LUT_2[21630] = 32'b11111111111111110010101010011010;
assign LUT_2[21631] = 32'b11111111111111101111100010110011;
assign LUT_2[21632] = 32'b00000000000000000101101110010010;
assign LUT_2[21633] = 32'b00000000000000000010100110101011;
assign LUT_2[21634] = 32'b00000000000000001100100111001110;
assign LUT_2[21635] = 32'b00000000000000001001011111100111;
assign LUT_2[21636] = 32'b00000000000000000010001011111010;
assign LUT_2[21637] = 32'b11111111111111111111000100010011;
assign LUT_2[21638] = 32'b00000000000000001001000100110110;
assign LUT_2[21639] = 32'b00000000000000000101111101001111;
assign LUT_2[21640] = 32'b00000000000000000000011111101111;
assign LUT_2[21641] = 32'b11111111111111111101011000001000;
assign LUT_2[21642] = 32'b00000000000000000111011000101011;
assign LUT_2[21643] = 32'b00000000000000000100010001000100;
assign LUT_2[21644] = 32'b11111111111111111100111101010111;
assign LUT_2[21645] = 32'b11111111111111111001110101110000;
assign LUT_2[21646] = 32'b00000000000000000011110110010011;
assign LUT_2[21647] = 32'b00000000000000000000101110101100;
assign LUT_2[21648] = 32'b00000000000000000000010010011100;
assign LUT_2[21649] = 32'b11111111111111111101001010110101;
assign LUT_2[21650] = 32'b00000000000000000111001011011000;
assign LUT_2[21651] = 32'b00000000000000000100000011110001;
assign LUT_2[21652] = 32'b11111111111111111100110000000100;
assign LUT_2[21653] = 32'b11111111111111111001101000011101;
assign LUT_2[21654] = 32'b00000000000000000011101001000000;
assign LUT_2[21655] = 32'b00000000000000000000100001011001;
assign LUT_2[21656] = 32'b11111111111111111011000011111001;
assign LUT_2[21657] = 32'b11111111111111110111111100010010;
assign LUT_2[21658] = 32'b00000000000000000001111100110101;
assign LUT_2[21659] = 32'b11111111111111111110110101001110;
assign LUT_2[21660] = 32'b11111111111111110111100001100001;
assign LUT_2[21661] = 32'b11111111111111110100011001111010;
assign LUT_2[21662] = 32'b11111111111111111110011010011101;
assign LUT_2[21663] = 32'b11111111111111111011010010110110;
assign LUT_2[21664] = 32'b00000000000000000110001001111011;
assign LUT_2[21665] = 32'b00000000000000000011000010010100;
assign LUT_2[21666] = 32'b00000000000000001101000010110111;
assign LUT_2[21667] = 32'b00000000000000001001111011010000;
assign LUT_2[21668] = 32'b00000000000000000010100111100011;
assign LUT_2[21669] = 32'b11111111111111111111011111111100;
assign LUT_2[21670] = 32'b00000000000000001001100000011111;
assign LUT_2[21671] = 32'b00000000000000000110011000111000;
assign LUT_2[21672] = 32'b00000000000000000000111011011000;
assign LUT_2[21673] = 32'b11111111111111111101110011110001;
assign LUT_2[21674] = 32'b00000000000000000111110100010100;
assign LUT_2[21675] = 32'b00000000000000000100101100101101;
assign LUT_2[21676] = 32'b11111111111111111101011001000000;
assign LUT_2[21677] = 32'b11111111111111111010010001011001;
assign LUT_2[21678] = 32'b00000000000000000100010001111100;
assign LUT_2[21679] = 32'b00000000000000000001001010010101;
assign LUT_2[21680] = 32'b00000000000000000000101110000101;
assign LUT_2[21681] = 32'b11111111111111111101100110011110;
assign LUT_2[21682] = 32'b00000000000000000111100111000001;
assign LUT_2[21683] = 32'b00000000000000000100011111011010;
assign LUT_2[21684] = 32'b11111111111111111101001011101101;
assign LUT_2[21685] = 32'b11111111111111111010000100000110;
assign LUT_2[21686] = 32'b00000000000000000100000100101001;
assign LUT_2[21687] = 32'b00000000000000000000111101000010;
assign LUT_2[21688] = 32'b11111111111111111011011111100010;
assign LUT_2[21689] = 32'b11111111111111111000010111111011;
assign LUT_2[21690] = 32'b00000000000000000010011000011110;
assign LUT_2[21691] = 32'b11111111111111111111010000110111;
assign LUT_2[21692] = 32'b11111111111111110111111101001010;
assign LUT_2[21693] = 32'b11111111111111110100110101100011;
assign LUT_2[21694] = 32'b11111111111111111110110110000110;
assign LUT_2[21695] = 32'b11111111111111111011101110011111;
assign LUT_2[21696] = 32'b11111111111111111101110110110101;
assign LUT_2[21697] = 32'b11111111111111111010101111001110;
assign LUT_2[21698] = 32'b00000000000000000100101111110001;
assign LUT_2[21699] = 32'b00000000000000000001101000001010;
assign LUT_2[21700] = 32'b11111111111111111010010100011101;
assign LUT_2[21701] = 32'b11111111111111110111001100110110;
assign LUT_2[21702] = 32'b00000000000000000001001101011001;
assign LUT_2[21703] = 32'b11111111111111111110000101110010;
assign LUT_2[21704] = 32'b11111111111111111000101000010010;
assign LUT_2[21705] = 32'b11111111111111110101100000101011;
assign LUT_2[21706] = 32'b11111111111111111111100001001110;
assign LUT_2[21707] = 32'b11111111111111111100011001100111;
assign LUT_2[21708] = 32'b11111111111111110101000101111010;
assign LUT_2[21709] = 32'b11111111111111110001111110010011;
assign LUT_2[21710] = 32'b11111111111111111011111110110110;
assign LUT_2[21711] = 32'b11111111111111111000110111001111;
assign LUT_2[21712] = 32'b11111111111111111000011010111111;
assign LUT_2[21713] = 32'b11111111111111110101010011011000;
assign LUT_2[21714] = 32'b11111111111111111111010011111011;
assign LUT_2[21715] = 32'b11111111111111111100001100010100;
assign LUT_2[21716] = 32'b11111111111111110100111000100111;
assign LUT_2[21717] = 32'b11111111111111110001110001000000;
assign LUT_2[21718] = 32'b11111111111111111011110001100011;
assign LUT_2[21719] = 32'b11111111111111111000101001111100;
assign LUT_2[21720] = 32'b11111111111111110011001100011100;
assign LUT_2[21721] = 32'b11111111111111110000000100110101;
assign LUT_2[21722] = 32'b11111111111111111010000101011000;
assign LUT_2[21723] = 32'b11111111111111110110111101110001;
assign LUT_2[21724] = 32'b11111111111111101111101010000100;
assign LUT_2[21725] = 32'b11111111111111101100100010011101;
assign LUT_2[21726] = 32'b11111111111111110110100011000000;
assign LUT_2[21727] = 32'b11111111111111110011011011011001;
assign LUT_2[21728] = 32'b11111111111111111110010010011110;
assign LUT_2[21729] = 32'b11111111111111111011001010110111;
assign LUT_2[21730] = 32'b00000000000000000101001011011010;
assign LUT_2[21731] = 32'b00000000000000000010000011110011;
assign LUT_2[21732] = 32'b11111111111111111010110000000110;
assign LUT_2[21733] = 32'b11111111111111110111101000011111;
assign LUT_2[21734] = 32'b00000000000000000001101001000010;
assign LUT_2[21735] = 32'b11111111111111111110100001011011;
assign LUT_2[21736] = 32'b11111111111111111001000011111011;
assign LUT_2[21737] = 32'b11111111111111110101111100010100;
assign LUT_2[21738] = 32'b11111111111111111111111100110111;
assign LUT_2[21739] = 32'b11111111111111111100110101010000;
assign LUT_2[21740] = 32'b11111111111111110101100001100011;
assign LUT_2[21741] = 32'b11111111111111110010011001111100;
assign LUT_2[21742] = 32'b11111111111111111100011010011111;
assign LUT_2[21743] = 32'b11111111111111111001010010111000;
assign LUT_2[21744] = 32'b11111111111111111000110110101000;
assign LUT_2[21745] = 32'b11111111111111110101101111000001;
assign LUT_2[21746] = 32'b11111111111111111111101111100100;
assign LUT_2[21747] = 32'b11111111111111111100100111111101;
assign LUT_2[21748] = 32'b11111111111111110101010100010000;
assign LUT_2[21749] = 32'b11111111111111110010001100101001;
assign LUT_2[21750] = 32'b11111111111111111100001101001100;
assign LUT_2[21751] = 32'b11111111111111111001000101100101;
assign LUT_2[21752] = 32'b11111111111111110011101000000101;
assign LUT_2[21753] = 32'b11111111111111110000100000011110;
assign LUT_2[21754] = 32'b11111111111111111010100001000001;
assign LUT_2[21755] = 32'b11111111111111110111011001011010;
assign LUT_2[21756] = 32'b11111111111111110000000101101101;
assign LUT_2[21757] = 32'b11111111111111101100111110000110;
assign LUT_2[21758] = 32'b11111111111111110110111110101001;
assign LUT_2[21759] = 32'b11111111111111110011110111000010;
assign LUT_2[21760] = 32'b00000000000000000101011000101001;
assign LUT_2[21761] = 32'b00000000000000000010010001000010;
assign LUT_2[21762] = 32'b00000000000000001100010001100101;
assign LUT_2[21763] = 32'b00000000000000001001001001111110;
assign LUT_2[21764] = 32'b00000000000000000001110110010001;
assign LUT_2[21765] = 32'b11111111111111111110101110101010;
assign LUT_2[21766] = 32'b00000000000000001000101111001101;
assign LUT_2[21767] = 32'b00000000000000000101100111100110;
assign LUT_2[21768] = 32'b00000000000000000000001010000110;
assign LUT_2[21769] = 32'b11111111111111111101000010011111;
assign LUT_2[21770] = 32'b00000000000000000111000011000010;
assign LUT_2[21771] = 32'b00000000000000000011111011011011;
assign LUT_2[21772] = 32'b11111111111111111100100111101110;
assign LUT_2[21773] = 32'b11111111111111111001100000000111;
assign LUT_2[21774] = 32'b00000000000000000011100000101010;
assign LUT_2[21775] = 32'b00000000000000000000011001000011;
assign LUT_2[21776] = 32'b11111111111111111111111100110011;
assign LUT_2[21777] = 32'b11111111111111111100110101001100;
assign LUT_2[21778] = 32'b00000000000000000110110101101111;
assign LUT_2[21779] = 32'b00000000000000000011101110001000;
assign LUT_2[21780] = 32'b11111111111111111100011010011011;
assign LUT_2[21781] = 32'b11111111111111111001010010110100;
assign LUT_2[21782] = 32'b00000000000000000011010011010111;
assign LUT_2[21783] = 32'b00000000000000000000001011110000;
assign LUT_2[21784] = 32'b11111111111111111010101110010000;
assign LUT_2[21785] = 32'b11111111111111110111100110101001;
assign LUT_2[21786] = 32'b00000000000000000001100111001100;
assign LUT_2[21787] = 32'b11111111111111111110011111100101;
assign LUT_2[21788] = 32'b11111111111111110111001011111000;
assign LUT_2[21789] = 32'b11111111111111110100000100010001;
assign LUT_2[21790] = 32'b11111111111111111110000100110100;
assign LUT_2[21791] = 32'b11111111111111111010111101001101;
assign LUT_2[21792] = 32'b00000000000000000101110100010010;
assign LUT_2[21793] = 32'b00000000000000000010101100101011;
assign LUT_2[21794] = 32'b00000000000000001100101101001110;
assign LUT_2[21795] = 32'b00000000000000001001100101100111;
assign LUT_2[21796] = 32'b00000000000000000010010001111010;
assign LUT_2[21797] = 32'b11111111111111111111001010010011;
assign LUT_2[21798] = 32'b00000000000000001001001010110110;
assign LUT_2[21799] = 32'b00000000000000000110000011001111;
assign LUT_2[21800] = 32'b00000000000000000000100101101111;
assign LUT_2[21801] = 32'b11111111111111111101011110001000;
assign LUT_2[21802] = 32'b00000000000000000111011110101011;
assign LUT_2[21803] = 32'b00000000000000000100010111000100;
assign LUT_2[21804] = 32'b11111111111111111101000011010111;
assign LUT_2[21805] = 32'b11111111111111111001111011110000;
assign LUT_2[21806] = 32'b00000000000000000011111100010011;
assign LUT_2[21807] = 32'b00000000000000000000110100101100;
assign LUT_2[21808] = 32'b00000000000000000000011000011100;
assign LUT_2[21809] = 32'b11111111111111111101010000110101;
assign LUT_2[21810] = 32'b00000000000000000111010001011000;
assign LUT_2[21811] = 32'b00000000000000000100001001110001;
assign LUT_2[21812] = 32'b11111111111111111100110110000100;
assign LUT_2[21813] = 32'b11111111111111111001101110011101;
assign LUT_2[21814] = 32'b00000000000000000011101111000000;
assign LUT_2[21815] = 32'b00000000000000000000100111011001;
assign LUT_2[21816] = 32'b11111111111111111011001001111001;
assign LUT_2[21817] = 32'b11111111111111111000000010010010;
assign LUT_2[21818] = 32'b00000000000000000010000010110101;
assign LUT_2[21819] = 32'b11111111111111111110111011001110;
assign LUT_2[21820] = 32'b11111111111111110111100111100001;
assign LUT_2[21821] = 32'b11111111111111110100011111111010;
assign LUT_2[21822] = 32'b11111111111111111110100000011101;
assign LUT_2[21823] = 32'b11111111111111111011011000110110;
assign LUT_2[21824] = 32'b11111111111111111101100001001100;
assign LUT_2[21825] = 32'b11111111111111111010011001100101;
assign LUT_2[21826] = 32'b00000000000000000100011010001000;
assign LUT_2[21827] = 32'b00000000000000000001010010100001;
assign LUT_2[21828] = 32'b11111111111111111001111110110100;
assign LUT_2[21829] = 32'b11111111111111110110110111001101;
assign LUT_2[21830] = 32'b00000000000000000000110111110000;
assign LUT_2[21831] = 32'b11111111111111111101110000001001;
assign LUT_2[21832] = 32'b11111111111111111000010010101001;
assign LUT_2[21833] = 32'b11111111111111110101001011000010;
assign LUT_2[21834] = 32'b11111111111111111111001011100101;
assign LUT_2[21835] = 32'b11111111111111111100000011111110;
assign LUT_2[21836] = 32'b11111111111111110100110000010001;
assign LUT_2[21837] = 32'b11111111111111110001101000101010;
assign LUT_2[21838] = 32'b11111111111111111011101001001101;
assign LUT_2[21839] = 32'b11111111111111111000100001100110;
assign LUT_2[21840] = 32'b11111111111111111000000101010110;
assign LUT_2[21841] = 32'b11111111111111110100111101101111;
assign LUT_2[21842] = 32'b11111111111111111110111110010010;
assign LUT_2[21843] = 32'b11111111111111111011110110101011;
assign LUT_2[21844] = 32'b11111111111111110100100010111110;
assign LUT_2[21845] = 32'b11111111111111110001011011010111;
assign LUT_2[21846] = 32'b11111111111111111011011011111010;
assign LUT_2[21847] = 32'b11111111111111111000010100010011;
assign LUT_2[21848] = 32'b11111111111111110010110110110011;
assign LUT_2[21849] = 32'b11111111111111101111101111001100;
assign LUT_2[21850] = 32'b11111111111111111001101111101111;
assign LUT_2[21851] = 32'b11111111111111110110101000001000;
assign LUT_2[21852] = 32'b11111111111111101111010100011011;
assign LUT_2[21853] = 32'b11111111111111101100001100110100;
assign LUT_2[21854] = 32'b11111111111111110110001101010111;
assign LUT_2[21855] = 32'b11111111111111110011000101110000;
assign LUT_2[21856] = 32'b11111111111111111101111100110101;
assign LUT_2[21857] = 32'b11111111111111111010110101001110;
assign LUT_2[21858] = 32'b00000000000000000100110101110001;
assign LUT_2[21859] = 32'b00000000000000000001101110001010;
assign LUT_2[21860] = 32'b11111111111111111010011010011101;
assign LUT_2[21861] = 32'b11111111111111110111010010110110;
assign LUT_2[21862] = 32'b00000000000000000001010011011001;
assign LUT_2[21863] = 32'b11111111111111111110001011110010;
assign LUT_2[21864] = 32'b11111111111111111000101110010010;
assign LUT_2[21865] = 32'b11111111111111110101100110101011;
assign LUT_2[21866] = 32'b11111111111111111111100111001110;
assign LUT_2[21867] = 32'b11111111111111111100011111100111;
assign LUT_2[21868] = 32'b11111111111111110101001011111010;
assign LUT_2[21869] = 32'b11111111111111110010000100010011;
assign LUT_2[21870] = 32'b11111111111111111100000100110110;
assign LUT_2[21871] = 32'b11111111111111111000111101001111;
assign LUT_2[21872] = 32'b11111111111111111000100000111111;
assign LUT_2[21873] = 32'b11111111111111110101011001011000;
assign LUT_2[21874] = 32'b11111111111111111111011001111011;
assign LUT_2[21875] = 32'b11111111111111111100010010010100;
assign LUT_2[21876] = 32'b11111111111111110100111110100111;
assign LUT_2[21877] = 32'b11111111111111110001110111000000;
assign LUT_2[21878] = 32'b11111111111111111011110111100011;
assign LUT_2[21879] = 32'b11111111111111111000101111111100;
assign LUT_2[21880] = 32'b11111111111111110011010010011100;
assign LUT_2[21881] = 32'b11111111111111110000001010110101;
assign LUT_2[21882] = 32'b11111111111111111010001011011000;
assign LUT_2[21883] = 32'b11111111111111110111000011110001;
assign LUT_2[21884] = 32'b11111111111111101111110000000100;
assign LUT_2[21885] = 32'b11111111111111101100101000011101;
assign LUT_2[21886] = 32'b11111111111111110110101001000000;
assign LUT_2[21887] = 32'b11111111111111110011100001011001;
assign LUT_2[21888] = 32'b00000000000000001001101100111000;
assign LUT_2[21889] = 32'b00000000000000000110100101010001;
assign LUT_2[21890] = 32'b00000000000000010000100101110100;
assign LUT_2[21891] = 32'b00000000000000001101011110001101;
assign LUT_2[21892] = 32'b00000000000000000110001010100000;
assign LUT_2[21893] = 32'b00000000000000000011000010111001;
assign LUT_2[21894] = 32'b00000000000000001101000011011100;
assign LUT_2[21895] = 32'b00000000000000001001111011110101;
assign LUT_2[21896] = 32'b00000000000000000100011110010101;
assign LUT_2[21897] = 32'b00000000000000000001010110101110;
assign LUT_2[21898] = 32'b00000000000000001011010111010001;
assign LUT_2[21899] = 32'b00000000000000001000001111101010;
assign LUT_2[21900] = 32'b00000000000000000000111011111101;
assign LUT_2[21901] = 32'b11111111111111111101110100010110;
assign LUT_2[21902] = 32'b00000000000000000111110100111001;
assign LUT_2[21903] = 32'b00000000000000000100101101010010;
assign LUT_2[21904] = 32'b00000000000000000100010001000010;
assign LUT_2[21905] = 32'b00000000000000000001001001011011;
assign LUT_2[21906] = 32'b00000000000000001011001001111110;
assign LUT_2[21907] = 32'b00000000000000001000000010010111;
assign LUT_2[21908] = 32'b00000000000000000000101110101010;
assign LUT_2[21909] = 32'b11111111111111111101100111000011;
assign LUT_2[21910] = 32'b00000000000000000111100111100110;
assign LUT_2[21911] = 32'b00000000000000000100011111111111;
assign LUT_2[21912] = 32'b11111111111111111111000010011111;
assign LUT_2[21913] = 32'b11111111111111111011111010111000;
assign LUT_2[21914] = 32'b00000000000000000101111011011011;
assign LUT_2[21915] = 32'b00000000000000000010110011110100;
assign LUT_2[21916] = 32'b11111111111111111011100000000111;
assign LUT_2[21917] = 32'b11111111111111111000011000100000;
assign LUT_2[21918] = 32'b00000000000000000010011001000011;
assign LUT_2[21919] = 32'b11111111111111111111010001011100;
assign LUT_2[21920] = 32'b00000000000000001010001000100001;
assign LUT_2[21921] = 32'b00000000000000000111000000111010;
assign LUT_2[21922] = 32'b00000000000000010001000001011101;
assign LUT_2[21923] = 32'b00000000000000001101111001110110;
assign LUT_2[21924] = 32'b00000000000000000110100110001001;
assign LUT_2[21925] = 32'b00000000000000000011011110100010;
assign LUT_2[21926] = 32'b00000000000000001101011111000101;
assign LUT_2[21927] = 32'b00000000000000001010010111011110;
assign LUT_2[21928] = 32'b00000000000000000100111001111110;
assign LUT_2[21929] = 32'b00000000000000000001110010010111;
assign LUT_2[21930] = 32'b00000000000000001011110010111010;
assign LUT_2[21931] = 32'b00000000000000001000101011010011;
assign LUT_2[21932] = 32'b00000000000000000001010111100110;
assign LUT_2[21933] = 32'b11111111111111111110001111111111;
assign LUT_2[21934] = 32'b00000000000000001000010000100010;
assign LUT_2[21935] = 32'b00000000000000000101001000111011;
assign LUT_2[21936] = 32'b00000000000000000100101100101011;
assign LUT_2[21937] = 32'b00000000000000000001100101000100;
assign LUT_2[21938] = 32'b00000000000000001011100101100111;
assign LUT_2[21939] = 32'b00000000000000001000011110000000;
assign LUT_2[21940] = 32'b00000000000000000001001010010011;
assign LUT_2[21941] = 32'b11111111111111111110000010101100;
assign LUT_2[21942] = 32'b00000000000000001000000011001111;
assign LUT_2[21943] = 32'b00000000000000000100111011101000;
assign LUT_2[21944] = 32'b11111111111111111111011110001000;
assign LUT_2[21945] = 32'b11111111111111111100010110100001;
assign LUT_2[21946] = 32'b00000000000000000110010111000100;
assign LUT_2[21947] = 32'b00000000000000000011001111011101;
assign LUT_2[21948] = 32'b11111111111111111011111011110000;
assign LUT_2[21949] = 32'b11111111111111111000110100001001;
assign LUT_2[21950] = 32'b00000000000000000010110100101100;
assign LUT_2[21951] = 32'b11111111111111111111101101000101;
assign LUT_2[21952] = 32'b00000000000000000001110101011011;
assign LUT_2[21953] = 32'b11111111111111111110101101110100;
assign LUT_2[21954] = 32'b00000000000000001000101110010111;
assign LUT_2[21955] = 32'b00000000000000000101100110110000;
assign LUT_2[21956] = 32'b11111111111111111110010011000011;
assign LUT_2[21957] = 32'b11111111111111111011001011011100;
assign LUT_2[21958] = 32'b00000000000000000101001011111111;
assign LUT_2[21959] = 32'b00000000000000000010000100011000;
assign LUT_2[21960] = 32'b11111111111111111100100110111000;
assign LUT_2[21961] = 32'b11111111111111111001011111010001;
assign LUT_2[21962] = 32'b00000000000000000011011111110100;
assign LUT_2[21963] = 32'b00000000000000000000011000001101;
assign LUT_2[21964] = 32'b11111111111111111001000100100000;
assign LUT_2[21965] = 32'b11111111111111110101111100111001;
assign LUT_2[21966] = 32'b11111111111111111111111101011100;
assign LUT_2[21967] = 32'b11111111111111111100110101110101;
assign LUT_2[21968] = 32'b11111111111111111100011001100101;
assign LUT_2[21969] = 32'b11111111111111111001010001111110;
assign LUT_2[21970] = 32'b00000000000000000011010010100001;
assign LUT_2[21971] = 32'b00000000000000000000001010111010;
assign LUT_2[21972] = 32'b11111111111111111000110111001101;
assign LUT_2[21973] = 32'b11111111111111110101101111100110;
assign LUT_2[21974] = 32'b11111111111111111111110000001001;
assign LUT_2[21975] = 32'b11111111111111111100101000100010;
assign LUT_2[21976] = 32'b11111111111111110111001011000010;
assign LUT_2[21977] = 32'b11111111111111110100000011011011;
assign LUT_2[21978] = 32'b11111111111111111110000011111110;
assign LUT_2[21979] = 32'b11111111111111111010111100010111;
assign LUT_2[21980] = 32'b11111111111111110011101000101010;
assign LUT_2[21981] = 32'b11111111111111110000100001000011;
assign LUT_2[21982] = 32'b11111111111111111010100001100110;
assign LUT_2[21983] = 32'b11111111111111110111011001111111;
assign LUT_2[21984] = 32'b00000000000000000010010001000100;
assign LUT_2[21985] = 32'b11111111111111111111001001011101;
assign LUT_2[21986] = 32'b00000000000000001001001010000000;
assign LUT_2[21987] = 32'b00000000000000000110000010011001;
assign LUT_2[21988] = 32'b11111111111111111110101110101100;
assign LUT_2[21989] = 32'b11111111111111111011100111000101;
assign LUT_2[21990] = 32'b00000000000000000101100111101000;
assign LUT_2[21991] = 32'b00000000000000000010100000000001;
assign LUT_2[21992] = 32'b11111111111111111101000010100001;
assign LUT_2[21993] = 32'b11111111111111111001111010111010;
assign LUT_2[21994] = 32'b00000000000000000011111011011101;
assign LUT_2[21995] = 32'b00000000000000000000110011110110;
assign LUT_2[21996] = 32'b11111111111111111001100000001001;
assign LUT_2[21997] = 32'b11111111111111110110011000100010;
assign LUT_2[21998] = 32'b00000000000000000000011001000101;
assign LUT_2[21999] = 32'b11111111111111111101010001011110;
assign LUT_2[22000] = 32'b11111111111111111100110101001110;
assign LUT_2[22001] = 32'b11111111111111111001101101100111;
assign LUT_2[22002] = 32'b00000000000000000011101110001010;
assign LUT_2[22003] = 32'b00000000000000000000100110100011;
assign LUT_2[22004] = 32'b11111111111111111001010010110110;
assign LUT_2[22005] = 32'b11111111111111110110001011001111;
assign LUT_2[22006] = 32'b00000000000000000000001011110010;
assign LUT_2[22007] = 32'b11111111111111111101000100001011;
assign LUT_2[22008] = 32'b11111111111111110111100110101011;
assign LUT_2[22009] = 32'b11111111111111110100011111000100;
assign LUT_2[22010] = 32'b11111111111111111110011111100111;
assign LUT_2[22011] = 32'b11111111111111111011011000000000;
assign LUT_2[22012] = 32'b11111111111111110100000100010011;
assign LUT_2[22013] = 32'b11111111111111110000111100101100;
assign LUT_2[22014] = 32'b11111111111111111010111101001111;
assign LUT_2[22015] = 32'b11111111111111110111110101101000;
assign LUT_2[22016] = 32'b00000000000000000110001011110101;
assign LUT_2[22017] = 32'b00000000000000000011000100001110;
assign LUT_2[22018] = 32'b00000000000000001101000100110001;
assign LUT_2[22019] = 32'b00000000000000001001111101001010;
assign LUT_2[22020] = 32'b00000000000000000010101001011101;
assign LUT_2[22021] = 32'b11111111111111111111100001110110;
assign LUT_2[22022] = 32'b00000000000000001001100010011001;
assign LUT_2[22023] = 32'b00000000000000000110011010110010;
assign LUT_2[22024] = 32'b00000000000000000000111101010010;
assign LUT_2[22025] = 32'b11111111111111111101110101101011;
assign LUT_2[22026] = 32'b00000000000000000111110110001110;
assign LUT_2[22027] = 32'b00000000000000000100101110100111;
assign LUT_2[22028] = 32'b11111111111111111101011010111010;
assign LUT_2[22029] = 32'b11111111111111111010010011010011;
assign LUT_2[22030] = 32'b00000000000000000100010011110110;
assign LUT_2[22031] = 32'b00000000000000000001001100001111;
assign LUT_2[22032] = 32'b00000000000000000000101111111111;
assign LUT_2[22033] = 32'b11111111111111111101101000011000;
assign LUT_2[22034] = 32'b00000000000000000111101000111011;
assign LUT_2[22035] = 32'b00000000000000000100100001010100;
assign LUT_2[22036] = 32'b11111111111111111101001101100111;
assign LUT_2[22037] = 32'b11111111111111111010000110000000;
assign LUT_2[22038] = 32'b00000000000000000100000110100011;
assign LUT_2[22039] = 32'b00000000000000000000111110111100;
assign LUT_2[22040] = 32'b11111111111111111011100001011100;
assign LUT_2[22041] = 32'b11111111111111111000011001110101;
assign LUT_2[22042] = 32'b00000000000000000010011010011000;
assign LUT_2[22043] = 32'b11111111111111111111010010110001;
assign LUT_2[22044] = 32'b11111111111111110111111111000100;
assign LUT_2[22045] = 32'b11111111111111110100110111011101;
assign LUT_2[22046] = 32'b11111111111111111110111000000000;
assign LUT_2[22047] = 32'b11111111111111111011110000011001;
assign LUT_2[22048] = 32'b00000000000000000110100111011110;
assign LUT_2[22049] = 32'b00000000000000000011011111110111;
assign LUT_2[22050] = 32'b00000000000000001101100000011010;
assign LUT_2[22051] = 32'b00000000000000001010011000110011;
assign LUT_2[22052] = 32'b00000000000000000011000101000110;
assign LUT_2[22053] = 32'b11111111111111111111111101011111;
assign LUT_2[22054] = 32'b00000000000000001001111110000010;
assign LUT_2[22055] = 32'b00000000000000000110110110011011;
assign LUT_2[22056] = 32'b00000000000000000001011000111011;
assign LUT_2[22057] = 32'b11111111111111111110010001010100;
assign LUT_2[22058] = 32'b00000000000000001000010001110111;
assign LUT_2[22059] = 32'b00000000000000000101001010010000;
assign LUT_2[22060] = 32'b11111111111111111101110110100011;
assign LUT_2[22061] = 32'b11111111111111111010101110111100;
assign LUT_2[22062] = 32'b00000000000000000100101111011111;
assign LUT_2[22063] = 32'b00000000000000000001100111111000;
assign LUT_2[22064] = 32'b00000000000000000001001011101000;
assign LUT_2[22065] = 32'b11111111111111111110000100000001;
assign LUT_2[22066] = 32'b00000000000000001000000100100100;
assign LUT_2[22067] = 32'b00000000000000000100111100111101;
assign LUT_2[22068] = 32'b11111111111111111101101001010000;
assign LUT_2[22069] = 32'b11111111111111111010100001101001;
assign LUT_2[22070] = 32'b00000000000000000100100010001100;
assign LUT_2[22071] = 32'b00000000000000000001011010100101;
assign LUT_2[22072] = 32'b11111111111111111011111101000101;
assign LUT_2[22073] = 32'b11111111111111111000110101011110;
assign LUT_2[22074] = 32'b00000000000000000010110110000001;
assign LUT_2[22075] = 32'b11111111111111111111101110011010;
assign LUT_2[22076] = 32'b11111111111111111000011010101101;
assign LUT_2[22077] = 32'b11111111111111110101010011000110;
assign LUT_2[22078] = 32'b11111111111111111111010011101001;
assign LUT_2[22079] = 32'b11111111111111111100001100000010;
assign LUT_2[22080] = 32'b11111111111111111110010100011000;
assign LUT_2[22081] = 32'b11111111111111111011001100110001;
assign LUT_2[22082] = 32'b00000000000000000101001101010100;
assign LUT_2[22083] = 32'b00000000000000000010000101101101;
assign LUT_2[22084] = 32'b11111111111111111010110010000000;
assign LUT_2[22085] = 32'b11111111111111110111101010011001;
assign LUT_2[22086] = 32'b00000000000000000001101010111100;
assign LUT_2[22087] = 32'b11111111111111111110100011010101;
assign LUT_2[22088] = 32'b11111111111111111001000101110101;
assign LUT_2[22089] = 32'b11111111111111110101111110001110;
assign LUT_2[22090] = 32'b11111111111111111111111110110001;
assign LUT_2[22091] = 32'b11111111111111111100110111001010;
assign LUT_2[22092] = 32'b11111111111111110101100011011101;
assign LUT_2[22093] = 32'b11111111111111110010011011110110;
assign LUT_2[22094] = 32'b11111111111111111100011100011001;
assign LUT_2[22095] = 32'b11111111111111111001010100110010;
assign LUT_2[22096] = 32'b11111111111111111000111000100010;
assign LUT_2[22097] = 32'b11111111111111110101110000111011;
assign LUT_2[22098] = 32'b11111111111111111111110001011110;
assign LUT_2[22099] = 32'b11111111111111111100101001110111;
assign LUT_2[22100] = 32'b11111111111111110101010110001010;
assign LUT_2[22101] = 32'b11111111111111110010001110100011;
assign LUT_2[22102] = 32'b11111111111111111100001111000110;
assign LUT_2[22103] = 32'b11111111111111111001000111011111;
assign LUT_2[22104] = 32'b11111111111111110011101001111111;
assign LUT_2[22105] = 32'b11111111111111110000100010011000;
assign LUT_2[22106] = 32'b11111111111111111010100010111011;
assign LUT_2[22107] = 32'b11111111111111110111011011010100;
assign LUT_2[22108] = 32'b11111111111111110000000111100111;
assign LUT_2[22109] = 32'b11111111111111101101000000000000;
assign LUT_2[22110] = 32'b11111111111111110111000000100011;
assign LUT_2[22111] = 32'b11111111111111110011111000111100;
assign LUT_2[22112] = 32'b11111111111111111110110000000001;
assign LUT_2[22113] = 32'b11111111111111111011101000011010;
assign LUT_2[22114] = 32'b00000000000000000101101000111101;
assign LUT_2[22115] = 32'b00000000000000000010100001010110;
assign LUT_2[22116] = 32'b11111111111111111011001101101001;
assign LUT_2[22117] = 32'b11111111111111111000000110000010;
assign LUT_2[22118] = 32'b00000000000000000010000110100101;
assign LUT_2[22119] = 32'b11111111111111111110111110111110;
assign LUT_2[22120] = 32'b11111111111111111001100001011110;
assign LUT_2[22121] = 32'b11111111111111110110011001110111;
assign LUT_2[22122] = 32'b00000000000000000000011010011010;
assign LUT_2[22123] = 32'b11111111111111111101010010110011;
assign LUT_2[22124] = 32'b11111111111111110101111111000110;
assign LUT_2[22125] = 32'b11111111111111110010110111011111;
assign LUT_2[22126] = 32'b11111111111111111100111000000010;
assign LUT_2[22127] = 32'b11111111111111111001110000011011;
assign LUT_2[22128] = 32'b11111111111111111001010100001011;
assign LUT_2[22129] = 32'b11111111111111110110001100100100;
assign LUT_2[22130] = 32'b00000000000000000000001101000111;
assign LUT_2[22131] = 32'b11111111111111111101000101100000;
assign LUT_2[22132] = 32'b11111111111111110101110001110011;
assign LUT_2[22133] = 32'b11111111111111110010101010001100;
assign LUT_2[22134] = 32'b11111111111111111100101010101111;
assign LUT_2[22135] = 32'b11111111111111111001100011001000;
assign LUT_2[22136] = 32'b11111111111111110100000101101000;
assign LUT_2[22137] = 32'b11111111111111110000111110000001;
assign LUT_2[22138] = 32'b11111111111111111010111110100100;
assign LUT_2[22139] = 32'b11111111111111110111110110111101;
assign LUT_2[22140] = 32'b11111111111111110000100011010000;
assign LUT_2[22141] = 32'b11111111111111101101011011101001;
assign LUT_2[22142] = 32'b11111111111111110111011100001100;
assign LUT_2[22143] = 32'b11111111111111110100010100100101;
assign LUT_2[22144] = 32'b00000000000000001010100000000100;
assign LUT_2[22145] = 32'b00000000000000000111011000011101;
assign LUT_2[22146] = 32'b00000000000000010001011001000000;
assign LUT_2[22147] = 32'b00000000000000001110010001011001;
assign LUT_2[22148] = 32'b00000000000000000110111101101100;
assign LUT_2[22149] = 32'b00000000000000000011110110000101;
assign LUT_2[22150] = 32'b00000000000000001101110110101000;
assign LUT_2[22151] = 32'b00000000000000001010101111000001;
assign LUT_2[22152] = 32'b00000000000000000101010001100001;
assign LUT_2[22153] = 32'b00000000000000000010001001111010;
assign LUT_2[22154] = 32'b00000000000000001100001010011101;
assign LUT_2[22155] = 32'b00000000000000001001000010110110;
assign LUT_2[22156] = 32'b00000000000000000001101111001001;
assign LUT_2[22157] = 32'b11111111111111111110100111100010;
assign LUT_2[22158] = 32'b00000000000000001000101000000101;
assign LUT_2[22159] = 32'b00000000000000000101100000011110;
assign LUT_2[22160] = 32'b00000000000000000101000100001110;
assign LUT_2[22161] = 32'b00000000000000000001111100100111;
assign LUT_2[22162] = 32'b00000000000000001011111101001010;
assign LUT_2[22163] = 32'b00000000000000001000110101100011;
assign LUT_2[22164] = 32'b00000000000000000001100001110110;
assign LUT_2[22165] = 32'b11111111111111111110011010001111;
assign LUT_2[22166] = 32'b00000000000000001000011010110010;
assign LUT_2[22167] = 32'b00000000000000000101010011001011;
assign LUT_2[22168] = 32'b11111111111111111111110101101011;
assign LUT_2[22169] = 32'b11111111111111111100101110000100;
assign LUT_2[22170] = 32'b00000000000000000110101110100111;
assign LUT_2[22171] = 32'b00000000000000000011100111000000;
assign LUT_2[22172] = 32'b11111111111111111100010011010011;
assign LUT_2[22173] = 32'b11111111111111111001001011101100;
assign LUT_2[22174] = 32'b00000000000000000011001100001111;
assign LUT_2[22175] = 32'b00000000000000000000000100101000;
assign LUT_2[22176] = 32'b00000000000000001010111011101101;
assign LUT_2[22177] = 32'b00000000000000000111110100000110;
assign LUT_2[22178] = 32'b00000000000000010001110100101001;
assign LUT_2[22179] = 32'b00000000000000001110101101000010;
assign LUT_2[22180] = 32'b00000000000000000111011001010101;
assign LUT_2[22181] = 32'b00000000000000000100010001101110;
assign LUT_2[22182] = 32'b00000000000000001110010010010001;
assign LUT_2[22183] = 32'b00000000000000001011001010101010;
assign LUT_2[22184] = 32'b00000000000000000101101101001010;
assign LUT_2[22185] = 32'b00000000000000000010100101100011;
assign LUT_2[22186] = 32'b00000000000000001100100110000110;
assign LUT_2[22187] = 32'b00000000000000001001011110011111;
assign LUT_2[22188] = 32'b00000000000000000010001010110010;
assign LUT_2[22189] = 32'b11111111111111111111000011001011;
assign LUT_2[22190] = 32'b00000000000000001001000011101110;
assign LUT_2[22191] = 32'b00000000000000000101111100000111;
assign LUT_2[22192] = 32'b00000000000000000101011111110111;
assign LUT_2[22193] = 32'b00000000000000000010011000010000;
assign LUT_2[22194] = 32'b00000000000000001100011000110011;
assign LUT_2[22195] = 32'b00000000000000001001010001001100;
assign LUT_2[22196] = 32'b00000000000000000001111101011111;
assign LUT_2[22197] = 32'b11111111111111111110110101111000;
assign LUT_2[22198] = 32'b00000000000000001000110110011011;
assign LUT_2[22199] = 32'b00000000000000000101101110110100;
assign LUT_2[22200] = 32'b00000000000000000000010001010100;
assign LUT_2[22201] = 32'b11111111111111111101001001101101;
assign LUT_2[22202] = 32'b00000000000000000111001010010000;
assign LUT_2[22203] = 32'b00000000000000000100000010101001;
assign LUT_2[22204] = 32'b11111111111111111100101110111100;
assign LUT_2[22205] = 32'b11111111111111111001100111010101;
assign LUT_2[22206] = 32'b00000000000000000011100111111000;
assign LUT_2[22207] = 32'b00000000000000000000100000010001;
assign LUT_2[22208] = 32'b00000000000000000010101000100111;
assign LUT_2[22209] = 32'b11111111111111111111100001000000;
assign LUT_2[22210] = 32'b00000000000000001001100001100011;
assign LUT_2[22211] = 32'b00000000000000000110011001111100;
assign LUT_2[22212] = 32'b11111111111111111111000110001111;
assign LUT_2[22213] = 32'b11111111111111111011111110101000;
assign LUT_2[22214] = 32'b00000000000000000101111111001011;
assign LUT_2[22215] = 32'b00000000000000000010110111100100;
assign LUT_2[22216] = 32'b11111111111111111101011010000100;
assign LUT_2[22217] = 32'b11111111111111111010010010011101;
assign LUT_2[22218] = 32'b00000000000000000100010011000000;
assign LUT_2[22219] = 32'b00000000000000000001001011011001;
assign LUT_2[22220] = 32'b11111111111111111001110111101100;
assign LUT_2[22221] = 32'b11111111111111110110110000000101;
assign LUT_2[22222] = 32'b00000000000000000000110000101000;
assign LUT_2[22223] = 32'b11111111111111111101101001000001;
assign LUT_2[22224] = 32'b11111111111111111101001100110001;
assign LUT_2[22225] = 32'b11111111111111111010000101001010;
assign LUT_2[22226] = 32'b00000000000000000100000101101101;
assign LUT_2[22227] = 32'b00000000000000000000111110000110;
assign LUT_2[22228] = 32'b11111111111111111001101010011001;
assign LUT_2[22229] = 32'b11111111111111110110100010110010;
assign LUT_2[22230] = 32'b00000000000000000000100011010101;
assign LUT_2[22231] = 32'b11111111111111111101011011101110;
assign LUT_2[22232] = 32'b11111111111111110111111110001110;
assign LUT_2[22233] = 32'b11111111111111110100110110100111;
assign LUT_2[22234] = 32'b11111111111111111110110111001010;
assign LUT_2[22235] = 32'b11111111111111111011101111100011;
assign LUT_2[22236] = 32'b11111111111111110100011011110110;
assign LUT_2[22237] = 32'b11111111111111110001010100001111;
assign LUT_2[22238] = 32'b11111111111111111011010100110010;
assign LUT_2[22239] = 32'b11111111111111111000001101001011;
assign LUT_2[22240] = 32'b00000000000000000011000100010000;
assign LUT_2[22241] = 32'b11111111111111111111111100101001;
assign LUT_2[22242] = 32'b00000000000000001001111101001100;
assign LUT_2[22243] = 32'b00000000000000000110110101100101;
assign LUT_2[22244] = 32'b11111111111111111111100001111000;
assign LUT_2[22245] = 32'b11111111111111111100011010010001;
assign LUT_2[22246] = 32'b00000000000000000110011010110100;
assign LUT_2[22247] = 32'b00000000000000000011010011001101;
assign LUT_2[22248] = 32'b11111111111111111101110101101101;
assign LUT_2[22249] = 32'b11111111111111111010101110000110;
assign LUT_2[22250] = 32'b00000000000000000100101110101001;
assign LUT_2[22251] = 32'b00000000000000000001100111000010;
assign LUT_2[22252] = 32'b11111111111111111010010011010101;
assign LUT_2[22253] = 32'b11111111111111110111001011101110;
assign LUT_2[22254] = 32'b00000000000000000001001100010001;
assign LUT_2[22255] = 32'b11111111111111111110000100101010;
assign LUT_2[22256] = 32'b11111111111111111101101000011010;
assign LUT_2[22257] = 32'b11111111111111111010100000110011;
assign LUT_2[22258] = 32'b00000000000000000100100001010110;
assign LUT_2[22259] = 32'b00000000000000000001011001101111;
assign LUT_2[22260] = 32'b11111111111111111010000110000010;
assign LUT_2[22261] = 32'b11111111111111110110111110011011;
assign LUT_2[22262] = 32'b00000000000000000000111110111110;
assign LUT_2[22263] = 32'b11111111111111111101110111010111;
assign LUT_2[22264] = 32'b11111111111111111000011001110111;
assign LUT_2[22265] = 32'b11111111111111110101010010010000;
assign LUT_2[22266] = 32'b11111111111111111111010010110011;
assign LUT_2[22267] = 32'b11111111111111111100001011001100;
assign LUT_2[22268] = 32'b11111111111111110100110111011111;
assign LUT_2[22269] = 32'b11111111111111110001101111111000;
assign LUT_2[22270] = 32'b11111111111111111011110000011011;
assign LUT_2[22271] = 32'b11111111111111111000101000110100;
assign LUT_2[22272] = 32'b00000000000000001010001010011011;
assign LUT_2[22273] = 32'b00000000000000000111000010110100;
assign LUT_2[22274] = 32'b00000000000000010001000011010111;
assign LUT_2[22275] = 32'b00000000000000001101111011110000;
assign LUT_2[22276] = 32'b00000000000000000110101000000011;
assign LUT_2[22277] = 32'b00000000000000000011100000011100;
assign LUT_2[22278] = 32'b00000000000000001101100000111111;
assign LUT_2[22279] = 32'b00000000000000001010011001011000;
assign LUT_2[22280] = 32'b00000000000000000100111011111000;
assign LUT_2[22281] = 32'b00000000000000000001110100010001;
assign LUT_2[22282] = 32'b00000000000000001011110100110100;
assign LUT_2[22283] = 32'b00000000000000001000101101001101;
assign LUT_2[22284] = 32'b00000000000000000001011001100000;
assign LUT_2[22285] = 32'b11111111111111111110010001111001;
assign LUT_2[22286] = 32'b00000000000000001000010010011100;
assign LUT_2[22287] = 32'b00000000000000000101001010110101;
assign LUT_2[22288] = 32'b00000000000000000100101110100101;
assign LUT_2[22289] = 32'b00000000000000000001100110111110;
assign LUT_2[22290] = 32'b00000000000000001011100111100001;
assign LUT_2[22291] = 32'b00000000000000001000011111111010;
assign LUT_2[22292] = 32'b00000000000000000001001100001101;
assign LUT_2[22293] = 32'b11111111111111111110000100100110;
assign LUT_2[22294] = 32'b00000000000000001000000101001001;
assign LUT_2[22295] = 32'b00000000000000000100111101100010;
assign LUT_2[22296] = 32'b11111111111111111111100000000010;
assign LUT_2[22297] = 32'b11111111111111111100011000011011;
assign LUT_2[22298] = 32'b00000000000000000110011000111110;
assign LUT_2[22299] = 32'b00000000000000000011010001010111;
assign LUT_2[22300] = 32'b11111111111111111011111101101010;
assign LUT_2[22301] = 32'b11111111111111111000110110000011;
assign LUT_2[22302] = 32'b00000000000000000010110110100110;
assign LUT_2[22303] = 32'b11111111111111111111101110111111;
assign LUT_2[22304] = 32'b00000000000000001010100110000100;
assign LUT_2[22305] = 32'b00000000000000000111011110011101;
assign LUT_2[22306] = 32'b00000000000000010001011111000000;
assign LUT_2[22307] = 32'b00000000000000001110010111011001;
assign LUT_2[22308] = 32'b00000000000000000111000011101100;
assign LUT_2[22309] = 32'b00000000000000000011111100000101;
assign LUT_2[22310] = 32'b00000000000000001101111100101000;
assign LUT_2[22311] = 32'b00000000000000001010110101000001;
assign LUT_2[22312] = 32'b00000000000000000101010111100001;
assign LUT_2[22313] = 32'b00000000000000000010001111111010;
assign LUT_2[22314] = 32'b00000000000000001100010000011101;
assign LUT_2[22315] = 32'b00000000000000001001001000110110;
assign LUT_2[22316] = 32'b00000000000000000001110101001001;
assign LUT_2[22317] = 32'b11111111111111111110101101100010;
assign LUT_2[22318] = 32'b00000000000000001000101110000101;
assign LUT_2[22319] = 32'b00000000000000000101100110011110;
assign LUT_2[22320] = 32'b00000000000000000101001010001110;
assign LUT_2[22321] = 32'b00000000000000000010000010100111;
assign LUT_2[22322] = 32'b00000000000000001100000011001010;
assign LUT_2[22323] = 32'b00000000000000001000111011100011;
assign LUT_2[22324] = 32'b00000000000000000001100111110110;
assign LUT_2[22325] = 32'b11111111111111111110100000001111;
assign LUT_2[22326] = 32'b00000000000000001000100000110010;
assign LUT_2[22327] = 32'b00000000000000000101011001001011;
assign LUT_2[22328] = 32'b11111111111111111111111011101011;
assign LUT_2[22329] = 32'b11111111111111111100110100000100;
assign LUT_2[22330] = 32'b00000000000000000110110100100111;
assign LUT_2[22331] = 32'b00000000000000000011101101000000;
assign LUT_2[22332] = 32'b11111111111111111100011001010011;
assign LUT_2[22333] = 32'b11111111111111111001010001101100;
assign LUT_2[22334] = 32'b00000000000000000011010010001111;
assign LUT_2[22335] = 32'b00000000000000000000001010101000;
assign LUT_2[22336] = 32'b00000000000000000010010010111110;
assign LUT_2[22337] = 32'b11111111111111111111001011010111;
assign LUT_2[22338] = 32'b00000000000000001001001011111010;
assign LUT_2[22339] = 32'b00000000000000000110000100010011;
assign LUT_2[22340] = 32'b11111111111111111110110000100110;
assign LUT_2[22341] = 32'b11111111111111111011101000111111;
assign LUT_2[22342] = 32'b00000000000000000101101001100010;
assign LUT_2[22343] = 32'b00000000000000000010100001111011;
assign LUT_2[22344] = 32'b11111111111111111101000100011011;
assign LUT_2[22345] = 32'b11111111111111111001111100110100;
assign LUT_2[22346] = 32'b00000000000000000011111101010111;
assign LUT_2[22347] = 32'b00000000000000000000110101110000;
assign LUT_2[22348] = 32'b11111111111111111001100010000011;
assign LUT_2[22349] = 32'b11111111111111110110011010011100;
assign LUT_2[22350] = 32'b00000000000000000000011010111111;
assign LUT_2[22351] = 32'b11111111111111111101010011011000;
assign LUT_2[22352] = 32'b11111111111111111100110111001000;
assign LUT_2[22353] = 32'b11111111111111111001101111100001;
assign LUT_2[22354] = 32'b00000000000000000011110000000100;
assign LUT_2[22355] = 32'b00000000000000000000101000011101;
assign LUT_2[22356] = 32'b11111111111111111001010100110000;
assign LUT_2[22357] = 32'b11111111111111110110001101001001;
assign LUT_2[22358] = 32'b00000000000000000000001101101100;
assign LUT_2[22359] = 32'b11111111111111111101000110000101;
assign LUT_2[22360] = 32'b11111111111111110111101000100101;
assign LUT_2[22361] = 32'b11111111111111110100100000111110;
assign LUT_2[22362] = 32'b11111111111111111110100001100001;
assign LUT_2[22363] = 32'b11111111111111111011011001111010;
assign LUT_2[22364] = 32'b11111111111111110100000110001101;
assign LUT_2[22365] = 32'b11111111111111110000111110100110;
assign LUT_2[22366] = 32'b11111111111111111010111111001001;
assign LUT_2[22367] = 32'b11111111111111110111110111100010;
assign LUT_2[22368] = 32'b00000000000000000010101110100111;
assign LUT_2[22369] = 32'b11111111111111111111100111000000;
assign LUT_2[22370] = 32'b00000000000000001001100111100011;
assign LUT_2[22371] = 32'b00000000000000000110011111111100;
assign LUT_2[22372] = 32'b11111111111111111111001100001111;
assign LUT_2[22373] = 32'b11111111111111111100000100101000;
assign LUT_2[22374] = 32'b00000000000000000110000101001011;
assign LUT_2[22375] = 32'b00000000000000000010111101100100;
assign LUT_2[22376] = 32'b11111111111111111101100000000100;
assign LUT_2[22377] = 32'b11111111111111111010011000011101;
assign LUT_2[22378] = 32'b00000000000000000100011001000000;
assign LUT_2[22379] = 32'b00000000000000000001010001011001;
assign LUT_2[22380] = 32'b11111111111111111001111101101100;
assign LUT_2[22381] = 32'b11111111111111110110110110000101;
assign LUT_2[22382] = 32'b00000000000000000000110110101000;
assign LUT_2[22383] = 32'b11111111111111111101101111000001;
assign LUT_2[22384] = 32'b11111111111111111101010010110001;
assign LUT_2[22385] = 32'b11111111111111111010001011001010;
assign LUT_2[22386] = 32'b00000000000000000100001011101101;
assign LUT_2[22387] = 32'b00000000000000000001000100000110;
assign LUT_2[22388] = 32'b11111111111111111001110000011001;
assign LUT_2[22389] = 32'b11111111111111110110101000110010;
assign LUT_2[22390] = 32'b00000000000000000000101001010101;
assign LUT_2[22391] = 32'b11111111111111111101100001101110;
assign LUT_2[22392] = 32'b11111111111111111000000100001110;
assign LUT_2[22393] = 32'b11111111111111110100111100100111;
assign LUT_2[22394] = 32'b11111111111111111110111101001010;
assign LUT_2[22395] = 32'b11111111111111111011110101100011;
assign LUT_2[22396] = 32'b11111111111111110100100001110110;
assign LUT_2[22397] = 32'b11111111111111110001011010001111;
assign LUT_2[22398] = 32'b11111111111111111011011010110010;
assign LUT_2[22399] = 32'b11111111111111111000010011001011;
assign LUT_2[22400] = 32'b00000000000000001110011110101010;
assign LUT_2[22401] = 32'b00000000000000001011010111000011;
assign LUT_2[22402] = 32'b00000000000000010101010111100110;
assign LUT_2[22403] = 32'b00000000000000010010001111111111;
assign LUT_2[22404] = 32'b00000000000000001010111100010010;
assign LUT_2[22405] = 32'b00000000000000000111110100101011;
assign LUT_2[22406] = 32'b00000000000000010001110101001110;
assign LUT_2[22407] = 32'b00000000000000001110101101100111;
assign LUT_2[22408] = 32'b00000000000000001001010000000111;
assign LUT_2[22409] = 32'b00000000000000000110001000100000;
assign LUT_2[22410] = 32'b00000000000000010000001001000011;
assign LUT_2[22411] = 32'b00000000000000001101000001011100;
assign LUT_2[22412] = 32'b00000000000000000101101101101111;
assign LUT_2[22413] = 32'b00000000000000000010100110001000;
assign LUT_2[22414] = 32'b00000000000000001100100110101011;
assign LUT_2[22415] = 32'b00000000000000001001011111000100;
assign LUT_2[22416] = 32'b00000000000000001001000010110100;
assign LUT_2[22417] = 32'b00000000000000000101111011001101;
assign LUT_2[22418] = 32'b00000000000000001111111011110000;
assign LUT_2[22419] = 32'b00000000000000001100110100001001;
assign LUT_2[22420] = 32'b00000000000000000101100000011100;
assign LUT_2[22421] = 32'b00000000000000000010011000110101;
assign LUT_2[22422] = 32'b00000000000000001100011001011000;
assign LUT_2[22423] = 32'b00000000000000001001010001110001;
assign LUT_2[22424] = 32'b00000000000000000011110100010001;
assign LUT_2[22425] = 32'b00000000000000000000101100101010;
assign LUT_2[22426] = 32'b00000000000000001010101101001101;
assign LUT_2[22427] = 32'b00000000000000000111100101100110;
assign LUT_2[22428] = 32'b00000000000000000000010001111001;
assign LUT_2[22429] = 32'b11111111111111111101001010010010;
assign LUT_2[22430] = 32'b00000000000000000111001010110101;
assign LUT_2[22431] = 32'b00000000000000000100000011001110;
assign LUT_2[22432] = 32'b00000000000000001110111010010011;
assign LUT_2[22433] = 32'b00000000000000001011110010101100;
assign LUT_2[22434] = 32'b00000000000000010101110011001111;
assign LUT_2[22435] = 32'b00000000000000010010101011101000;
assign LUT_2[22436] = 32'b00000000000000001011010111111011;
assign LUT_2[22437] = 32'b00000000000000001000010000010100;
assign LUT_2[22438] = 32'b00000000000000010010010000110111;
assign LUT_2[22439] = 32'b00000000000000001111001001010000;
assign LUT_2[22440] = 32'b00000000000000001001101011110000;
assign LUT_2[22441] = 32'b00000000000000000110100100001001;
assign LUT_2[22442] = 32'b00000000000000010000100100101100;
assign LUT_2[22443] = 32'b00000000000000001101011101000101;
assign LUT_2[22444] = 32'b00000000000000000110001001011000;
assign LUT_2[22445] = 32'b00000000000000000011000001110001;
assign LUT_2[22446] = 32'b00000000000000001101000010010100;
assign LUT_2[22447] = 32'b00000000000000001001111010101101;
assign LUT_2[22448] = 32'b00000000000000001001011110011101;
assign LUT_2[22449] = 32'b00000000000000000110010110110110;
assign LUT_2[22450] = 32'b00000000000000010000010111011001;
assign LUT_2[22451] = 32'b00000000000000001101001111110010;
assign LUT_2[22452] = 32'b00000000000000000101111100000101;
assign LUT_2[22453] = 32'b00000000000000000010110100011110;
assign LUT_2[22454] = 32'b00000000000000001100110101000001;
assign LUT_2[22455] = 32'b00000000000000001001101101011010;
assign LUT_2[22456] = 32'b00000000000000000100001111111010;
assign LUT_2[22457] = 32'b00000000000000000001001000010011;
assign LUT_2[22458] = 32'b00000000000000001011001000110110;
assign LUT_2[22459] = 32'b00000000000000001000000001001111;
assign LUT_2[22460] = 32'b00000000000000000000101101100010;
assign LUT_2[22461] = 32'b11111111111111111101100101111011;
assign LUT_2[22462] = 32'b00000000000000000111100110011110;
assign LUT_2[22463] = 32'b00000000000000000100011110110111;
assign LUT_2[22464] = 32'b00000000000000000110100111001101;
assign LUT_2[22465] = 32'b00000000000000000011011111100110;
assign LUT_2[22466] = 32'b00000000000000001101100000001001;
assign LUT_2[22467] = 32'b00000000000000001010011000100010;
assign LUT_2[22468] = 32'b00000000000000000011000100110101;
assign LUT_2[22469] = 32'b11111111111111111111111101001110;
assign LUT_2[22470] = 32'b00000000000000001001111101110001;
assign LUT_2[22471] = 32'b00000000000000000110110110001010;
assign LUT_2[22472] = 32'b00000000000000000001011000101010;
assign LUT_2[22473] = 32'b11111111111111111110010001000011;
assign LUT_2[22474] = 32'b00000000000000001000010001100110;
assign LUT_2[22475] = 32'b00000000000000000101001001111111;
assign LUT_2[22476] = 32'b11111111111111111101110110010010;
assign LUT_2[22477] = 32'b11111111111111111010101110101011;
assign LUT_2[22478] = 32'b00000000000000000100101111001110;
assign LUT_2[22479] = 32'b00000000000000000001100111100111;
assign LUT_2[22480] = 32'b00000000000000000001001011010111;
assign LUT_2[22481] = 32'b11111111111111111110000011110000;
assign LUT_2[22482] = 32'b00000000000000001000000100010011;
assign LUT_2[22483] = 32'b00000000000000000100111100101100;
assign LUT_2[22484] = 32'b11111111111111111101101000111111;
assign LUT_2[22485] = 32'b11111111111111111010100001011000;
assign LUT_2[22486] = 32'b00000000000000000100100001111011;
assign LUT_2[22487] = 32'b00000000000000000001011010010100;
assign LUT_2[22488] = 32'b11111111111111111011111100110100;
assign LUT_2[22489] = 32'b11111111111111111000110101001101;
assign LUT_2[22490] = 32'b00000000000000000010110101110000;
assign LUT_2[22491] = 32'b11111111111111111111101110001001;
assign LUT_2[22492] = 32'b11111111111111111000011010011100;
assign LUT_2[22493] = 32'b11111111111111110101010010110101;
assign LUT_2[22494] = 32'b11111111111111111111010011011000;
assign LUT_2[22495] = 32'b11111111111111111100001011110001;
assign LUT_2[22496] = 32'b00000000000000000111000010110110;
assign LUT_2[22497] = 32'b00000000000000000011111011001111;
assign LUT_2[22498] = 32'b00000000000000001101111011110010;
assign LUT_2[22499] = 32'b00000000000000001010110100001011;
assign LUT_2[22500] = 32'b00000000000000000011100000011110;
assign LUT_2[22501] = 32'b00000000000000000000011000110111;
assign LUT_2[22502] = 32'b00000000000000001010011001011010;
assign LUT_2[22503] = 32'b00000000000000000111010001110011;
assign LUT_2[22504] = 32'b00000000000000000001110100010011;
assign LUT_2[22505] = 32'b11111111111111111110101100101100;
assign LUT_2[22506] = 32'b00000000000000001000101101001111;
assign LUT_2[22507] = 32'b00000000000000000101100101101000;
assign LUT_2[22508] = 32'b11111111111111111110010001111011;
assign LUT_2[22509] = 32'b11111111111111111011001010010100;
assign LUT_2[22510] = 32'b00000000000000000101001010110111;
assign LUT_2[22511] = 32'b00000000000000000010000011010000;
assign LUT_2[22512] = 32'b00000000000000000001100111000000;
assign LUT_2[22513] = 32'b11111111111111111110011111011001;
assign LUT_2[22514] = 32'b00000000000000001000011111111100;
assign LUT_2[22515] = 32'b00000000000000000101011000010101;
assign LUT_2[22516] = 32'b11111111111111111110000100101000;
assign LUT_2[22517] = 32'b11111111111111111010111101000001;
assign LUT_2[22518] = 32'b00000000000000000100111101100100;
assign LUT_2[22519] = 32'b00000000000000000001110101111101;
assign LUT_2[22520] = 32'b11111111111111111100011000011101;
assign LUT_2[22521] = 32'b11111111111111111001010000110110;
assign LUT_2[22522] = 32'b00000000000000000011010001011001;
assign LUT_2[22523] = 32'b00000000000000000000001001110010;
assign LUT_2[22524] = 32'b11111111111111111000110110000101;
assign LUT_2[22525] = 32'b11111111111111110101101110011110;
assign LUT_2[22526] = 32'b11111111111111111111101111000001;
assign LUT_2[22527] = 32'b11111111111111111100100111011010;
assign LUT_2[22528] = 32'b11111111111111110110100011111010;
assign LUT_2[22529] = 32'b11111111111111110011011100010011;
assign LUT_2[22530] = 32'b11111111111111111101011100110110;
assign LUT_2[22531] = 32'b11111111111111111010010101001111;
assign LUT_2[22532] = 32'b11111111111111110011000001100010;
assign LUT_2[22533] = 32'b11111111111111101111111001111011;
assign LUT_2[22534] = 32'b11111111111111111001111010011110;
assign LUT_2[22535] = 32'b11111111111111110110110010110111;
assign LUT_2[22536] = 32'b11111111111111110001010101010111;
assign LUT_2[22537] = 32'b11111111111111101110001101110000;
assign LUT_2[22538] = 32'b11111111111111111000001110010011;
assign LUT_2[22539] = 32'b11111111111111110101000110101100;
assign LUT_2[22540] = 32'b11111111111111101101110010111111;
assign LUT_2[22541] = 32'b11111111111111101010101011011000;
assign LUT_2[22542] = 32'b11111111111111110100101011111011;
assign LUT_2[22543] = 32'b11111111111111110001100100010100;
assign LUT_2[22544] = 32'b11111111111111110001001000000100;
assign LUT_2[22545] = 32'b11111111111111101110000000011101;
assign LUT_2[22546] = 32'b11111111111111111000000001000000;
assign LUT_2[22547] = 32'b11111111111111110100111001011001;
assign LUT_2[22548] = 32'b11111111111111101101100101101100;
assign LUT_2[22549] = 32'b11111111111111101010011110000101;
assign LUT_2[22550] = 32'b11111111111111110100011110101000;
assign LUT_2[22551] = 32'b11111111111111110001010111000001;
assign LUT_2[22552] = 32'b11111111111111101011111001100001;
assign LUT_2[22553] = 32'b11111111111111101000110001111010;
assign LUT_2[22554] = 32'b11111111111111110010110010011101;
assign LUT_2[22555] = 32'b11111111111111101111101010110110;
assign LUT_2[22556] = 32'b11111111111111101000010111001001;
assign LUT_2[22557] = 32'b11111111111111100101001111100010;
assign LUT_2[22558] = 32'b11111111111111101111010000000101;
assign LUT_2[22559] = 32'b11111111111111101100001000011110;
assign LUT_2[22560] = 32'b11111111111111110110111111100011;
assign LUT_2[22561] = 32'b11111111111111110011110111111100;
assign LUT_2[22562] = 32'b11111111111111111101111000011111;
assign LUT_2[22563] = 32'b11111111111111111010110000111000;
assign LUT_2[22564] = 32'b11111111111111110011011101001011;
assign LUT_2[22565] = 32'b11111111111111110000010101100100;
assign LUT_2[22566] = 32'b11111111111111111010010110000111;
assign LUT_2[22567] = 32'b11111111111111110111001110100000;
assign LUT_2[22568] = 32'b11111111111111110001110001000000;
assign LUT_2[22569] = 32'b11111111111111101110101001011001;
assign LUT_2[22570] = 32'b11111111111111111000101001111100;
assign LUT_2[22571] = 32'b11111111111111110101100010010101;
assign LUT_2[22572] = 32'b11111111111111101110001110101000;
assign LUT_2[22573] = 32'b11111111111111101011000111000001;
assign LUT_2[22574] = 32'b11111111111111110101000111100100;
assign LUT_2[22575] = 32'b11111111111111110001111111111101;
assign LUT_2[22576] = 32'b11111111111111110001100011101101;
assign LUT_2[22577] = 32'b11111111111111101110011100000110;
assign LUT_2[22578] = 32'b11111111111111111000011100101001;
assign LUT_2[22579] = 32'b11111111111111110101010101000010;
assign LUT_2[22580] = 32'b11111111111111101110000001010101;
assign LUT_2[22581] = 32'b11111111111111101010111001101110;
assign LUT_2[22582] = 32'b11111111111111110100111010010001;
assign LUT_2[22583] = 32'b11111111111111110001110010101010;
assign LUT_2[22584] = 32'b11111111111111101100010101001010;
assign LUT_2[22585] = 32'b11111111111111101001001101100011;
assign LUT_2[22586] = 32'b11111111111111110011001110000110;
assign LUT_2[22587] = 32'b11111111111111110000000110011111;
assign LUT_2[22588] = 32'b11111111111111101000110010110010;
assign LUT_2[22589] = 32'b11111111111111100101101011001011;
assign LUT_2[22590] = 32'b11111111111111101111101011101110;
assign LUT_2[22591] = 32'b11111111111111101100100100000111;
assign LUT_2[22592] = 32'b11111111111111101110101100011101;
assign LUT_2[22593] = 32'b11111111111111101011100100110110;
assign LUT_2[22594] = 32'b11111111111111110101100101011001;
assign LUT_2[22595] = 32'b11111111111111110010011101110010;
assign LUT_2[22596] = 32'b11111111111111101011001010000101;
assign LUT_2[22597] = 32'b11111111111111101000000010011110;
assign LUT_2[22598] = 32'b11111111111111110010000011000001;
assign LUT_2[22599] = 32'b11111111111111101110111011011010;
assign LUT_2[22600] = 32'b11111111111111101001011101111010;
assign LUT_2[22601] = 32'b11111111111111100110010110010011;
assign LUT_2[22602] = 32'b11111111111111110000010110110110;
assign LUT_2[22603] = 32'b11111111111111101101001111001111;
assign LUT_2[22604] = 32'b11111111111111100101111011100010;
assign LUT_2[22605] = 32'b11111111111111100010110011111011;
assign LUT_2[22606] = 32'b11111111111111101100110100011110;
assign LUT_2[22607] = 32'b11111111111111101001101100110111;
assign LUT_2[22608] = 32'b11111111111111101001010000100111;
assign LUT_2[22609] = 32'b11111111111111100110001001000000;
assign LUT_2[22610] = 32'b11111111111111110000001001100011;
assign LUT_2[22611] = 32'b11111111111111101101000001111100;
assign LUT_2[22612] = 32'b11111111111111100101101110001111;
assign LUT_2[22613] = 32'b11111111111111100010100110101000;
assign LUT_2[22614] = 32'b11111111111111101100100111001011;
assign LUT_2[22615] = 32'b11111111111111101001011111100100;
assign LUT_2[22616] = 32'b11111111111111100100000010000100;
assign LUT_2[22617] = 32'b11111111111111100000111010011101;
assign LUT_2[22618] = 32'b11111111111111101010111011000000;
assign LUT_2[22619] = 32'b11111111111111100111110011011001;
assign LUT_2[22620] = 32'b11111111111111100000011111101100;
assign LUT_2[22621] = 32'b11111111111111011101011000000101;
assign LUT_2[22622] = 32'b11111111111111100111011000101000;
assign LUT_2[22623] = 32'b11111111111111100100010001000001;
assign LUT_2[22624] = 32'b11111111111111101111001000000110;
assign LUT_2[22625] = 32'b11111111111111101100000000011111;
assign LUT_2[22626] = 32'b11111111111111110110000001000010;
assign LUT_2[22627] = 32'b11111111111111110010111001011011;
assign LUT_2[22628] = 32'b11111111111111101011100101101110;
assign LUT_2[22629] = 32'b11111111111111101000011110000111;
assign LUT_2[22630] = 32'b11111111111111110010011110101010;
assign LUT_2[22631] = 32'b11111111111111101111010111000011;
assign LUT_2[22632] = 32'b11111111111111101001111001100011;
assign LUT_2[22633] = 32'b11111111111111100110110001111100;
assign LUT_2[22634] = 32'b11111111111111110000110010011111;
assign LUT_2[22635] = 32'b11111111111111101101101010111000;
assign LUT_2[22636] = 32'b11111111111111100110010111001011;
assign LUT_2[22637] = 32'b11111111111111100011001111100100;
assign LUT_2[22638] = 32'b11111111111111101101010000000111;
assign LUT_2[22639] = 32'b11111111111111101010001000100000;
assign LUT_2[22640] = 32'b11111111111111101001101100010000;
assign LUT_2[22641] = 32'b11111111111111100110100100101001;
assign LUT_2[22642] = 32'b11111111111111110000100101001100;
assign LUT_2[22643] = 32'b11111111111111101101011101100101;
assign LUT_2[22644] = 32'b11111111111111100110001001111000;
assign LUT_2[22645] = 32'b11111111111111100011000010010001;
assign LUT_2[22646] = 32'b11111111111111101101000010110100;
assign LUT_2[22647] = 32'b11111111111111101001111011001101;
assign LUT_2[22648] = 32'b11111111111111100100011101101101;
assign LUT_2[22649] = 32'b11111111111111100001010110000110;
assign LUT_2[22650] = 32'b11111111111111101011010110101001;
assign LUT_2[22651] = 32'b11111111111111101000001111000010;
assign LUT_2[22652] = 32'b11111111111111100000111011010101;
assign LUT_2[22653] = 32'b11111111111111011101110011101110;
assign LUT_2[22654] = 32'b11111111111111100111110100010001;
assign LUT_2[22655] = 32'b11111111111111100100101100101010;
assign LUT_2[22656] = 32'b11111111111111111010111000001001;
assign LUT_2[22657] = 32'b11111111111111110111110000100010;
assign LUT_2[22658] = 32'b00000000000000000001110001000101;
assign LUT_2[22659] = 32'b11111111111111111110101001011110;
assign LUT_2[22660] = 32'b11111111111111110111010101110001;
assign LUT_2[22661] = 32'b11111111111111110100001110001010;
assign LUT_2[22662] = 32'b11111111111111111110001110101101;
assign LUT_2[22663] = 32'b11111111111111111011000111000110;
assign LUT_2[22664] = 32'b11111111111111110101101001100110;
assign LUT_2[22665] = 32'b11111111111111110010100001111111;
assign LUT_2[22666] = 32'b11111111111111111100100010100010;
assign LUT_2[22667] = 32'b11111111111111111001011010111011;
assign LUT_2[22668] = 32'b11111111111111110010000111001110;
assign LUT_2[22669] = 32'b11111111111111101110111111100111;
assign LUT_2[22670] = 32'b11111111111111111001000000001010;
assign LUT_2[22671] = 32'b11111111111111110101111000100011;
assign LUT_2[22672] = 32'b11111111111111110101011100010011;
assign LUT_2[22673] = 32'b11111111111111110010010100101100;
assign LUT_2[22674] = 32'b11111111111111111100010101001111;
assign LUT_2[22675] = 32'b11111111111111111001001101101000;
assign LUT_2[22676] = 32'b11111111111111110001111001111011;
assign LUT_2[22677] = 32'b11111111111111101110110010010100;
assign LUT_2[22678] = 32'b11111111111111111000110010110111;
assign LUT_2[22679] = 32'b11111111111111110101101011010000;
assign LUT_2[22680] = 32'b11111111111111110000001101110000;
assign LUT_2[22681] = 32'b11111111111111101101000110001001;
assign LUT_2[22682] = 32'b11111111111111110111000110101100;
assign LUT_2[22683] = 32'b11111111111111110011111111000101;
assign LUT_2[22684] = 32'b11111111111111101100101011011000;
assign LUT_2[22685] = 32'b11111111111111101001100011110001;
assign LUT_2[22686] = 32'b11111111111111110011100100010100;
assign LUT_2[22687] = 32'b11111111111111110000011100101101;
assign LUT_2[22688] = 32'b11111111111111111011010011110010;
assign LUT_2[22689] = 32'b11111111111111111000001100001011;
assign LUT_2[22690] = 32'b00000000000000000010001100101110;
assign LUT_2[22691] = 32'b11111111111111111111000101000111;
assign LUT_2[22692] = 32'b11111111111111110111110001011010;
assign LUT_2[22693] = 32'b11111111111111110100101001110011;
assign LUT_2[22694] = 32'b11111111111111111110101010010110;
assign LUT_2[22695] = 32'b11111111111111111011100010101111;
assign LUT_2[22696] = 32'b11111111111111110110000101001111;
assign LUT_2[22697] = 32'b11111111111111110010111101101000;
assign LUT_2[22698] = 32'b11111111111111111100111110001011;
assign LUT_2[22699] = 32'b11111111111111111001110110100100;
assign LUT_2[22700] = 32'b11111111111111110010100010110111;
assign LUT_2[22701] = 32'b11111111111111101111011011010000;
assign LUT_2[22702] = 32'b11111111111111111001011011110011;
assign LUT_2[22703] = 32'b11111111111111110110010100001100;
assign LUT_2[22704] = 32'b11111111111111110101110111111100;
assign LUT_2[22705] = 32'b11111111111111110010110000010101;
assign LUT_2[22706] = 32'b11111111111111111100110000111000;
assign LUT_2[22707] = 32'b11111111111111111001101001010001;
assign LUT_2[22708] = 32'b11111111111111110010010101100100;
assign LUT_2[22709] = 32'b11111111111111101111001101111101;
assign LUT_2[22710] = 32'b11111111111111111001001110100000;
assign LUT_2[22711] = 32'b11111111111111110110000110111001;
assign LUT_2[22712] = 32'b11111111111111110000101001011001;
assign LUT_2[22713] = 32'b11111111111111101101100001110010;
assign LUT_2[22714] = 32'b11111111111111110111100010010101;
assign LUT_2[22715] = 32'b11111111111111110100011010101110;
assign LUT_2[22716] = 32'b11111111111111101101000111000001;
assign LUT_2[22717] = 32'b11111111111111101001111111011010;
assign LUT_2[22718] = 32'b11111111111111110011111111111101;
assign LUT_2[22719] = 32'b11111111111111110000111000010110;
assign LUT_2[22720] = 32'b11111111111111110011000000101100;
assign LUT_2[22721] = 32'b11111111111111101111111001000101;
assign LUT_2[22722] = 32'b11111111111111111001111001101000;
assign LUT_2[22723] = 32'b11111111111111110110110010000001;
assign LUT_2[22724] = 32'b11111111111111101111011110010100;
assign LUT_2[22725] = 32'b11111111111111101100010110101101;
assign LUT_2[22726] = 32'b11111111111111110110010111010000;
assign LUT_2[22727] = 32'b11111111111111110011001111101001;
assign LUT_2[22728] = 32'b11111111111111101101110010001001;
assign LUT_2[22729] = 32'b11111111111111101010101010100010;
assign LUT_2[22730] = 32'b11111111111111110100101011000101;
assign LUT_2[22731] = 32'b11111111111111110001100011011110;
assign LUT_2[22732] = 32'b11111111111111101010001111110001;
assign LUT_2[22733] = 32'b11111111111111100111001000001010;
assign LUT_2[22734] = 32'b11111111111111110001001000101101;
assign LUT_2[22735] = 32'b11111111111111101110000001000110;
assign LUT_2[22736] = 32'b11111111111111101101100100110110;
assign LUT_2[22737] = 32'b11111111111111101010011101001111;
assign LUT_2[22738] = 32'b11111111111111110100011101110010;
assign LUT_2[22739] = 32'b11111111111111110001010110001011;
assign LUT_2[22740] = 32'b11111111111111101010000010011110;
assign LUT_2[22741] = 32'b11111111111111100110111010110111;
assign LUT_2[22742] = 32'b11111111111111110000111011011010;
assign LUT_2[22743] = 32'b11111111111111101101110011110011;
assign LUT_2[22744] = 32'b11111111111111101000010110010011;
assign LUT_2[22745] = 32'b11111111111111100101001110101100;
assign LUT_2[22746] = 32'b11111111111111101111001111001111;
assign LUT_2[22747] = 32'b11111111111111101100000111101000;
assign LUT_2[22748] = 32'b11111111111111100100110011111011;
assign LUT_2[22749] = 32'b11111111111111100001101100010100;
assign LUT_2[22750] = 32'b11111111111111101011101100110111;
assign LUT_2[22751] = 32'b11111111111111101000100101010000;
assign LUT_2[22752] = 32'b11111111111111110011011100010101;
assign LUT_2[22753] = 32'b11111111111111110000010100101110;
assign LUT_2[22754] = 32'b11111111111111111010010101010001;
assign LUT_2[22755] = 32'b11111111111111110111001101101010;
assign LUT_2[22756] = 32'b11111111111111101111111001111101;
assign LUT_2[22757] = 32'b11111111111111101100110010010110;
assign LUT_2[22758] = 32'b11111111111111110110110010111001;
assign LUT_2[22759] = 32'b11111111111111110011101011010010;
assign LUT_2[22760] = 32'b11111111111111101110001101110010;
assign LUT_2[22761] = 32'b11111111111111101011000110001011;
assign LUT_2[22762] = 32'b11111111111111110101000110101110;
assign LUT_2[22763] = 32'b11111111111111110001111111000111;
assign LUT_2[22764] = 32'b11111111111111101010101011011010;
assign LUT_2[22765] = 32'b11111111111111100111100011110011;
assign LUT_2[22766] = 32'b11111111111111110001100100010110;
assign LUT_2[22767] = 32'b11111111111111101110011100101111;
assign LUT_2[22768] = 32'b11111111111111101110000000011111;
assign LUT_2[22769] = 32'b11111111111111101010111000111000;
assign LUT_2[22770] = 32'b11111111111111110100111001011011;
assign LUT_2[22771] = 32'b11111111111111110001110001110100;
assign LUT_2[22772] = 32'b11111111111111101010011110000111;
assign LUT_2[22773] = 32'b11111111111111100111010110100000;
assign LUT_2[22774] = 32'b11111111111111110001010111000011;
assign LUT_2[22775] = 32'b11111111111111101110001111011100;
assign LUT_2[22776] = 32'b11111111111111101000110001111100;
assign LUT_2[22777] = 32'b11111111111111100101101010010101;
assign LUT_2[22778] = 32'b11111111111111101111101010111000;
assign LUT_2[22779] = 32'b11111111111111101100100011010001;
assign LUT_2[22780] = 32'b11111111111111100101001111100100;
assign LUT_2[22781] = 32'b11111111111111100010000111111101;
assign LUT_2[22782] = 32'b11111111111111101100001000100000;
assign LUT_2[22783] = 32'b11111111111111101001000000111001;
assign LUT_2[22784] = 32'b11111111111111111010100010100000;
assign LUT_2[22785] = 32'b11111111111111110111011010111001;
assign LUT_2[22786] = 32'b00000000000000000001011011011100;
assign LUT_2[22787] = 32'b11111111111111111110010011110101;
assign LUT_2[22788] = 32'b11111111111111110111000000001000;
assign LUT_2[22789] = 32'b11111111111111110011111000100001;
assign LUT_2[22790] = 32'b11111111111111111101111001000100;
assign LUT_2[22791] = 32'b11111111111111111010110001011101;
assign LUT_2[22792] = 32'b11111111111111110101010011111101;
assign LUT_2[22793] = 32'b11111111111111110010001100010110;
assign LUT_2[22794] = 32'b11111111111111111100001100111001;
assign LUT_2[22795] = 32'b11111111111111111001000101010010;
assign LUT_2[22796] = 32'b11111111111111110001110001100101;
assign LUT_2[22797] = 32'b11111111111111101110101001111110;
assign LUT_2[22798] = 32'b11111111111111111000101010100001;
assign LUT_2[22799] = 32'b11111111111111110101100010111010;
assign LUT_2[22800] = 32'b11111111111111110101000110101010;
assign LUT_2[22801] = 32'b11111111111111110001111111000011;
assign LUT_2[22802] = 32'b11111111111111111011111111100110;
assign LUT_2[22803] = 32'b11111111111111111000110111111111;
assign LUT_2[22804] = 32'b11111111111111110001100100010010;
assign LUT_2[22805] = 32'b11111111111111101110011100101011;
assign LUT_2[22806] = 32'b11111111111111111000011101001110;
assign LUT_2[22807] = 32'b11111111111111110101010101100111;
assign LUT_2[22808] = 32'b11111111111111101111111000000111;
assign LUT_2[22809] = 32'b11111111111111101100110000100000;
assign LUT_2[22810] = 32'b11111111111111110110110001000011;
assign LUT_2[22811] = 32'b11111111111111110011101001011100;
assign LUT_2[22812] = 32'b11111111111111101100010101101111;
assign LUT_2[22813] = 32'b11111111111111101001001110001000;
assign LUT_2[22814] = 32'b11111111111111110011001110101011;
assign LUT_2[22815] = 32'b11111111111111110000000111000100;
assign LUT_2[22816] = 32'b11111111111111111010111110001001;
assign LUT_2[22817] = 32'b11111111111111110111110110100010;
assign LUT_2[22818] = 32'b00000000000000000001110111000101;
assign LUT_2[22819] = 32'b11111111111111111110101111011110;
assign LUT_2[22820] = 32'b11111111111111110111011011110001;
assign LUT_2[22821] = 32'b11111111111111110100010100001010;
assign LUT_2[22822] = 32'b11111111111111111110010100101101;
assign LUT_2[22823] = 32'b11111111111111111011001101000110;
assign LUT_2[22824] = 32'b11111111111111110101101111100110;
assign LUT_2[22825] = 32'b11111111111111110010100111111111;
assign LUT_2[22826] = 32'b11111111111111111100101000100010;
assign LUT_2[22827] = 32'b11111111111111111001100000111011;
assign LUT_2[22828] = 32'b11111111111111110010001101001110;
assign LUT_2[22829] = 32'b11111111111111101111000101100111;
assign LUT_2[22830] = 32'b11111111111111111001000110001010;
assign LUT_2[22831] = 32'b11111111111111110101111110100011;
assign LUT_2[22832] = 32'b11111111111111110101100010010011;
assign LUT_2[22833] = 32'b11111111111111110010011010101100;
assign LUT_2[22834] = 32'b11111111111111111100011011001111;
assign LUT_2[22835] = 32'b11111111111111111001010011101000;
assign LUT_2[22836] = 32'b11111111111111110001111111111011;
assign LUT_2[22837] = 32'b11111111111111101110111000010100;
assign LUT_2[22838] = 32'b11111111111111111000111000110111;
assign LUT_2[22839] = 32'b11111111111111110101110001010000;
assign LUT_2[22840] = 32'b11111111111111110000010011110000;
assign LUT_2[22841] = 32'b11111111111111101101001100001001;
assign LUT_2[22842] = 32'b11111111111111110111001100101100;
assign LUT_2[22843] = 32'b11111111111111110100000101000101;
assign LUT_2[22844] = 32'b11111111111111101100110001011000;
assign LUT_2[22845] = 32'b11111111111111101001101001110001;
assign LUT_2[22846] = 32'b11111111111111110011101010010100;
assign LUT_2[22847] = 32'b11111111111111110000100010101101;
assign LUT_2[22848] = 32'b11111111111111110010101011000011;
assign LUT_2[22849] = 32'b11111111111111101111100011011100;
assign LUT_2[22850] = 32'b11111111111111111001100011111111;
assign LUT_2[22851] = 32'b11111111111111110110011100011000;
assign LUT_2[22852] = 32'b11111111111111101111001000101011;
assign LUT_2[22853] = 32'b11111111111111101100000001000100;
assign LUT_2[22854] = 32'b11111111111111110110000001100111;
assign LUT_2[22855] = 32'b11111111111111110010111010000000;
assign LUT_2[22856] = 32'b11111111111111101101011100100000;
assign LUT_2[22857] = 32'b11111111111111101010010100111001;
assign LUT_2[22858] = 32'b11111111111111110100010101011100;
assign LUT_2[22859] = 32'b11111111111111110001001101110101;
assign LUT_2[22860] = 32'b11111111111111101001111010001000;
assign LUT_2[22861] = 32'b11111111111111100110110010100001;
assign LUT_2[22862] = 32'b11111111111111110000110011000100;
assign LUT_2[22863] = 32'b11111111111111101101101011011101;
assign LUT_2[22864] = 32'b11111111111111101101001111001101;
assign LUT_2[22865] = 32'b11111111111111101010000111100110;
assign LUT_2[22866] = 32'b11111111111111110100001000001001;
assign LUT_2[22867] = 32'b11111111111111110001000000100010;
assign LUT_2[22868] = 32'b11111111111111101001101100110101;
assign LUT_2[22869] = 32'b11111111111111100110100101001110;
assign LUT_2[22870] = 32'b11111111111111110000100101110001;
assign LUT_2[22871] = 32'b11111111111111101101011110001010;
assign LUT_2[22872] = 32'b11111111111111101000000000101010;
assign LUT_2[22873] = 32'b11111111111111100100111001000011;
assign LUT_2[22874] = 32'b11111111111111101110111001100110;
assign LUT_2[22875] = 32'b11111111111111101011110001111111;
assign LUT_2[22876] = 32'b11111111111111100100011110010010;
assign LUT_2[22877] = 32'b11111111111111100001010110101011;
assign LUT_2[22878] = 32'b11111111111111101011010111001110;
assign LUT_2[22879] = 32'b11111111111111101000001111100111;
assign LUT_2[22880] = 32'b11111111111111110011000110101100;
assign LUT_2[22881] = 32'b11111111111111101111111111000101;
assign LUT_2[22882] = 32'b11111111111111111001111111101000;
assign LUT_2[22883] = 32'b11111111111111110110111000000001;
assign LUT_2[22884] = 32'b11111111111111101111100100010100;
assign LUT_2[22885] = 32'b11111111111111101100011100101101;
assign LUT_2[22886] = 32'b11111111111111110110011101010000;
assign LUT_2[22887] = 32'b11111111111111110011010101101001;
assign LUT_2[22888] = 32'b11111111111111101101111000001001;
assign LUT_2[22889] = 32'b11111111111111101010110000100010;
assign LUT_2[22890] = 32'b11111111111111110100110001000101;
assign LUT_2[22891] = 32'b11111111111111110001101001011110;
assign LUT_2[22892] = 32'b11111111111111101010010101110001;
assign LUT_2[22893] = 32'b11111111111111100111001110001010;
assign LUT_2[22894] = 32'b11111111111111110001001110101101;
assign LUT_2[22895] = 32'b11111111111111101110000111000110;
assign LUT_2[22896] = 32'b11111111111111101101101010110110;
assign LUT_2[22897] = 32'b11111111111111101010100011001111;
assign LUT_2[22898] = 32'b11111111111111110100100011110010;
assign LUT_2[22899] = 32'b11111111111111110001011100001011;
assign LUT_2[22900] = 32'b11111111111111101010001000011110;
assign LUT_2[22901] = 32'b11111111111111100111000000110111;
assign LUT_2[22902] = 32'b11111111111111110001000001011010;
assign LUT_2[22903] = 32'b11111111111111101101111001110011;
assign LUT_2[22904] = 32'b11111111111111101000011100010011;
assign LUT_2[22905] = 32'b11111111111111100101010100101100;
assign LUT_2[22906] = 32'b11111111111111101111010101001111;
assign LUT_2[22907] = 32'b11111111111111101100001101101000;
assign LUT_2[22908] = 32'b11111111111111100100111001111011;
assign LUT_2[22909] = 32'b11111111111111100001110010010100;
assign LUT_2[22910] = 32'b11111111111111101011110010110111;
assign LUT_2[22911] = 32'b11111111111111101000101011010000;
assign LUT_2[22912] = 32'b11111111111111111110110110101111;
assign LUT_2[22913] = 32'b11111111111111111011101111001000;
assign LUT_2[22914] = 32'b00000000000000000101101111101011;
assign LUT_2[22915] = 32'b00000000000000000010101000000100;
assign LUT_2[22916] = 32'b11111111111111111011010100010111;
assign LUT_2[22917] = 32'b11111111111111111000001100110000;
assign LUT_2[22918] = 32'b00000000000000000010001101010011;
assign LUT_2[22919] = 32'b11111111111111111111000101101100;
assign LUT_2[22920] = 32'b11111111111111111001101000001100;
assign LUT_2[22921] = 32'b11111111111111110110100000100101;
assign LUT_2[22922] = 32'b00000000000000000000100001001000;
assign LUT_2[22923] = 32'b11111111111111111101011001100001;
assign LUT_2[22924] = 32'b11111111111111110110000101110100;
assign LUT_2[22925] = 32'b11111111111111110010111110001101;
assign LUT_2[22926] = 32'b11111111111111111100111110110000;
assign LUT_2[22927] = 32'b11111111111111111001110111001001;
assign LUT_2[22928] = 32'b11111111111111111001011010111001;
assign LUT_2[22929] = 32'b11111111111111110110010011010010;
assign LUT_2[22930] = 32'b00000000000000000000010011110101;
assign LUT_2[22931] = 32'b11111111111111111101001100001110;
assign LUT_2[22932] = 32'b11111111111111110101111000100001;
assign LUT_2[22933] = 32'b11111111111111110010110000111010;
assign LUT_2[22934] = 32'b11111111111111111100110001011101;
assign LUT_2[22935] = 32'b11111111111111111001101001110110;
assign LUT_2[22936] = 32'b11111111111111110100001100010110;
assign LUT_2[22937] = 32'b11111111111111110001000100101111;
assign LUT_2[22938] = 32'b11111111111111111011000101010010;
assign LUT_2[22939] = 32'b11111111111111110111111101101011;
assign LUT_2[22940] = 32'b11111111111111110000101001111110;
assign LUT_2[22941] = 32'b11111111111111101101100010010111;
assign LUT_2[22942] = 32'b11111111111111110111100010111010;
assign LUT_2[22943] = 32'b11111111111111110100011011010011;
assign LUT_2[22944] = 32'b11111111111111111111010010011000;
assign LUT_2[22945] = 32'b11111111111111111100001010110001;
assign LUT_2[22946] = 32'b00000000000000000110001011010100;
assign LUT_2[22947] = 32'b00000000000000000011000011101101;
assign LUT_2[22948] = 32'b11111111111111111011110000000000;
assign LUT_2[22949] = 32'b11111111111111111000101000011001;
assign LUT_2[22950] = 32'b00000000000000000010101000111100;
assign LUT_2[22951] = 32'b11111111111111111111100001010101;
assign LUT_2[22952] = 32'b11111111111111111010000011110101;
assign LUT_2[22953] = 32'b11111111111111110110111100001110;
assign LUT_2[22954] = 32'b00000000000000000000111100110001;
assign LUT_2[22955] = 32'b11111111111111111101110101001010;
assign LUT_2[22956] = 32'b11111111111111110110100001011101;
assign LUT_2[22957] = 32'b11111111111111110011011001110110;
assign LUT_2[22958] = 32'b11111111111111111101011010011001;
assign LUT_2[22959] = 32'b11111111111111111010010010110010;
assign LUT_2[22960] = 32'b11111111111111111001110110100010;
assign LUT_2[22961] = 32'b11111111111111110110101110111011;
assign LUT_2[22962] = 32'b00000000000000000000101111011110;
assign LUT_2[22963] = 32'b11111111111111111101100111110111;
assign LUT_2[22964] = 32'b11111111111111110110010100001010;
assign LUT_2[22965] = 32'b11111111111111110011001100100011;
assign LUT_2[22966] = 32'b11111111111111111101001101000110;
assign LUT_2[22967] = 32'b11111111111111111010000101011111;
assign LUT_2[22968] = 32'b11111111111111110100100111111111;
assign LUT_2[22969] = 32'b11111111111111110001100000011000;
assign LUT_2[22970] = 32'b11111111111111111011100000111011;
assign LUT_2[22971] = 32'b11111111111111111000011001010100;
assign LUT_2[22972] = 32'b11111111111111110001000101100111;
assign LUT_2[22973] = 32'b11111111111111101101111110000000;
assign LUT_2[22974] = 32'b11111111111111110111111110100011;
assign LUT_2[22975] = 32'b11111111111111110100110110111100;
assign LUT_2[22976] = 32'b11111111111111110110111111010010;
assign LUT_2[22977] = 32'b11111111111111110011110111101011;
assign LUT_2[22978] = 32'b11111111111111111101111000001110;
assign LUT_2[22979] = 32'b11111111111111111010110000100111;
assign LUT_2[22980] = 32'b11111111111111110011011100111010;
assign LUT_2[22981] = 32'b11111111111111110000010101010011;
assign LUT_2[22982] = 32'b11111111111111111010010101110110;
assign LUT_2[22983] = 32'b11111111111111110111001110001111;
assign LUT_2[22984] = 32'b11111111111111110001110000101111;
assign LUT_2[22985] = 32'b11111111111111101110101001001000;
assign LUT_2[22986] = 32'b11111111111111111000101001101011;
assign LUT_2[22987] = 32'b11111111111111110101100010000100;
assign LUT_2[22988] = 32'b11111111111111101110001110010111;
assign LUT_2[22989] = 32'b11111111111111101011000110110000;
assign LUT_2[22990] = 32'b11111111111111110101000111010011;
assign LUT_2[22991] = 32'b11111111111111110001111111101100;
assign LUT_2[22992] = 32'b11111111111111110001100011011100;
assign LUT_2[22993] = 32'b11111111111111101110011011110101;
assign LUT_2[22994] = 32'b11111111111111111000011100011000;
assign LUT_2[22995] = 32'b11111111111111110101010100110001;
assign LUT_2[22996] = 32'b11111111111111101110000001000100;
assign LUT_2[22997] = 32'b11111111111111101010111001011101;
assign LUT_2[22998] = 32'b11111111111111110100111010000000;
assign LUT_2[22999] = 32'b11111111111111110001110010011001;
assign LUT_2[23000] = 32'b11111111111111101100010100111001;
assign LUT_2[23001] = 32'b11111111111111101001001101010010;
assign LUT_2[23002] = 32'b11111111111111110011001101110101;
assign LUT_2[23003] = 32'b11111111111111110000000110001110;
assign LUT_2[23004] = 32'b11111111111111101000110010100001;
assign LUT_2[23005] = 32'b11111111111111100101101010111010;
assign LUT_2[23006] = 32'b11111111111111101111101011011101;
assign LUT_2[23007] = 32'b11111111111111101100100011110110;
assign LUT_2[23008] = 32'b11111111111111110111011010111011;
assign LUT_2[23009] = 32'b11111111111111110100010011010100;
assign LUT_2[23010] = 32'b11111111111111111110010011110111;
assign LUT_2[23011] = 32'b11111111111111111011001100010000;
assign LUT_2[23012] = 32'b11111111111111110011111000100011;
assign LUT_2[23013] = 32'b11111111111111110000110000111100;
assign LUT_2[23014] = 32'b11111111111111111010110001011111;
assign LUT_2[23015] = 32'b11111111111111110111101001111000;
assign LUT_2[23016] = 32'b11111111111111110010001100011000;
assign LUT_2[23017] = 32'b11111111111111101111000100110001;
assign LUT_2[23018] = 32'b11111111111111111001000101010100;
assign LUT_2[23019] = 32'b11111111111111110101111101101101;
assign LUT_2[23020] = 32'b11111111111111101110101010000000;
assign LUT_2[23021] = 32'b11111111111111101011100010011001;
assign LUT_2[23022] = 32'b11111111111111110101100010111100;
assign LUT_2[23023] = 32'b11111111111111110010011011010101;
assign LUT_2[23024] = 32'b11111111111111110001111111000101;
assign LUT_2[23025] = 32'b11111111111111101110110111011110;
assign LUT_2[23026] = 32'b11111111111111111000111000000001;
assign LUT_2[23027] = 32'b11111111111111110101110000011010;
assign LUT_2[23028] = 32'b11111111111111101110011100101101;
assign LUT_2[23029] = 32'b11111111111111101011010101000110;
assign LUT_2[23030] = 32'b11111111111111110101010101101001;
assign LUT_2[23031] = 32'b11111111111111110010001110000010;
assign LUT_2[23032] = 32'b11111111111111101100110000100010;
assign LUT_2[23033] = 32'b11111111111111101001101000111011;
assign LUT_2[23034] = 32'b11111111111111110011101001011110;
assign LUT_2[23035] = 32'b11111111111111110000100001110111;
assign LUT_2[23036] = 32'b11111111111111101001001110001010;
assign LUT_2[23037] = 32'b11111111111111100110000110100011;
assign LUT_2[23038] = 32'b11111111111111110000000111000110;
assign LUT_2[23039] = 32'b11111111111111101100111111011111;
assign LUT_2[23040] = 32'b11111111111111111011010101101100;
assign LUT_2[23041] = 32'b11111111111111111000001110000101;
assign LUT_2[23042] = 32'b00000000000000000010001110101000;
assign LUT_2[23043] = 32'b11111111111111111111000111000001;
assign LUT_2[23044] = 32'b11111111111111110111110011010100;
assign LUT_2[23045] = 32'b11111111111111110100101011101101;
assign LUT_2[23046] = 32'b11111111111111111110101100010000;
assign LUT_2[23047] = 32'b11111111111111111011100100101001;
assign LUT_2[23048] = 32'b11111111111111110110000111001001;
assign LUT_2[23049] = 32'b11111111111111110010111111100010;
assign LUT_2[23050] = 32'b11111111111111111101000000000101;
assign LUT_2[23051] = 32'b11111111111111111001111000011110;
assign LUT_2[23052] = 32'b11111111111111110010100100110001;
assign LUT_2[23053] = 32'b11111111111111101111011101001010;
assign LUT_2[23054] = 32'b11111111111111111001011101101101;
assign LUT_2[23055] = 32'b11111111111111110110010110000110;
assign LUT_2[23056] = 32'b11111111111111110101111001110110;
assign LUT_2[23057] = 32'b11111111111111110010110010001111;
assign LUT_2[23058] = 32'b11111111111111111100110010110010;
assign LUT_2[23059] = 32'b11111111111111111001101011001011;
assign LUT_2[23060] = 32'b11111111111111110010010111011110;
assign LUT_2[23061] = 32'b11111111111111101111001111110111;
assign LUT_2[23062] = 32'b11111111111111111001010000011010;
assign LUT_2[23063] = 32'b11111111111111110110001000110011;
assign LUT_2[23064] = 32'b11111111111111110000101011010011;
assign LUT_2[23065] = 32'b11111111111111101101100011101100;
assign LUT_2[23066] = 32'b11111111111111110111100100001111;
assign LUT_2[23067] = 32'b11111111111111110100011100101000;
assign LUT_2[23068] = 32'b11111111111111101101001000111011;
assign LUT_2[23069] = 32'b11111111111111101010000001010100;
assign LUT_2[23070] = 32'b11111111111111110100000001110111;
assign LUT_2[23071] = 32'b11111111111111110000111010010000;
assign LUT_2[23072] = 32'b11111111111111111011110001010101;
assign LUT_2[23073] = 32'b11111111111111111000101001101110;
assign LUT_2[23074] = 32'b00000000000000000010101010010001;
assign LUT_2[23075] = 32'b11111111111111111111100010101010;
assign LUT_2[23076] = 32'b11111111111111111000001110111101;
assign LUT_2[23077] = 32'b11111111111111110101000111010110;
assign LUT_2[23078] = 32'b11111111111111111111000111111001;
assign LUT_2[23079] = 32'b11111111111111111100000000010010;
assign LUT_2[23080] = 32'b11111111111111110110100010110010;
assign LUT_2[23081] = 32'b11111111111111110011011011001011;
assign LUT_2[23082] = 32'b11111111111111111101011011101110;
assign LUT_2[23083] = 32'b11111111111111111010010100000111;
assign LUT_2[23084] = 32'b11111111111111110011000000011010;
assign LUT_2[23085] = 32'b11111111111111101111111000110011;
assign LUT_2[23086] = 32'b11111111111111111001111001010110;
assign LUT_2[23087] = 32'b11111111111111110110110001101111;
assign LUT_2[23088] = 32'b11111111111111110110010101011111;
assign LUT_2[23089] = 32'b11111111111111110011001101111000;
assign LUT_2[23090] = 32'b11111111111111111101001110011011;
assign LUT_2[23091] = 32'b11111111111111111010000110110100;
assign LUT_2[23092] = 32'b11111111111111110010110011000111;
assign LUT_2[23093] = 32'b11111111111111101111101011100000;
assign LUT_2[23094] = 32'b11111111111111111001101100000011;
assign LUT_2[23095] = 32'b11111111111111110110100100011100;
assign LUT_2[23096] = 32'b11111111111111110001000110111100;
assign LUT_2[23097] = 32'b11111111111111101101111111010101;
assign LUT_2[23098] = 32'b11111111111111110111111111111000;
assign LUT_2[23099] = 32'b11111111111111110100111000010001;
assign LUT_2[23100] = 32'b11111111111111101101100100100100;
assign LUT_2[23101] = 32'b11111111111111101010011100111101;
assign LUT_2[23102] = 32'b11111111111111110100011101100000;
assign LUT_2[23103] = 32'b11111111111111110001010101111001;
assign LUT_2[23104] = 32'b11111111111111110011011110001111;
assign LUT_2[23105] = 32'b11111111111111110000010110101000;
assign LUT_2[23106] = 32'b11111111111111111010010111001011;
assign LUT_2[23107] = 32'b11111111111111110111001111100100;
assign LUT_2[23108] = 32'b11111111111111101111111011110111;
assign LUT_2[23109] = 32'b11111111111111101100110100010000;
assign LUT_2[23110] = 32'b11111111111111110110110100110011;
assign LUT_2[23111] = 32'b11111111111111110011101101001100;
assign LUT_2[23112] = 32'b11111111111111101110001111101100;
assign LUT_2[23113] = 32'b11111111111111101011001000000101;
assign LUT_2[23114] = 32'b11111111111111110101001000101000;
assign LUT_2[23115] = 32'b11111111111111110010000001000001;
assign LUT_2[23116] = 32'b11111111111111101010101101010100;
assign LUT_2[23117] = 32'b11111111111111100111100101101101;
assign LUT_2[23118] = 32'b11111111111111110001100110010000;
assign LUT_2[23119] = 32'b11111111111111101110011110101001;
assign LUT_2[23120] = 32'b11111111111111101110000010011001;
assign LUT_2[23121] = 32'b11111111111111101010111010110010;
assign LUT_2[23122] = 32'b11111111111111110100111011010101;
assign LUT_2[23123] = 32'b11111111111111110001110011101110;
assign LUT_2[23124] = 32'b11111111111111101010100000000001;
assign LUT_2[23125] = 32'b11111111111111100111011000011010;
assign LUT_2[23126] = 32'b11111111111111110001011000111101;
assign LUT_2[23127] = 32'b11111111111111101110010001010110;
assign LUT_2[23128] = 32'b11111111111111101000110011110110;
assign LUT_2[23129] = 32'b11111111111111100101101100001111;
assign LUT_2[23130] = 32'b11111111111111101111101100110010;
assign LUT_2[23131] = 32'b11111111111111101100100101001011;
assign LUT_2[23132] = 32'b11111111111111100101010001011110;
assign LUT_2[23133] = 32'b11111111111111100010001001110111;
assign LUT_2[23134] = 32'b11111111111111101100001010011010;
assign LUT_2[23135] = 32'b11111111111111101001000010110011;
assign LUT_2[23136] = 32'b11111111111111110011111001111000;
assign LUT_2[23137] = 32'b11111111111111110000110010010001;
assign LUT_2[23138] = 32'b11111111111111111010110010110100;
assign LUT_2[23139] = 32'b11111111111111110111101011001101;
assign LUT_2[23140] = 32'b11111111111111110000010111100000;
assign LUT_2[23141] = 32'b11111111111111101101001111111001;
assign LUT_2[23142] = 32'b11111111111111110111010000011100;
assign LUT_2[23143] = 32'b11111111111111110100001000110101;
assign LUT_2[23144] = 32'b11111111111111101110101011010101;
assign LUT_2[23145] = 32'b11111111111111101011100011101110;
assign LUT_2[23146] = 32'b11111111111111110101100100010001;
assign LUT_2[23147] = 32'b11111111111111110010011100101010;
assign LUT_2[23148] = 32'b11111111111111101011001000111101;
assign LUT_2[23149] = 32'b11111111111111101000000001010110;
assign LUT_2[23150] = 32'b11111111111111110010000001111001;
assign LUT_2[23151] = 32'b11111111111111101110111010010010;
assign LUT_2[23152] = 32'b11111111111111101110011110000010;
assign LUT_2[23153] = 32'b11111111111111101011010110011011;
assign LUT_2[23154] = 32'b11111111111111110101010110111110;
assign LUT_2[23155] = 32'b11111111111111110010001111010111;
assign LUT_2[23156] = 32'b11111111111111101010111011101010;
assign LUT_2[23157] = 32'b11111111111111100111110100000011;
assign LUT_2[23158] = 32'b11111111111111110001110100100110;
assign LUT_2[23159] = 32'b11111111111111101110101100111111;
assign LUT_2[23160] = 32'b11111111111111101001001111011111;
assign LUT_2[23161] = 32'b11111111111111100110000111111000;
assign LUT_2[23162] = 32'b11111111111111110000001000011011;
assign LUT_2[23163] = 32'b11111111111111101101000000110100;
assign LUT_2[23164] = 32'b11111111111111100101101101000111;
assign LUT_2[23165] = 32'b11111111111111100010100101100000;
assign LUT_2[23166] = 32'b11111111111111101100100110000011;
assign LUT_2[23167] = 32'b11111111111111101001011110011100;
assign LUT_2[23168] = 32'b11111111111111111111101001111011;
assign LUT_2[23169] = 32'b11111111111111111100100010010100;
assign LUT_2[23170] = 32'b00000000000000000110100010110111;
assign LUT_2[23171] = 32'b00000000000000000011011011010000;
assign LUT_2[23172] = 32'b11111111111111111100000111100011;
assign LUT_2[23173] = 32'b11111111111111111000111111111100;
assign LUT_2[23174] = 32'b00000000000000000011000000011111;
assign LUT_2[23175] = 32'b11111111111111111111111000111000;
assign LUT_2[23176] = 32'b11111111111111111010011011011000;
assign LUT_2[23177] = 32'b11111111111111110111010011110001;
assign LUT_2[23178] = 32'b00000000000000000001010100010100;
assign LUT_2[23179] = 32'b11111111111111111110001100101101;
assign LUT_2[23180] = 32'b11111111111111110110111001000000;
assign LUT_2[23181] = 32'b11111111111111110011110001011001;
assign LUT_2[23182] = 32'b11111111111111111101110001111100;
assign LUT_2[23183] = 32'b11111111111111111010101010010101;
assign LUT_2[23184] = 32'b11111111111111111010001110000101;
assign LUT_2[23185] = 32'b11111111111111110111000110011110;
assign LUT_2[23186] = 32'b00000000000000000001000111000001;
assign LUT_2[23187] = 32'b11111111111111111101111111011010;
assign LUT_2[23188] = 32'b11111111111111110110101011101101;
assign LUT_2[23189] = 32'b11111111111111110011100100000110;
assign LUT_2[23190] = 32'b11111111111111111101100100101001;
assign LUT_2[23191] = 32'b11111111111111111010011101000010;
assign LUT_2[23192] = 32'b11111111111111110100111111100010;
assign LUT_2[23193] = 32'b11111111111111110001110111111011;
assign LUT_2[23194] = 32'b11111111111111111011111000011110;
assign LUT_2[23195] = 32'b11111111111111111000110000110111;
assign LUT_2[23196] = 32'b11111111111111110001011101001010;
assign LUT_2[23197] = 32'b11111111111111101110010101100011;
assign LUT_2[23198] = 32'b11111111111111111000010110000110;
assign LUT_2[23199] = 32'b11111111111111110101001110011111;
assign LUT_2[23200] = 32'b00000000000000000000000101100100;
assign LUT_2[23201] = 32'b11111111111111111100111101111101;
assign LUT_2[23202] = 32'b00000000000000000110111110100000;
assign LUT_2[23203] = 32'b00000000000000000011110110111001;
assign LUT_2[23204] = 32'b11111111111111111100100011001100;
assign LUT_2[23205] = 32'b11111111111111111001011011100101;
assign LUT_2[23206] = 32'b00000000000000000011011100001000;
assign LUT_2[23207] = 32'b00000000000000000000010100100001;
assign LUT_2[23208] = 32'b11111111111111111010110111000001;
assign LUT_2[23209] = 32'b11111111111111110111101111011010;
assign LUT_2[23210] = 32'b00000000000000000001101111111101;
assign LUT_2[23211] = 32'b11111111111111111110101000010110;
assign LUT_2[23212] = 32'b11111111111111110111010100101001;
assign LUT_2[23213] = 32'b11111111111111110100001101000010;
assign LUT_2[23214] = 32'b11111111111111111110001101100101;
assign LUT_2[23215] = 32'b11111111111111111011000101111110;
assign LUT_2[23216] = 32'b11111111111111111010101001101110;
assign LUT_2[23217] = 32'b11111111111111110111100010000111;
assign LUT_2[23218] = 32'b00000000000000000001100010101010;
assign LUT_2[23219] = 32'b11111111111111111110011011000011;
assign LUT_2[23220] = 32'b11111111111111110111000111010110;
assign LUT_2[23221] = 32'b11111111111111110011111111101111;
assign LUT_2[23222] = 32'b11111111111111111110000000010010;
assign LUT_2[23223] = 32'b11111111111111111010111000101011;
assign LUT_2[23224] = 32'b11111111111111110101011011001011;
assign LUT_2[23225] = 32'b11111111111111110010010011100100;
assign LUT_2[23226] = 32'b11111111111111111100010100000111;
assign LUT_2[23227] = 32'b11111111111111111001001100100000;
assign LUT_2[23228] = 32'b11111111111111110001111000110011;
assign LUT_2[23229] = 32'b11111111111111101110110001001100;
assign LUT_2[23230] = 32'b11111111111111111000110001101111;
assign LUT_2[23231] = 32'b11111111111111110101101010001000;
assign LUT_2[23232] = 32'b11111111111111110111110010011110;
assign LUT_2[23233] = 32'b11111111111111110100101010110111;
assign LUT_2[23234] = 32'b11111111111111111110101011011010;
assign LUT_2[23235] = 32'b11111111111111111011100011110011;
assign LUT_2[23236] = 32'b11111111111111110100010000000110;
assign LUT_2[23237] = 32'b11111111111111110001001000011111;
assign LUT_2[23238] = 32'b11111111111111111011001001000010;
assign LUT_2[23239] = 32'b11111111111111111000000001011011;
assign LUT_2[23240] = 32'b11111111111111110010100011111011;
assign LUT_2[23241] = 32'b11111111111111101111011100010100;
assign LUT_2[23242] = 32'b11111111111111111001011100110111;
assign LUT_2[23243] = 32'b11111111111111110110010101010000;
assign LUT_2[23244] = 32'b11111111111111101111000001100011;
assign LUT_2[23245] = 32'b11111111111111101011111001111100;
assign LUT_2[23246] = 32'b11111111111111110101111010011111;
assign LUT_2[23247] = 32'b11111111111111110010110010111000;
assign LUT_2[23248] = 32'b11111111111111110010010110101000;
assign LUT_2[23249] = 32'b11111111111111101111001111000001;
assign LUT_2[23250] = 32'b11111111111111111001001111100100;
assign LUT_2[23251] = 32'b11111111111111110110000111111101;
assign LUT_2[23252] = 32'b11111111111111101110110100010000;
assign LUT_2[23253] = 32'b11111111111111101011101100101001;
assign LUT_2[23254] = 32'b11111111111111110101101101001100;
assign LUT_2[23255] = 32'b11111111111111110010100101100101;
assign LUT_2[23256] = 32'b11111111111111101101001000000101;
assign LUT_2[23257] = 32'b11111111111111101010000000011110;
assign LUT_2[23258] = 32'b11111111111111110100000001000001;
assign LUT_2[23259] = 32'b11111111111111110000111001011010;
assign LUT_2[23260] = 32'b11111111111111101001100101101101;
assign LUT_2[23261] = 32'b11111111111111100110011110000110;
assign LUT_2[23262] = 32'b11111111111111110000011110101001;
assign LUT_2[23263] = 32'b11111111111111101101010111000010;
assign LUT_2[23264] = 32'b11111111111111111000001110000111;
assign LUT_2[23265] = 32'b11111111111111110101000110100000;
assign LUT_2[23266] = 32'b11111111111111111111000111000011;
assign LUT_2[23267] = 32'b11111111111111111011111111011100;
assign LUT_2[23268] = 32'b11111111111111110100101011101111;
assign LUT_2[23269] = 32'b11111111111111110001100100001000;
assign LUT_2[23270] = 32'b11111111111111111011100100101011;
assign LUT_2[23271] = 32'b11111111111111111000011101000100;
assign LUT_2[23272] = 32'b11111111111111110010111111100100;
assign LUT_2[23273] = 32'b11111111111111101111110111111101;
assign LUT_2[23274] = 32'b11111111111111111001111000100000;
assign LUT_2[23275] = 32'b11111111111111110110110000111001;
assign LUT_2[23276] = 32'b11111111111111101111011101001100;
assign LUT_2[23277] = 32'b11111111111111101100010101100101;
assign LUT_2[23278] = 32'b11111111111111110110010110001000;
assign LUT_2[23279] = 32'b11111111111111110011001110100001;
assign LUT_2[23280] = 32'b11111111111111110010110010010001;
assign LUT_2[23281] = 32'b11111111111111101111101010101010;
assign LUT_2[23282] = 32'b11111111111111111001101011001101;
assign LUT_2[23283] = 32'b11111111111111110110100011100110;
assign LUT_2[23284] = 32'b11111111111111101111001111111001;
assign LUT_2[23285] = 32'b11111111111111101100001000010010;
assign LUT_2[23286] = 32'b11111111111111110110001000110101;
assign LUT_2[23287] = 32'b11111111111111110011000001001110;
assign LUT_2[23288] = 32'b11111111111111101101100011101110;
assign LUT_2[23289] = 32'b11111111111111101010011100000111;
assign LUT_2[23290] = 32'b11111111111111110100011100101010;
assign LUT_2[23291] = 32'b11111111111111110001010101000011;
assign LUT_2[23292] = 32'b11111111111111101010000001010110;
assign LUT_2[23293] = 32'b11111111111111100110111001101111;
assign LUT_2[23294] = 32'b11111111111111110000111010010010;
assign LUT_2[23295] = 32'b11111111111111101101110010101011;
assign LUT_2[23296] = 32'b11111111111111111111010100010010;
assign LUT_2[23297] = 32'b11111111111111111100001100101011;
assign LUT_2[23298] = 32'b00000000000000000110001101001110;
assign LUT_2[23299] = 32'b00000000000000000011000101100111;
assign LUT_2[23300] = 32'b11111111111111111011110001111010;
assign LUT_2[23301] = 32'b11111111111111111000101010010011;
assign LUT_2[23302] = 32'b00000000000000000010101010110110;
assign LUT_2[23303] = 32'b11111111111111111111100011001111;
assign LUT_2[23304] = 32'b11111111111111111010000101101111;
assign LUT_2[23305] = 32'b11111111111111110110111110001000;
assign LUT_2[23306] = 32'b00000000000000000000111110101011;
assign LUT_2[23307] = 32'b11111111111111111101110111000100;
assign LUT_2[23308] = 32'b11111111111111110110100011010111;
assign LUT_2[23309] = 32'b11111111111111110011011011110000;
assign LUT_2[23310] = 32'b11111111111111111101011100010011;
assign LUT_2[23311] = 32'b11111111111111111010010100101100;
assign LUT_2[23312] = 32'b11111111111111111001111000011100;
assign LUT_2[23313] = 32'b11111111111111110110110000110101;
assign LUT_2[23314] = 32'b00000000000000000000110001011000;
assign LUT_2[23315] = 32'b11111111111111111101101001110001;
assign LUT_2[23316] = 32'b11111111111111110110010110000100;
assign LUT_2[23317] = 32'b11111111111111110011001110011101;
assign LUT_2[23318] = 32'b11111111111111111101001111000000;
assign LUT_2[23319] = 32'b11111111111111111010000111011001;
assign LUT_2[23320] = 32'b11111111111111110100101001111001;
assign LUT_2[23321] = 32'b11111111111111110001100010010010;
assign LUT_2[23322] = 32'b11111111111111111011100010110101;
assign LUT_2[23323] = 32'b11111111111111111000011011001110;
assign LUT_2[23324] = 32'b11111111111111110001000111100001;
assign LUT_2[23325] = 32'b11111111111111101101111111111010;
assign LUT_2[23326] = 32'b11111111111111111000000000011101;
assign LUT_2[23327] = 32'b11111111111111110100111000110110;
assign LUT_2[23328] = 32'b11111111111111111111101111111011;
assign LUT_2[23329] = 32'b11111111111111111100101000010100;
assign LUT_2[23330] = 32'b00000000000000000110101000110111;
assign LUT_2[23331] = 32'b00000000000000000011100001010000;
assign LUT_2[23332] = 32'b11111111111111111100001101100011;
assign LUT_2[23333] = 32'b11111111111111111001000101111100;
assign LUT_2[23334] = 32'b00000000000000000011000110011111;
assign LUT_2[23335] = 32'b11111111111111111111111110111000;
assign LUT_2[23336] = 32'b11111111111111111010100001011000;
assign LUT_2[23337] = 32'b11111111111111110111011001110001;
assign LUT_2[23338] = 32'b00000000000000000001011010010100;
assign LUT_2[23339] = 32'b11111111111111111110010010101101;
assign LUT_2[23340] = 32'b11111111111111110110111111000000;
assign LUT_2[23341] = 32'b11111111111111110011110111011001;
assign LUT_2[23342] = 32'b11111111111111111101110111111100;
assign LUT_2[23343] = 32'b11111111111111111010110000010101;
assign LUT_2[23344] = 32'b11111111111111111010010100000101;
assign LUT_2[23345] = 32'b11111111111111110111001100011110;
assign LUT_2[23346] = 32'b00000000000000000001001101000001;
assign LUT_2[23347] = 32'b11111111111111111110000101011010;
assign LUT_2[23348] = 32'b11111111111111110110110001101101;
assign LUT_2[23349] = 32'b11111111111111110011101010000110;
assign LUT_2[23350] = 32'b11111111111111111101101010101001;
assign LUT_2[23351] = 32'b11111111111111111010100011000010;
assign LUT_2[23352] = 32'b11111111111111110101000101100010;
assign LUT_2[23353] = 32'b11111111111111110001111101111011;
assign LUT_2[23354] = 32'b11111111111111111011111110011110;
assign LUT_2[23355] = 32'b11111111111111111000110110110111;
assign LUT_2[23356] = 32'b11111111111111110001100011001010;
assign LUT_2[23357] = 32'b11111111111111101110011011100011;
assign LUT_2[23358] = 32'b11111111111111111000011100000110;
assign LUT_2[23359] = 32'b11111111111111110101010100011111;
assign LUT_2[23360] = 32'b11111111111111110111011100110101;
assign LUT_2[23361] = 32'b11111111111111110100010101001110;
assign LUT_2[23362] = 32'b11111111111111111110010101110001;
assign LUT_2[23363] = 32'b11111111111111111011001110001010;
assign LUT_2[23364] = 32'b11111111111111110011111010011101;
assign LUT_2[23365] = 32'b11111111111111110000110010110110;
assign LUT_2[23366] = 32'b11111111111111111010110011011001;
assign LUT_2[23367] = 32'b11111111111111110111101011110010;
assign LUT_2[23368] = 32'b11111111111111110010001110010010;
assign LUT_2[23369] = 32'b11111111111111101111000110101011;
assign LUT_2[23370] = 32'b11111111111111111001000111001110;
assign LUT_2[23371] = 32'b11111111111111110101111111100111;
assign LUT_2[23372] = 32'b11111111111111101110101011111010;
assign LUT_2[23373] = 32'b11111111111111101011100100010011;
assign LUT_2[23374] = 32'b11111111111111110101100100110110;
assign LUT_2[23375] = 32'b11111111111111110010011101001111;
assign LUT_2[23376] = 32'b11111111111111110010000000111111;
assign LUT_2[23377] = 32'b11111111111111101110111001011000;
assign LUT_2[23378] = 32'b11111111111111111000111001111011;
assign LUT_2[23379] = 32'b11111111111111110101110010010100;
assign LUT_2[23380] = 32'b11111111111111101110011110100111;
assign LUT_2[23381] = 32'b11111111111111101011010111000000;
assign LUT_2[23382] = 32'b11111111111111110101010111100011;
assign LUT_2[23383] = 32'b11111111111111110010001111111100;
assign LUT_2[23384] = 32'b11111111111111101100110010011100;
assign LUT_2[23385] = 32'b11111111111111101001101010110101;
assign LUT_2[23386] = 32'b11111111111111110011101011011000;
assign LUT_2[23387] = 32'b11111111111111110000100011110001;
assign LUT_2[23388] = 32'b11111111111111101001010000000100;
assign LUT_2[23389] = 32'b11111111111111100110001000011101;
assign LUT_2[23390] = 32'b11111111111111110000001001000000;
assign LUT_2[23391] = 32'b11111111111111101101000001011001;
assign LUT_2[23392] = 32'b11111111111111110111111000011110;
assign LUT_2[23393] = 32'b11111111111111110100110000110111;
assign LUT_2[23394] = 32'b11111111111111111110110001011010;
assign LUT_2[23395] = 32'b11111111111111111011101001110011;
assign LUT_2[23396] = 32'b11111111111111110100010110000110;
assign LUT_2[23397] = 32'b11111111111111110001001110011111;
assign LUT_2[23398] = 32'b11111111111111111011001111000010;
assign LUT_2[23399] = 32'b11111111111111111000000111011011;
assign LUT_2[23400] = 32'b11111111111111110010101001111011;
assign LUT_2[23401] = 32'b11111111111111101111100010010100;
assign LUT_2[23402] = 32'b11111111111111111001100010110111;
assign LUT_2[23403] = 32'b11111111111111110110011011010000;
assign LUT_2[23404] = 32'b11111111111111101111000111100011;
assign LUT_2[23405] = 32'b11111111111111101011111111111100;
assign LUT_2[23406] = 32'b11111111111111110110000000011111;
assign LUT_2[23407] = 32'b11111111111111110010111000111000;
assign LUT_2[23408] = 32'b11111111111111110010011100101000;
assign LUT_2[23409] = 32'b11111111111111101111010101000001;
assign LUT_2[23410] = 32'b11111111111111111001010101100100;
assign LUT_2[23411] = 32'b11111111111111110110001101111101;
assign LUT_2[23412] = 32'b11111111111111101110111010010000;
assign LUT_2[23413] = 32'b11111111111111101011110010101001;
assign LUT_2[23414] = 32'b11111111111111110101110011001100;
assign LUT_2[23415] = 32'b11111111111111110010101011100101;
assign LUT_2[23416] = 32'b11111111111111101101001110000101;
assign LUT_2[23417] = 32'b11111111111111101010000110011110;
assign LUT_2[23418] = 32'b11111111111111110100000111000001;
assign LUT_2[23419] = 32'b11111111111111110000111111011010;
assign LUT_2[23420] = 32'b11111111111111101001101011101101;
assign LUT_2[23421] = 32'b11111111111111100110100100000110;
assign LUT_2[23422] = 32'b11111111111111110000100100101001;
assign LUT_2[23423] = 32'b11111111111111101101011101000010;
assign LUT_2[23424] = 32'b00000000000000000011101000100001;
assign LUT_2[23425] = 32'b00000000000000000000100000111010;
assign LUT_2[23426] = 32'b00000000000000001010100001011101;
assign LUT_2[23427] = 32'b00000000000000000111011001110110;
assign LUT_2[23428] = 32'b00000000000000000000000110001001;
assign LUT_2[23429] = 32'b11111111111111111100111110100010;
assign LUT_2[23430] = 32'b00000000000000000110111111000101;
assign LUT_2[23431] = 32'b00000000000000000011110111011110;
assign LUT_2[23432] = 32'b11111111111111111110011001111110;
assign LUT_2[23433] = 32'b11111111111111111011010010010111;
assign LUT_2[23434] = 32'b00000000000000000101010010111010;
assign LUT_2[23435] = 32'b00000000000000000010001011010011;
assign LUT_2[23436] = 32'b11111111111111111010110111100110;
assign LUT_2[23437] = 32'b11111111111111110111101111111111;
assign LUT_2[23438] = 32'b00000000000000000001110000100010;
assign LUT_2[23439] = 32'b11111111111111111110101000111011;
assign LUT_2[23440] = 32'b11111111111111111110001100101011;
assign LUT_2[23441] = 32'b11111111111111111011000101000100;
assign LUT_2[23442] = 32'b00000000000000000101000101100111;
assign LUT_2[23443] = 32'b00000000000000000001111110000000;
assign LUT_2[23444] = 32'b11111111111111111010101010010011;
assign LUT_2[23445] = 32'b11111111111111110111100010101100;
assign LUT_2[23446] = 32'b00000000000000000001100011001111;
assign LUT_2[23447] = 32'b11111111111111111110011011101000;
assign LUT_2[23448] = 32'b11111111111111111000111110001000;
assign LUT_2[23449] = 32'b11111111111111110101110110100001;
assign LUT_2[23450] = 32'b11111111111111111111110111000100;
assign LUT_2[23451] = 32'b11111111111111111100101111011101;
assign LUT_2[23452] = 32'b11111111111111110101011011110000;
assign LUT_2[23453] = 32'b11111111111111110010010100001001;
assign LUT_2[23454] = 32'b11111111111111111100010100101100;
assign LUT_2[23455] = 32'b11111111111111111001001101000101;
assign LUT_2[23456] = 32'b00000000000000000100000100001010;
assign LUT_2[23457] = 32'b00000000000000000000111100100011;
assign LUT_2[23458] = 32'b00000000000000001010111101000110;
assign LUT_2[23459] = 32'b00000000000000000111110101011111;
assign LUT_2[23460] = 32'b00000000000000000000100001110010;
assign LUT_2[23461] = 32'b11111111111111111101011010001011;
assign LUT_2[23462] = 32'b00000000000000000111011010101110;
assign LUT_2[23463] = 32'b00000000000000000100010011000111;
assign LUT_2[23464] = 32'b11111111111111111110110101100111;
assign LUT_2[23465] = 32'b11111111111111111011101110000000;
assign LUT_2[23466] = 32'b00000000000000000101101110100011;
assign LUT_2[23467] = 32'b00000000000000000010100110111100;
assign LUT_2[23468] = 32'b11111111111111111011010011001111;
assign LUT_2[23469] = 32'b11111111111111111000001011101000;
assign LUT_2[23470] = 32'b00000000000000000010001100001011;
assign LUT_2[23471] = 32'b11111111111111111111000100100100;
assign LUT_2[23472] = 32'b11111111111111111110101000010100;
assign LUT_2[23473] = 32'b11111111111111111011100000101101;
assign LUT_2[23474] = 32'b00000000000000000101100001010000;
assign LUT_2[23475] = 32'b00000000000000000010011001101001;
assign LUT_2[23476] = 32'b11111111111111111011000101111100;
assign LUT_2[23477] = 32'b11111111111111110111111110010101;
assign LUT_2[23478] = 32'b00000000000000000001111110111000;
assign LUT_2[23479] = 32'b11111111111111111110110111010001;
assign LUT_2[23480] = 32'b11111111111111111001011001110001;
assign LUT_2[23481] = 32'b11111111111111110110010010001010;
assign LUT_2[23482] = 32'b00000000000000000000010010101101;
assign LUT_2[23483] = 32'b11111111111111111101001011000110;
assign LUT_2[23484] = 32'b11111111111111110101110111011001;
assign LUT_2[23485] = 32'b11111111111111110010101111110010;
assign LUT_2[23486] = 32'b11111111111111111100110000010101;
assign LUT_2[23487] = 32'b11111111111111111001101000101110;
assign LUT_2[23488] = 32'b11111111111111111011110001000100;
assign LUT_2[23489] = 32'b11111111111111111000101001011101;
assign LUT_2[23490] = 32'b00000000000000000010101010000000;
assign LUT_2[23491] = 32'b11111111111111111111100010011001;
assign LUT_2[23492] = 32'b11111111111111111000001110101100;
assign LUT_2[23493] = 32'b11111111111111110101000111000101;
assign LUT_2[23494] = 32'b11111111111111111111000111101000;
assign LUT_2[23495] = 32'b11111111111111111100000000000001;
assign LUT_2[23496] = 32'b11111111111111110110100010100001;
assign LUT_2[23497] = 32'b11111111111111110011011010111010;
assign LUT_2[23498] = 32'b11111111111111111101011011011101;
assign LUT_2[23499] = 32'b11111111111111111010010011110110;
assign LUT_2[23500] = 32'b11111111111111110011000000001001;
assign LUT_2[23501] = 32'b11111111111111101111111000100010;
assign LUT_2[23502] = 32'b11111111111111111001111001000101;
assign LUT_2[23503] = 32'b11111111111111110110110001011110;
assign LUT_2[23504] = 32'b11111111111111110110010101001110;
assign LUT_2[23505] = 32'b11111111111111110011001101100111;
assign LUT_2[23506] = 32'b11111111111111111101001110001010;
assign LUT_2[23507] = 32'b11111111111111111010000110100011;
assign LUT_2[23508] = 32'b11111111111111110010110010110110;
assign LUT_2[23509] = 32'b11111111111111101111101011001111;
assign LUT_2[23510] = 32'b11111111111111111001101011110010;
assign LUT_2[23511] = 32'b11111111111111110110100100001011;
assign LUT_2[23512] = 32'b11111111111111110001000110101011;
assign LUT_2[23513] = 32'b11111111111111101101111111000100;
assign LUT_2[23514] = 32'b11111111111111110111111111100111;
assign LUT_2[23515] = 32'b11111111111111110100111000000000;
assign LUT_2[23516] = 32'b11111111111111101101100100010011;
assign LUT_2[23517] = 32'b11111111111111101010011100101100;
assign LUT_2[23518] = 32'b11111111111111110100011101001111;
assign LUT_2[23519] = 32'b11111111111111110001010101101000;
assign LUT_2[23520] = 32'b11111111111111111100001100101101;
assign LUT_2[23521] = 32'b11111111111111111001000101000110;
assign LUT_2[23522] = 32'b00000000000000000011000101101001;
assign LUT_2[23523] = 32'b11111111111111111111111110000010;
assign LUT_2[23524] = 32'b11111111111111111000101010010101;
assign LUT_2[23525] = 32'b11111111111111110101100010101110;
assign LUT_2[23526] = 32'b11111111111111111111100011010001;
assign LUT_2[23527] = 32'b11111111111111111100011011101010;
assign LUT_2[23528] = 32'b11111111111111110110111110001010;
assign LUT_2[23529] = 32'b11111111111111110011110110100011;
assign LUT_2[23530] = 32'b11111111111111111101110111000110;
assign LUT_2[23531] = 32'b11111111111111111010101111011111;
assign LUT_2[23532] = 32'b11111111111111110011011011110010;
assign LUT_2[23533] = 32'b11111111111111110000010100001011;
assign LUT_2[23534] = 32'b11111111111111111010010100101110;
assign LUT_2[23535] = 32'b11111111111111110111001101000111;
assign LUT_2[23536] = 32'b11111111111111110110110000110111;
assign LUT_2[23537] = 32'b11111111111111110011101001010000;
assign LUT_2[23538] = 32'b11111111111111111101101001110011;
assign LUT_2[23539] = 32'b11111111111111111010100010001100;
assign LUT_2[23540] = 32'b11111111111111110011001110011111;
assign LUT_2[23541] = 32'b11111111111111110000000110111000;
assign LUT_2[23542] = 32'b11111111111111111010000111011011;
assign LUT_2[23543] = 32'b11111111111111110110111111110100;
assign LUT_2[23544] = 32'b11111111111111110001100010010100;
assign LUT_2[23545] = 32'b11111111111111101110011010101101;
assign LUT_2[23546] = 32'b11111111111111111000011011010000;
assign LUT_2[23547] = 32'b11111111111111110101010011101001;
assign LUT_2[23548] = 32'b11111111111111101101111111111100;
assign LUT_2[23549] = 32'b11111111111111101010111000010101;
assign LUT_2[23550] = 32'b11111111111111110100111000111000;
assign LUT_2[23551] = 32'b11111111111111110001110001010001;
assign LUT_2[23552] = 32'b11111111111111111101001111111111;
assign LUT_2[23553] = 32'b11111111111111111010001000011000;
assign LUT_2[23554] = 32'b00000000000000000100001000111011;
assign LUT_2[23555] = 32'b00000000000000000001000001010100;
assign LUT_2[23556] = 32'b11111111111111111001101101100111;
assign LUT_2[23557] = 32'b11111111111111110110100110000000;
assign LUT_2[23558] = 32'b00000000000000000000100110100011;
assign LUT_2[23559] = 32'b11111111111111111101011110111100;
assign LUT_2[23560] = 32'b11111111111111111000000001011100;
assign LUT_2[23561] = 32'b11111111111111110100111001110101;
assign LUT_2[23562] = 32'b11111111111111111110111010011000;
assign LUT_2[23563] = 32'b11111111111111111011110010110001;
assign LUT_2[23564] = 32'b11111111111111110100011111000100;
assign LUT_2[23565] = 32'b11111111111111110001010111011101;
assign LUT_2[23566] = 32'b11111111111111111011011000000000;
assign LUT_2[23567] = 32'b11111111111111111000010000011001;
assign LUT_2[23568] = 32'b11111111111111110111110100001001;
assign LUT_2[23569] = 32'b11111111111111110100101100100010;
assign LUT_2[23570] = 32'b11111111111111111110101101000101;
assign LUT_2[23571] = 32'b11111111111111111011100101011110;
assign LUT_2[23572] = 32'b11111111111111110100010001110001;
assign LUT_2[23573] = 32'b11111111111111110001001010001010;
assign LUT_2[23574] = 32'b11111111111111111011001010101101;
assign LUT_2[23575] = 32'b11111111111111111000000011000110;
assign LUT_2[23576] = 32'b11111111111111110010100101100110;
assign LUT_2[23577] = 32'b11111111111111101111011101111111;
assign LUT_2[23578] = 32'b11111111111111111001011110100010;
assign LUT_2[23579] = 32'b11111111111111110110010110111011;
assign LUT_2[23580] = 32'b11111111111111101111000011001110;
assign LUT_2[23581] = 32'b11111111111111101011111011100111;
assign LUT_2[23582] = 32'b11111111111111110101111100001010;
assign LUT_2[23583] = 32'b11111111111111110010110100100011;
assign LUT_2[23584] = 32'b11111111111111111101101011101000;
assign LUT_2[23585] = 32'b11111111111111111010100100000001;
assign LUT_2[23586] = 32'b00000000000000000100100100100100;
assign LUT_2[23587] = 32'b00000000000000000001011100111101;
assign LUT_2[23588] = 32'b11111111111111111010001001010000;
assign LUT_2[23589] = 32'b11111111111111110111000001101001;
assign LUT_2[23590] = 32'b00000000000000000001000010001100;
assign LUT_2[23591] = 32'b11111111111111111101111010100101;
assign LUT_2[23592] = 32'b11111111111111111000011101000101;
assign LUT_2[23593] = 32'b11111111111111110101010101011110;
assign LUT_2[23594] = 32'b11111111111111111111010110000001;
assign LUT_2[23595] = 32'b11111111111111111100001110011010;
assign LUT_2[23596] = 32'b11111111111111110100111010101101;
assign LUT_2[23597] = 32'b11111111111111110001110011000110;
assign LUT_2[23598] = 32'b11111111111111111011110011101001;
assign LUT_2[23599] = 32'b11111111111111111000101100000010;
assign LUT_2[23600] = 32'b11111111111111111000001111110010;
assign LUT_2[23601] = 32'b11111111111111110101001000001011;
assign LUT_2[23602] = 32'b11111111111111111111001000101110;
assign LUT_2[23603] = 32'b11111111111111111100000001000111;
assign LUT_2[23604] = 32'b11111111111111110100101101011010;
assign LUT_2[23605] = 32'b11111111111111110001100101110011;
assign LUT_2[23606] = 32'b11111111111111111011100110010110;
assign LUT_2[23607] = 32'b11111111111111111000011110101111;
assign LUT_2[23608] = 32'b11111111111111110011000001001111;
assign LUT_2[23609] = 32'b11111111111111101111111001101000;
assign LUT_2[23610] = 32'b11111111111111111001111010001011;
assign LUT_2[23611] = 32'b11111111111111110110110010100100;
assign LUT_2[23612] = 32'b11111111111111101111011110110111;
assign LUT_2[23613] = 32'b11111111111111101100010111010000;
assign LUT_2[23614] = 32'b11111111111111110110010111110011;
assign LUT_2[23615] = 32'b11111111111111110011010000001100;
assign LUT_2[23616] = 32'b11111111111111110101011000100010;
assign LUT_2[23617] = 32'b11111111111111110010010000111011;
assign LUT_2[23618] = 32'b11111111111111111100010001011110;
assign LUT_2[23619] = 32'b11111111111111111001001001110111;
assign LUT_2[23620] = 32'b11111111111111110001110110001010;
assign LUT_2[23621] = 32'b11111111111111101110101110100011;
assign LUT_2[23622] = 32'b11111111111111111000101111000110;
assign LUT_2[23623] = 32'b11111111111111110101100111011111;
assign LUT_2[23624] = 32'b11111111111111110000001001111111;
assign LUT_2[23625] = 32'b11111111111111101101000010011000;
assign LUT_2[23626] = 32'b11111111111111110111000010111011;
assign LUT_2[23627] = 32'b11111111111111110011111011010100;
assign LUT_2[23628] = 32'b11111111111111101100100111100111;
assign LUT_2[23629] = 32'b11111111111111101001100000000000;
assign LUT_2[23630] = 32'b11111111111111110011100000100011;
assign LUT_2[23631] = 32'b11111111111111110000011000111100;
assign LUT_2[23632] = 32'b11111111111111101111111100101100;
assign LUT_2[23633] = 32'b11111111111111101100110101000101;
assign LUT_2[23634] = 32'b11111111111111110110110101101000;
assign LUT_2[23635] = 32'b11111111111111110011101110000001;
assign LUT_2[23636] = 32'b11111111111111101100011010010100;
assign LUT_2[23637] = 32'b11111111111111101001010010101101;
assign LUT_2[23638] = 32'b11111111111111110011010011010000;
assign LUT_2[23639] = 32'b11111111111111110000001011101001;
assign LUT_2[23640] = 32'b11111111111111101010101110001001;
assign LUT_2[23641] = 32'b11111111111111100111100110100010;
assign LUT_2[23642] = 32'b11111111111111110001100111000101;
assign LUT_2[23643] = 32'b11111111111111101110011111011110;
assign LUT_2[23644] = 32'b11111111111111100111001011110001;
assign LUT_2[23645] = 32'b11111111111111100100000100001010;
assign LUT_2[23646] = 32'b11111111111111101110000100101101;
assign LUT_2[23647] = 32'b11111111111111101010111101000110;
assign LUT_2[23648] = 32'b11111111111111110101110100001011;
assign LUT_2[23649] = 32'b11111111111111110010101100100100;
assign LUT_2[23650] = 32'b11111111111111111100101101000111;
assign LUT_2[23651] = 32'b11111111111111111001100101100000;
assign LUT_2[23652] = 32'b11111111111111110010010001110011;
assign LUT_2[23653] = 32'b11111111111111101111001010001100;
assign LUT_2[23654] = 32'b11111111111111111001001010101111;
assign LUT_2[23655] = 32'b11111111111111110110000011001000;
assign LUT_2[23656] = 32'b11111111111111110000100101101000;
assign LUT_2[23657] = 32'b11111111111111101101011110000001;
assign LUT_2[23658] = 32'b11111111111111110111011110100100;
assign LUT_2[23659] = 32'b11111111111111110100010110111101;
assign LUT_2[23660] = 32'b11111111111111101101000011010000;
assign LUT_2[23661] = 32'b11111111111111101001111011101001;
assign LUT_2[23662] = 32'b11111111111111110011111100001100;
assign LUT_2[23663] = 32'b11111111111111110000110100100101;
assign LUT_2[23664] = 32'b11111111111111110000011000010101;
assign LUT_2[23665] = 32'b11111111111111101101010000101110;
assign LUT_2[23666] = 32'b11111111111111110111010001010001;
assign LUT_2[23667] = 32'b11111111111111110100001001101010;
assign LUT_2[23668] = 32'b11111111111111101100110101111101;
assign LUT_2[23669] = 32'b11111111111111101001101110010110;
assign LUT_2[23670] = 32'b11111111111111110011101110111001;
assign LUT_2[23671] = 32'b11111111111111110000100111010010;
assign LUT_2[23672] = 32'b11111111111111101011001001110010;
assign LUT_2[23673] = 32'b11111111111111101000000010001011;
assign LUT_2[23674] = 32'b11111111111111110010000010101110;
assign LUT_2[23675] = 32'b11111111111111101110111011000111;
assign LUT_2[23676] = 32'b11111111111111100111100111011010;
assign LUT_2[23677] = 32'b11111111111111100100011111110011;
assign LUT_2[23678] = 32'b11111111111111101110100000010110;
assign LUT_2[23679] = 32'b11111111111111101011011000101111;
assign LUT_2[23680] = 32'b00000000000000000001100100001110;
assign LUT_2[23681] = 32'b11111111111111111110011100100111;
assign LUT_2[23682] = 32'b00000000000000001000011101001010;
assign LUT_2[23683] = 32'b00000000000000000101010101100011;
assign LUT_2[23684] = 32'b11111111111111111110000001110110;
assign LUT_2[23685] = 32'b11111111111111111010111010001111;
assign LUT_2[23686] = 32'b00000000000000000100111010110010;
assign LUT_2[23687] = 32'b00000000000000000001110011001011;
assign LUT_2[23688] = 32'b11111111111111111100010101101011;
assign LUT_2[23689] = 32'b11111111111111111001001110000100;
assign LUT_2[23690] = 32'b00000000000000000011001110100111;
assign LUT_2[23691] = 32'b00000000000000000000000111000000;
assign LUT_2[23692] = 32'b11111111111111111000110011010011;
assign LUT_2[23693] = 32'b11111111111111110101101011101100;
assign LUT_2[23694] = 32'b11111111111111111111101100001111;
assign LUT_2[23695] = 32'b11111111111111111100100100101000;
assign LUT_2[23696] = 32'b11111111111111111100001000011000;
assign LUT_2[23697] = 32'b11111111111111111001000000110001;
assign LUT_2[23698] = 32'b00000000000000000011000001010100;
assign LUT_2[23699] = 32'b11111111111111111111111001101101;
assign LUT_2[23700] = 32'b11111111111111111000100110000000;
assign LUT_2[23701] = 32'b11111111111111110101011110011001;
assign LUT_2[23702] = 32'b11111111111111111111011110111100;
assign LUT_2[23703] = 32'b11111111111111111100010111010101;
assign LUT_2[23704] = 32'b11111111111111110110111001110101;
assign LUT_2[23705] = 32'b11111111111111110011110010001110;
assign LUT_2[23706] = 32'b11111111111111111101110010110001;
assign LUT_2[23707] = 32'b11111111111111111010101011001010;
assign LUT_2[23708] = 32'b11111111111111110011010111011101;
assign LUT_2[23709] = 32'b11111111111111110000001111110110;
assign LUT_2[23710] = 32'b11111111111111111010010000011001;
assign LUT_2[23711] = 32'b11111111111111110111001000110010;
assign LUT_2[23712] = 32'b00000000000000000001111111110111;
assign LUT_2[23713] = 32'b11111111111111111110111000010000;
assign LUT_2[23714] = 32'b00000000000000001000111000110011;
assign LUT_2[23715] = 32'b00000000000000000101110001001100;
assign LUT_2[23716] = 32'b11111111111111111110011101011111;
assign LUT_2[23717] = 32'b11111111111111111011010101111000;
assign LUT_2[23718] = 32'b00000000000000000101010110011011;
assign LUT_2[23719] = 32'b00000000000000000010001110110100;
assign LUT_2[23720] = 32'b11111111111111111100110001010100;
assign LUT_2[23721] = 32'b11111111111111111001101001101101;
assign LUT_2[23722] = 32'b00000000000000000011101010010000;
assign LUT_2[23723] = 32'b00000000000000000000100010101001;
assign LUT_2[23724] = 32'b11111111111111111001001110111100;
assign LUT_2[23725] = 32'b11111111111111110110000111010101;
assign LUT_2[23726] = 32'b00000000000000000000000111111000;
assign LUT_2[23727] = 32'b11111111111111111101000000010001;
assign LUT_2[23728] = 32'b11111111111111111100100100000001;
assign LUT_2[23729] = 32'b11111111111111111001011100011010;
assign LUT_2[23730] = 32'b00000000000000000011011100111101;
assign LUT_2[23731] = 32'b00000000000000000000010101010110;
assign LUT_2[23732] = 32'b11111111111111111001000001101001;
assign LUT_2[23733] = 32'b11111111111111110101111010000010;
assign LUT_2[23734] = 32'b11111111111111111111111010100101;
assign LUT_2[23735] = 32'b11111111111111111100110010111110;
assign LUT_2[23736] = 32'b11111111111111110111010101011110;
assign LUT_2[23737] = 32'b11111111111111110100001101110111;
assign LUT_2[23738] = 32'b11111111111111111110001110011010;
assign LUT_2[23739] = 32'b11111111111111111011000110110011;
assign LUT_2[23740] = 32'b11111111111111110011110011000110;
assign LUT_2[23741] = 32'b11111111111111110000101011011111;
assign LUT_2[23742] = 32'b11111111111111111010101100000010;
assign LUT_2[23743] = 32'b11111111111111110111100100011011;
assign LUT_2[23744] = 32'b11111111111111111001101100110001;
assign LUT_2[23745] = 32'b11111111111111110110100101001010;
assign LUT_2[23746] = 32'b00000000000000000000100101101101;
assign LUT_2[23747] = 32'b11111111111111111101011110000110;
assign LUT_2[23748] = 32'b11111111111111110110001010011001;
assign LUT_2[23749] = 32'b11111111111111110011000010110010;
assign LUT_2[23750] = 32'b11111111111111111101000011010101;
assign LUT_2[23751] = 32'b11111111111111111001111011101110;
assign LUT_2[23752] = 32'b11111111111111110100011110001110;
assign LUT_2[23753] = 32'b11111111111111110001010110100111;
assign LUT_2[23754] = 32'b11111111111111111011010111001010;
assign LUT_2[23755] = 32'b11111111111111111000001111100011;
assign LUT_2[23756] = 32'b11111111111111110000111011110110;
assign LUT_2[23757] = 32'b11111111111111101101110100001111;
assign LUT_2[23758] = 32'b11111111111111110111110100110010;
assign LUT_2[23759] = 32'b11111111111111110100101101001011;
assign LUT_2[23760] = 32'b11111111111111110100010000111011;
assign LUT_2[23761] = 32'b11111111111111110001001001010100;
assign LUT_2[23762] = 32'b11111111111111111011001001110111;
assign LUT_2[23763] = 32'b11111111111111111000000010010000;
assign LUT_2[23764] = 32'b11111111111111110000101110100011;
assign LUT_2[23765] = 32'b11111111111111101101100110111100;
assign LUT_2[23766] = 32'b11111111111111110111100111011111;
assign LUT_2[23767] = 32'b11111111111111110100011111111000;
assign LUT_2[23768] = 32'b11111111111111101111000010011000;
assign LUT_2[23769] = 32'b11111111111111101011111010110001;
assign LUT_2[23770] = 32'b11111111111111110101111011010100;
assign LUT_2[23771] = 32'b11111111111111110010110011101101;
assign LUT_2[23772] = 32'b11111111111111101011100000000000;
assign LUT_2[23773] = 32'b11111111111111101000011000011001;
assign LUT_2[23774] = 32'b11111111111111110010011000111100;
assign LUT_2[23775] = 32'b11111111111111101111010001010101;
assign LUT_2[23776] = 32'b11111111111111111010001000011010;
assign LUT_2[23777] = 32'b11111111111111110111000000110011;
assign LUT_2[23778] = 32'b00000000000000000001000001010110;
assign LUT_2[23779] = 32'b11111111111111111101111001101111;
assign LUT_2[23780] = 32'b11111111111111110110100110000010;
assign LUT_2[23781] = 32'b11111111111111110011011110011011;
assign LUT_2[23782] = 32'b11111111111111111101011110111110;
assign LUT_2[23783] = 32'b11111111111111111010010111010111;
assign LUT_2[23784] = 32'b11111111111111110100111001110111;
assign LUT_2[23785] = 32'b11111111111111110001110010010000;
assign LUT_2[23786] = 32'b11111111111111111011110010110011;
assign LUT_2[23787] = 32'b11111111111111111000101011001100;
assign LUT_2[23788] = 32'b11111111111111110001010111011111;
assign LUT_2[23789] = 32'b11111111111111101110001111111000;
assign LUT_2[23790] = 32'b11111111111111111000010000011011;
assign LUT_2[23791] = 32'b11111111111111110101001000110100;
assign LUT_2[23792] = 32'b11111111111111110100101100100100;
assign LUT_2[23793] = 32'b11111111111111110001100100111101;
assign LUT_2[23794] = 32'b11111111111111111011100101100000;
assign LUT_2[23795] = 32'b11111111111111111000011101111001;
assign LUT_2[23796] = 32'b11111111111111110001001010001100;
assign LUT_2[23797] = 32'b11111111111111101110000010100101;
assign LUT_2[23798] = 32'b11111111111111111000000011001000;
assign LUT_2[23799] = 32'b11111111111111110100111011100001;
assign LUT_2[23800] = 32'b11111111111111101111011110000001;
assign LUT_2[23801] = 32'b11111111111111101100010110011010;
assign LUT_2[23802] = 32'b11111111111111110110010110111101;
assign LUT_2[23803] = 32'b11111111111111110011001111010110;
assign LUT_2[23804] = 32'b11111111111111101011111011101001;
assign LUT_2[23805] = 32'b11111111111111101000110100000010;
assign LUT_2[23806] = 32'b11111111111111110010110100100101;
assign LUT_2[23807] = 32'b11111111111111101111101100111110;
assign LUT_2[23808] = 32'b00000000000000000001001110100101;
assign LUT_2[23809] = 32'b11111111111111111110000110111110;
assign LUT_2[23810] = 32'b00000000000000001000000111100001;
assign LUT_2[23811] = 32'b00000000000000000100111111111010;
assign LUT_2[23812] = 32'b11111111111111111101101100001101;
assign LUT_2[23813] = 32'b11111111111111111010100100100110;
assign LUT_2[23814] = 32'b00000000000000000100100101001001;
assign LUT_2[23815] = 32'b00000000000000000001011101100010;
assign LUT_2[23816] = 32'b11111111111111111100000000000010;
assign LUT_2[23817] = 32'b11111111111111111000111000011011;
assign LUT_2[23818] = 32'b00000000000000000010111000111110;
assign LUT_2[23819] = 32'b11111111111111111111110001010111;
assign LUT_2[23820] = 32'b11111111111111111000011101101010;
assign LUT_2[23821] = 32'b11111111111111110101010110000011;
assign LUT_2[23822] = 32'b11111111111111111111010110100110;
assign LUT_2[23823] = 32'b11111111111111111100001110111111;
assign LUT_2[23824] = 32'b11111111111111111011110010101111;
assign LUT_2[23825] = 32'b11111111111111111000101011001000;
assign LUT_2[23826] = 32'b00000000000000000010101011101011;
assign LUT_2[23827] = 32'b11111111111111111111100100000100;
assign LUT_2[23828] = 32'b11111111111111111000010000010111;
assign LUT_2[23829] = 32'b11111111111111110101001000110000;
assign LUT_2[23830] = 32'b11111111111111111111001001010011;
assign LUT_2[23831] = 32'b11111111111111111100000001101100;
assign LUT_2[23832] = 32'b11111111111111110110100100001100;
assign LUT_2[23833] = 32'b11111111111111110011011100100101;
assign LUT_2[23834] = 32'b11111111111111111101011101001000;
assign LUT_2[23835] = 32'b11111111111111111010010101100001;
assign LUT_2[23836] = 32'b11111111111111110011000001110100;
assign LUT_2[23837] = 32'b11111111111111101111111010001101;
assign LUT_2[23838] = 32'b11111111111111111001111010110000;
assign LUT_2[23839] = 32'b11111111111111110110110011001001;
assign LUT_2[23840] = 32'b00000000000000000001101010001110;
assign LUT_2[23841] = 32'b11111111111111111110100010100111;
assign LUT_2[23842] = 32'b00000000000000001000100011001010;
assign LUT_2[23843] = 32'b00000000000000000101011011100011;
assign LUT_2[23844] = 32'b11111111111111111110000111110110;
assign LUT_2[23845] = 32'b11111111111111111011000000001111;
assign LUT_2[23846] = 32'b00000000000000000101000000110010;
assign LUT_2[23847] = 32'b00000000000000000001111001001011;
assign LUT_2[23848] = 32'b11111111111111111100011011101011;
assign LUT_2[23849] = 32'b11111111111111111001010100000100;
assign LUT_2[23850] = 32'b00000000000000000011010100100111;
assign LUT_2[23851] = 32'b00000000000000000000001101000000;
assign LUT_2[23852] = 32'b11111111111111111000111001010011;
assign LUT_2[23853] = 32'b11111111111111110101110001101100;
assign LUT_2[23854] = 32'b11111111111111111111110010001111;
assign LUT_2[23855] = 32'b11111111111111111100101010101000;
assign LUT_2[23856] = 32'b11111111111111111100001110011000;
assign LUT_2[23857] = 32'b11111111111111111001000110110001;
assign LUT_2[23858] = 32'b00000000000000000011000111010100;
assign LUT_2[23859] = 32'b11111111111111111111111111101101;
assign LUT_2[23860] = 32'b11111111111111111000101100000000;
assign LUT_2[23861] = 32'b11111111111111110101100100011001;
assign LUT_2[23862] = 32'b11111111111111111111100100111100;
assign LUT_2[23863] = 32'b11111111111111111100011101010101;
assign LUT_2[23864] = 32'b11111111111111110110111111110101;
assign LUT_2[23865] = 32'b11111111111111110011111000001110;
assign LUT_2[23866] = 32'b11111111111111111101111000110001;
assign LUT_2[23867] = 32'b11111111111111111010110001001010;
assign LUT_2[23868] = 32'b11111111111111110011011101011101;
assign LUT_2[23869] = 32'b11111111111111110000010101110110;
assign LUT_2[23870] = 32'b11111111111111111010010110011001;
assign LUT_2[23871] = 32'b11111111111111110111001110110010;
assign LUT_2[23872] = 32'b11111111111111111001010111001000;
assign LUT_2[23873] = 32'b11111111111111110110001111100001;
assign LUT_2[23874] = 32'b00000000000000000000010000000100;
assign LUT_2[23875] = 32'b11111111111111111101001000011101;
assign LUT_2[23876] = 32'b11111111111111110101110100110000;
assign LUT_2[23877] = 32'b11111111111111110010101101001001;
assign LUT_2[23878] = 32'b11111111111111111100101101101100;
assign LUT_2[23879] = 32'b11111111111111111001100110000101;
assign LUT_2[23880] = 32'b11111111111111110100001000100101;
assign LUT_2[23881] = 32'b11111111111111110001000000111110;
assign LUT_2[23882] = 32'b11111111111111111011000001100001;
assign LUT_2[23883] = 32'b11111111111111110111111001111010;
assign LUT_2[23884] = 32'b11111111111111110000100110001101;
assign LUT_2[23885] = 32'b11111111111111101101011110100110;
assign LUT_2[23886] = 32'b11111111111111110111011111001001;
assign LUT_2[23887] = 32'b11111111111111110100010111100010;
assign LUT_2[23888] = 32'b11111111111111110011111011010010;
assign LUT_2[23889] = 32'b11111111111111110000110011101011;
assign LUT_2[23890] = 32'b11111111111111111010110100001110;
assign LUT_2[23891] = 32'b11111111111111110111101100100111;
assign LUT_2[23892] = 32'b11111111111111110000011000111010;
assign LUT_2[23893] = 32'b11111111111111101101010001010011;
assign LUT_2[23894] = 32'b11111111111111110111010001110110;
assign LUT_2[23895] = 32'b11111111111111110100001010001111;
assign LUT_2[23896] = 32'b11111111111111101110101100101111;
assign LUT_2[23897] = 32'b11111111111111101011100101001000;
assign LUT_2[23898] = 32'b11111111111111110101100101101011;
assign LUT_2[23899] = 32'b11111111111111110010011110000100;
assign LUT_2[23900] = 32'b11111111111111101011001010010111;
assign LUT_2[23901] = 32'b11111111111111101000000010110000;
assign LUT_2[23902] = 32'b11111111111111110010000011010011;
assign LUT_2[23903] = 32'b11111111111111101110111011101100;
assign LUT_2[23904] = 32'b11111111111111111001110010110001;
assign LUT_2[23905] = 32'b11111111111111110110101011001010;
assign LUT_2[23906] = 32'b00000000000000000000101011101101;
assign LUT_2[23907] = 32'b11111111111111111101100100000110;
assign LUT_2[23908] = 32'b11111111111111110110010000011001;
assign LUT_2[23909] = 32'b11111111111111110011001000110010;
assign LUT_2[23910] = 32'b11111111111111111101001001010101;
assign LUT_2[23911] = 32'b11111111111111111010000001101110;
assign LUT_2[23912] = 32'b11111111111111110100100100001110;
assign LUT_2[23913] = 32'b11111111111111110001011100100111;
assign LUT_2[23914] = 32'b11111111111111111011011101001010;
assign LUT_2[23915] = 32'b11111111111111111000010101100011;
assign LUT_2[23916] = 32'b11111111111111110001000001110110;
assign LUT_2[23917] = 32'b11111111111111101101111010001111;
assign LUT_2[23918] = 32'b11111111111111110111111010110010;
assign LUT_2[23919] = 32'b11111111111111110100110011001011;
assign LUT_2[23920] = 32'b11111111111111110100010110111011;
assign LUT_2[23921] = 32'b11111111111111110001001111010100;
assign LUT_2[23922] = 32'b11111111111111111011001111110111;
assign LUT_2[23923] = 32'b11111111111111111000001000010000;
assign LUT_2[23924] = 32'b11111111111111110000110100100011;
assign LUT_2[23925] = 32'b11111111111111101101101100111100;
assign LUT_2[23926] = 32'b11111111111111110111101101011111;
assign LUT_2[23927] = 32'b11111111111111110100100101111000;
assign LUT_2[23928] = 32'b11111111111111101111001000011000;
assign LUT_2[23929] = 32'b11111111111111101100000000110001;
assign LUT_2[23930] = 32'b11111111111111110110000001010100;
assign LUT_2[23931] = 32'b11111111111111110010111001101101;
assign LUT_2[23932] = 32'b11111111111111101011100110000000;
assign LUT_2[23933] = 32'b11111111111111101000011110011001;
assign LUT_2[23934] = 32'b11111111111111110010011110111100;
assign LUT_2[23935] = 32'b11111111111111101111010111010101;
assign LUT_2[23936] = 32'b00000000000000000101100010110100;
assign LUT_2[23937] = 32'b00000000000000000010011011001101;
assign LUT_2[23938] = 32'b00000000000000001100011011110000;
assign LUT_2[23939] = 32'b00000000000000001001010100001001;
assign LUT_2[23940] = 32'b00000000000000000010000000011100;
assign LUT_2[23941] = 32'b11111111111111111110111000110101;
assign LUT_2[23942] = 32'b00000000000000001000111001011000;
assign LUT_2[23943] = 32'b00000000000000000101110001110001;
assign LUT_2[23944] = 32'b00000000000000000000010100010001;
assign LUT_2[23945] = 32'b11111111111111111101001100101010;
assign LUT_2[23946] = 32'b00000000000000000111001101001101;
assign LUT_2[23947] = 32'b00000000000000000100000101100110;
assign LUT_2[23948] = 32'b11111111111111111100110001111001;
assign LUT_2[23949] = 32'b11111111111111111001101010010010;
assign LUT_2[23950] = 32'b00000000000000000011101010110101;
assign LUT_2[23951] = 32'b00000000000000000000100011001110;
assign LUT_2[23952] = 32'b00000000000000000000000110111110;
assign LUT_2[23953] = 32'b11111111111111111100111111010111;
assign LUT_2[23954] = 32'b00000000000000000110111111111010;
assign LUT_2[23955] = 32'b00000000000000000011111000010011;
assign LUT_2[23956] = 32'b11111111111111111100100100100110;
assign LUT_2[23957] = 32'b11111111111111111001011100111111;
assign LUT_2[23958] = 32'b00000000000000000011011101100010;
assign LUT_2[23959] = 32'b00000000000000000000010101111011;
assign LUT_2[23960] = 32'b11111111111111111010111000011011;
assign LUT_2[23961] = 32'b11111111111111110111110000110100;
assign LUT_2[23962] = 32'b00000000000000000001110001010111;
assign LUT_2[23963] = 32'b11111111111111111110101001110000;
assign LUT_2[23964] = 32'b11111111111111110111010110000011;
assign LUT_2[23965] = 32'b11111111111111110100001110011100;
assign LUT_2[23966] = 32'b11111111111111111110001110111111;
assign LUT_2[23967] = 32'b11111111111111111011000111011000;
assign LUT_2[23968] = 32'b00000000000000000101111110011101;
assign LUT_2[23969] = 32'b00000000000000000010110110110110;
assign LUT_2[23970] = 32'b00000000000000001100110111011001;
assign LUT_2[23971] = 32'b00000000000000001001101111110010;
assign LUT_2[23972] = 32'b00000000000000000010011100000101;
assign LUT_2[23973] = 32'b11111111111111111111010100011110;
assign LUT_2[23974] = 32'b00000000000000001001010101000001;
assign LUT_2[23975] = 32'b00000000000000000110001101011010;
assign LUT_2[23976] = 32'b00000000000000000000101111111010;
assign LUT_2[23977] = 32'b11111111111111111101101000010011;
assign LUT_2[23978] = 32'b00000000000000000111101000110110;
assign LUT_2[23979] = 32'b00000000000000000100100001001111;
assign LUT_2[23980] = 32'b11111111111111111101001101100010;
assign LUT_2[23981] = 32'b11111111111111111010000101111011;
assign LUT_2[23982] = 32'b00000000000000000100000110011110;
assign LUT_2[23983] = 32'b00000000000000000000111110110111;
assign LUT_2[23984] = 32'b00000000000000000000100010100111;
assign LUT_2[23985] = 32'b11111111111111111101011011000000;
assign LUT_2[23986] = 32'b00000000000000000111011011100011;
assign LUT_2[23987] = 32'b00000000000000000100010011111100;
assign LUT_2[23988] = 32'b11111111111111111101000000001111;
assign LUT_2[23989] = 32'b11111111111111111001111000101000;
assign LUT_2[23990] = 32'b00000000000000000011111001001011;
assign LUT_2[23991] = 32'b00000000000000000000110001100100;
assign LUT_2[23992] = 32'b11111111111111111011010100000100;
assign LUT_2[23993] = 32'b11111111111111111000001100011101;
assign LUT_2[23994] = 32'b00000000000000000010001101000000;
assign LUT_2[23995] = 32'b11111111111111111111000101011001;
assign LUT_2[23996] = 32'b11111111111111110111110001101100;
assign LUT_2[23997] = 32'b11111111111111110100101010000101;
assign LUT_2[23998] = 32'b11111111111111111110101010101000;
assign LUT_2[23999] = 32'b11111111111111111011100011000001;
assign LUT_2[24000] = 32'b11111111111111111101101011010111;
assign LUT_2[24001] = 32'b11111111111111111010100011110000;
assign LUT_2[24002] = 32'b00000000000000000100100100010011;
assign LUT_2[24003] = 32'b00000000000000000001011100101100;
assign LUT_2[24004] = 32'b11111111111111111010001000111111;
assign LUT_2[24005] = 32'b11111111111111110111000001011000;
assign LUT_2[24006] = 32'b00000000000000000001000001111011;
assign LUT_2[24007] = 32'b11111111111111111101111010010100;
assign LUT_2[24008] = 32'b11111111111111111000011100110100;
assign LUT_2[24009] = 32'b11111111111111110101010101001101;
assign LUT_2[24010] = 32'b11111111111111111111010101110000;
assign LUT_2[24011] = 32'b11111111111111111100001110001001;
assign LUT_2[24012] = 32'b11111111111111110100111010011100;
assign LUT_2[24013] = 32'b11111111111111110001110010110101;
assign LUT_2[24014] = 32'b11111111111111111011110011011000;
assign LUT_2[24015] = 32'b11111111111111111000101011110001;
assign LUT_2[24016] = 32'b11111111111111111000001111100001;
assign LUT_2[24017] = 32'b11111111111111110101000111111010;
assign LUT_2[24018] = 32'b11111111111111111111001000011101;
assign LUT_2[24019] = 32'b11111111111111111100000000110110;
assign LUT_2[24020] = 32'b11111111111111110100101101001001;
assign LUT_2[24021] = 32'b11111111111111110001100101100010;
assign LUT_2[24022] = 32'b11111111111111111011100110000101;
assign LUT_2[24023] = 32'b11111111111111111000011110011110;
assign LUT_2[24024] = 32'b11111111111111110011000000111110;
assign LUT_2[24025] = 32'b11111111111111101111111001010111;
assign LUT_2[24026] = 32'b11111111111111111001111001111010;
assign LUT_2[24027] = 32'b11111111111111110110110010010011;
assign LUT_2[24028] = 32'b11111111111111101111011110100110;
assign LUT_2[24029] = 32'b11111111111111101100010110111111;
assign LUT_2[24030] = 32'b11111111111111110110010111100010;
assign LUT_2[24031] = 32'b11111111111111110011001111111011;
assign LUT_2[24032] = 32'b11111111111111111110000111000000;
assign LUT_2[24033] = 32'b11111111111111111010111111011001;
assign LUT_2[24034] = 32'b00000000000000000100111111111100;
assign LUT_2[24035] = 32'b00000000000000000001111000010101;
assign LUT_2[24036] = 32'b11111111111111111010100100101000;
assign LUT_2[24037] = 32'b11111111111111110111011101000001;
assign LUT_2[24038] = 32'b00000000000000000001011101100100;
assign LUT_2[24039] = 32'b11111111111111111110010101111101;
assign LUT_2[24040] = 32'b11111111111111111000111000011101;
assign LUT_2[24041] = 32'b11111111111111110101110000110110;
assign LUT_2[24042] = 32'b11111111111111111111110001011001;
assign LUT_2[24043] = 32'b11111111111111111100101001110010;
assign LUT_2[24044] = 32'b11111111111111110101010110000101;
assign LUT_2[24045] = 32'b11111111111111110010001110011110;
assign LUT_2[24046] = 32'b11111111111111111100001111000001;
assign LUT_2[24047] = 32'b11111111111111111001000111011010;
assign LUT_2[24048] = 32'b11111111111111111000101011001010;
assign LUT_2[24049] = 32'b11111111111111110101100011100011;
assign LUT_2[24050] = 32'b11111111111111111111100100000110;
assign LUT_2[24051] = 32'b11111111111111111100011100011111;
assign LUT_2[24052] = 32'b11111111111111110101001000110010;
assign LUT_2[24053] = 32'b11111111111111110010000001001011;
assign LUT_2[24054] = 32'b11111111111111111100000001101110;
assign LUT_2[24055] = 32'b11111111111111111000111010000111;
assign LUT_2[24056] = 32'b11111111111111110011011100100111;
assign LUT_2[24057] = 32'b11111111111111110000010101000000;
assign LUT_2[24058] = 32'b11111111111111111010010101100011;
assign LUT_2[24059] = 32'b11111111111111110111001101111100;
assign LUT_2[24060] = 32'b11111111111111101111111010001111;
assign LUT_2[24061] = 32'b11111111111111101100110010101000;
assign LUT_2[24062] = 32'b11111111111111110110110011001011;
assign LUT_2[24063] = 32'b11111111111111110011101011100100;
assign LUT_2[24064] = 32'b00000000000000000010000001110001;
assign LUT_2[24065] = 32'b11111111111111111110111010001010;
assign LUT_2[24066] = 32'b00000000000000001000111010101101;
assign LUT_2[24067] = 32'b00000000000000000101110011000110;
assign LUT_2[24068] = 32'b11111111111111111110011111011001;
assign LUT_2[24069] = 32'b11111111111111111011010111110010;
assign LUT_2[24070] = 32'b00000000000000000101011000010101;
assign LUT_2[24071] = 32'b00000000000000000010010000101110;
assign LUT_2[24072] = 32'b11111111111111111100110011001110;
assign LUT_2[24073] = 32'b11111111111111111001101011100111;
assign LUT_2[24074] = 32'b00000000000000000011101100001010;
assign LUT_2[24075] = 32'b00000000000000000000100100100011;
assign LUT_2[24076] = 32'b11111111111111111001010000110110;
assign LUT_2[24077] = 32'b11111111111111110110001001001111;
assign LUT_2[24078] = 32'b00000000000000000000001001110010;
assign LUT_2[24079] = 32'b11111111111111111101000010001011;
assign LUT_2[24080] = 32'b11111111111111111100100101111011;
assign LUT_2[24081] = 32'b11111111111111111001011110010100;
assign LUT_2[24082] = 32'b00000000000000000011011110110111;
assign LUT_2[24083] = 32'b00000000000000000000010111010000;
assign LUT_2[24084] = 32'b11111111111111111001000011100011;
assign LUT_2[24085] = 32'b11111111111111110101111011111100;
assign LUT_2[24086] = 32'b11111111111111111111111100011111;
assign LUT_2[24087] = 32'b11111111111111111100110100111000;
assign LUT_2[24088] = 32'b11111111111111110111010111011000;
assign LUT_2[24089] = 32'b11111111111111110100001111110001;
assign LUT_2[24090] = 32'b11111111111111111110010000010100;
assign LUT_2[24091] = 32'b11111111111111111011001000101101;
assign LUT_2[24092] = 32'b11111111111111110011110101000000;
assign LUT_2[24093] = 32'b11111111111111110000101101011001;
assign LUT_2[24094] = 32'b11111111111111111010101101111100;
assign LUT_2[24095] = 32'b11111111111111110111100110010101;
assign LUT_2[24096] = 32'b00000000000000000010011101011010;
assign LUT_2[24097] = 32'b11111111111111111111010101110011;
assign LUT_2[24098] = 32'b00000000000000001001010110010110;
assign LUT_2[24099] = 32'b00000000000000000110001110101111;
assign LUT_2[24100] = 32'b11111111111111111110111011000010;
assign LUT_2[24101] = 32'b11111111111111111011110011011011;
assign LUT_2[24102] = 32'b00000000000000000101110011111110;
assign LUT_2[24103] = 32'b00000000000000000010101100010111;
assign LUT_2[24104] = 32'b11111111111111111101001110110111;
assign LUT_2[24105] = 32'b11111111111111111010000111010000;
assign LUT_2[24106] = 32'b00000000000000000100000111110011;
assign LUT_2[24107] = 32'b00000000000000000001000000001100;
assign LUT_2[24108] = 32'b11111111111111111001101100011111;
assign LUT_2[24109] = 32'b11111111111111110110100100111000;
assign LUT_2[24110] = 32'b00000000000000000000100101011011;
assign LUT_2[24111] = 32'b11111111111111111101011101110100;
assign LUT_2[24112] = 32'b11111111111111111101000001100100;
assign LUT_2[24113] = 32'b11111111111111111001111001111101;
assign LUT_2[24114] = 32'b00000000000000000011111010100000;
assign LUT_2[24115] = 32'b00000000000000000000110010111001;
assign LUT_2[24116] = 32'b11111111111111111001011111001100;
assign LUT_2[24117] = 32'b11111111111111110110010111100101;
assign LUT_2[24118] = 32'b00000000000000000000011000001000;
assign LUT_2[24119] = 32'b11111111111111111101010000100001;
assign LUT_2[24120] = 32'b11111111111111110111110011000001;
assign LUT_2[24121] = 32'b11111111111111110100101011011010;
assign LUT_2[24122] = 32'b11111111111111111110101011111101;
assign LUT_2[24123] = 32'b11111111111111111011100100010110;
assign LUT_2[24124] = 32'b11111111111111110100010000101001;
assign LUT_2[24125] = 32'b11111111111111110001001001000010;
assign LUT_2[24126] = 32'b11111111111111111011001001100101;
assign LUT_2[24127] = 32'b11111111111111111000000001111110;
assign LUT_2[24128] = 32'b11111111111111111010001010010100;
assign LUT_2[24129] = 32'b11111111111111110111000010101101;
assign LUT_2[24130] = 32'b00000000000000000001000011010000;
assign LUT_2[24131] = 32'b11111111111111111101111011101001;
assign LUT_2[24132] = 32'b11111111111111110110100111111100;
assign LUT_2[24133] = 32'b11111111111111110011100000010101;
assign LUT_2[24134] = 32'b11111111111111111101100000111000;
assign LUT_2[24135] = 32'b11111111111111111010011001010001;
assign LUT_2[24136] = 32'b11111111111111110100111011110001;
assign LUT_2[24137] = 32'b11111111111111110001110100001010;
assign LUT_2[24138] = 32'b11111111111111111011110100101101;
assign LUT_2[24139] = 32'b11111111111111111000101101000110;
assign LUT_2[24140] = 32'b11111111111111110001011001011001;
assign LUT_2[24141] = 32'b11111111111111101110010001110010;
assign LUT_2[24142] = 32'b11111111111111111000010010010101;
assign LUT_2[24143] = 32'b11111111111111110101001010101110;
assign LUT_2[24144] = 32'b11111111111111110100101110011110;
assign LUT_2[24145] = 32'b11111111111111110001100110110111;
assign LUT_2[24146] = 32'b11111111111111111011100111011010;
assign LUT_2[24147] = 32'b11111111111111111000011111110011;
assign LUT_2[24148] = 32'b11111111111111110001001100000110;
assign LUT_2[24149] = 32'b11111111111111101110000100011111;
assign LUT_2[24150] = 32'b11111111111111111000000101000010;
assign LUT_2[24151] = 32'b11111111111111110100111101011011;
assign LUT_2[24152] = 32'b11111111111111101111011111111011;
assign LUT_2[24153] = 32'b11111111111111101100011000010100;
assign LUT_2[24154] = 32'b11111111111111110110011000110111;
assign LUT_2[24155] = 32'b11111111111111110011010001010000;
assign LUT_2[24156] = 32'b11111111111111101011111101100011;
assign LUT_2[24157] = 32'b11111111111111101000110101111100;
assign LUT_2[24158] = 32'b11111111111111110010110110011111;
assign LUT_2[24159] = 32'b11111111111111101111101110111000;
assign LUT_2[24160] = 32'b11111111111111111010100101111101;
assign LUT_2[24161] = 32'b11111111111111110111011110010110;
assign LUT_2[24162] = 32'b00000000000000000001011110111001;
assign LUT_2[24163] = 32'b11111111111111111110010111010010;
assign LUT_2[24164] = 32'b11111111111111110111000011100101;
assign LUT_2[24165] = 32'b11111111111111110011111011111110;
assign LUT_2[24166] = 32'b11111111111111111101111100100001;
assign LUT_2[24167] = 32'b11111111111111111010110100111010;
assign LUT_2[24168] = 32'b11111111111111110101010111011010;
assign LUT_2[24169] = 32'b11111111111111110010001111110011;
assign LUT_2[24170] = 32'b11111111111111111100010000010110;
assign LUT_2[24171] = 32'b11111111111111111001001000101111;
assign LUT_2[24172] = 32'b11111111111111110001110101000010;
assign LUT_2[24173] = 32'b11111111111111101110101101011011;
assign LUT_2[24174] = 32'b11111111111111111000101101111110;
assign LUT_2[24175] = 32'b11111111111111110101100110010111;
assign LUT_2[24176] = 32'b11111111111111110101001010000111;
assign LUT_2[24177] = 32'b11111111111111110010000010100000;
assign LUT_2[24178] = 32'b11111111111111111100000011000011;
assign LUT_2[24179] = 32'b11111111111111111000111011011100;
assign LUT_2[24180] = 32'b11111111111111110001100111101111;
assign LUT_2[24181] = 32'b11111111111111101110100000001000;
assign LUT_2[24182] = 32'b11111111111111111000100000101011;
assign LUT_2[24183] = 32'b11111111111111110101011001000100;
assign LUT_2[24184] = 32'b11111111111111101111111011100100;
assign LUT_2[24185] = 32'b11111111111111101100110011111101;
assign LUT_2[24186] = 32'b11111111111111110110110100100000;
assign LUT_2[24187] = 32'b11111111111111110011101100111001;
assign LUT_2[24188] = 32'b11111111111111101100011001001100;
assign LUT_2[24189] = 32'b11111111111111101001010001100101;
assign LUT_2[24190] = 32'b11111111111111110011010010001000;
assign LUT_2[24191] = 32'b11111111111111110000001010100001;
assign LUT_2[24192] = 32'b00000000000000000110010110000000;
assign LUT_2[24193] = 32'b00000000000000000011001110011001;
assign LUT_2[24194] = 32'b00000000000000001101001110111100;
assign LUT_2[24195] = 32'b00000000000000001010000111010101;
assign LUT_2[24196] = 32'b00000000000000000010110011101000;
assign LUT_2[24197] = 32'b11111111111111111111101100000001;
assign LUT_2[24198] = 32'b00000000000000001001101100100100;
assign LUT_2[24199] = 32'b00000000000000000110100100111101;
assign LUT_2[24200] = 32'b00000000000000000001000111011101;
assign LUT_2[24201] = 32'b11111111111111111101111111110110;
assign LUT_2[24202] = 32'b00000000000000001000000000011001;
assign LUT_2[24203] = 32'b00000000000000000100111000110010;
assign LUT_2[24204] = 32'b11111111111111111101100101000101;
assign LUT_2[24205] = 32'b11111111111111111010011101011110;
assign LUT_2[24206] = 32'b00000000000000000100011110000001;
assign LUT_2[24207] = 32'b00000000000000000001010110011010;
assign LUT_2[24208] = 32'b00000000000000000000111010001010;
assign LUT_2[24209] = 32'b11111111111111111101110010100011;
assign LUT_2[24210] = 32'b00000000000000000111110011000110;
assign LUT_2[24211] = 32'b00000000000000000100101011011111;
assign LUT_2[24212] = 32'b11111111111111111101010111110010;
assign LUT_2[24213] = 32'b11111111111111111010010000001011;
assign LUT_2[24214] = 32'b00000000000000000100010000101110;
assign LUT_2[24215] = 32'b00000000000000000001001001000111;
assign LUT_2[24216] = 32'b11111111111111111011101011100111;
assign LUT_2[24217] = 32'b11111111111111111000100100000000;
assign LUT_2[24218] = 32'b00000000000000000010100100100011;
assign LUT_2[24219] = 32'b11111111111111111111011100111100;
assign LUT_2[24220] = 32'b11111111111111111000001001001111;
assign LUT_2[24221] = 32'b11111111111111110101000001101000;
assign LUT_2[24222] = 32'b11111111111111111111000010001011;
assign LUT_2[24223] = 32'b11111111111111111011111010100100;
assign LUT_2[24224] = 32'b00000000000000000110110001101001;
assign LUT_2[24225] = 32'b00000000000000000011101010000010;
assign LUT_2[24226] = 32'b00000000000000001101101010100101;
assign LUT_2[24227] = 32'b00000000000000001010100010111110;
assign LUT_2[24228] = 32'b00000000000000000011001111010001;
assign LUT_2[24229] = 32'b00000000000000000000000111101010;
assign LUT_2[24230] = 32'b00000000000000001010001000001101;
assign LUT_2[24231] = 32'b00000000000000000111000000100110;
assign LUT_2[24232] = 32'b00000000000000000001100011000110;
assign LUT_2[24233] = 32'b11111111111111111110011011011111;
assign LUT_2[24234] = 32'b00000000000000001000011100000010;
assign LUT_2[24235] = 32'b00000000000000000101010100011011;
assign LUT_2[24236] = 32'b11111111111111111110000000101110;
assign LUT_2[24237] = 32'b11111111111111111010111001000111;
assign LUT_2[24238] = 32'b00000000000000000100111001101010;
assign LUT_2[24239] = 32'b00000000000000000001110010000011;
assign LUT_2[24240] = 32'b00000000000000000001010101110011;
assign LUT_2[24241] = 32'b11111111111111111110001110001100;
assign LUT_2[24242] = 32'b00000000000000001000001110101111;
assign LUT_2[24243] = 32'b00000000000000000101000111001000;
assign LUT_2[24244] = 32'b11111111111111111101110011011011;
assign LUT_2[24245] = 32'b11111111111111111010101011110100;
assign LUT_2[24246] = 32'b00000000000000000100101100010111;
assign LUT_2[24247] = 32'b00000000000000000001100100110000;
assign LUT_2[24248] = 32'b11111111111111111100000111010000;
assign LUT_2[24249] = 32'b11111111111111111000111111101001;
assign LUT_2[24250] = 32'b00000000000000000011000000001100;
assign LUT_2[24251] = 32'b11111111111111111111111000100101;
assign LUT_2[24252] = 32'b11111111111111111000100100111000;
assign LUT_2[24253] = 32'b11111111111111110101011101010001;
assign LUT_2[24254] = 32'b11111111111111111111011101110100;
assign LUT_2[24255] = 32'b11111111111111111100010110001101;
assign LUT_2[24256] = 32'b11111111111111111110011110100011;
assign LUT_2[24257] = 32'b11111111111111111011010110111100;
assign LUT_2[24258] = 32'b00000000000000000101010111011111;
assign LUT_2[24259] = 32'b00000000000000000010001111111000;
assign LUT_2[24260] = 32'b11111111111111111010111100001011;
assign LUT_2[24261] = 32'b11111111111111110111110100100100;
assign LUT_2[24262] = 32'b00000000000000000001110101000111;
assign LUT_2[24263] = 32'b11111111111111111110101101100000;
assign LUT_2[24264] = 32'b11111111111111111001010000000000;
assign LUT_2[24265] = 32'b11111111111111110110001000011001;
assign LUT_2[24266] = 32'b00000000000000000000001000111100;
assign LUT_2[24267] = 32'b11111111111111111101000001010101;
assign LUT_2[24268] = 32'b11111111111111110101101101101000;
assign LUT_2[24269] = 32'b11111111111111110010100110000001;
assign LUT_2[24270] = 32'b11111111111111111100100110100100;
assign LUT_2[24271] = 32'b11111111111111111001011110111101;
assign LUT_2[24272] = 32'b11111111111111111001000010101101;
assign LUT_2[24273] = 32'b11111111111111110101111011000110;
assign LUT_2[24274] = 32'b11111111111111111111111011101001;
assign LUT_2[24275] = 32'b11111111111111111100110100000010;
assign LUT_2[24276] = 32'b11111111111111110101100000010101;
assign LUT_2[24277] = 32'b11111111111111110010011000101110;
assign LUT_2[24278] = 32'b11111111111111111100011001010001;
assign LUT_2[24279] = 32'b11111111111111111001010001101010;
assign LUT_2[24280] = 32'b11111111111111110011110100001010;
assign LUT_2[24281] = 32'b11111111111111110000101100100011;
assign LUT_2[24282] = 32'b11111111111111111010101101000110;
assign LUT_2[24283] = 32'b11111111111111110111100101011111;
assign LUT_2[24284] = 32'b11111111111111110000010001110010;
assign LUT_2[24285] = 32'b11111111111111101101001010001011;
assign LUT_2[24286] = 32'b11111111111111110111001010101110;
assign LUT_2[24287] = 32'b11111111111111110100000011000111;
assign LUT_2[24288] = 32'b11111111111111111110111010001100;
assign LUT_2[24289] = 32'b11111111111111111011110010100101;
assign LUT_2[24290] = 32'b00000000000000000101110011001000;
assign LUT_2[24291] = 32'b00000000000000000010101011100001;
assign LUT_2[24292] = 32'b11111111111111111011010111110100;
assign LUT_2[24293] = 32'b11111111111111111000010000001101;
assign LUT_2[24294] = 32'b00000000000000000010010000110000;
assign LUT_2[24295] = 32'b11111111111111111111001001001001;
assign LUT_2[24296] = 32'b11111111111111111001101011101001;
assign LUT_2[24297] = 32'b11111111111111110110100100000010;
assign LUT_2[24298] = 32'b00000000000000000000100100100101;
assign LUT_2[24299] = 32'b11111111111111111101011100111110;
assign LUT_2[24300] = 32'b11111111111111110110001001010001;
assign LUT_2[24301] = 32'b11111111111111110011000001101010;
assign LUT_2[24302] = 32'b11111111111111111101000010001101;
assign LUT_2[24303] = 32'b11111111111111111001111010100110;
assign LUT_2[24304] = 32'b11111111111111111001011110010110;
assign LUT_2[24305] = 32'b11111111111111110110010110101111;
assign LUT_2[24306] = 32'b00000000000000000000010111010010;
assign LUT_2[24307] = 32'b11111111111111111101001111101011;
assign LUT_2[24308] = 32'b11111111111111110101111011111110;
assign LUT_2[24309] = 32'b11111111111111110010110100010111;
assign LUT_2[24310] = 32'b11111111111111111100110100111010;
assign LUT_2[24311] = 32'b11111111111111111001101101010011;
assign LUT_2[24312] = 32'b11111111111111110100001111110011;
assign LUT_2[24313] = 32'b11111111111111110001001000001100;
assign LUT_2[24314] = 32'b11111111111111111011001000101111;
assign LUT_2[24315] = 32'b11111111111111111000000001001000;
assign LUT_2[24316] = 32'b11111111111111110000101101011011;
assign LUT_2[24317] = 32'b11111111111111101101100101110100;
assign LUT_2[24318] = 32'b11111111111111110111100110010111;
assign LUT_2[24319] = 32'b11111111111111110100011110110000;
assign LUT_2[24320] = 32'b00000000000000000110000000010111;
assign LUT_2[24321] = 32'b00000000000000000010111000110000;
assign LUT_2[24322] = 32'b00000000000000001100111001010011;
assign LUT_2[24323] = 32'b00000000000000001001110001101100;
assign LUT_2[24324] = 32'b00000000000000000010011101111111;
assign LUT_2[24325] = 32'b11111111111111111111010110011000;
assign LUT_2[24326] = 32'b00000000000000001001010110111011;
assign LUT_2[24327] = 32'b00000000000000000110001111010100;
assign LUT_2[24328] = 32'b00000000000000000000110001110100;
assign LUT_2[24329] = 32'b11111111111111111101101010001101;
assign LUT_2[24330] = 32'b00000000000000000111101010110000;
assign LUT_2[24331] = 32'b00000000000000000100100011001001;
assign LUT_2[24332] = 32'b11111111111111111101001111011100;
assign LUT_2[24333] = 32'b11111111111111111010000111110101;
assign LUT_2[24334] = 32'b00000000000000000100001000011000;
assign LUT_2[24335] = 32'b00000000000000000001000000110001;
assign LUT_2[24336] = 32'b00000000000000000000100100100001;
assign LUT_2[24337] = 32'b11111111111111111101011100111010;
assign LUT_2[24338] = 32'b00000000000000000111011101011101;
assign LUT_2[24339] = 32'b00000000000000000100010101110110;
assign LUT_2[24340] = 32'b11111111111111111101000010001001;
assign LUT_2[24341] = 32'b11111111111111111001111010100010;
assign LUT_2[24342] = 32'b00000000000000000011111011000101;
assign LUT_2[24343] = 32'b00000000000000000000110011011110;
assign LUT_2[24344] = 32'b11111111111111111011010101111110;
assign LUT_2[24345] = 32'b11111111111111111000001110010111;
assign LUT_2[24346] = 32'b00000000000000000010001110111010;
assign LUT_2[24347] = 32'b11111111111111111111000111010011;
assign LUT_2[24348] = 32'b11111111111111110111110011100110;
assign LUT_2[24349] = 32'b11111111111111110100101011111111;
assign LUT_2[24350] = 32'b11111111111111111110101100100010;
assign LUT_2[24351] = 32'b11111111111111111011100100111011;
assign LUT_2[24352] = 32'b00000000000000000110011100000000;
assign LUT_2[24353] = 32'b00000000000000000011010100011001;
assign LUT_2[24354] = 32'b00000000000000001101010100111100;
assign LUT_2[24355] = 32'b00000000000000001010001101010101;
assign LUT_2[24356] = 32'b00000000000000000010111001101000;
assign LUT_2[24357] = 32'b11111111111111111111110010000001;
assign LUT_2[24358] = 32'b00000000000000001001110010100100;
assign LUT_2[24359] = 32'b00000000000000000110101010111101;
assign LUT_2[24360] = 32'b00000000000000000001001101011101;
assign LUT_2[24361] = 32'b11111111111111111110000101110110;
assign LUT_2[24362] = 32'b00000000000000001000000110011001;
assign LUT_2[24363] = 32'b00000000000000000100111110110010;
assign LUT_2[24364] = 32'b11111111111111111101101011000101;
assign LUT_2[24365] = 32'b11111111111111111010100011011110;
assign LUT_2[24366] = 32'b00000000000000000100100100000001;
assign LUT_2[24367] = 32'b00000000000000000001011100011010;
assign LUT_2[24368] = 32'b00000000000000000001000000001010;
assign LUT_2[24369] = 32'b11111111111111111101111000100011;
assign LUT_2[24370] = 32'b00000000000000000111111001000110;
assign LUT_2[24371] = 32'b00000000000000000100110001011111;
assign LUT_2[24372] = 32'b11111111111111111101011101110010;
assign LUT_2[24373] = 32'b11111111111111111010010110001011;
assign LUT_2[24374] = 32'b00000000000000000100010110101110;
assign LUT_2[24375] = 32'b00000000000000000001001111000111;
assign LUT_2[24376] = 32'b11111111111111111011110001100111;
assign LUT_2[24377] = 32'b11111111111111111000101010000000;
assign LUT_2[24378] = 32'b00000000000000000010101010100011;
assign LUT_2[24379] = 32'b11111111111111111111100010111100;
assign LUT_2[24380] = 32'b11111111111111111000001111001111;
assign LUT_2[24381] = 32'b11111111111111110101000111101000;
assign LUT_2[24382] = 32'b11111111111111111111001000001011;
assign LUT_2[24383] = 32'b11111111111111111100000000100100;
assign LUT_2[24384] = 32'b11111111111111111110001000111010;
assign LUT_2[24385] = 32'b11111111111111111011000001010011;
assign LUT_2[24386] = 32'b00000000000000000101000001110110;
assign LUT_2[24387] = 32'b00000000000000000001111010001111;
assign LUT_2[24388] = 32'b11111111111111111010100110100010;
assign LUT_2[24389] = 32'b11111111111111110111011110111011;
assign LUT_2[24390] = 32'b00000000000000000001011111011110;
assign LUT_2[24391] = 32'b11111111111111111110010111110111;
assign LUT_2[24392] = 32'b11111111111111111000111010010111;
assign LUT_2[24393] = 32'b11111111111111110101110010110000;
assign LUT_2[24394] = 32'b11111111111111111111110011010011;
assign LUT_2[24395] = 32'b11111111111111111100101011101100;
assign LUT_2[24396] = 32'b11111111111111110101010111111111;
assign LUT_2[24397] = 32'b11111111111111110010010000011000;
assign LUT_2[24398] = 32'b11111111111111111100010000111011;
assign LUT_2[24399] = 32'b11111111111111111001001001010100;
assign LUT_2[24400] = 32'b11111111111111111000101101000100;
assign LUT_2[24401] = 32'b11111111111111110101100101011101;
assign LUT_2[24402] = 32'b11111111111111111111100110000000;
assign LUT_2[24403] = 32'b11111111111111111100011110011001;
assign LUT_2[24404] = 32'b11111111111111110101001010101100;
assign LUT_2[24405] = 32'b11111111111111110010000011000101;
assign LUT_2[24406] = 32'b11111111111111111100000011101000;
assign LUT_2[24407] = 32'b11111111111111111000111100000001;
assign LUT_2[24408] = 32'b11111111111111110011011110100001;
assign LUT_2[24409] = 32'b11111111111111110000010110111010;
assign LUT_2[24410] = 32'b11111111111111111010010111011101;
assign LUT_2[24411] = 32'b11111111111111110111001111110110;
assign LUT_2[24412] = 32'b11111111111111101111111100001001;
assign LUT_2[24413] = 32'b11111111111111101100110100100010;
assign LUT_2[24414] = 32'b11111111111111110110110101000101;
assign LUT_2[24415] = 32'b11111111111111110011101101011110;
assign LUT_2[24416] = 32'b11111111111111111110100100100011;
assign LUT_2[24417] = 32'b11111111111111111011011100111100;
assign LUT_2[24418] = 32'b00000000000000000101011101011111;
assign LUT_2[24419] = 32'b00000000000000000010010101111000;
assign LUT_2[24420] = 32'b11111111111111111011000010001011;
assign LUT_2[24421] = 32'b11111111111111110111111010100100;
assign LUT_2[24422] = 32'b00000000000000000001111011000111;
assign LUT_2[24423] = 32'b11111111111111111110110011100000;
assign LUT_2[24424] = 32'b11111111111111111001010110000000;
assign LUT_2[24425] = 32'b11111111111111110110001110011001;
assign LUT_2[24426] = 32'b00000000000000000000001110111100;
assign LUT_2[24427] = 32'b11111111111111111101000111010101;
assign LUT_2[24428] = 32'b11111111111111110101110011101000;
assign LUT_2[24429] = 32'b11111111111111110010101100000001;
assign LUT_2[24430] = 32'b11111111111111111100101100100100;
assign LUT_2[24431] = 32'b11111111111111111001100100111101;
assign LUT_2[24432] = 32'b11111111111111111001001000101101;
assign LUT_2[24433] = 32'b11111111111111110110000001000110;
assign LUT_2[24434] = 32'b00000000000000000000000001101001;
assign LUT_2[24435] = 32'b11111111111111111100111010000010;
assign LUT_2[24436] = 32'b11111111111111110101100110010101;
assign LUT_2[24437] = 32'b11111111111111110010011110101110;
assign LUT_2[24438] = 32'b11111111111111111100011111010001;
assign LUT_2[24439] = 32'b11111111111111111001010111101010;
assign LUT_2[24440] = 32'b11111111111111110011111010001010;
assign LUT_2[24441] = 32'b11111111111111110000110010100011;
assign LUT_2[24442] = 32'b11111111111111111010110011000110;
assign LUT_2[24443] = 32'b11111111111111110111101011011111;
assign LUT_2[24444] = 32'b11111111111111110000010111110010;
assign LUT_2[24445] = 32'b11111111111111101101010000001011;
assign LUT_2[24446] = 32'b11111111111111110111010000101110;
assign LUT_2[24447] = 32'b11111111111111110100001001000111;
assign LUT_2[24448] = 32'b00000000000000001010010100100110;
assign LUT_2[24449] = 32'b00000000000000000111001100111111;
assign LUT_2[24450] = 32'b00000000000000010001001101100010;
assign LUT_2[24451] = 32'b00000000000000001110000101111011;
assign LUT_2[24452] = 32'b00000000000000000110110010001110;
assign LUT_2[24453] = 32'b00000000000000000011101010100111;
assign LUT_2[24454] = 32'b00000000000000001101101011001010;
assign LUT_2[24455] = 32'b00000000000000001010100011100011;
assign LUT_2[24456] = 32'b00000000000000000101000110000011;
assign LUT_2[24457] = 32'b00000000000000000001111110011100;
assign LUT_2[24458] = 32'b00000000000000001011111110111111;
assign LUT_2[24459] = 32'b00000000000000001000110111011000;
assign LUT_2[24460] = 32'b00000000000000000001100011101011;
assign LUT_2[24461] = 32'b11111111111111111110011100000100;
assign LUT_2[24462] = 32'b00000000000000001000011100100111;
assign LUT_2[24463] = 32'b00000000000000000101010101000000;
assign LUT_2[24464] = 32'b00000000000000000100111000110000;
assign LUT_2[24465] = 32'b00000000000000000001110001001001;
assign LUT_2[24466] = 32'b00000000000000001011110001101100;
assign LUT_2[24467] = 32'b00000000000000001000101010000101;
assign LUT_2[24468] = 32'b00000000000000000001010110011000;
assign LUT_2[24469] = 32'b11111111111111111110001110110001;
assign LUT_2[24470] = 32'b00000000000000001000001111010100;
assign LUT_2[24471] = 32'b00000000000000000101000111101101;
assign LUT_2[24472] = 32'b11111111111111111111101010001101;
assign LUT_2[24473] = 32'b11111111111111111100100010100110;
assign LUT_2[24474] = 32'b00000000000000000110100011001001;
assign LUT_2[24475] = 32'b00000000000000000011011011100010;
assign LUT_2[24476] = 32'b11111111111111111100000111110101;
assign LUT_2[24477] = 32'b11111111111111111001000000001110;
assign LUT_2[24478] = 32'b00000000000000000011000000110001;
assign LUT_2[24479] = 32'b11111111111111111111111001001010;
assign LUT_2[24480] = 32'b00000000000000001010110000001111;
assign LUT_2[24481] = 32'b00000000000000000111101000101000;
assign LUT_2[24482] = 32'b00000000000000010001101001001011;
assign LUT_2[24483] = 32'b00000000000000001110100001100100;
assign LUT_2[24484] = 32'b00000000000000000111001101110111;
assign LUT_2[24485] = 32'b00000000000000000100000110010000;
assign LUT_2[24486] = 32'b00000000000000001110000110110011;
assign LUT_2[24487] = 32'b00000000000000001010111111001100;
assign LUT_2[24488] = 32'b00000000000000000101100001101100;
assign LUT_2[24489] = 32'b00000000000000000010011010000101;
assign LUT_2[24490] = 32'b00000000000000001100011010101000;
assign LUT_2[24491] = 32'b00000000000000001001010011000001;
assign LUT_2[24492] = 32'b00000000000000000001111111010100;
assign LUT_2[24493] = 32'b11111111111111111110110111101101;
assign LUT_2[24494] = 32'b00000000000000001000111000010000;
assign LUT_2[24495] = 32'b00000000000000000101110000101001;
assign LUT_2[24496] = 32'b00000000000000000101010100011001;
assign LUT_2[24497] = 32'b00000000000000000010001100110010;
assign LUT_2[24498] = 32'b00000000000000001100001101010101;
assign LUT_2[24499] = 32'b00000000000000001001000101101110;
assign LUT_2[24500] = 32'b00000000000000000001110010000001;
assign LUT_2[24501] = 32'b11111111111111111110101010011010;
assign LUT_2[24502] = 32'b00000000000000001000101010111101;
assign LUT_2[24503] = 32'b00000000000000000101100011010110;
assign LUT_2[24504] = 32'b00000000000000000000000101110110;
assign LUT_2[24505] = 32'b11111111111111111100111110001111;
assign LUT_2[24506] = 32'b00000000000000000110111110110010;
assign LUT_2[24507] = 32'b00000000000000000011110111001011;
assign LUT_2[24508] = 32'b11111111111111111100100011011110;
assign LUT_2[24509] = 32'b11111111111111111001011011110111;
assign LUT_2[24510] = 32'b00000000000000000011011100011010;
assign LUT_2[24511] = 32'b00000000000000000000010100110011;
assign LUT_2[24512] = 32'b00000000000000000010011101001001;
assign LUT_2[24513] = 32'b11111111111111111111010101100010;
assign LUT_2[24514] = 32'b00000000000000001001010110000101;
assign LUT_2[24515] = 32'b00000000000000000110001110011110;
assign LUT_2[24516] = 32'b11111111111111111110111010110001;
assign LUT_2[24517] = 32'b11111111111111111011110011001010;
assign LUT_2[24518] = 32'b00000000000000000101110011101101;
assign LUT_2[24519] = 32'b00000000000000000010101100000110;
assign LUT_2[24520] = 32'b11111111111111111101001110100110;
assign LUT_2[24521] = 32'b11111111111111111010000110111111;
assign LUT_2[24522] = 32'b00000000000000000100000111100010;
assign LUT_2[24523] = 32'b00000000000000000000111111111011;
assign LUT_2[24524] = 32'b11111111111111111001101100001110;
assign LUT_2[24525] = 32'b11111111111111110110100100100111;
assign LUT_2[24526] = 32'b00000000000000000000100101001010;
assign LUT_2[24527] = 32'b11111111111111111101011101100011;
assign LUT_2[24528] = 32'b11111111111111111101000001010011;
assign LUT_2[24529] = 32'b11111111111111111001111001101100;
assign LUT_2[24530] = 32'b00000000000000000011111010001111;
assign LUT_2[24531] = 32'b00000000000000000000110010101000;
assign LUT_2[24532] = 32'b11111111111111111001011110111011;
assign LUT_2[24533] = 32'b11111111111111110110010111010100;
assign LUT_2[24534] = 32'b00000000000000000000010111110111;
assign LUT_2[24535] = 32'b11111111111111111101010000010000;
assign LUT_2[24536] = 32'b11111111111111110111110010110000;
assign LUT_2[24537] = 32'b11111111111111110100101011001001;
assign LUT_2[24538] = 32'b11111111111111111110101011101100;
assign LUT_2[24539] = 32'b11111111111111111011100100000101;
assign LUT_2[24540] = 32'b11111111111111110100010000011000;
assign LUT_2[24541] = 32'b11111111111111110001001000110001;
assign LUT_2[24542] = 32'b11111111111111111011001001010100;
assign LUT_2[24543] = 32'b11111111111111111000000001101101;
assign LUT_2[24544] = 32'b00000000000000000010111000110010;
assign LUT_2[24545] = 32'b11111111111111111111110001001011;
assign LUT_2[24546] = 32'b00000000000000001001110001101110;
assign LUT_2[24547] = 32'b00000000000000000110101010000111;
assign LUT_2[24548] = 32'b11111111111111111111010110011010;
assign LUT_2[24549] = 32'b11111111111111111100001110110011;
assign LUT_2[24550] = 32'b00000000000000000110001111010110;
assign LUT_2[24551] = 32'b00000000000000000011000111101111;
assign LUT_2[24552] = 32'b11111111111111111101101010001111;
assign LUT_2[24553] = 32'b11111111111111111010100010101000;
assign LUT_2[24554] = 32'b00000000000000000100100011001011;
assign LUT_2[24555] = 32'b00000000000000000001011011100100;
assign LUT_2[24556] = 32'b11111111111111111010000111110111;
assign LUT_2[24557] = 32'b11111111111111110111000000010000;
assign LUT_2[24558] = 32'b00000000000000000001000000110011;
assign LUT_2[24559] = 32'b11111111111111111101111001001100;
assign LUT_2[24560] = 32'b11111111111111111101011100111100;
assign LUT_2[24561] = 32'b11111111111111111010010101010101;
assign LUT_2[24562] = 32'b00000000000000000100010101111000;
assign LUT_2[24563] = 32'b00000000000000000001001110010001;
assign LUT_2[24564] = 32'b11111111111111111001111010100100;
assign LUT_2[24565] = 32'b11111111111111110110110010111101;
assign LUT_2[24566] = 32'b00000000000000000000110011100000;
assign LUT_2[24567] = 32'b11111111111111111101101011111001;
assign LUT_2[24568] = 32'b11111111111111111000001110011001;
assign LUT_2[24569] = 32'b11111111111111110101000110110010;
assign LUT_2[24570] = 32'b11111111111111111111000111010101;
assign LUT_2[24571] = 32'b11111111111111111011111111101110;
assign LUT_2[24572] = 32'b11111111111111110100101100000001;
assign LUT_2[24573] = 32'b11111111111111110001100100011010;
assign LUT_2[24574] = 32'b11111111111111111011100100111101;
assign LUT_2[24575] = 32'b11111111111111111000011101010110;
assign LUT_2[24576] = 32'b11111111111111110100111111110001;
assign LUT_2[24577] = 32'b11111111111111110001111000001010;
assign LUT_2[24578] = 32'b11111111111111111011111000101101;
assign LUT_2[24579] = 32'b11111111111111111000110001000110;
assign LUT_2[24580] = 32'b11111111111111110001011101011001;
assign LUT_2[24581] = 32'b11111111111111101110010101110010;
assign LUT_2[24582] = 32'b11111111111111111000010110010101;
assign LUT_2[24583] = 32'b11111111111111110101001110101110;
assign LUT_2[24584] = 32'b11111111111111101111110001001110;
assign LUT_2[24585] = 32'b11111111111111101100101001100111;
assign LUT_2[24586] = 32'b11111111111111110110101010001010;
assign LUT_2[24587] = 32'b11111111111111110011100010100011;
assign LUT_2[24588] = 32'b11111111111111101100001110110110;
assign LUT_2[24589] = 32'b11111111111111101001000111001111;
assign LUT_2[24590] = 32'b11111111111111110011000111110010;
assign LUT_2[24591] = 32'b11111111111111110000000000001011;
assign LUT_2[24592] = 32'b11111111111111101111100011111011;
assign LUT_2[24593] = 32'b11111111111111101100011100010100;
assign LUT_2[24594] = 32'b11111111111111110110011100110111;
assign LUT_2[24595] = 32'b11111111111111110011010101010000;
assign LUT_2[24596] = 32'b11111111111111101100000001100011;
assign LUT_2[24597] = 32'b11111111111111101000111001111100;
assign LUT_2[24598] = 32'b11111111111111110010111010011111;
assign LUT_2[24599] = 32'b11111111111111101111110010111000;
assign LUT_2[24600] = 32'b11111111111111101010010101011000;
assign LUT_2[24601] = 32'b11111111111111100111001101110001;
assign LUT_2[24602] = 32'b11111111111111110001001110010100;
assign LUT_2[24603] = 32'b11111111111111101110000110101101;
assign LUT_2[24604] = 32'b11111111111111100110110011000000;
assign LUT_2[24605] = 32'b11111111111111100011101011011001;
assign LUT_2[24606] = 32'b11111111111111101101101011111100;
assign LUT_2[24607] = 32'b11111111111111101010100100010101;
assign LUT_2[24608] = 32'b11111111111111110101011011011010;
assign LUT_2[24609] = 32'b11111111111111110010010011110011;
assign LUT_2[24610] = 32'b11111111111111111100010100010110;
assign LUT_2[24611] = 32'b11111111111111111001001100101111;
assign LUT_2[24612] = 32'b11111111111111110001111001000010;
assign LUT_2[24613] = 32'b11111111111111101110110001011011;
assign LUT_2[24614] = 32'b11111111111111111000110001111110;
assign LUT_2[24615] = 32'b11111111111111110101101010010111;
assign LUT_2[24616] = 32'b11111111111111110000001100110111;
assign LUT_2[24617] = 32'b11111111111111101101000101010000;
assign LUT_2[24618] = 32'b11111111111111110111000101110011;
assign LUT_2[24619] = 32'b11111111111111110011111110001100;
assign LUT_2[24620] = 32'b11111111111111101100101010011111;
assign LUT_2[24621] = 32'b11111111111111101001100010111000;
assign LUT_2[24622] = 32'b11111111111111110011100011011011;
assign LUT_2[24623] = 32'b11111111111111110000011011110100;
assign LUT_2[24624] = 32'b11111111111111101111111111100100;
assign LUT_2[24625] = 32'b11111111111111101100110111111101;
assign LUT_2[24626] = 32'b11111111111111110110111000100000;
assign LUT_2[24627] = 32'b11111111111111110011110000111001;
assign LUT_2[24628] = 32'b11111111111111101100011101001100;
assign LUT_2[24629] = 32'b11111111111111101001010101100101;
assign LUT_2[24630] = 32'b11111111111111110011010110001000;
assign LUT_2[24631] = 32'b11111111111111110000001110100001;
assign LUT_2[24632] = 32'b11111111111111101010110001000001;
assign LUT_2[24633] = 32'b11111111111111100111101001011010;
assign LUT_2[24634] = 32'b11111111111111110001101001111101;
assign LUT_2[24635] = 32'b11111111111111101110100010010110;
assign LUT_2[24636] = 32'b11111111111111100111001110101001;
assign LUT_2[24637] = 32'b11111111111111100100000111000010;
assign LUT_2[24638] = 32'b11111111111111101110000111100101;
assign LUT_2[24639] = 32'b11111111111111101010111111111110;
assign LUT_2[24640] = 32'b11111111111111101101001000010100;
assign LUT_2[24641] = 32'b11111111111111101010000000101101;
assign LUT_2[24642] = 32'b11111111111111110100000001010000;
assign LUT_2[24643] = 32'b11111111111111110000111001101001;
assign LUT_2[24644] = 32'b11111111111111101001100101111100;
assign LUT_2[24645] = 32'b11111111111111100110011110010101;
assign LUT_2[24646] = 32'b11111111111111110000011110111000;
assign LUT_2[24647] = 32'b11111111111111101101010111010001;
assign LUT_2[24648] = 32'b11111111111111100111111001110001;
assign LUT_2[24649] = 32'b11111111111111100100110010001010;
assign LUT_2[24650] = 32'b11111111111111101110110010101101;
assign LUT_2[24651] = 32'b11111111111111101011101011000110;
assign LUT_2[24652] = 32'b11111111111111100100010111011001;
assign LUT_2[24653] = 32'b11111111111111100001001111110010;
assign LUT_2[24654] = 32'b11111111111111101011010000010101;
assign LUT_2[24655] = 32'b11111111111111101000001000101110;
assign LUT_2[24656] = 32'b11111111111111100111101100011110;
assign LUT_2[24657] = 32'b11111111111111100100100100110111;
assign LUT_2[24658] = 32'b11111111111111101110100101011010;
assign LUT_2[24659] = 32'b11111111111111101011011101110011;
assign LUT_2[24660] = 32'b11111111111111100100001010000110;
assign LUT_2[24661] = 32'b11111111111111100001000010011111;
assign LUT_2[24662] = 32'b11111111111111101011000011000010;
assign LUT_2[24663] = 32'b11111111111111100111111011011011;
assign LUT_2[24664] = 32'b11111111111111100010011101111011;
assign LUT_2[24665] = 32'b11111111111111011111010110010100;
assign LUT_2[24666] = 32'b11111111111111101001010110110111;
assign LUT_2[24667] = 32'b11111111111111100110001111010000;
assign LUT_2[24668] = 32'b11111111111111011110111011100011;
assign LUT_2[24669] = 32'b11111111111111011011110011111100;
assign LUT_2[24670] = 32'b11111111111111100101110100011111;
assign LUT_2[24671] = 32'b11111111111111100010101100111000;
assign LUT_2[24672] = 32'b11111111111111101101100011111101;
assign LUT_2[24673] = 32'b11111111111111101010011100010110;
assign LUT_2[24674] = 32'b11111111111111110100011100111001;
assign LUT_2[24675] = 32'b11111111111111110001010101010010;
assign LUT_2[24676] = 32'b11111111111111101010000001100101;
assign LUT_2[24677] = 32'b11111111111111100110111001111110;
assign LUT_2[24678] = 32'b11111111111111110000111010100001;
assign LUT_2[24679] = 32'b11111111111111101101110010111010;
assign LUT_2[24680] = 32'b11111111111111101000010101011010;
assign LUT_2[24681] = 32'b11111111111111100101001101110011;
assign LUT_2[24682] = 32'b11111111111111101111001110010110;
assign LUT_2[24683] = 32'b11111111111111101100000110101111;
assign LUT_2[24684] = 32'b11111111111111100100110011000010;
assign LUT_2[24685] = 32'b11111111111111100001101011011011;
assign LUT_2[24686] = 32'b11111111111111101011101011111110;
assign LUT_2[24687] = 32'b11111111111111101000100100010111;
assign LUT_2[24688] = 32'b11111111111111101000001000000111;
assign LUT_2[24689] = 32'b11111111111111100101000000100000;
assign LUT_2[24690] = 32'b11111111111111101111000001000011;
assign LUT_2[24691] = 32'b11111111111111101011111001011100;
assign LUT_2[24692] = 32'b11111111111111100100100101101111;
assign LUT_2[24693] = 32'b11111111111111100001011110001000;
assign LUT_2[24694] = 32'b11111111111111101011011110101011;
assign LUT_2[24695] = 32'b11111111111111101000010111000100;
assign LUT_2[24696] = 32'b11111111111111100010111001100100;
assign LUT_2[24697] = 32'b11111111111111011111110001111101;
assign LUT_2[24698] = 32'b11111111111111101001110010100000;
assign LUT_2[24699] = 32'b11111111111111100110101010111001;
assign LUT_2[24700] = 32'b11111111111111011111010111001100;
assign LUT_2[24701] = 32'b11111111111111011100001111100101;
assign LUT_2[24702] = 32'b11111111111111100110010000001000;
assign LUT_2[24703] = 32'b11111111111111100011001000100001;
assign LUT_2[24704] = 32'b11111111111111111001010100000000;
assign LUT_2[24705] = 32'b11111111111111110110001100011001;
assign LUT_2[24706] = 32'b00000000000000000000001100111100;
assign LUT_2[24707] = 32'b11111111111111111101000101010101;
assign LUT_2[24708] = 32'b11111111111111110101110001101000;
assign LUT_2[24709] = 32'b11111111111111110010101010000001;
assign LUT_2[24710] = 32'b11111111111111111100101010100100;
assign LUT_2[24711] = 32'b11111111111111111001100010111101;
assign LUT_2[24712] = 32'b11111111111111110100000101011101;
assign LUT_2[24713] = 32'b11111111111111110000111101110110;
assign LUT_2[24714] = 32'b11111111111111111010111110011001;
assign LUT_2[24715] = 32'b11111111111111110111110110110010;
assign LUT_2[24716] = 32'b11111111111111110000100011000101;
assign LUT_2[24717] = 32'b11111111111111101101011011011110;
assign LUT_2[24718] = 32'b11111111111111110111011100000001;
assign LUT_2[24719] = 32'b11111111111111110100010100011010;
assign LUT_2[24720] = 32'b11111111111111110011111000001010;
assign LUT_2[24721] = 32'b11111111111111110000110000100011;
assign LUT_2[24722] = 32'b11111111111111111010110001000110;
assign LUT_2[24723] = 32'b11111111111111110111101001011111;
assign LUT_2[24724] = 32'b11111111111111110000010101110010;
assign LUT_2[24725] = 32'b11111111111111101101001110001011;
assign LUT_2[24726] = 32'b11111111111111110111001110101110;
assign LUT_2[24727] = 32'b11111111111111110100000111000111;
assign LUT_2[24728] = 32'b11111111111111101110101001100111;
assign LUT_2[24729] = 32'b11111111111111101011100010000000;
assign LUT_2[24730] = 32'b11111111111111110101100010100011;
assign LUT_2[24731] = 32'b11111111111111110010011010111100;
assign LUT_2[24732] = 32'b11111111111111101011000111001111;
assign LUT_2[24733] = 32'b11111111111111100111111111101000;
assign LUT_2[24734] = 32'b11111111111111110010000000001011;
assign LUT_2[24735] = 32'b11111111111111101110111000100100;
assign LUT_2[24736] = 32'b11111111111111111001101111101001;
assign LUT_2[24737] = 32'b11111111111111110110101000000010;
assign LUT_2[24738] = 32'b00000000000000000000101000100101;
assign LUT_2[24739] = 32'b11111111111111111101100000111110;
assign LUT_2[24740] = 32'b11111111111111110110001101010001;
assign LUT_2[24741] = 32'b11111111111111110011000101101010;
assign LUT_2[24742] = 32'b11111111111111111101000110001101;
assign LUT_2[24743] = 32'b11111111111111111001111110100110;
assign LUT_2[24744] = 32'b11111111111111110100100001000110;
assign LUT_2[24745] = 32'b11111111111111110001011001011111;
assign LUT_2[24746] = 32'b11111111111111111011011010000010;
assign LUT_2[24747] = 32'b11111111111111111000010010011011;
assign LUT_2[24748] = 32'b11111111111111110000111110101110;
assign LUT_2[24749] = 32'b11111111111111101101110111000111;
assign LUT_2[24750] = 32'b11111111111111110111110111101010;
assign LUT_2[24751] = 32'b11111111111111110100110000000011;
assign LUT_2[24752] = 32'b11111111111111110100010011110011;
assign LUT_2[24753] = 32'b11111111111111110001001100001100;
assign LUT_2[24754] = 32'b11111111111111111011001100101111;
assign LUT_2[24755] = 32'b11111111111111111000000101001000;
assign LUT_2[24756] = 32'b11111111111111110000110001011011;
assign LUT_2[24757] = 32'b11111111111111101101101001110100;
assign LUT_2[24758] = 32'b11111111111111110111101010010111;
assign LUT_2[24759] = 32'b11111111111111110100100010110000;
assign LUT_2[24760] = 32'b11111111111111101111000101010000;
assign LUT_2[24761] = 32'b11111111111111101011111101101001;
assign LUT_2[24762] = 32'b11111111111111110101111110001100;
assign LUT_2[24763] = 32'b11111111111111110010110110100101;
assign LUT_2[24764] = 32'b11111111111111101011100010111000;
assign LUT_2[24765] = 32'b11111111111111101000011011010001;
assign LUT_2[24766] = 32'b11111111111111110010011011110100;
assign LUT_2[24767] = 32'b11111111111111101111010100001101;
assign LUT_2[24768] = 32'b11111111111111110001011100100011;
assign LUT_2[24769] = 32'b11111111111111101110010100111100;
assign LUT_2[24770] = 32'b11111111111111111000010101011111;
assign LUT_2[24771] = 32'b11111111111111110101001101111000;
assign LUT_2[24772] = 32'b11111111111111101101111010001011;
assign LUT_2[24773] = 32'b11111111111111101010110010100100;
assign LUT_2[24774] = 32'b11111111111111110100110011000111;
assign LUT_2[24775] = 32'b11111111111111110001101011100000;
assign LUT_2[24776] = 32'b11111111111111101100001110000000;
assign LUT_2[24777] = 32'b11111111111111101001000110011001;
assign LUT_2[24778] = 32'b11111111111111110011000110111100;
assign LUT_2[24779] = 32'b11111111111111101111111111010101;
assign LUT_2[24780] = 32'b11111111111111101000101011101000;
assign LUT_2[24781] = 32'b11111111111111100101100100000001;
assign LUT_2[24782] = 32'b11111111111111101111100100100100;
assign LUT_2[24783] = 32'b11111111111111101100011100111101;
assign LUT_2[24784] = 32'b11111111111111101100000000101101;
assign LUT_2[24785] = 32'b11111111111111101000111001000110;
assign LUT_2[24786] = 32'b11111111111111110010111001101001;
assign LUT_2[24787] = 32'b11111111111111101111110010000010;
assign LUT_2[24788] = 32'b11111111111111101000011110010101;
assign LUT_2[24789] = 32'b11111111111111100101010110101110;
assign LUT_2[24790] = 32'b11111111111111101111010111010001;
assign LUT_2[24791] = 32'b11111111111111101100001111101010;
assign LUT_2[24792] = 32'b11111111111111100110110010001010;
assign LUT_2[24793] = 32'b11111111111111100011101010100011;
assign LUT_2[24794] = 32'b11111111111111101101101011000110;
assign LUT_2[24795] = 32'b11111111111111101010100011011111;
assign LUT_2[24796] = 32'b11111111111111100011001111110010;
assign LUT_2[24797] = 32'b11111111111111100000001000001011;
assign LUT_2[24798] = 32'b11111111111111101010001000101110;
assign LUT_2[24799] = 32'b11111111111111100111000001000111;
assign LUT_2[24800] = 32'b11111111111111110001111000001100;
assign LUT_2[24801] = 32'b11111111111111101110110000100101;
assign LUT_2[24802] = 32'b11111111111111111000110001001000;
assign LUT_2[24803] = 32'b11111111111111110101101001100001;
assign LUT_2[24804] = 32'b11111111111111101110010101110100;
assign LUT_2[24805] = 32'b11111111111111101011001110001101;
assign LUT_2[24806] = 32'b11111111111111110101001110110000;
assign LUT_2[24807] = 32'b11111111111111110010000111001001;
assign LUT_2[24808] = 32'b11111111111111101100101001101001;
assign LUT_2[24809] = 32'b11111111111111101001100010000010;
assign LUT_2[24810] = 32'b11111111111111110011100010100101;
assign LUT_2[24811] = 32'b11111111111111110000011010111110;
assign LUT_2[24812] = 32'b11111111111111101001000111010001;
assign LUT_2[24813] = 32'b11111111111111100101111111101010;
assign LUT_2[24814] = 32'b11111111111111110000000000001101;
assign LUT_2[24815] = 32'b11111111111111101100111000100110;
assign LUT_2[24816] = 32'b11111111111111101100011100010110;
assign LUT_2[24817] = 32'b11111111111111101001010100101111;
assign LUT_2[24818] = 32'b11111111111111110011010101010010;
assign LUT_2[24819] = 32'b11111111111111110000001101101011;
assign LUT_2[24820] = 32'b11111111111111101000111001111110;
assign LUT_2[24821] = 32'b11111111111111100101110010010111;
assign LUT_2[24822] = 32'b11111111111111101111110010111010;
assign LUT_2[24823] = 32'b11111111111111101100101011010011;
assign LUT_2[24824] = 32'b11111111111111100111001101110011;
assign LUT_2[24825] = 32'b11111111111111100100000110001100;
assign LUT_2[24826] = 32'b11111111111111101110000110101111;
assign LUT_2[24827] = 32'b11111111111111101010111111001000;
assign LUT_2[24828] = 32'b11111111111111100011101011011011;
assign LUT_2[24829] = 32'b11111111111111100000100011110100;
assign LUT_2[24830] = 32'b11111111111111101010100100010111;
assign LUT_2[24831] = 32'b11111111111111100111011100110000;
assign LUT_2[24832] = 32'b11111111111111111000111110010111;
assign LUT_2[24833] = 32'b11111111111111110101110110110000;
assign LUT_2[24834] = 32'b11111111111111111111110111010011;
assign LUT_2[24835] = 32'b11111111111111111100101111101100;
assign LUT_2[24836] = 32'b11111111111111110101011011111111;
assign LUT_2[24837] = 32'b11111111111111110010010100011000;
assign LUT_2[24838] = 32'b11111111111111111100010100111011;
assign LUT_2[24839] = 32'b11111111111111111001001101010100;
assign LUT_2[24840] = 32'b11111111111111110011101111110100;
assign LUT_2[24841] = 32'b11111111111111110000101000001101;
assign LUT_2[24842] = 32'b11111111111111111010101000110000;
assign LUT_2[24843] = 32'b11111111111111110111100001001001;
assign LUT_2[24844] = 32'b11111111111111110000001101011100;
assign LUT_2[24845] = 32'b11111111111111101101000101110101;
assign LUT_2[24846] = 32'b11111111111111110111000110011000;
assign LUT_2[24847] = 32'b11111111111111110011111110110001;
assign LUT_2[24848] = 32'b11111111111111110011100010100001;
assign LUT_2[24849] = 32'b11111111111111110000011010111010;
assign LUT_2[24850] = 32'b11111111111111111010011011011101;
assign LUT_2[24851] = 32'b11111111111111110111010011110110;
assign LUT_2[24852] = 32'b11111111111111110000000000001001;
assign LUT_2[24853] = 32'b11111111111111101100111000100010;
assign LUT_2[24854] = 32'b11111111111111110110111001000101;
assign LUT_2[24855] = 32'b11111111111111110011110001011110;
assign LUT_2[24856] = 32'b11111111111111101110010011111110;
assign LUT_2[24857] = 32'b11111111111111101011001100010111;
assign LUT_2[24858] = 32'b11111111111111110101001100111010;
assign LUT_2[24859] = 32'b11111111111111110010000101010011;
assign LUT_2[24860] = 32'b11111111111111101010110001100110;
assign LUT_2[24861] = 32'b11111111111111100111101001111111;
assign LUT_2[24862] = 32'b11111111111111110001101010100010;
assign LUT_2[24863] = 32'b11111111111111101110100010111011;
assign LUT_2[24864] = 32'b11111111111111111001011010000000;
assign LUT_2[24865] = 32'b11111111111111110110010010011001;
assign LUT_2[24866] = 32'b00000000000000000000010010111100;
assign LUT_2[24867] = 32'b11111111111111111101001011010101;
assign LUT_2[24868] = 32'b11111111111111110101110111101000;
assign LUT_2[24869] = 32'b11111111111111110010110000000001;
assign LUT_2[24870] = 32'b11111111111111111100110000100100;
assign LUT_2[24871] = 32'b11111111111111111001101000111101;
assign LUT_2[24872] = 32'b11111111111111110100001011011101;
assign LUT_2[24873] = 32'b11111111111111110001000011110110;
assign LUT_2[24874] = 32'b11111111111111111011000100011001;
assign LUT_2[24875] = 32'b11111111111111110111111100110010;
assign LUT_2[24876] = 32'b11111111111111110000101001000101;
assign LUT_2[24877] = 32'b11111111111111101101100001011110;
assign LUT_2[24878] = 32'b11111111111111110111100010000001;
assign LUT_2[24879] = 32'b11111111111111110100011010011010;
assign LUT_2[24880] = 32'b11111111111111110011111110001010;
assign LUT_2[24881] = 32'b11111111111111110000110110100011;
assign LUT_2[24882] = 32'b11111111111111111010110111000110;
assign LUT_2[24883] = 32'b11111111111111110111101111011111;
assign LUT_2[24884] = 32'b11111111111111110000011011110010;
assign LUT_2[24885] = 32'b11111111111111101101010100001011;
assign LUT_2[24886] = 32'b11111111111111110111010100101110;
assign LUT_2[24887] = 32'b11111111111111110100001101000111;
assign LUT_2[24888] = 32'b11111111111111101110101111100111;
assign LUT_2[24889] = 32'b11111111111111101011101000000000;
assign LUT_2[24890] = 32'b11111111111111110101101000100011;
assign LUT_2[24891] = 32'b11111111111111110010100000111100;
assign LUT_2[24892] = 32'b11111111111111101011001101001111;
assign LUT_2[24893] = 32'b11111111111111101000000101101000;
assign LUT_2[24894] = 32'b11111111111111110010000110001011;
assign LUT_2[24895] = 32'b11111111111111101110111110100100;
assign LUT_2[24896] = 32'b11111111111111110001000110111010;
assign LUT_2[24897] = 32'b11111111111111101101111111010011;
assign LUT_2[24898] = 32'b11111111111111110111111111110110;
assign LUT_2[24899] = 32'b11111111111111110100111000001111;
assign LUT_2[24900] = 32'b11111111111111101101100100100010;
assign LUT_2[24901] = 32'b11111111111111101010011100111011;
assign LUT_2[24902] = 32'b11111111111111110100011101011110;
assign LUT_2[24903] = 32'b11111111111111110001010101110111;
assign LUT_2[24904] = 32'b11111111111111101011111000010111;
assign LUT_2[24905] = 32'b11111111111111101000110000110000;
assign LUT_2[24906] = 32'b11111111111111110010110001010011;
assign LUT_2[24907] = 32'b11111111111111101111101001101100;
assign LUT_2[24908] = 32'b11111111111111101000010101111111;
assign LUT_2[24909] = 32'b11111111111111100101001110011000;
assign LUT_2[24910] = 32'b11111111111111101111001110111011;
assign LUT_2[24911] = 32'b11111111111111101100000111010100;
assign LUT_2[24912] = 32'b11111111111111101011101011000100;
assign LUT_2[24913] = 32'b11111111111111101000100011011101;
assign LUT_2[24914] = 32'b11111111111111110010100100000000;
assign LUT_2[24915] = 32'b11111111111111101111011100011001;
assign LUT_2[24916] = 32'b11111111111111101000001000101100;
assign LUT_2[24917] = 32'b11111111111111100101000001000101;
assign LUT_2[24918] = 32'b11111111111111101111000001101000;
assign LUT_2[24919] = 32'b11111111111111101011111010000001;
assign LUT_2[24920] = 32'b11111111111111100110011100100001;
assign LUT_2[24921] = 32'b11111111111111100011010100111010;
assign LUT_2[24922] = 32'b11111111111111101101010101011101;
assign LUT_2[24923] = 32'b11111111111111101010001101110110;
assign LUT_2[24924] = 32'b11111111111111100010111010001001;
assign LUT_2[24925] = 32'b11111111111111011111110010100010;
assign LUT_2[24926] = 32'b11111111111111101001110011000101;
assign LUT_2[24927] = 32'b11111111111111100110101011011110;
assign LUT_2[24928] = 32'b11111111111111110001100010100011;
assign LUT_2[24929] = 32'b11111111111111101110011010111100;
assign LUT_2[24930] = 32'b11111111111111111000011011011111;
assign LUT_2[24931] = 32'b11111111111111110101010011111000;
assign LUT_2[24932] = 32'b11111111111111101110000000001011;
assign LUT_2[24933] = 32'b11111111111111101010111000100100;
assign LUT_2[24934] = 32'b11111111111111110100111001000111;
assign LUT_2[24935] = 32'b11111111111111110001110001100000;
assign LUT_2[24936] = 32'b11111111111111101100010100000000;
assign LUT_2[24937] = 32'b11111111111111101001001100011001;
assign LUT_2[24938] = 32'b11111111111111110011001100111100;
assign LUT_2[24939] = 32'b11111111111111110000000101010101;
assign LUT_2[24940] = 32'b11111111111111101000110001101000;
assign LUT_2[24941] = 32'b11111111111111100101101010000001;
assign LUT_2[24942] = 32'b11111111111111101111101010100100;
assign LUT_2[24943] = 32'b11111111111111101100100010111101;
assign LUT_2[24944] = 32'b11111111111111101100000110101101;
assign LUT_2[24945] = 32'b11111111111111101000111111000110;
assign LUT_2[24946] = 32'b11111111111111110010111111101001;
assign LUT_2[24947] = 32'b11111111111111101111111000000010;
assign LUT_2[24948] = 32'b11111111111111101000100100010101;
assign LUT_2[24949] = 32'b11111111111111100101011100101110;
assign LUT_2[24950] = 32'b11111111111111101111011101010001;
assign LUT_2[24951] = 32'b11111111111111101100010101101010;
assign LUT_2[24952] = 32'b11111111111111100110111000001010;
assign LUT_2[24953] = 32'b11111111111111100011110000100011;
assign LUT_2[24954] = 32'b11111111111111101101110001000110;
assign LUT_2[24955] = 32'b11111111111111101010101001011111;
assign LUT_2[24956] = 32'b11111111111111100011010101110010;
assign LUT_2[24957] = 32'b11111111111111100000001110001011;
assign LUT_2[24958] = 32'b11111111111111101010001110101110;
assign LUT_2[24959] = 32'b11111111111111100111000111000111;
assign LUT_2[24960] = 32'b11111111111111111101010010100110;
assign LUT_2[24961] = 32'b11111111111111111010001010111111;
assign LUT_2[24962] = 32'b00000000000000000100001011100010;
assign LUT_2[24963] = 32'b00000000000000000001000011111011;
assign LUT_2[24964] = 32'b11111111111111111001110000001110;
assign LUT_2[24965] = 32'b11111111111111110110101000100111;
assign LUT_2[24966] = 32'b00000000000000000000101001001010;
assign LUT_2[24967] = 32'b11111111111111111101100001100011;
assign LUT_2[24968] = 32'b11111111111111111000000100000011;
assign LUT_2[24969] = 32'b11111111111111110100111100011100;
assign LUT_2[24970] = 32'b11111111111111111110111100111111;
assign LUT_2[24971] = 32'b11111111111111111011110101011000;
assign LUT_2[24972] = 32'b11111111111111110100100001101011;
assign LUT_2[24973] = 32'b11111111111111110001011010000100;
assign LUT_2[24974] = 32'b11111111111111111011011010100111;
assign LUT_2[24975] = 32'b11111111111111111000010011000000;
assign LUT_2[24976] = 32'b11111111111111110111110110110000;
assign LUT_2[24977] = 32'b11111111111111110100101111001001;
assign LUT_2[24978] = 32'b11111111111111111110101111101100;
assign LUT_2[24979] = 32'b11111111111111111011101000000101;
assign LUT_2[24980] = 32'b11111111111111110100010100011000;
assign LUT_2[24981] = 32'b11111111111111110001001100110001;
assign LUT_2[24982] = 32'b11111111111111111011001101010100;
assign LUT_2[24983] = 32'b11111111111111111000000101101101;
assign LUT_2[24984] = 32'b11111111111111110010101000001101;
assign LUT_2[24985] = 32'b11111111111111101111100000100110;
assign LUT_2[24986] = 32'b11111111111111111001100001001001;
assign LUT_2[24987] = 32'b11111111111111110110011001100010;
assign LUT_2[24988] = 32'b11111111111111101111000101110101;
assign LUT_2[24989] = 32'b11111111111111101011111110001110;
assign LUT_2[24990] = 32'b11111111111111110101111110110001;
assign LUT_2[24991] = 32'b11111111111111110010110111001010;
assign LUT_2[24992] = 32'b11111111111111111101101110001111;
assign LUT_2[24993] = 32'b11111111111111111010100110101000;
assign LUT_2[24994] = 32'b00000000000000000100100111001011;
assign LUT_2[24995] = 32'b00000000000000000001011111100100;
assign LUT_2[24996] = 32'b11111111111111111010001011110111;
assign LUT_2[24997] = 32'b11111111111111110111000100010000;
assign LUT_2[24998] = 32'b00000000000000000001000100110011;
assign LUT_2[24999] = 32'b11111111111111111101111101001100;
assign LUT_2[25000] = 32'b11111111111111111000011111101100;
assign LUT_2[25001] = 32'b11111111111111110101011000000101;
assign LUT_2[25002] = 32'b11111111111111111111011000101000;
assign LUT_2[25003] = 32'b11111111111111111100010001000001;
assign LUT_2[25004] = 32'b11111111111111110100111101010100;
assign LUT_2[25005] = 32'b11111111111111110001110101101101;
assign LUT_2[25006] = 32'b11111111111111111011110110010000;
assign LUT_2[25007] = 32'b11111111111111111000101110101001;
assign LUT_2[25008] = 32'b11111111111111111000010010011001;
assign LUT_2[25009] = 32'b11111111111111110101001010110010;
assign LUT_2[25010] = 32'b11111111111111111111001011010101;
assign LUT_2[25011] = 32'b11111111111111111100000011101110;
assign LUT_2[25012] = 32'b11111111111111110100110000000001;
assign LUT_2[25013] = 32'b11111111111111110001101000011010;
assign LUT_2[25014] = 32'b11111111111111111011101000111101;
assign LUT_2[25015] = 32'b11111111111111111000100001010110;
assign LUT_2[25016] = 32'b11111111111111110011000011110110;
assign LUT_2[25017] = 32'b11111111111111101111111100001111;
assign LUT_2[25018] = 32'b11111111111111111001111100110010;
assign LUT_2[25019] = 32'b11111111111111110110110101001011;
assign LUT_2[25020] = 32'b11111111111111101111100001011110;
assign LUT_2[25021] = 32'b11111111111111101100011001110111;
assign LUT_2[25022] = 32'b11111111111111110110011010011010;
assign LUT_2[25023] = 32'b11111111111111110011010010110011;
assign LUT_2[25024] = 32'b11111111111111110101011011001001;
assign LUT_2[25025] = 32'b11111111111111110010010011100010;
assign LUT_2[25026] = 32'b11111111111111111100010100000101;
assign LUT_2[25027] = 32'b11111111111111111001001100011110;
assign LUT_2[25028] = 32'b11111111111111110001111000110001;
assign LUT_2[25029] = 32'b11111111111111101110110001001010;
assign LUT_2[25030] = 32'b11111111111111111000110001101101;
assign LUT_2[25031] = 32'b11111111111111110101101010000110;
assign LUT_2[25032] = 32'b11111111111111110000001100100110;
assign LUT_2[25033] = 32'b11111111111111101101000100111111;
assign LUT_2[25034] = 32'b11111111111111110111000101100010;
assign LUT_2[25035] = 32'b11111111111111110011111101111011;
assign LUT_2[25036] = 32'b11111111111111101100101010001110;
assign LUT_2[25037] = 32'b11111111111111101001100010100111;
assign LUT_2[25038] = 32'b11111111111111110011100011001010;
assign LUT_2[25039] = 32'b11111111111111110000011011100011;
assign LUT_2[25040] = 32'b11111111111111101111111111010011;
assign LUT_2[25041] = 32'b11111111111111101100110111101100;
assign LUT_2[25042] = 32'b11111111111111110110111000001111;
assign LUT_2[25043] = 32'b11111111111111110011110000101000;
assign LUT_2[25044] = 32'b11111111111111101100011100111011;
assign LUT_2[25045] = 32'b11111111111111101001010101010100;
assign LUT_2[25046] = 32'b11111111111111110011010101110111;
assign LUT_2[25047] = 32'b11111111111111110000001110010000;
assign LUT_2[25048] = 32'b11111111111111101010110000110000;
assign LUT_2[25049] = 32'b11111111111111100111101001001001;
assign LUT_2[25050] = 32'b11111111111111110001101001101100;
assign LUT_2[25051] = 32'b11111111111111101110100010000101;
assign LUT_2[25052] = 32'b11111111111111100111001110011000;
assign LUT_2[25053] = 32'b11111111111111100100000110110001;
assign LUT_2[25054] = 32'b11111111111111101110000111010100;
assign LUT_2[25055] = 32'b11111111111111101010111111101101;
assign LUT_2[25056] = 32'b11111111111111110101110110110010;
assign LUT_2[25057] = 32'b11111111111111110010101111001011;
assign LUT_2[25058] = 32'b11111111111111111100101111101110;
assign LUT_2[25059] = 32'b11111111111111111001101000000111;
assign LUT_2[25060] = 32'b11111111111111110010010100011010;
assign LUT_2[25061] = 32'b11111111111111101111001100110011;
assign LUT_2[25062] = 32'b11111111111111111001001101010110;
assign LUT_2[25063] = 32'b11111111111111110110000101101111;
assign LUT_2[25064] = 32'b11111111111111110000101000001111;
assign LUT_2[25065] = 32'b11111111111111101101100000101000;
assign LUT_2[25066] = 32'b11111111111111110111100001001011;
assign LUT_2[25067] = 32'b11111111111111110100011001100100;
assign LUT_2[25068] = 32'b11111111111111101101000101110111;
assign LUT_2[25069] = 32'b11111111111111101001111110010000;
assign LUT_2[25070] = 32'b11111111111111110011111110110011;
assign LUT_2[25071] = 32'b11111111111111110000110111001100;
assign LUT_2[25072] = 32'b11111111111111110000011010111100;
assign LUT_2[25073] = 32'b11111111111111101101010011010101;
assign LUT_2[25074] = 32'b11111111111111110111010011111000;
assign LUT_2[25075] = 32'b11111111111111110100001100010001;
assign LUT_2[25076] = 32'b11111111111111101100111000100100;
assign LUT_2[25077] = 32'b11111111111111101001110000111101;
assign LUT_2[25078] = 32'b11111111111111110011110001100000;
assign LUT_2[25079] = 32'b11111111111111110000101001111001;
assign LUT_2[25080] = 32'b11111111111111101011001100011001;
assign LUT_2[25081] = 32'b11111111111111101000000100110010;
assign LUT_2[25082] = 32'b11111111111111110010000101010101;
assign LUT_2[25083] = 32'b11111111111111101110111101101110;
assign LUT_2[25084] = 32'b11111111111111100111101010000001;
assign LUT_2[25085] = 32'b11111111111111100100100010011010;
assign LUT_2[25086] = 32'b11111111111111101110100010111101;
assign LUT_2[25087] = 32'b11111111111111101011011011010110;
assign LUT_2[25088] = 32'b11111111111111111001110001100011;
assign LUT_2[25089] = 32'b11111111111111110110101001111100;
assign LUT_2[25090] = 32'b00000000000000000000101010011111;
assign LUT_2[25091] = 32'b11111111111111111101100010111000;
assign LUT_2[25092] = 32'b11111111111111110110001111001011;
assign LUT_2[25093] = 32'b11111111111111110011000111100100;
assign LUT_2[25094] = 32'b11111111111111111101001000000111;
assign LUT_2[25095] = 32'b11111111111111111010000000100000;
assign LUT_2[25096] = 32'b11111111111111110100100011000000;
assign LUT_2[25097] = 32'b11111111111111110001011011011001;
assign LUT_2[25098] = 32'b11111111111111111011011011111100;
assign LUT_2[25099] = 32'b11111111111111111000010100010101;
assign LUT_2[25100] = 32'b11111111111111110001000000101000;
assign LUT_2[25101] = 32'b11111111111111101101111001000001;
assign LUT_2[25102] = 32'b11111111111111110111111001100100;
assign LUT_2[25103] = 32'b11111111111111110100110001111101;
assign LUT_2[25104] = 32'b11111111111111110100010101101101;
assign LUT_2[25105] = 32'b11111111111111110001001110000110;
assign LUT_2[25106] = 32'b11111111111111111011001110101001;
assign LUT_2[25107] = 32'b11111111111111111000000111000010;
assign LUT_2[25108] = 32'b11111111111111110000110011010101;
assign LUT_2[25109] = 32'b11111111111111101101101011101110;
assign LUT_2[25110] = 32'b11111111111111110111101100010001;
assign LUT_2[25111] = 32'b11111111111111110100100100101010;
assign LUT_2[25112] = 32'b11111111111111101111000111001010;
assign LUT_2[25113] = 32'b11111111111111101011111111100011;
assign LUT_2[25114] = 32'b11111111111111110110000000000110;
assign LUT_2[25115] = 32'b11111111111111110010111000011111;
assign LUT_2[25116] = 32'b11111111111111101011100100110010;
assign LUT_2[25117] = 32'b11111111111111101000011101001011;
assign LUT_2[25118] = 32'b11111111111111110010011101101110;
assign LUT_2[25119] = 32'b11111111111111101111010110000111;
assign LUT_2[25120] = 32'b11111111111111111010001101001100;
assign LUT_2[25121] = 32'b11111111111111110111000101100101;
assign LUT_2[25122] = 32'b00000000000000000001000110001000;
assign LUT_2[25123] = 32'b11111111111111111101111110100001;
assign LUT_2[25124] = 32'b11111111111111110110101010110100;
assign LUT_2[25125] = 32'b11111111111111110011100011001101;
assign LUT_2[25126] = 32'b11111111111111111101100011110000;
assign LUT_2[25127] = 32'b11111111111111111010011100001001;
assign LUT_2[25128] = 32'b11111111111111110100111110101001;
assign LUT_2[25129] = 32'b11111111111111110001110111000010;
assign LUT_2[25130] = 32'b11111111111111111011110111100101;
assign LUT_2[25131] = 32'b11111111111111111000101111111110;
assign LUT_2[25132] = 32'b11111111111111110001011100010001;
assign LUT_2[25133] = 32'b11111111111111101110010100101010;
assign LUT_2[25134] = 32'b11111111111111111000010101001101;
assign LUT_2[25135] = 32'b11111111111111110101001101100110;
assign LUT_2[25136] = 32'b11111111111111110100110001010110;
assign LUT_2[25137] = 32'b11111111111111110001101001101111;
assign LUT_2[25138] = 32'b11111111111111111011101010010010;
assign LUT_2[25139] = 32'b11111111111111111000100010101011;
assign LUT_2[25140] = 32'b11111111111111110001001110111110;
assign LUT_2[25141] = 32'b11111111111111101110000111010111;
assign LUT_2[25142] = 32'b11111111111111111000000111111010;
assign LUT_2[25143] = 32'b11111111111111110101000000010011;
assign LUT_2[25144] = 32'b11111111111111101111100010110011;
assign LUT_2[25145] = 32'b11111111111111101100011011001100;
assign LUT_2[25146] = 32'b11111111111111110110011011101111;
assign LUT_2[25147] = 32'b11111111111111110011010100001000;
assign LUT_2[25148] = 32'b11111111111111101100000000011011;
assign LUT_2[25149] = 32'b11111111111111101000111000110100;
assign LUT_2[25150] = 32'b11111111111111110010111001010111;
assign LUT_2[25151] = 32'b11111111111111101111110001110000;
assign LUT_2[25152] = 32'b11111111111111110001111010000110;
assign LUT_2[25153] = 32'b11111111111111101110110010011111;
assign LUT_2[25154] = 32'b11111111111111111000110011000010;
assign LUT_2[25155] = 32'b11111111111111110101101011011011;
assign LUT_2[25156] = 32'b11111111111111101110010111101110;
assign LUT_2[25157] = 32'b11111111111111101011010000000111;
assign LUT_2[25158] = 32'b11111111111111110101010000101010;
assign LUT_2[25159] = 32'b11111111111111110010001001000011;
assign LUT_2[25160] = 32'b11111111111111101100101011100011;
assign LUT_2[25161] = 32'b11111111111111101001100011111100;
assign LUT_2[25162] = 32'b11111111111111110011100100011111;
assign LUT_2[25163] = 32'b11111111111111110000011100111000;
assign LUT_2[25164] = 32'b11111111111111101001001001001011;
assign LUT_2[25165] = 32'b11111111111111100110000001100100;
assign LUT_2[25166] = 32'b11111111111111110000000010000111;
assign LUT_2[25167] = 32'b11111111111111101100111010100000;
assign LUT_2[25168] = 32'b11111111111111101100011110010000;
assign LUT_2[25169] = 32'b11111111111111101001010110101001;
assign LUT_2[25170] = 32'b11111111111111110011010111001100;
assign LUT_2[25171] = 32'b11111111111111110000001111100101;
assign LUT_2[25172] = 32'b11111111111111101000111011111000;
assign LUT_2[25173] = 32'b11111111111111100101110100010001;
assign LUT_2[25174] = 32'b11111111111111101111110100110100;
assign LUT_2[25175] = 32'b11111111111111101100101101001101;
assign LUT_2[25176] = 32'b11111111111111100111001111101101;
assign LUT_2[25177] = 32'b11111111111111100100001000000110;
assign LUT_2[25178] = 32'b11111111111111101110001000101001;
assign LUT_2[25179] = 32'b11111111111111101011000001000010;
assign LUT_2[25180] = 32'b11111111111111100011101101010101;
assign LUT_2[25181] = 32'b11111111111111100000100101101110;
assign LUT_2[25182] = 32'b11111111111111101010100110010001;
assign LUT_2[25183] = 32'b11111111111111100111011110101010;
assign LUT_2[25184] = 32'b11111111111111110010010101101111;
assign LUT_2[25185] = 32'b11111111111111101111001110001000;
assign LUT_2[25186] = 32'b11111111111111111001001110101011;
assign LUT_2[25187] = 32'b11111111111111110110000111000100;
assign LUT_2[25188] = 32'b11111111111111101110110011010111;
assign LUT_2[25189] = 32'b11111111111111101011101011110000;
assign LUT_2[25190] = 32'b11111111111111110101101100010011;
assign LUT_2[25191] = 32'b11111111111111110010100100101100;
assign LUT_2[25192] = 32'b11111111111111101101000111001100;
assign LUT_2[25193] = 32'b11111111111111101001111111100101;
assign LUT_2[25194] = 32'b11111111111111110100000000001000;
assign LUT_2[25195] = 32'b11111111111111110000111000100001;
assign LUT_2[25196] = 32'b11111111111111101001100100110100;
assign LUT_2[25197] = 32'b11111111111111100110011101001101;
assign LUT_2[25198] = 32'b11111111111111110000011101110000;
assign LUT_2[25199] = 32'b11111111111111101101010110001001;
assign LUT_2[25200] = 32'b11111111111111101100111001111001;
assign LUT_2[25201] = 32'b11111111111111101001110010010010;
assign LUT_2[25202] = 32'b11111111111111110011110010110101;
assign LUT_2[25203] = 32'b11111111111111110000101011001110;
assign LUT_2[25204] = 32'b11111111111111101001010111100001;
assign LUT_2[25205] = 32'b11111111111111100110001111111010;
assign LUT_2[25206] = 32'b11111111111111110000010000011101;
assign LUT_2[25207] = 32'b11111111111111101101001000110110;
assign LUT_2[25208] = 32'b11111111111111100111101011010110;
assign LUT_2[25209] = 32'b11111111111111100100100011101111;
assign LUT_2[25210] = 32'b11111111111111101110100100010010;
assign LUT_2[25211] = 32'b11111111111111101011011100101011;
assign LUT_2[25212] = 32'b11111111111111100100001000111110;
assign LUT_2[25213] = 32'b11111111111111100001000001010111;
assign LUT_2[25214] = 32'b11111111111111101011000001111010;
assign LUT_2[25215] = 32'b11111111111111100111111010010011;
assign LUT_2[25216] = 32'b11111111111111111110000101110010;
assign LUT_2[25217] = 32'b11111111111111111010111110001011;
assign LUT_2[25218] = 32'b00000000000000000100111110101110;
assign LUT_2[25219] = 32'b00000000000000000001110111000111;
assign LUT_2[25220] = 32'b11111111111111111010100011011010;
assign LUT_2[25221] = 32'b11111111111111110111011011110011;
assign LUT_2[25222] = 32'b00000000000000000001011100010110;
assign LUT_2[25223] = 32'b11111111111111111110010100101111;
assign LUT_2[25224] = 32'b11111111111111111000110111001111;
assign LUT_2[25225] = 32'b11111111111111110101101111101000;
assign LUT_2[25226] = 32'b11111111111111111111110000001011;
assign LUT_2[25227] = 32'b11111111111111111100101000100100;
assign LUT_2[25228] = 32'b11111111111111110101010100110111;
assign LUT_2[25229] = 32'b11111111111111110010001101010000;
assign LUT_2[25230] = 32'b11111111111111111100001101110011;
assign LUT_2[25231] = 32'b11111111111111111001000110001100;
assign LUT_2[25232] = 32'b11111111111111111000101001111100;
assign LUT_2[25233] = 32'b11111111111111110101100010010101;
assign LUT_2[25234] = 32'b11111111111111111111100010111000;
assign LUT_2[25235] = 32'b11111111111111111100011011010001;
assign LUT_2[25236] = 32'b11111111111111110101000111100100;
assign LUT_2[25237] = 32'b11111111111111110001111111111101;
assign LUT_2[25238] = 32'b11111111111111111100000000100000;
assign LUT_2[25239] = 32'b11111111111111111000111000111001;
assign LUT_2[25240] = 32'b11111111111111110011011011011001;
assign LUT_2[25241] = 32'b11111111111111110000010011110010;
assign LUT_2[25242] = 32'b11111111111111111010010100010101;
assign LUT_2[25243] = 32'b11111111111111110111001100101110;
assign LUT_2[25244] = 32'b11111111111111101111111001000001;
assign LUT_2[25245] = 32'b11111111111111101100110001011010;
assign LUT_2[25246] = 32'b11111111111111110110110001111101;
assign LUT_2[25247] = 32'b11111111111111110011101010010110;
assign LUT_2[25248] = 32'b11111111111111111110100001011011;
assign LUT_2[25249] = 32'b11111111111111111011011001110100;
assign LUT_2[25250] = 32'b00000000000000000101011010010111;
assign LUT_2[25251] = 32'b00000000000000000010010010110000;
assign LUT_2[25252] = 32'b11111111111111111010111111000011;
assign LUT_2[25253] = 32'b11111111111111110111110111011100;
assign LUT_2[25254] = 32'b00000000000000000001110111111111;
assign LUT_2[25255] = 32'b11111111111111111110110000011000;
assign LUT_2[25256] = 32'b11111111111111111001010010111000;
assign LUT_2[25257] = 32'b11111111111111110110001011010001;
assign LUT_2[25258] = 32'b00000000000000000000001011110100;
assign LUT_2[25259] = 32'b11111111111111111101000100001101;
assign LUT_2[25260] = 32'b11111111111111110101110000100000;
assign LUT_2[25261] = 32'b11111111111111110010101000111001;
assign LUT_2[25262] = 32'b11111111111111111100101001011100;
assign LUT_2[25263] = 32'b11111111111111111001100001110101;
assign LUT_2[25264] = 32'b11111111111111111001000101100101;
assign LUT_2[25265] = 32'b11111111111111110101111101111110;
assign LUT_2[25266] = 32'b11111111111111111111111110100001;
assign LUT_2[25267] = 32'b11111111111111111100110110111010;
assign LUT_2[25268] = 32'b11111111111111110101100011001101;
assign LUT_2[25269] = 32'b11111111111111110010011011100110;
assign LUT_2[25270] = 32'b11111111111111111100011100001001;
assign LUT_2[25271] = 32'b11111111111111111001010100100010;
assign LUT_2[25272] = 32'b11111111111111110011110111000010;
assign LUT_2[25273] = 32'b11111111111111110000101111011011;
assign LUT_2[25274] = 32'b11111111111111111010101111111110;
assign LUT_2[25275] = 32'b11111111111111110111101000010111;
assign LUT_2[25276] = 32'b11111111111111110000010100101010;
assign LUT_2[25277] = 32'b11111111111111101101001101000011;
assign LUT_2[25278] = 32'b11111111111111110111001101100110;
assign LUT_2[25279] = 32'b11111111111111110100000101111111;
assign LUT_2[25280] = 32'b11111111111111110110001110010101;
assign LUT_2[25281] = 32'b11111111111111110011000110101110;
assign LUT_2[25282] = 32'b11111111111111111101000111010001;
assign LUT_2[25283] = 32'b11111111111111111001111111101010;
assign LUT_2[25284] = 32'b11111111111111110010101011111101;
assign LUT_2[25285] = 32'b11111111111111101111100100010110;
assign LUT_2[25286] = 32'b11111111111111111001100100111001;
assign LUT_2[25287] = 32'b11111111111111110110011101010010;
assign LUT_2[25288] = 32'b11111111111111110000111111110010;
assign LUT_2[25289] = 32'b11111111111111101101111000001011;
assign LUT_2[25290] = 32'b11111111111111110111111000101110;
assign LUT_2[25291] = 32'b11111111111111110100110001000111;
assign LUT_2[25292] = 32'b11111111111111101101011101011010;
assign LUT_2[25293] = 32'b11111111111111101010010101110011;
assign LUT_2[25294] = 32'b11111111111111110100010110010110;
assign LUT_2[25295] = 32'b11111111111111110001001110101111;
assign LUT_2[25296] = 32'b11111111111111110000110010011111;
assign LUT_2[25297] = 32'b11111111111111101101101010111000;
assign LUT_2[25298] = 32'b11111111111111110111101011011011;
assign LUT_2[25299] = 32'b11111111111111110100100011110100;
assign LUT_2[25300] = 32'b11111111111111101101010000000111;
assign LUT_2[25301] = 32'b11111111111111101010001000100000;
assign LUT_2[25302] = 32'b11111111111111110100001001000011;
assign LUT_2[25303] = 32'b11111111111111110001000001011100;
assign LUT_2[25304] = 32'b11111111111111101011100011111100;
assign LUT_2[25305] = 32'b11111111111111101000011100010101;
assign LUT_2[25306] = 32'b11111111111111110010011100111000;
assign LUT_2[25307] = 32'b11111111111111101111010101010001;
assign LUT_2[25308] = 32'b11111111111111101000000001100100;
assign LUT_2[25309] = 32'b11111111111111100100111001111101;
assign LUT_2[25310] = 32'b11111111111111101110111010100000;
assign LUT_2[25311] = 32'b11111111111111101011110010111001;
assign LUT_2[25312] = 32'b11111111111111110110101001111110;
assign LUT_2[25313] = 32'b11111111111111110011100010010111;
assign LUT_2[25314] = 32'b11111111111111111101100010111010;
assign LUT_2[25315] = 32'b11111111111111111010011011010011;
assign LUT_2[25316] = 32'b11111111111111110011000111100110;
assign LUT_2[25317] = 32'b11111111111111101111111111111111;
assign LUT_2[25318] = 32'b11111111111111111010000000100010;
assign LUT_2[25319] = 32'b11111111111111110110111000111011;
assign LUT_2[25320] = 32'b11111111111111110001011011011011;
assign LUT_2[25321] = 32'b11111111111111101110010011110100;
assign LUT_2[25322] = 32'b11111111111111111000010100010111;
assign LUT_2[25323] = 32'b11111111111111110101001100110000;
assign LUT_2[25324] = 32'b11111111111111101101111001000011;
assign LUT_2[25325] = 32'b11111111111111101010110001011100;
assign LUT_2[25326] = 32'b11111111111111110100110001111111;
assign LUT_2[25327] = 32'b11111111111111110001101010011000;
assign LUT_2[25328] = 32'b11111111111111110001001110001000;
assign LUT_2[25329] = 32'b11111111111111101110000110100001;
assign LUT_2[25330] = 32'b11111111111111111000000111000100;
assign LUT_2[25331] = 32'b11111111111111110100111111011101;
assign LUT_2[25332] = 32'b11111111111111101101101011110000;
assign LUT_2[25333] = 32'b11111111111111101010100100001001;
assign LUT_2[25334] = 32'b11111111111111110100100100101100;
assign LUT_2[25335] = 32'b11111111111111110001011101000101;
assign LUT_2[25336] = 32'b11111111111111101011111111100101;
assign LUT_2[25337] = 32'b11111111111111101000110111111110;
assign LUT_2[25338] = 32'b11111111111111110010111000100001;
assign LUT_2[25339] = 32'b11111111111111101111110000111010;
assign LUT_2[25340] = 32'b11111111111111101000011101001101;
assign LUT_2[25341] = 32'b11111111111111100101010101100110;
assign LUT_2[25342] = 32'b11111111111111101111010110001001;
assign LUT_2[25343] = 32'b11111111111111101100001110100010;
assign LUT_2[25344] = 32'b11111111111111111101110000001001;
assign LUT_2[25345] = 32'b11111111111111111010101000100010;
assign LUT_2[25346] = 32'b00000000000000000100101001000101;
assign LUT_2[25347] = 32'b00000000000000000001100001011110;
assign LUT_2[25348] = 32'b11111111111111111010001101110001;
assign LUT_2[25349] = 32'b11111111111111110111000110001010;
assign LUT_2[25350] = 32'b00000000000000000001000110101101;
assign LUT_2[25351] = 32'b11111111111111111101111111000110;
assign LUT_2[25352] = 32'b11111111111111111000100001100110;
assign LUT_2[25353] = 32'b11111111111111110101011001111111;
assign LUT_2[25354] = 32'b11111111111111111111011010100010;
assign LUT_2[25355] = 32'b11111111111111111100010010111011;
assign LUT_2[25356] = 32'b11111111111111110100111111001110;
assign LUT_2[25357] = 32'b11111111111111110001110111100111;
assign LUT_2[25358] = 32'b11111111111111111011111000001010;
assign LUT_2[25359] = 32'b11111111111111111000110000100011;
assign LUT_2[25360] = 32'b11111111111111111000010100010011;
assign LUT_2[25361] = 32'b11111111111111110101001100101100;
assign LUT_2[25362] = 32'b11111111111111111111001101001111;
assign LUT_2[25363] = 32'b11111111111111111100000101101000;
assign LUT_2[25364] = 32'b11111111111111110100110001111011;
assign LUT_2[25365] = 32'b11111111111111110001101010010100;
assign LUT_2[25366] = 32'b11111111111111111011101010110111;
assign LUT_2[25367] = 32'b11111111111111111000100011010000;
assign LUT_2[25368] = 32'b11111111111111110011000101110000;
assign LUT_2[25369] = 32'b11111111111111101111111110001001;
assign LUT_2[25370] = 32'b11111111111111111001111110101100;
assign LUT_2[25371] = 32'b11111111111111110110110111000101;
assign LUT_2[25372] = 32'b11111111111111101111100011011000;
assign LUT_2[25373] = 32'b11111111111111101100011011110001;
assign LUT_2[25374] = 32'b11111111111111110110011100010100;
assign LUT_2[25375] = 32'b11111111111111110011010100101101;
assign LUT_2[25376] = 32'b11111111111111111110001011110010;
assign LUT_2[25377] = 32'b11111111111111111011000100001011;
assign LUT_2[25378] = 32'b00000000000000000101000100101110;
assign LUT_2[25379] = 32'b00000000000000000001111101000111;
assign LUT_2[25380] = 32'b11111111111111111010101001011010;
assign LUT_2[25381] = 32'b11111111111111110111100001110011;
assign LUT_2[25382] = 32'b00000000000000000001100010010110;
assign LUT_2[25383] = 32'b11111111111111111110011010101111;
assign LUT_2[25384] = 32'b11111111111111111000111101001111;
assign LUT_2[25385] = 32'b11111111111111110101110101101000;
assign LUT_2[25386] = 32'b11111111111111111111110110001011;
assign LUT_2[25387] = 32'b11111111111111111100101110100100;
assign LUT_2[25388] = 32'b11111111111111110101011010110111;
assign LUT_2[25389] = 32'b11111111111111110010010011010000;
assign LUT_2[25390] = 32'b11111111111111111100010011110011;
assign LUT_2[25391] = 32'b11111111111111111001001100001100;
assign LUT_2[25392] = 32'b11111111111111111000101111111100;
assign LUT_2[25393] = 32'b11111111111111110101101000010101;
assign LUT_2[25394] = 32'b11111111111111111111101000111000;
assign LUT_2[25395] = 32'b11111111111111111100100001010001;
assign LUT_2[25396] = 32'b11111111111111110101001101100100;
assign LUT_2[25397] = 32'b11111111111111110010000101111101;
assign LUT_2[25398] = 32'b11111111111111111100000110100000;
assign LUT_2[25399] = 32'b11111111111111111000111110111001;
assign LUT_2[25400] = 32'b11111111111111110011100001011001;
assign LUT_2[25401] = 32'b11111111111111110000011001110010;
assign LUT_2[25402] = 32'b11111111111111111010011010010101;
assign LUT_2[25403] = 32'b11111111111111110111010010101110;
assign LUT_2[25404] = 32'b11111111111111101111111111000001;
assign LUT_2[25405] = 32'b11111111111111101100110111011010;
assign LUT_2[25406] = 32'b11111111111111110110110111111101;
assign LUT_2[25407] = 32'b11111111111111110011110000010110;
assign LUT_2[25408] = 32'b11111111111111110101111000101100;
assign LUT_2[25409] = 32'b11111111111111110010110001000101;
assign LUT_2[25410] = 32'b11111111111111111100110001101000;
assign LUT_2[25411] = 32'b11111111111111111001101010000001;
assign LUT_2[25412] = 32'b11111111111111110010010110010100;
assign LUT_2[25413] = 32'b11111111111111101111001110101101;
assign LUT_2[25414] = 32'b11111111111111111001001111010000;
assign LUT_2[25415] = 32'b11111111111111110110000111101001;
assign LUT_2[25416] = 32'b11111111111111110000101010001001;
assign LUT_2[25417] = 32'b11111111111111101101100010100010;
assign LUT_2[25418] = 32'b11111111111111110111100011000101;
assign LUT_2[25419] = 32'b11111111111111110100011011011110;
assign LUT_2[25420] = 32'b11111111111111101101000111110001;
assign LUT_2[25421] = 32'b11111111111111101010000000001010;
assign LUT_2[25422] = 32'b11111111111111110100000000101101;
assign LUT_2[25423] = 32'b11111111111111110000111001000110;
assign LUT_2[25424] = 32'b11111111111111110000011100110110;
assign LUT_2[25425] = 32'b11111111111111101101010101001111;
assign LUT_2[25426] = 32'b11111111111111110111010101110010;
assign LUT_2[25427] = 32'b11111111111111110100001110001011;
assign LUT_2[25428] = 32'b11111111111111101100111010011110;
assign LUT_2[25429] = 32'b11111111111111101001110010110111;
assign LUT_2[25430] = 32'b11111111111111110011110011011010;
assign LUT_2[25431] = 32'b11111111111111110000101011110011;
assign LUT_2[25432] = 32'b11111111111111101011001110010011;
assign LUT_2[25433] = 32'b11111111111111101000000110101100;
assign LUT_2[25434] = 32'b11111111111111110010000111001111;
assign LUT_2[25435] = 32'b11111111111111101110111111101000;
assign LUT_2[25436] = 32'b11111111111111100111101011111011;
assign LUT_2[25437] = 32'b11111111111111100100100100010100;
assign LUT_2[25438] = 32'b11111111111111101110100100110111;
assign LUT_2[25439] = 32'b11111111111111101011011101010000;
assign LUT_2[25440] = 32'b11111111111111110110010100010101;
assign LUT_2[25441] = 32'b11111111111111110011001100101110;
assign LUT_2[25442] = 32'b11111111111111111101001101010001;
assign LUT_2[25443] = 32'b11111111111111111010000101101010;
assign LUT_2[25444] = 32'b11111111111111110010110001111101;
assign LUT_2[25445] = 32'b11111111111111101111101010010110;
assign LUT_2[25446] = 32'b11111111111111111001101010111001;
assign LUT_2[25447] = 32'b11111111111111110110100011010010;
assign LUT_2[25448] = 32'b11111111111111110001000101110010;
assign LUT_2[25449] = 32'b11111111111111101101111110001011;
assign LUT_2[25450] = 32'b11111111111111110111111110101110;
assign LUT_2[25451] = 32'b11111111111111110100110111000111;
assign LUT_2[25452] = 32'b11111111111111101101100011011010;
assign LUT_2[25453] = 32'b11111111111111101010011011110011;
assign LUT_2[25454] = 32'b11111111111111110100011100010110;
assign LUT_2[25455] = 32'b11111111111111110001010100101111;
assign LUT_2[25456] = 32'b11111111111111110000111000011111;
assign LUT_2[25457] = 32'b11111111111111101101110000111000;
assign LUT_2[25458] = 32'b11111111111111110111110001011011;
assign LUT_2[25459] = 32'b11111111111111110100101001110100;
assign LUT_2[25460] = 32'b11111111111111101101010110000111;
assign LUT_2[25461] = 32'b11111111111111101010001110100000;
assign LUT_2[25462] = 32'b11111111111111110100001111000011;
assign LUT_2[25463] = 32'b11111111111111110001000111011100;
assign LUT_2[25464] = 32'b11111111111111101011101001111100;
assign LUT_2[25465] = 32'b11111111111111101000100010010101;
assign LUT_2[25466] = 32'b11111111111111110010100010111000;
assign LUT_2[25467] = 32'b11111111111111101111011011010001;
assign LUT_2[25468] = 32'b11111111111111101000000111100100;
assign LUT_2[25469] = 32'b11111111111111100100111111111101;
assign LUT_2[25470] = 32'b11111111111111101111000000100000;
assign LUT_2[25471] = 32'b11111111111111101011111000111001;
assign LUT_2[25472] = 32'b00000000000000000010000100011000;
assign LUT_2[25473] = 32'b11111111111111111110111100110001;
assign LUT_2[25474] = 32'b00000000000000001000111101010100;
assign LUT_2[25475] = 32'b00000000000000000101110101101101;
assign LUT_2[25476] = 32'b11111111111111111110100010000000;
assign LUT_2[25477] = 32'b11111111111111111011011010011001;
assign LUT_2[25478] = 32'b00000000000000000101011010111100;
assign LUT_2[25479] = 32'b00000000000000000010010011010101;
assign LUT_2[25480] = 32'b11111111111111111100110101110101;
assign LUT_2[25481] = 32'b11111111111111111001101110001110;
assign LUT_2[25482] = 32'b00000000000000000011101110110001;
assign LUT_2[25483] = 32'b00000000000000000000100111001010;
assign LUT_2[25484] = 32'b11111111111111111001010011011101;
assign LUT_2[25485] = 32'b11111111111111110110001011110110;
assign LUT_2[25486] = 32'b00000000000000000000001100011001;
assign LUT_2[25487] = 32'b11111111111111111101000100110010;
assign LUT_2[25488] = 32'b11111111111111111100101000100010;
assign LUT_2[25489] = 32'b11111111111111111001100000111011;
assign LUT_2[25490] = 32'b00000000000000000011100001011110;
assign LUT_2[25491] = 32'b00000000000000000000011001110111;
assign LUT_2[25492] = 32'b11111111111111111001000110001010;
assign LUT_2[25493] = 32'b11111111111111110101111110100011;
assign LUT_2[25494] = 32'b11111111111111111111111111000110;
assign LUT_2[25495] = 32'b11111111111111111100110111011111;
assign LUT_2[25496] = 32'b11111111111111110111011001111111;
assign LUT_2[25497] = 32'b11111111111111110100010010011000;
assign LUT_2[25498] = 32'b11111111111111111110010010111011;
assign LUT_2[25499] = 32'b11111111111111111011001011010100;
assign LUT_2[25500] = 32'b11111111111111110011110111100111;
assign LUT_2[25501] = 32'b11111111111111110000110000000000;
assign LUT_2[25502] = 32'b11111111111111111010110000100011;
assign LUT_2[25503] = 32'b11111111111111110111101000111100;
assign LUT_2[25504] = 32'b00000000000000000010100000000001;
assign LUT_2[25505] = 32'b11111111111111111111011000011010;
assign LUT_2[25506] = 32'b00000000000000001001011000111101;
assign LUT_2[25507] = 32'b00000000000000000110010001010110;
assign LUT_2[25508] = 32'b11111111111111111110111101101001;
assign LUT_2[25509] = 32'b11111111111111111011110110000010;
assign LUT_2[25510] = 32'b00000000000000000101110110100101;
assign LUT_2[25511] = 32'b00000000000000000010101110111110;
assign LUT_2[25512] = 32'b11111111111111111101010001011110;
assign LUT_2[25513] = 32'b11111111111111111010001001110111;
assign LUT_2[25514] = 32'b00000000000000000100001010011010;
assign LUT_2[25515] = 32'b00000000000000000001000010110011;
assign LUT_2[25516] = 32'b11111111111111111001101111000110;
assign LUT_2[25517] = 32'b11111111111111110110100111011111;
assign LUT_2[25518] = 32'b00000000000000000000101000000010;
assign LUT_2[25519] = 32'b11111111111111111101100000011011;
assign LUT_2[25520] = 32'b11111111111111111101000100001011;
assign LUT_2[25521] = 32'b11111111111111111001111100100100;
assign LUT_2[25522] = 32'b00000000000000000011111101000111;
assign LUT_2[25523] = 32'b00000000000000000000110101100000;
assign LUT_2[25524] = 32'b11111111111111111001100001110011;
assign LUT_2[25525] = 32'b11111111111111110110011010001100;
assign LUT_2[25526] = 32'b00000000000000000000011010101111;
assign LUT_2[25527] = 32'b11111111111111111101010011001000;
assign LUT_2[25528] = 32'b11111111111111110111110101101000;
assign LUT_2[25529] = 32'b11111111111111110100101110000001;
assign LUT_2[25530] = 32'b11111111111111111110101110100100;
assign LUT_2[25531] = 32'b11111111111111111011100110111101;
assign LUT_2[25532] = 32'b11111111111111110100010011010000;
assign LUT_2[25533] = 32'b11111111111111110001001011101001;
assign LUT_2[25534] = 32'b11111111111111111011001100001100;
assign LUT_2[25535] = 32'b11111111111111111000000100100101;
assign LUT_2[25536] = 32'b11111111111111111010001100111011;
assign LUT_2[25537] = 32'b11111111111111110111000101010100;
assign LUT_2[25538] = 32'b00000000000000000001000101110111;
assign LUT_2[25539] = 32'b11111111111111111101111110010000;
assign LUT_2[25540] = 32'b11111111111111110110101010100011;
assign LUT_2[25541] = 32'b11111111111111110011100010111100;
assign LUT_2[25542] = 32'b11111111111111111101100011011111;
assign LUT_2[25543] = 32'b11111111111111111010011011111000;
assign LUT_2[25544] = 32'b11111111111111110100111110011000;
assign LUT_2[25545] = 32'b11111111111111110001110110110001;
assign LUT_2[25546] = 32'b11111111111111111011110111010100;
assign LUT_2[25547] = 32'b11111111111111111000101111101101;
assign LUT_2[25548] = 32'b11111111111111110001011100000000;
assign LUT_2[25549] = 32'b11111111111111101110010100011001;
assign LUT_2[25550] = 32'b11111111111111111000010100111100;
assign LUT_2[25551] = 32'b11111111111111110101001101010101;
assign LUT_2[25552] = 32'b11111111111111110100110001000101;
assign LUT_2[25553] = 32'b11111111111111110001101001011110;
assign LUT_2[25554] = 32'b11111111111111111011101010000001;
assign LUT_2[25555] = 32'b11111111111111111000100010011010;
assign LUT_2[25556] = 32'b11111111111111110001001110101101;
assign LUT_2[25557] = 32'b11111111111111101110000111000110;
assign LUT_2[25558] = 32'b11111111111111111000000111101001;
assign LUT_2[25559] = 32'b11111111111111110101000000000010;
assign LUT_2[25560] = 32'b11111111111111101111100010100010;
assign LUT_2[25561] = 32'b11111111111111101100011010111011;
assign LUT_2[25562] = 32'b11111111111111110110011011011110;
assign LUT_2[25563] = 32'b11111111111111110011010011110111;
assign LUT_2[25564] = 32'b11111111111111101100000000001010;
assign LUT_2[25565] = 32'b11111111111111101000111000100011;
assign LUT_2[25566] = 32'b11111111111111110010111001000110;
assign LUT_2[25567] = 32'b11111111111111101111110001011111;
assign LUT_2[25568] = 32'b11111111111111111010101000100100;
assign LUT_2[25569] = 32'b11111111111111110111100000111101;
assign LUT_2[25570] = 32'b00000000000000000001100001100000;
assign LUT_2[25571] = 32'b11111111111111111110011001111001;
assign LUT_2[25572] = 32'b11111111111111110111000110001100;
assign LUT_2[25573] = 32'b11111111111111110011111110100101;
assign LUT_2[25574] = 32'b11111111111111111101111111001000;
assign LUT_2[25575] = 32'b11111111111111111010110111100001;
assign LUT_2[25576] = 32'b11111111111111110101011010000001;
assign LUT_2[25577] = 32'b11111111111111110010010010011010;
assign LUT_2[25578] = 32'b11111111111111111100010010111101;
assign LUT_2[25579] = 32'b11111111111111111001001011010110;
assign LUT_2[25580] = 32'b11111111111111110001110111101001;
assign LUT_2[25581] = 32'b11111111111111101110110000000010;
assign LUT_2[25582] = 32'b11111111111111111000110000100101;
assign LUT_2[25583] = 32'b11111111111111110101101000111110;
assign LUT_2[25584] = 32'b11111111111111110101001100101110;
assign LUT_2[25585] = 32'b11111111111111110010000101000111;
assign LUT_2[25586] = 32'b11111111111111111100000101101010;
assign LUT_2[25587] = 32'b11111111111111111000111110000011;
assign LUT_2[25588] = 32'b11111111111111110001101010010110;
assign LUT_2[25589] = 32'b11111111111111101110100010101111;
assign LUT_2[25590] = 32'b11111111111111111000100011010010;
assign LUT_2[25591] = 32'b11111111111111110101011011101011;
assign LUT_2[25592] = 32'b11111111111111101111111110001011;
assign LUT_2[25593] = 32'b11111111111111101100110110100100;
assign LUT_2[25594] = 32'b11111111111111110110110111000111;
assign LUT_2[25595] = 32'b11111111111111110011101111100000;
assign LUT_2[25596] = 32'b11111111111111101100011011110011;
assign LUT_2[25597] = 32'b11111111111111101001010100001100;
assign LUT_2[25598] = 32'b11111111111111110011010100101111;
assign LUT_2[25599] = 32'b11111111111111110000001101001000;
assign LUT_2[25600] = 32'b11111111111111111011101011110110;
assign LUT_2[25601] = 32'b11111111111111111000100100001111;
assign LUT_2[25602] = 32'b00000000000000000010100100110010;
assign LUT_2[25603] = 32'b11111111111111111111011101001011;
assign LUT_2[25604] = 32'b11111111111111111000001001011110;
assign LUT_2[25605] = 32'b11111111111111110101000001110111;
assign LUT_2[25606] = 32'b11111111111111111111000010011010;
assign LUT_2[25607] = 32'b11111111111111111011111010110011;
assign LUT_2[25608] = 32'b11111111111111110110011101010011;
assign LUT_2[25609] = 32'b11111111111111110011010101101100;
assign LUT_2[25610] = 32'b11111111111111111101010110001111;
assign LUT_2[25611] = 32'b11111111111111111010001110101000;
assign LUT_2[25612] = 32'b11111111111111110010111010111011;
assign LUT_2[25613] = 32'b11111111111111101111110011010100;
assign LUT_2[25614] = 32'b11111111111111111001110011110111;
assign LUT_2[25615] = 32'b11111111111111110110101100010000;
assign LUT_2[25616] = 32'b11111111111111110110010000000000;
assign LUT_2[25617] = 32'b11111111111111110011001000011001;
assign LUT_2[25618] = 32'b11111111111111111101001000111100;
assign LUT_2[25619] = 32'b11111111111111111010000001010101;
assign LUT_2[25620] = 32'b11111111111111110010101101101000;
assign LUT_2[25621] = 32'b11111111111111101111100110000001;
assign LUT_2[25622] = 32'b11111111111111111001100110100100;
assign LUT_2[25623] = 32'b11111111111111110110011110111101;
assign LUT_2[25624] = 32'b11111111111111110001000001011101;
assign LUT_2[25625] = 32'b11111111111111101101111001110110;
assign LUT_2[25626] = 32'b11111111111111110111111010011001;
assign LUT_2[25627] = 32'b11111111111111110100110010110010;
assign LUT_2[25628] = 32'b11111111111111101101011111000101;
assign LUT_2[25629] = 32'b11111111111111101010010111011110;
assign LUT_2[25630] = 32'b11111111111111110100011000000001;
assign LUT_2[25631] = 32'b11111111111111110001010000011010;
assign LUT_2[25632] = 32'b11111111111111111100000111011111;
assign LUT_2[25633] = 32'b11111111111111111000111111111000;
assign LUT_2[25634] = 32'b00000000000000000011000000011011;
assign LUT_2[25635] = 32'b11111111111111111111111000110100;
assign LUT_2[25636] = 32'b11111111111111111000100101000111;
assign LUT_2[25637] = 32'b11111111111111110101011101100000;
assign LUT_2[25638] = 32'b11111111111111111111011110000011;
assign LUT_2[25639] = 32'b11111111111111111100010110011100;
assign LUT_2[25640] = 32'b11111111111111110110111000111100;
assign LUT_2[25641] = 32'b11111111111111110011110001010101;
assign LUT_2[25642] = 32'b11111111111111111101110001111000;
assign LUT_2[25643] = 32'b11111111111111111010101010010001;
assign LUT_2[25644] = 32'b11111111111111110011010110100100;
assign LUT_2[25645] = 32'b11111111111111110000001110111101;
assign LUT_2[25646] = 32'b11111111111111111010001111100000;
assign LUT_2[25647] = 32'b11111111111111110111000111111001;
assign LUT_2[25648] = 32'b11111111111111110110101011101001;
assign LUT_2[25649] = 32'b11111111111111110011100100000010;
assign LUT_2[25650] = 32'b11111111111111111101100100100101;
assign LUT_2[25651] = 32'b11111111111111111010011100111110;
assign LUT_2[25652] = 32'b11111111111111110011001001010001;
assign LUT_2[25653] = 32'b11111111111111110000000001101010;
assign LUT_2[25654] = 32'b11111111111111111010000010001101;
assign LUT_2[25655] = 32'b11111111111111110110111010100110;
assign LUT_2[25656] = 32'b11111111111111110001011101000110;
assign LUT_2[25657] = 32'b11111111111111101110010101011111;
assign LUT_2[25658] = 32'b11111111111111111000010110000010;
assign LUT_2[25659] = 32'b11111111111111110101001110011011;
assign LUT_2[25660] = 32'b11111111111111101101111010101110;
assign LUT_2[25661] = 32'b11111111111111101010110011000111;
assign LUT_2[25662] = 32'b11111111111111110100110011101010;
assign LUT_2[25663] = 32'b11111111111111110001101100000011;
assign LUT_2[25664] = 32'b11111111111111110011110100011001;
assign LUT_2[25665] = 32'b11111111111111110000101100110010;
assign LUT_2[25666] = 32'b11111111111111111010101101010101;
assign LUT_2[25667] = 32'b11111111111111110111100101101110;
assign LUT_2[25668] = 32'b11111111111111110000010010000001;
assign LUT_2[25669] = 32'b11111111111111101101001010011010;
assign LUT_2[25670] = 32'b11111111111111110111001010111101;
assign LUT_2[25671] = 32'b11111111111111110100000011010110;
assign LUT_2[25672] = 32'b11111111111111101110100101110110;
assign LUT_2[25673] = 32'b11111111111111101011011110001111;
assign LUT_2[25674] = 32'b11111111111111110101011110110010;
assign LUT_2[25675] = 32'b11111111111111110010010111001011;
assign LUT_2[25676] = 32'b11111111111111101011000011011110;
assign LUT_2[25677] = 32'b11111111111111100111111011110111;
assign LUT_2[25678] = 32'b11111111111111110001111100011010;
assign LUT_2[25679] = 32'b11111111111111101110110100110011;
assign LUT_2[25680] = 32'b11111111111111101110011000100011;
assign LUT_2[25681] = 32'b11111111111111101011010000111100;
assign LUT_2[25682] = 32'b11111111111111110101010001011111;
assign LUT_2[25683] = 32'b11111111111111110010001001111000;
assign LUT_2[25684] = 32'b11111111111111101010110110001011;
assign LUT_2[25685] = 32'b11111111111111100111101110100100;
assign LUT_2[25686] = 32'b11111111111111110001101111000111;
assign LUT_2[25687] = 32'b11111111111111101110100111100000;
assign LUT_2[25688] = 32'b11111111111111101001001010000000;
assign LUT_2[25689] = 32'b11111111111111100110000010011001;
assign LUT_2[25690] = 32'b11111111111111110000000010111100;
assign LUT_2[25691] = 32'b11111111111111101100111011010101;
assign LUT_2[25692] = 32'b11111111111111100101100111101000;
assign LUT_2[25693] = 32'b11111111111111100010100000000001;
assign LUT_2[25694] = 32'b11111111111111101100100000100100;
assign LUT_2[25695] = 32'b11111111111111101001011000111101;
assign LUT_2[25696] = 32'b11111111111111110100010000000010;
assign LUT_2[25697] = 32'b11111111111111110001001000011011;
assign LUT_2[25698] = 32'b11111111111111111011001000111110;
assign LUT_2[25699] = 32'b11111111111111111000000001010111;
assign LUT_2[25700] = 32'b11111111111111110000101101101010;
assign LUT_2[25701] = 32'b11111111111111101101100110000011;
assign LUT_2[25702] = 32'b11111111111111110111100110100110;
assign LUT_2[25703] = 32'b11111111111111110100011110111111;
assign LUT_2[25704] = 32'b11111111111111101111000001011111;
assign LUT_2[25705] = 32'b11111111111111101011111001111000;
assign LUT_2[25706] = 32'b11111111111111110101111010011011;
assign LUT_2[25707] = 32'b11111111111111110010110010110100;
assign LUT_2[25708] = 32'b11111111111111101011011111000111;
assign LUT_2[25709] = 32'b11111111111111101000010111100000;
assign LUT_2[25710] = 32'b11111111111111110010011000000011;
assign LUT_2[25711] = 32'b11111111111111101111010000011100;
assign LUT_2[25712] = 32'b11111111111111101110110100001100;
assign LUT_2[25713] = 32'b11111111111111101011101100100101;
assign LUT_2[25714] = 32'b11111111111111110101101101001000;
assign LUT_2[25715] = 32'b11111111111111110010100101100001;
assign LUT_2[25716] = 32'b11111111111111101011010001110100;
assign LUT_2[25717] = 32'b11111111111111101000001010001101;
assign LUT_2[25718] = 32'b11111111111111110010001010110000;
assign LUT_2[25719] = 32'b11111111111111101111000011001001;
assign LUT_2[25720] = 32'b11111111111111101001100101101001;
assign LUT_2[25721] = 32'b11111111111111100110011110000010;
assign LUT_2[25722] = 32'b11111111111111110000011110100101;
assign LUT_2[25723] = 32'b11111111111111101101010110111110;
assign LUT_2[25724] = 32'b11111111111111100110000011010001;
assign LUT_2[25725] = 32'b11111111111111100010111011101010;
assign LUT_2[25726] = 32'b11111111111111101100111100001101;
assign LUT_2[25727] = 32'b11111111111111101001110100100110;
assign LUT_2[25728] = 32'b00000000000000000000000000000101;
assign LUT_2[25729] = 32'b11111111111111111100111000011110;
assign LUT_2[25730] = 32'b00000000000000000110111001000001;
assign LUT_2[25731] = 32'b00000000000000000011110001011010;
assign LUT_2[25732] = 32'b11111111111111111100011101101101;
assign LUT_2[25733] = 32'b11111111111111111001010110000110;
assign LUT_2[25734] = 32'b00000000000000000011010110101001;
assign LUT_2[25735] = 32'b00000000000000000000001111000010;
assign LUT_2[25736] = 32'b11111111111111111010110001100010;
assign LUT_2[25737] = 32'b11111111111111110111101001111011;
assign LUT_2[25738] = 32'b00000000000000000001101010011110;
assign LUT_2[25739] = 32'b11111111111111111110100010110111;
assign LUT_2[25740] = 32'b11111111111111110111001111001010;
assign LUT_2[25741] = 32'b11111111111111110100000111100011;
assign LUT_2[25742] = 32'b11111111111111111110001000000110;
assign LUT_2[25743] = 32'b11111111111111111011000000011111;
assign LUT_2[25744] = 32'b11111111111111111010100100001111;
assign LUT_2[25745] = 32'b11111111111111110111011100101000;
assign LUT_2[25746] = 32'b00000000000000000001011101001011;
assign LUT_2[25747] = 32'b11111111111111111110010101100100;
assign LUT_2[25748] = 32'b11111111111111110111000001110111;
assign LUT_2[25749] = 32'b11111111111111110011111010010000;
assign LUT_2[25750] = 32'b11111111111111111101111010110011;
assign LUT_2[25751] = 32'b11111111111111111010110011001100;
assign LUT_2[25752] = 32'b11111111111111110101010101101100;
assign LUT_2[25753] = 32'b11111111111111110010001110000101;
assign LUT_2[25754] = 32'b11111111111111111100001110101000;
assign LUT_2[25755] = 32'b11111111111111111001000111000001;
assign LUT_2[25756] = 32'b11111111111111110001110011010100;
assign LUT_2[25757] = 32'b11111111111111101110101011101101;
assign LUT_2[25758] = 32'b11111111111111111000101100010000;
assign LUT_2[25759] = 32'b11111111111111110101100100101001;
assign LUT_2[25760] = 32'b00000000000000000000011011101110;
assign LUT_2[25761] = 32'b11111111111111111101010100000111;
assign LUT_2[25762] = 32'b00000000000000000111010100101010;
assign LUT_2[25763] = 32'b00000000000000000100001101000011;
assign LUT_2[25764] = 32'b11111111111111111100111001010110;
assign LUT_2[25765] = 32'b11111111111111111001110001101111;
assign LUT_2[25766] = 32'b00000000000000000011110010010010;
assign LUT_2[25767] = 32'b00000000000000000000101010101011;
assign LUT_2[25768] = 32'b11111111111111111011001101001011;
assign LUT_2[25769] = 32'b11111111111111111000000101100100;
assign LUT_2[25770] = 32'b00000000000000000010000110000111;
assign LUT_2[25771] = 32'b11111111111111111110111110100000;
assign LUT_2[25772] = 32'b11111111111111110111101010110011;
assign LUT_2[25773] = 32'b11111111111111110100100011001100;
assign LUT_2[25774] = 32'b11111111111111111110100011101111;
assign LUT_2[25775] = 32'b11111111111111111011011100001000;
assign LUT_2[25776] = 32'b11111111111111111010111111111000;
assign LUT_2[25777] = 32'b11111111111111110111111000010001;
assign LUT_2[25778] = 32'b00000000000000000001111000110100;
assign LUT_2[25779] = 32'b11111111111111111110110001001101;
assign LUT_2[25780] = 32'b11111111111111110111011101100000;
assign LUT_2[25781] = 32'b11111111111111110100010101111001;
assign LUT_2[25782] = 32'b11111111111111111110010110011100;
assign LUT_2[25783] = 32'b11111111111111111011001110110101;
assign LUT_2[25784] = 32'b11111111111111110101110001010101;
assign LUT_2[25785] = 32'b11111111111111110010101001101110;
assign LUT_2[25786] = 32'b11111111111111111100101010010001;
assign LUT_2[25787] = 32'b11111111111111111001100010101010;
assign LUT_2[25788] = 32'b11111111111111110010001110111101;
assign LUT_2[25789] = 32'b11111111111111101111000111010110;
assign LUT_2[25790] = 32'b11111111111111111001000111111001;
assign LUT_2[25791] = 32'b11111111111111110110000000010010;
assign LUT_2[25792] = 32'b11111111111111111000001000101000;
assign LUT_2[25793] = 32'b11111111111111110101000001000001;
assign LUT_2[25794] = 32'b11111111111111111111000001100100;
assign LUT_2[25795] = 32'b11111111111111111011111001111101;
assign LUT_2[25796] = 32'b11111111111111110100100110010000;
assign LUT_2[25797] = 32'b11111111111111110001011110101001;
assign LUT_2[25798] = 32'b11111111111111111011011111001100;
assign LUT_2[25799] = 32'b11111111111111111000010111100101;
assign LUT_2[25800] = 32'b11111111111111110010111010000101;
assign LUT_2[25801] = 32'b11111111111111101111110010011110;
assign LUT_2[25802] = 32'b11111111111111111001110011000001;
assign LUT_2[25803] = 32'b11111111111111110110101011011010;
assign LUT_2[25804] = 32'b11111111111111101111010111101101;
assign LUT_2[25805] = 32'b11111111111111101100010000000110;
assign LUT_2[25806] = 32'b11111111111111110110010000101001;
assign LUT_2[25807] = 32'b11111111111111110011001001000010;
assign LUT_2[25808] = 32'b11111111111111110010101100110010;
assign LUT_2[25809] = 32'b11111111111111101111100101001011;
assign LUT_2[25810] = 32'b11111111111111111001100101101110;
assign LUT_2[25811] = 32'b11111111111111110110011110000111;
assign LUT_2[25812] = 32'b11111111111111101111001010011010;
assign LUT_2[25813] = 32'b11111111111111101100000010110011;
assign LUT_2[25814] = 32'b11111111111111110110000011010110;
assign LUT_2[25815] = 32'b11111111111111110010111011101111;
assign LUT_2[25816] = 32'b11111111111111101101011110001111;
assign LUT_2[25817] = 32'b11111111111111101010010110101000;
assign LUT_2[25818] = 32'b11111111111111110100010111001011;
assign LUT_2[25819] = 32'b11111111111111110001001111100100;
assign LUT_2[25820] = 32'b11111111111111101001111011110111;
assign LUT_2[25821] = 32'b11111111111111100110110100010000;
assign LUT_2[25822] = 32'b11111111111111110000110100110011;
assign LUT_2[25823] = 32'b11111111111111101101101101001100;
assign LUT_2[25824] = 32'b11111111111111111000100100010001;
assign LUT_2[25825] = 32'b11111111111111110101011100101010;
assign LUT_2[25826] = 32'b11111111111111111111011101001101;
assign LUT_2[25827] = 32'b11111111111111111100010101100110;
assign LUT_2[25828] = 32'b11111111111111110101000001111001;
assign LUT_2[25829] = 32'b11111111111111110001111010010010;
assign LUT_2[25830] = 32'b11111111111111111011111010110101;
assign LUT_2[25831] = 32'b11111111111111111000110011001110;
assign LUT_2[25832] = 32'b11111111111111110011010101101110;
assign LUT_2[25833] = 32'b11111111111111110000001110000111;
assign LUT_2[25834] = 32'b11111111111111111010001110101010;
assign LUT_2[25835] = 32'b11111111111111110111000111000011;
assign LUT_2[25836] = 32'b11111111111111101111110011010110;
assign LUT_2[25837] = 32'b11111111111111101100101011101111;
assign LUT_2[25838] = 32'b11111111111111110110101100010010;
assign LUT_2[25839] = 32'b11111111111111110011100100101011;
assign LUT_2[25840] = 32'b11111111111111110011001000011011;
assign LUT_2[25841] = 32'b11111111111111110000000000110100;
assign LUT_2[25842] = 32'b11111111111111111010000001010111;
assign LUT_2[25843] = 32'b11111111111111110110111001110000;
assign LUT_2[25844] = 32'b11111111111111101111100110000011;
assign LUT_2[25845] = 32'b11111111111111101100011110011100;
assign LUT_2[25846] = 32'b11111111111111110110011110111111;
assign LUT_2[25847] = 32'b11111111111111110011010111011000;
assign LUT_2[25848] = 32'b11111111111111101101111001111000;
assign LUT_2[25849] = 32'b11111111111111101010110010010001;
assign LUT_2[25850] = 32'b11111111111111110100110010110100;
assign LUT_2[25851] = 32'b11111111111111110001101011001101;
assign LUT_2[25852] = 32'b11111111111111101010010111100000;
assign LUT_2[25853] = 32'b11111111111111100111001111111001;
assign LUT_2[25854] = 32'b11111111111111110001010000011100;
assign LUT_2[25855] = 32'b11111111111111101110001000110101;
assign LUT_2[25856] = 32'b11111111111111111111101010011100;
assign LUT_2[25857] = 32'b11111111111111111100100010110101;
assign LUT_2[25858] = 32'b00000000000000000110100011011000;
assign LUT_2[25859] = 32'b00000000000000000011011011110001;
assign LUT_2[25860] = 32'b11111111111111111100001000000100;
assign LUT_2[25861] = 32'b11111111111111111001000000011101;
assign LUT_2[25862] = 32'b00000000000000000011000001000000;
assign LUT_2[25863] = 32'b11111111111111111111111001011001;
assign LUT_2[25864] = 32'b11111111111111111010011011111001;
assign LUT_2[25865] = 32'b11111111111111110111010100010010;
assign LUT_2[25866] = 32'b00000000000000000001010100110101;
assign LUT_2[25867] = 32'b11111111111111111110001101001110;
assign LUT_2[25868] = 32'b11111111111111110110111001100001;
assign LUT_2[25869] = 32'b11111111111111110011110001111010;
assign LUT_2[25870] = 32'b11111111111111111101110010011101;
assign LUT_2[25871] = 32'b11111111111111111010101010110110;
assign LUT_2[25872] = 32'b11111111111111111010001110100110;
assign LUT_2[25873] = 32'b11111111111111110111000110111111;
assign LUT_2[25874] = 32'b00000000000000000001000111100010;
assign LUT_2[25875] = 32'b11111111111111111101111111111011;
assign LUT_2[25876] = 32'b11111111111111110110101100001110;
assign LUT_2[25877] = 32'b11111111111111110011100100100111;
assign LUT_2[25878] = 32'b11111111111111111101100101001010;
assign LUT_2[25879] = 32'b11111111111111111010011101100011;
assign LUT_2[25880] = 32'b11111111111111110101000000000011;
assign LUT_2[25881] = 32'b11111111111111110001111000011100;
assign LUT_2[25882] = 32'b11111111111111111011111000111111;
assign LUT_2[25883] = 32'b11111111111111111000110001011000;
assign LUT_2[25884] = 32'b11111111111111110001011101101011;
assign LUT_2[25885] = 32'b11111111111111101110010110000100;
assign LUT_2[25886] = 32'b11111111111111111000010110100111;
assign LUT_2[25887] = 32'b11111111111111110101001111000000;
assign LUT_2[25888] = 32'b00000000000000000000000110000101;
assign LUT_2[25889] = 32'b11111111111111111100111110011110;
assign LUT_2[25890] = 32'b00000000000000000110111111000001;
assign LUT_2[25891] = 32'b00000000000000000011110111011010;
assign LUT_2[25892] = 32'b11111111111111111100100011101101;
assign LUT_2[25893] = 32'b11111111111111111001011100000110;
assign LUT_2[25894] = 32'b00000000000000000011011100101001;
assign LUT_2[25895] = 32'b00000000000000000000010101000010;
assign LUT_2[25896] = 32'b11111111111111111010110111100010;
assign LUT_2[25897] = 32'b11111111111111110111101111111011;
assign LUT_2[25898] = 32'b00000000000000000001110000011110;
assign LUT_2[25899] = 32'b11111111111111111110101000110111;
assign LUT_2[25900] = 32'b11111111111111110111010101001010;
assign LUT_2[25901] = 32'b11111111111111110100001101100011;
assign LUT_2[25902] = 32'b11111111111111111110001110000110;
assign LUT_2[25903] = 32'b11111111111111111011000110011111;
assign LUT_2[25904] = 32'b11111111111111111010101010001111;
assign LUT_2[25905] = 32'b11111111111111110111100010101000;
assign LUT_2[25906] = 32'b00000000000000000001100011001011;
assign LUT_2[25907] = 32'b11111111111111111110011011100100;
assign LUT_2[25908] = 32'b11111111111111110111000111110111;
assign LUT_2[25909] = 32'b11111111111111110100000000010000;
assign LUT_2[25910] = 32'b11111111111111111110000000110011;
assign LUT_2[25911] = 32'b11111111111111111010111001001100;
assign LUT_2[25912] = 32'b11111111111111110101011011101100;
assign LUT_2[25913] = 32'b11111111111111110010010100000101;
assign LUT_2[25914] = 32'b11111111111111111100010100101000;
assign LUT_2[25915] = 32'b11111111111111111001001101000001;
assign LUT_2[25916] = 32'b11111111111111110001111001010100;
assign LUT_2[25917] = 32'b11111111111111101110110001101101;
assign LUT_2[25918] = 32'b11111111111111111000110010010000;
assign LUT_2[25919] = 32'b11111111111111110101101010101001;
assign LUT_2[25920] = 32'b11111111111111110111110010111111;
assign LUT_2[25921] = 32'b11111111111111110100101011011000;
assign LUT_2[25922] = 32'b11111111111111111110101011111011;
assign LUT_2[25923] = 32'b11111111111111111011100100010100;
assign LUT_2[25924] = 32'b11111111111111110100010000100111;
assign LUT_2[25925] = 32'b11111111111111110001001001000000;
assign LUT_2[25926] = 32'b11111111111111111011001001100011;
assign LUT_2[25927] = 32'b11111111111111111000000001111100;
assign LUT_2[25928] = 32'b11111111111111110010100100011100;
assign LUT_2[25929] = 32'b11111111111111101111011100110101;
assign LUT_2[25930] = 32'b11111111111111111001011101011000;
assign LUT_2[25931] = 32'b11111111111111110110010101110001;
assign LUT_2[25932] = 32'b11111111111111101111000010000100;
assign LUT_2[25933] = 32'b11111111111111101011111010011101;
assign LUT_2[25934] = 32'b11111111111111110101111011000000;
assign LUT_2[25935] = 32'b11111111111111110010110011011001;
assign LUT_2[25936] = 32'b11111111111111110010010111001001;
assign LUT_2[25937] = 32'b11111111111111101111001111100010;
assign LUT_2[25938] = 32'b11111111111111111001010000000101;
assign LUT_2[25939] = 32'b11111111111111110110001000011110;
assign LUT_2[25940] = 32'b11111111111111101110110100110001;
assign LUT_2[25941] = 32'b11111111111111101011101101001010;
assign LUT_2[25942] = 32'b11111111111111110101101101101101;
assign LUT_2[25943] = 32'b11111111111111110010100110000110;
assign LUT_2[25944] = 32'b11111111111111101101001000100110;
assign LUT_2[25945] = 32'b11111111111111101010000000111111;
assign LUT_2[25946] = 32'b11111111111111110100000001100010;
assign LUT_2[25947] = 32'b11111111111111110000111001111011;
assign LUT_2[25948] = 32'b11111111111111101001100110001110;
assign LUT_2[25949] = 32'b11111111111111100110011110100111;
assign LUT_2[25950] = 32'b11111111111111110000011111001010;
assign LUT_2[25951] = 32'b11111111111111101101010111100011;
assign LUT_2[25952] = 32'b11111111111111111000001110101000;
assign LUT_2[25953] = 32'b11111111111111110101000111000001;
assign LUT_2[25954] = 32'b11111111111111111111000111100100;
assign LUT_2[25955] = 32'b11111111111111111011111111111101;
assign LUT_2[25956] = 32'b11111111111111110100101100010000;
assign LUT_2[25957] = 32'b11111111111111110001100100101001;
assign LUT_2[25958] = 32'b11111111111111111011100101001100;
assign LUT_2[25959] = 32'b11111111111111111000011101100101;
assign LUT_2[25960] = 32'b11111111111111110011000000000101;
assign LUT_2[25961] = 32'b11111111111111101111111000011110;
assign LUT_2[25962] = 32'b11111111111111111001111001000001;
assign LUT_2[25963] = 32'b11111111111111110110110001011010;
assign LUT_2[25964] = 32'b11111111111111101111011101101101;
assign LUT_2[25965] = 32'b11111111111111101100010110000110;
assign LUT_2[25966] = 32'b11111111111111110110010110101001;
assign LUT_2[25967] = 32'b11111111111111110011001111000010;
assign LUT_2[25968] = 32'b11111111111111110010110010110010;
assign LUT_2[25969] = 32'b11111111111111101111101011001011;
assign LUT_2[25970] = 32'b11111111111111111001101011101110;
assign LUT_2[25971] = 32'b11111111111111110110100100000111;
assign LUT_2[25972] = 32'b11111111111111101111010000011010;
assign LUT_2[25973] = 32'b11111111111111101100001000110011;
assign LUT_2[25974] = 32'b11111111111111110110001001010110;
assign LUT_2[25975] = 32'b11111111111111110011000001101111;
assign LUT_2[25976] = 32'b11111111111111101101100100001111;
assign LUT_2[25977] = 32'b11111111111111101010011100101000;
assign LUT_2[25978] = 32'b11111111111111110100011101001011;
assign LUT_2[25979] = 32'b11111111111111110001010101100100;
assign LUT_2[25980] = 32'b11111111111111101010000001110111;
assign LUT_2[25981] = 32'b11111111111111100110111010010000;
assign LUT_2[25982] = 32'b11111111111111110000111010110011;
assign LUT_2[25983] = 32'b11111111111111101101110011001100;
assign LUT_2[25984] = 32'b00000000000000000011111110101011;
assign LUT_2[25985] = 32'b00000000000000000000110111000100;
assign LUT_2[25986] = 32'b00000000000000001010110111100111;
assign LUT_2[25987] = 32'b00000000000000000111110000000000;
assign LUT_2[25988] = 32'b00000000000000000000011100010011;
assign LUT_2[25989] = 32'b11111111111111111101010100101100;
assign LUT_2[25990] = 32'b00000000000000000111010101001111;
assign LUT_2[25991] = 32'b00000000000000000100001101101000;
assign LUT_2[25992] = 32'b11111111111111111110110000001000;
assign LUT_2[25993] = 32'b11111111111111111011101000100001;
assign LUT_2[25994] = 32'b00000000000000000101101001000100;
assign LUT_2[25995] = 32'b00000000000000000010100001011101;
assign LUT_2[25996] = 32'b11111111111111111011001101110000;
assign LUT_2[25997] = 32'b11111111111111111000000110001001;
assign LUT_2[25998] = 32'b00000000000000000010000110101100;
assign LUT_2[25999] = 32'b11111111111111111110111111000101;
assign LUT_2[26000] = 32'b11111111111111111110100010110101;
assign LUT_2[26001] = 32'b11111111111111111011011011001110;
assign LUT_2[26002] = 32'b00000000000000000101011011110001;
assign LUT_2[26003] = 32'b00000000000000000010010100001010;
assign LUT_2[26004] = 32'b11111111111111111011000000011101;
assign LUT_2[26005] = 32'b11111111111111110111111000110110;
assign LUT_2[26006] = 32'b00000000000000000001111001011001;
assign LUT_2[26007] = 32'b11111111111111111110110001110010;
assign LUT_2[26008] = 32'b11111111111111111001010100010010;
assign LUT_2[26009] = 32'b11111111111111110110001100101011;
assign LUT_2[26010] = 32'b00000000000000000000001101001110;
assign LUT_2[26011] = 32'b11111111111111111101000101100111;
assign LUT_2[26012] = 32'b11111111111111110101110001111010;
assign LUT_2[26013] = 32'b11111111111111110010101010010011;
assign LUT_2[26014] = 32'b11111111111111111100101010110110;
assign LUT_2[26015] = 32'b11111111111111111001100011001111;
assign LUT_2[26016] = 32'b00000000000000000100011010010100;
assign LUT_2[26017] = 32'b00000000000000000001010010101101;
assign LUT_2[26018] = 32'b00000000000000001011010011010000;
assign LUT_2[26019] = 32'b00000000000000001000001011101001;
assign LUT_2[26020] = 32'b00000000000000000000110111111100;
assign LUT_2[26021] = 32'b11111111111111111101110000010101;
assign LUT_2[26022] = 32'b00000000000000000111110000111000;
assign LUT_2[26023] = 32'b00000000000000000100101001010001;
assign LUT_2[26024] = 32'b11111111111111111111001011110001;
assign LUT_2[26025] = 32'b11111111111111111100000100001010;
assign LUT_2[26026] = 32'b00000000000000000110000100101101;
assign LUT_2[26027] = 32'b00000000000000000010111101000110;
assign LUT_2[26028] = 32'b11111111111111111011101001011001;
assign LUT_2[26029] = 32'b11111111111111111000100001110010;
assign LUT_2[26030] = 32'b00000000000000000010100010010101;
assign LUT_2[26031] = 32'b11111111111111111111011010101110;
assign LUT_2[26032] = 32'b11111111111111111110111110011110;
assign LUT_2[26033] = 32'b11111111111111111011110110110111;
assign LUT_2[26034] = 32'b00000000000000000101110111011010;
assign LUT_2[26035] = 32'b00000000000000000010101111110011;
assign LUT_2[26036] = 32'b11111111111111111011011100000110;
assign LUT_2[26037] = 32'b11111111111111111000010100011111;
assign LUT_2[26038] = 32'b00000000000000000010010101000010;
assign LUT_2[26039] = 32'b11111111111111111111001101011011;
assign LUT_2[26040] = 32'b11111111111111111001101111111011;
assign LUT_2[26041] = 32'b11111111111111110110101000010100;
assign LUT_2[26042] = 32'b00000000000000000000101000110111;
assign LUT_2[26043] = 32'b11111111111111111101100001010000;
assign LUT_2[26044] = 32'b11111111111111110110001101100011;
assign LUT_2[26045] = 32'b11111111111111110011000101111100;
assign LUT_2[26046] = 32'b11111111111111111101000110011111;
assign LUT_2[26047] = 32'b11111111111111111001111110111000;
assign LUT_2[26048] = 32'b11111111111111111100000111001110;
assign LUT_2[26049] = 32'b11111111111111111000111111100111;
assign LUT_2[26050] = 32'b00000000000000000011000000001010;
assign LUT_2[26051] = 32'b11111111111111111111111000100011;
assign LUT_2[26052] = 32'b11111111111111111000100100110110;
assign LUT_2[26053] = 32'b11111111111111110101011101001111;
assign LUT_2[26054] = 32'b11111111111111111111011101110010;
assign LUT_2[26055] = 32'b11111111111111111100010110001011;
assign LUT_2[26056] = 32'b11111111111111110110111000101011;
assign LUT_2[26057] = 32'b11111111111111110011110001000100;
assign LUT_2[26058] = 32'b11111111111111111101110001100111;
assign LUT_2[26059] = 32'b11111111111111111010101010000000;
assign LUT_2[26060] = 32'b11111111111111110011010110010011;
assign LUT_2[26061] = 32'b11111111111111110000001110101100;
assign LUT_2[26062] = 32'b11111111111111111010001111001111;
assign LUT_2[26063] = 32'b11111111111111110111000111101000;
assign LUT_2[26064] = 32'b11111111111111110110101011011000;
assign LUT_2[26065] = 32'b11111111111111110011100011110001;
assign LUT_2[26066] = 32'b11111111111111111101100100010100;
assign LUT_2[26067] = 32'b11111111111111111010011100101101;
assign LUT_2[26068] = 32'b11111111111111110011001001000000;
assign LUT_2[26069] = 32'b11111111111111110000000001011001;
assign LUT_2[26070] = 32'b11111111111111111010000001111100;
assign LUT_2[26071] = 32'b11111111111111110110111010010101;
assign LUT_2[26072] = 32'b11111111111111110001011100110101;
assign LUT_2[26073] = 32'b11111111111111101110010101001110;
assign LUT_2[26074] = 32'b11111111111111111000010101110001;
assign LUT_2[26075] = 32'b11111111111111110101001110001010;
assign LUT_2[26076] = 32'b11111111111111101101111010011101;
assign LUT_2[26077] = 32'b11111111111111101010110010110110;
assign LUT_2[26078] = 32'b11111111111111110100110011011001;
assign LUT_2[26079] = 32'b11111111111111110001101011110010;
assign LUT_2[26080] = 32'b11111111111111111100100010110111;
assign LUT_2[26081] = 32'b11111111111111111001011011010000;
assign LUT_2[26082] = 32'b00000000000000000011011011110011;
assign LUT_2[26083] = 32'b00000000000000000000010100001100;
assign LUT_2[26084] = 32'b11111111111111111001000000011111;
assign LUT_2[26085] = 32'b11111111111111110101111000111000;
assign LUT_2[26086] = 32'b11111111111111111111111001011011;
assign LUT_2[26087] = 32'b11111111111111111100110001110100;
assign LUT_2[26088] = 32'b11111111111111110111010100010100;
assign LUT_2[26089] = 32'b11111111111111110100001100101101;
assign LUT_2[26090] = 32'b11111111111111111110001101010000;
assign LUT_2[26091] = 32'b11111111111111111011000101101001;
assign LUT_2[26092] = 32'b11111111111111110011110001111100;
assign LUT_2[26093] = 32'b11111111111111110000101010010101;
assign LUT_2[26094] = 32'b11111111111111111010101010111000;
assign LUT_2[26095] = 32'b11111111111111110111100011010001;
assign LUT_2[26096] = 32'b11111111111111110111000111000001;
assign LUT_2[26097] = 32'b11111111111111110011111111011010;
assign LUT_2[26098] = 32'b11111111111111111101111111111101;
assign LUT_2[26099] = 32'b11111111111111111010111000010110;
assign LUT_2[26100] = 32'b11111111111111110011100100101001;
assign LUT_2[26101] = 32'b11111111111111110000011101000010;
assign LUT_2[26102] = 32'b11111111111111111010011101100101;
assign LUT_2[26103] = 32'b11111111111111110111010101111110;
assign LUT_2[26104] = 32'b11111111111111110001111000011110;
assign LUT_2[26105] = 32'b11111111111111101110110000110111;
assign LUT_2[26106] = 32'b11111111111111111000110001011010;
assign LUT_2[26107] = 32'b11111111111111110101101001110011;
assign LUT_2[26108] = 32'b11111111111111101110010110000110;
assign LUT_2[26109] = 32'b11111111111111101011001110011111;
assign LUT_2[26110] = 32'b11111111111111110101001111000010;
assign LUT_2[26111] = 32'b11111111111111110010000111011011;
assign LUT_2[26112] = 32'b00000000000000000000011101101000;
assign LUT_2[26113] = 32'b11111111111111111101010110000001;
assign LUT_2[26114] = 32'b00000000000000000111010110100100;
assign LUT_2[26115] = 32'b00000000000000000100001110111101;
assign LUT_2[26116] = 32'b11111111111111111100111011010000;
assign LUT_2[26117] = 32'b11111111111111111001110011101001;
assign LUT_2[26118] = 32'b00000000000000000011110100001100;
assign LUT_2[26119] = 32'b00000000000000000000101100100101;
assign LUT_2[26120] = 32'b11111111111111111011001111000101;
assign LUT_2[26121] = 32'b11111111111111111000000111011110;
assign LUT_2[26122] = 32'b00000000000000000010001000000001;
assign LUT_2[26123] = 32'b11111111111111111111000000011010;
assign LUT_2[26124] = 32'b11111111111111110111101100101101;
assign LUT_2[26125] = 32'b11111111111111110100100101000110;
assign LUT_2[26126] = 32'b11111111111111111110100101101001;
assign LUT_2[26127] = 32'b11111111111111111011011110000010;
assign LUT_2[26128] = 32'b11111111111111111011000001110010;
assign LUT_2[26129] = 32'b11111111111111110111111010001011;
assign LUT_2[26130] = 32'b00000000000000000001111010101110;
assign LUT_2[26131] = 32'b11111111111111111110110011000111;
assign LUT_2[26132] = 32'b11111111111111110111011111011010;
assign LUT_2[26133] = 32'b11111111111111110100010111110011;
assign LUT_2[26134] = 32'b11111111111111111110011000010110;
assign LUT_2[26135] = 32'b11111111111111111011010000101111;
assign LUT_2[26136] = 32'b11111111111111110101110011001111;
assign LUT_2[26137] = 32'b11111111111111110010101011101000;
assign LUT_2[26138] = 32'b11111111111111111100101100001011;
assign LUT_2[26139] = 32'b11111111111111111001100100100100;
assign LUT_2[26140] = 32'b11111111111111110010010000110111;
assign LUT_2[26141] = 32'b11111111111111101111001001010000;
assign LUT_2[26142] = 32'b11111111111111111001001001110011;
assign LUT_2[26143] = 32'b11111111111111110110000010001100;
assign LUT_2[26144] = 32'b00000000000000000000111001010001;
assign LUT_2[26145] = 32'b11111111111111111101110001101010;
assign LUT_2[26146] = 32'b00000000000000000111110010001101;
assign LUT_2[26147] = 32'b00000000000000000100101010100110;
assign LUT_2[26148] = 32'b11111111111111111101010110111001;
assign LUT_2[26149] = 32'b11111111111111111010001111010010;
assign LUT_2[26150] = 32'b00000000000000000100001111110101;
assign LUT_2[26151] = 32'b00000000000000000001001000001110;
assign LUT_2[26152] = 32'b11111111111111111011101010101110;
assign LUT_2[26153] = 32'b11111111111111111000100011000111;
assign LUT_2[26154] = 32'b00000000000000000010100011101010;
assign LUT_2[26155] = 32'b11111111111111111111011100000011;
assign LUT_2[26156] = 32'b11111111111111111000001000010110;
assign LUT_2[26157] = 32'b11111111111111110101000000101111;
assign LUT_2[26158] = 32'b11111111111111111111000001010010;
assign LUT_2[26159] = 32'b11111111111111111011111001101011;
assign LUT_2[26160] = 32'b11111111111111111011011101011011;
assign LUT_2[26161] = 32'b11111111111111111000010101110100;
assign LUT_2[26162] = 32'b00000000000000000010010110010111;
assign LUT_2[26163] = 32'b11111111111111111111001110110000;
assign LUT_2[26164] = 32'b11111111111111110111111011000011;
assign LUT_2[26165] = 32'b11111111111111110100110011011100;
assign LUT_2[26166] = 32'b11111111111111111110110011111111;
assign LUT_2[26167] = 32'b11111111111111111011101100011000;
assign LUT_2[26168] = 32'b11111111111111110110001110111000;
assign LUT_2[26169] = 32'b11111111111111110011000111010001;
assign LUT_2[26170] = 32'b11111111111111111101000111110100;
assign LUT_2[26171] = 32'b11111111111111111010000000001101;
assign LUT_2[26172] = 32'b11111111111111110010101100100000;
assign LUT_2[26173] = 32'b11111111111111101111100100111001;
assign LUT_2[26174] = 32'b11111111111111111001100101011100;
assign LUT_2[26175] = 32'b11111111111111110110011101110101;
assign LUT_2[26176] = 32'b11111111111111111000100110001011;
assign LUT_2[26177] = 32'b11111111111111110101011110100100;
assign LUT_2[26178] = 32'b11111111111111111111011111000111;
assign LUT_2[26179] = 32'b11111111111111111100010111100000;
assign LUT_2[26180] = 32'b11111111111111110101000011110011;
assign LUT_2[26181] = 32'b11111111111111110001111100001100;
assign LUT_2[26182] = 32'b11111111111111111011111100101111;
assign LUT_2[26183] = 32'b11111111111111111000110101001000;
assign LUT_2[26184] = 32'b11111111111111110011010111101000;
assign LUT_2[26185] = 32'b11111111111111110000010000000001;
assign LUT_2[26186] = 32'b11111111111111111010010000100100;
assign LUT_2[26187] = 32'b11111111111111110111001000111101;
assign LUT_2[26188] = 32'b11111111111111101111110101010000;
assign LUT_2[26189] = 32'b11111111111111101100101101101001;
assign LUT_2[26190] = 32'b11111111111111110110101110001100;
assign LUT_2[26191] = 32'b11111111111111110011100110100101;
assign LUT_2[26192] = 32'b11111111111111110011001010010101;
assign LUT_2[26193] = 32'b11111111111111110000000010101110;
assign LUT_2[26194] = 32'b11111111111111111010000011010001;
assign LUT_2[26195] = 32'b11111111111111110110111011101010;
assign LUT_2[26196] = 32'b11111111111111101111100111111101;
assign LUT_2[26197] = 32'b11111111111111101100100000010110;
assign LUT_2[26198] = 32'b11111111111111110110100000111001;
assign LUT_2[26199] = 32'b11111111111111110011011001010010;
assign LUT_2[26200] = 32'b11111111111111101101111011110010;
assign LUT_2[26201] = 32'b11111111111111101010110100001011;
assign LUT_2[26202] = 32'b11111111111111110100110100101110;
assign LUT_2[26203] = 32'b11111111111111110001101101000111;
assign LUT_2[26204] = 32'b11111111111111101010011001011010;
assign LUT_2[26205] = 32'b11111111111111100111010001110011;
assign LUT_2[26206] = 32'b11111111111111110001010010010110;
assign LUT_2[26207] = 32'b11111111111111101110001010101111;
assign LUT_2[26208] = 32'b11111111111111111001000001110100;
assign LUT_2[26209] = 32'b11111111111111110101111010001101;
assign LUT_2[26210] = 32'b11111111111111111111111010110000;
assign LUT_2[26211] = 32'b11111111111111111100110011001001;
assign LUT_2[26212] = 32'b11111111111111110101011111011100;
assign LUT_2[26213] = 32'b11111111111111110010010111110101;
assign LUT_2[26214] = 32'b11111111111111111100011000011000;
assign LUT_2[26215] = 32'b11111111111111111001010000110001;
assign LUT_2[26216] = 32'b11111111111111110011110011010001;
assign LUT_2[26217] = 32'b11111111111111110000101011101010;
assign LUT_2[26218] = 32'b11111111111111111010101100001101;
assign LUT_2[26219] = 32'b11111111111111110111100100100110;
assign LUT_2[26220] = 32'b11111111111111110000010000111001;
assign LUT_2[26221] = 32'b11111111111111101101001001010010;
assign LUT_2[26222] = 32'b11111111111111110111001001110101;
assign LUT_2[26223] = 32'b11111111111111110100000010001110;
assign LUT_2[26224] = 32'b11111111111111110011100101111110;
assign LUT_2[26225] = 32'b11111111111111110000011110010111;
assign LUT_2[26226] = 32'b11111111111111111010011110111010;
assign LUT_2[26227] = 32'b11111111111111110111010111010011;
assign LUT_2[26228] = 32'b11111111111111110000000011100110;
assign LUT_2[26229] = 32'b11111111111111101100111011111111;
assign LUT_2[26230] = 32'b11111111111111110110111100100010;
assign LUT_2[26231] = 32'b11111111111111110011110100111011;
assign LUT_2[26232] = 32'b11111111111111101110010111011011;
assign LUT_2[26233] = 32'b11111111111111101011001111110100;
assign LUT_2[26234] = 32'b11111111111111110101010000010111;
assign LUT_2[26235] = 32'b11111111111111110010001000110000;
assign LUT_2[26236] = 32'b11111111111111101010110101000011;
assign LUT_2[26237] = 32'b11111111111111100111101101011100;
assign LUT_2[26238] = 32'b11111111111111110001101101111111;
assign LUT_2[26239] = 32'b11111111111111101110100110011000;
assign LUT_2[26240] = 32'b00000000000000000100110001110111;
assign LUT_2[26241] = 32'b00000000000000000001101010010000;
assign LUT_2[26242] = 32'b00000000000000001011101010110011;
assign LUT_2[26243] = 32'b00000000000000001000100011001100;
assign LUT_2[26244] = 32'b00000000000000000001001111011111;
assign LUT_2[26245] = 32'b11111111111111111110000111111000;
assign LUT_2[26246] = 32'b00000000000000001000001000011011;
assign LUT_2[26247] = 32'b00000000000000000101000000110100;
assign LUT_2[26248] = 32'b11111111111111111111100011010100;
assign LUT_2[26249] = 32'b11111111111111111100011011101101;
assign LUT_2[26250] = 32'b00000000000000000110011100010000;
assign LUT_2[26251] = 32'b00000000000000000011010100101001;
assign LUT_2[26252] = 32'b11111111111111111100000000111100;
assign LUT_2[26253] = 32'b11111111111111111000111001010101;
assign LUT_2[26254] = 32'b00000000000000000010111001111000;
assign LUT_2[26255] = 32'b11111111111111111111110010010001;
assign LUT_2[26256] = 32'b11111111111111111111010110000001;
assign LUT_2[26257] = 32'b11111111111111111100001110011010;
assign LUT_2[26258] = 32'b00000000000000000110001110111101;
assign LUT_2[26259] = 32'b00000000000000000011000111010110;
assign LUT_2[26260] = 32'b11111111111111111011110011101001;
assign LUT_2[26261] = 32'b11111111111111111000101100000010;
assign LUT_2[26262] = 32'b00000000000000000010101100100101;
assign LUT_2[26263] = 32'b11111111111111111111100100111110;
assign LUT_2[26264] = 32'b11111111111111111010000111011110;
assign LUT_2[26265] = 32'b11111111111111110110111111110111;
assign LUT_2[26266] = 32'b00000000000000000001000000011010;
assign LUT_2[26267] = 32'b11111111111111111101111000110011;
assign LUT_2[26268] = 32'b11111111111111110110100101000110;
assign LUT_2[26269] = 32'b11111111111111110011011101011111;
assign LUT_2[26270] = 32'b11111111111111111101011110000010;
assign LUT_2[26271] = 32'b11111111111111111010010110011011;
assign LUT_2[26272] = 32'b00000000000000000101001101100000;
assign LUT_2[26273] = 32'b00000000000000000010000101111001;
assign LUT_2[26274] = 32'b00000000000000001100000110011100;
assign LUT_2[26275] = 32'b00000000000000001000111110110101;
assign LUT_2[26276] = 32'b00000000000000000001101011001000;
assign LUT_2[26277] = 32'b11111111111111111110100011100001;
assign LUT_2[26278] = 32'b00000000000000001000100100000100;
assign LUT_2[26279] = 32'b00000000000000000101011100011101;
assign LUT_2[26280] = 32'b11111111111111111111111110111101;
assign LUT_2[26281] = 32'b11111111111111111100110111010110;
assign LUT_2[26282] = 32'b00000000000000000110110111111001;
assign LUT_2[26283] = 32'b00000000000000000011110000010010;
assign LUT_2[26284] = 32'b11111111111111111100011100100101;
assign LUT_2[26285] = 32'b11111111111111111001010100111110;
assign LUT_2[26286] = 32'b00000000000000000011010101100001;
assign LUT_2[26287] = 32'b00000000000000000000001101111010;
assign LUT_2[26288] = 32'b11111111111111111111110001101010;
assign LUT_2[26289] = 32'b11111111111111111100101010000011;
assign LUT_2[26290] = 32'b00000000000000000110101010100110;
assign LUT_2[26291] = 32'b00000000000000000011100010111111;
assign LUT_2[26292] = 32'b11111111111111111100001111010010;
assign LUT_2[26293] = 32'b11111111111111111001000111101011;
assign LUT_2[26294] = 32'b00000000000000000011001000001110;
assign LUT_2[26295] = 32'b00000000000000000000000000100111;
assign LUT_2[26296] = 32'b11111111111111111010100011000111;
assign LUT_2[26297] = 32'b11111111111111110111011011100000;
assign LUT_2[26298] = 32'b00000000000000000001011100000011;
assign LUT_2[26299] = 32'b11111111111111111110010100011100;
assign LUT_2[26300] = 32'b11111111111111110111000000101111;
assign LUT_2[26301] = 32'b11111111111111110011111001001000;
assign LUT_2[26302] = 32'b11111111111111111101111001101011;
assign LUT_2[26303] = 32'b11111111111111111010110010000100;
assign LUT_2[26304] = 32'b11111111111111111100111010011010;
assign LUT_2[26305] = 32'b11111111111111111001110010110011;
assign LUT_2[26306] = 32'b00000000000000000011110011010110;
assign LUT_2[26307] = 32'b00000000000000000000101011101111;
assign LUT_2[26308] = 32'b11111111111111111001011000000010;
assign LUT_2[26309] = 32'b11111111111111110110010000011011;
assign LUT_2[26310] = 32'b00000000000000000000010000111110;
assign LUT_2[26311] = 32'b11111111111111111101001001010111;
assign LUT_2[26312] = 32'b11111111111111110111101011110111;
assign LUT_2[26313] = 32'b11111111111111110100100100010000;
assign LUT_2[26314] = 32'b11111111111111111110100100110011;
assign LUT_2[26315] = 32'b11111111111111111011011101001100;
assign LUT_2[26316] = 32'b11111111111111110100001001011111;
assign LUT_2[26317] = 32'b11111111111111110001000001111000;
assign LUT_2[26318] = 32'b11111111111111111011000010011011;
assign LUT_2[26319] = 32'b11111111111111110111111010110100;
assign LUT_2[26320] = 32'b11111111111111110111011110100100;
assign LUT_2[26321] = 32'b11111111111111110100010110111101;
assign LUT_2[26322] = 32'b11111111111111111110010111100000;
assign LUT_2[26323] = 32'b11111111111111111011001111111001;
assign LUT_2[26324] = 32'b11111111111111110011111100001100;
assign LUT_2[26325] = 32'b11111111111111110000110100100101;
assign LUT_2[26326] = 32'b11111111111111111010110101001000;
assign LUT_2[26327] = 32'b11111111111111110111101101100001;
assign LUT_2[26328] = 32'b11111111111111110010010000000001;
assign LUT_2[26329] = 32'b11111111111111101111001000011010;
assign LUT_2[26330] = 32'b11111111111111111001001000111101;
assign LUT_2[26331] = 32'b11111111111111110110000001010110;
assign LUT_2[26332] = 32'b11111111111111101110101101101001;
assign LUT_2[26333] = 32'b11111111111111101011100110000010;
assign LUT_2[26334] = 32'b11111111111111110101100110100101;
assign LUT_2[26335] = 32'b11111111111111110010011110111110;
assign LUT_2[26336] = 32'b11111111111111111101010110000011;
assign LUT_2[26337] = 32'b11111111111111111010001110011100;
assign LUT_2[26338] = 32'b00000000000000000100001110111111;
assign LUT_2[26339] = 32'b00000000000000000001000111011000;
assign LUT_2[26340] = 32'b11111111111111111001110011101011;
assign LUT_2[26341] = 32'b11111111111111110110101100000100;
assign LUT_2[26342] = 32'b00000000000000000000101100100111;
assign LUT_2[26343] = 32'b11111111111111111101100101000000;
assign LUT_2[26344] = 32'b11111111111111111000000111100000;
assign LUT_2[26345] = 32'b11111111111111110100111111111001;
assign LUT_2[26346] = 32'b11111111111111111111000000011100;
assign LUT_2[26347] = 32'b11111111111111111011111000110101;
assign LUT_2[26348] = 32'b11111111111111110100100101001000;
assign LUT_2[26349] = 32'b11111111111111110001011101100001;
assign LUT_2[26350] = 32'b11111111111111111011011110000100;
assign LUT_2[26351] = 32'b11111111111111111000010110011101;
assign LUT_2[26352] = 32'b11111111111111110111111010001101;
assign LUT_2[26353] = 32'b11111111111111110100110010100110;
assign LUT_2[26354] = 32'b11111111111111111110110011001001;
assign LUT_2[26355] = 32'b11111111111111111011101011100010;
assign LUT_2[26356] = 32'b11111111111111110100010111110101;
assign LUT_2[26357] = 32'b11111111111111110001010000001110;
assign LUT_2[26358] = 32'b11111111111111111011010000110001;
assign LUT_2[26359] = 32'b11111111111111111000001001001010;
assign LUT_2[26360] = 32'b11111111111111110010101011101010;
assign LUT_2[26361] = 32'b11111111111111101111100100000011;
assign LUT_2[26362] = 32'b11111111111111111001100100100110;
assign LUT_2[26363] = 32'b11111111111111110110011100111111;
assign LUT_2[26364] = 32'b11111111111111101111001001010010;
assign LUT_2[26365] = 32'b11111111111111101100000001101011;
assign LUT_2[26366] = 32'b11111111111111110110000010001110;
assign LUT_2[26367] = 32'b11111111111111110010111010100111;
assign LUT_2[26368] = 32'b00000000000000000100011100001110;
assign LUT_2[26369] = 32'b00000000000000000001010100100111;
assign LUT_2[26370] = 32'b00000000000000001011010101001010;
assign LUT_2[26371] = 32'b00000000000000001000001101100011;
assign LUT_2[26372] = 32'b00000000000000000000111001110110;
assign LUT_2[26373] = 32'b11111111111111111101110010001111;
assign LUT_2[26374] = 32'b00000000000000000111110010110010;
assign LUT_2[26375] = 32'b00000000000000000100101011001011;
assign LUT_2[26376] = 32'b11111111111111111111001101101011;
assign LUT_2[26377] = 32'b11111111111111111100000110000100;
assign LUT_2[26378] = 32'b00000000000000000110000110100111;
assign LUT_2[26379] = 32'b00000000000000000010111111000000;
assign LUT_2[26380] = 32'b11111111111111111011101011010011;
assign LUT_2[26381] = 32'b11111111111111111000100011101100;
assign LUT_2[26382] = 32'b00000000000000000010100100001111;
assign LUT_2[26383] = 32'b11111111111111111111011100101000;
assign LUT_2[26384] = 32'b11111111111111111111000000011000;
assign LUT_2[26385] = 32'b11111111111111111011111000110001;
assign LUT_2[26386] = 32'b00000000000000000101111001010100;
assign LUT_2[26387] = 32'b00000000000000000010110001101101;
assign LUT_2[26388] = 32'b11111111111111111011011110000000;
assign LUT_2[26389] = 32'b11111111111111111000010110011001;
assign LUT_2[26390] = 32'b00000000000000000010010110111100;
assign LUT_2[26391] = 32'b11111111111111111111001111010101;
assign LUT_2[26392] = 32'b11111111111111111001110001110101;
assign LUT_2[26393] = 32'b11111111111111110110101010001110;
assign LUT_2[26394] = 32'b00000000000000000000101010110001;
assign LUT_2[26395] = 32'b11111111111111111101100011001010;
assign LUT_2[26396] = 32'b11111111111111110110001111011101;
assign LUT_2[26397] = 32'b11111111111111110011000111110110;
assign LUT_2[26398] = 32'b11111111111111111101001000011001;
assign LUT_2[26399] = 32'b11111111111111111010000000110010;
assign LUT_2[26400] = 32'b00000000000000000100110111110111;
assign LUT_2[26401] = 32'b00000000000000000001110000010000;
assign LUT_2[26402] = 32'b00000000000000001011110000110011;
assign LUT_2[26403] = 32'b00000000000000001000101001001100;
assign LUT_2[26404] = 32'b00000000000000000001010101011111;
assign LUT_2[26405] = 32'b11111111111111111110001101111000;
assign LUT_2[26406] = 32'b00000000000000001000001110011011;
assign LUT_2[26407] = 32'b00000000000000000101000110110100;
assign LUT_2[26408] = 32'b11111111111111111111101001010100;
assign LUT_2[26409] = 32'b11111111111111111100100001101101;
assign LUT_2[26410] = 32'b00000000000000000110100010010000;
assign LUT_2[26411] = 32'b00000000000000000011011010101001;
assign LUT_2[26412] = 32'b11111111111111111100000110111100;
assign LUT_2[26413] = 32'b11111111111111111000111111010101;
assign LUT_2[26414] = 32'b00000000000000000010111111111000;
assign LUT_2[26415] = 32'b11111111111111111111111000010001;
assign LUT_2[26416] = 32'b11111111111111111111011100000001;
assign LUT_2[26417] = 32'b11111111111111111100010100011010;
assign LUT_2[26418] = 32'b00000000000000000110010100111101;
assign LUT_2[26419] = 32'b00000000000000000011001101010110;
assign LUT_2[26420] = 32'b11111111111111111011111001101001;
assign LUT_2[26421] = 32'b11111111111111111000110010000010;
assign LUT_2[26422] = 32'b00000000000000000010110010100101;
assign LUT_2[26423] = 32'b11111111111111111111101010111110;
assign LUT_2[26424] = 32'b11111111111111111010001101011110;
assign LUT_2[26425] = 32'b11111111111111110111000101110111;
assign LUT_2[26426] = 32'b00000000000000000001000110011010;
assign LUT_2[26427] = 32'b11111111111111111101111110110011;
assign LUT_2[26428] = 32'b11111111111111110110101011000110;
assign LUT_2[26429] = 32'b11111111111111110011100011011111;
assign LUT_2[26430] = 32'b11111111111111111101100100000010;
assign LUT_2[26431] = 32'b11111111111111111010011100011011;
assign LUT_2[26432] = 32'b11111111111111111100100100110001;
assign LUT_2[26433] = 32'b11111111111111111001011101001010;
assign LUT_2[26434] = 32'b00000000000000000011011101101101;
assign LUT_2[26435] = 32'b00000000000000000000010110000110;
assign LUT_2[26436] = 32'b11111111111111111001000010011001;
assign LUT_2[26437] = 32'b11111111111111110101111010110010;
assign LUT_2[26438] = 32'b11111111111111111111111011010101;
assign LUT_2[26439] = 32'b11111111111111111100110011101110;
assign LUT_2[26440] = 32'b11111111111111110111010110001110;
assign LUT_2[26441] = 32'b11111111111111110100001110100111;
assign LUT_2[26442] = 32'b11111111111111111110001111001010;
assign LUT_2[26443] = 32'b11111111111111111011000111100011;
assign LUT_2[26444] = 32'b11111111111111110011110011110110;
assign LUT_2[26445] = 32'b11111111111111110000101100001111;
assign LUT_2[26446] = 32'b11111111111111111010101100110010;
assign LUT_2[26447] = 32'b11111111111111110111100101001011;
assign LUT_2[26448] = 32'b11111111111111110111001000111011;
assign LUT_2[26449] = 32'b11111111111111110100000001010100;
assign LUT_2[26450] = 32'b11111111111111111110000001110111;
assign LUT_2[26451] = 32'b11111111111111111010111010010000;
assign LUT_2[26452] = 32'b11111111111111110011100110100011;
assign LUT_2[26453] = 32'b11111111111111110000011110111100;
assign LUT_2[26454] = 32'b11111111111111111010011111011111;
assign LUT_2[26455] = 32'b11111111111111110111010111111000;
assign LUT_2[26456] = 32'b11111111111111110001111010011000;
assign LUT_2[26457] = 32'b11111111111111101110110010110001;
assign LUT_2[26458] = 32'b11111111111111111000110011010100;
assign LUT_2[26459] = 32'b11111111111111110101101011101101;
assign LUT_2[26460] = 32'b11111111111111101110011000000000;
assign LUT_2[26461] = 32'b11111111111111101011010000011001;
assign LUT_2[26462] = 32'b11111111111111110101010000111100;
assign LUT_2[26463] = 32'b11111111111111110010001001010101;
assign LUT_2[26464] = 32'b11111111111111111101000000011010;
assign LUT_2[26465] = 32'b11111111111111111001111000110011;
assign LUT_2[26466] = 32'b00000000000000000011111001010110;
assign LUT_2[26467] = 32'b00000000000000000000110001101111;
assign LUT_2[26468] = 32'b11111111111111111001011110000010;
assign LUT_2[26469] = 32'b11111111111111110110010110011011;
assign LUT_2[26470] = 32'b00000000000000000000010110111110;
assign LUT_2[26471] = 32'b11111111111111111101001111010111;
assign LUT_2[26472] = 32'b11111111111111110111110001110111;
assign LUT_2[26473] = 32'b11111111111111110100101010010000;
assign LUT_2[26474] = 32'b11111111111111111110101010110011;
assign LUT_2[26475] = 32'b11111111111111111011100011001100;
assign LUT_2[26476] = 32'b11111111111111110100001111011111;
assign LUT_2[26477] = 32'b11111111111111110001000111111000;
assign LUT_2[26478] = 32'b11111111111111111011001000011011;
assign LUT_2[26479] = 32'b11111111111111111000000000110100;
assign LUT_2[26480] = 32'b11111111111111110111100100100100;
assign LUT_2[26481] = 32'b11111111111111110100011100111101;
assign LUT_2[26482] = 32'b11111111111111111110011101100000;
assign LUT_2[26483] = 32'b11111111111111111011010101111001;
assign LUT_2[26484] = 32'b11111111111111110100000010001100;
assign LUT_2[26485] = 32'b11111111111111110000111010100101;
assign LUT_2[26486] = 32'b11111111111111111010111011001000;
assign LUT_2[26487] = 32'b11111111111111110111110011100001;
assign LUT_2[26488] = 32'b11111111111111110010010110000001;
assign LUT_2[26489] = 32'b11111111111111101111001110011010;
assign LUT_2[26490] = 32'b11111111111111111001001110111101;
assign LUT_2[26491] = 32'b11111111111111110110000111010110;
assign LUT_2[26492] = 32'b11111111111111101110110011101001;
assign LUT_2[26493] = 32'b11111111111111101011101100000010;
assign LUT_2[26494] = 32'b11111111111111110101101100100101;
assign LUT_2[26495] = 32'b11111111111111110010100100111110;
assign LUT_2[26496] = 32'b00000000000000001000110000011101;
assign LUT_2[26497] = 32'b00000000000000000101101000110110;
assign LUT_2[26498] = 32'b00000000000000001111101001011001;
assign LUT_2[26499] = 32'b00000000000000001100100001110010;
assign LUT_2[26500] = 32'b00000000000000000101001110000101;
assign LUT_2[26501] = 32'b00000000000000000010000110011110;
assign LUT_2[26502] = 32'b00000000000000001100000111000001;
assign LUT_2[26503] = 32'b00000000000000001000111111011010;
assign LUT_2[26504] = 32'b00000000000000000011100001111010;
assign LUT_2[26505] = 32'b00000000000000000000011010010011;
assign LUT_2[26506] = 32'b00000000000000001010011010110110;
assign LUT_2[26507] = 32'b00000000000000000111010011001111;
assign LUT_2[26508] = 32'b11111111111111111111111111100010;
assign LUT_2[26509] = 32'b11111111111111111100110111111011;
assign LUT_2[26510] = 32'b00000000000000000110111000011110;
assign LUT_2[26511] = 32'b00000000000000000011110000110111;
assign LUT_2[26512] = 32'b00000000000000000011010100100111;
assign LUT_2[26513] = 32'b00000000000000000000001101000000;
assign LUT_2[26514] = 32'b00000000000000001010001101100011;
assign LUT_2[26515] = 32'b00000000000000000111000101111100;
assign LUT_2[26516] = 32'b11111111111111111111110010001111;
assign LUT_2[26517] = 32'b11111111111111111100101010101000;
assign LUT_2[26518] = 32'b00000000000000000110101011001011;
assign LUT_2[26519] = 32'b00000000000000000011100011100100;
assign LUT_2[26520] = 32'b11111111111111111110000110000100;
assign LUT_2[26521] = 32'b11111111111111111010111110011101;
assign LUT_2[26522] = 32'b00000000000000000100111111000000;
assign LUT_2[26523] = 32'b00000000000000000001110111011001;
assign LUT_2[26524] = 32'b11111111111111111010100011101100;
assign LUT_2[26525] = 32'b11111111111111110111011100000101;
assign LUT_2[26526] = 32'b00000000000000000001011100101000;
assign LUT_2[26527] = 32'b11111111111111111110010101000001;
assign LUT_2[26528] = 32'b00000000000000001001001100000110;
assign LUT_2[26529] = 32'b00000000000000000110000100011111;
assign LUT_2[26530] = 32'b00000000000000010000000101000010;
assign LUT_2[26531] = 32'b00000000000000001100111101011011;
assign LUT_2[26532] = 32'b00000000000000000101101001101110;
assign LUT_2[26533] = 32'b00000000000000000010100010000111;
assign LUT_2[26534] = 32'b00000000000000001100100010101010;
assign LUT_2[26535] = 32'b00000000000000001001011011000011;
assign LUT_2[26536] = 32'b00000000000000000011111101100011;
assign LUT_2[26537] = 32'b00000000000000000000110101111100;
assign LUT_2[26538] = 32'b00000000000000001010110110011111;
assign LUT_2[26539] = 32'b00000000000000000111101110111000;
assign LUT_2[26540] = 32'b00000000000000000000011011001011;
assign LUT_2[26541] = 32'b11111111111111111101010011100100;
assign LUT_2[26542] = 32'b00000000000000000111010100000111;
assign LUT_2[26543] = 32'b00000000000000000100001100100000;
assign LUT_2[26544] = 32'b00000000000000000011110000010000;
assign LUT_2[26545] = 32'b00000000000000000000101000101001;
assign LUT_2[26546] = 32'b00000000000000001010101001001100;
assign LUT_2[26547] = 32'b00000000000000000111100001100101;
assign LUT_2[26548] = 32'b00000000000000000000001101111000;
assign LUT_2[26549] = 32'b11111111111111111101000110010001;
assign LUT_2[26550] = 32'b00000000000000000111000110110100;
assign LUT_2[26551] = 32'b00000000000000000011111111001101;
assign LUT_2[26552] = 32'b11111111111111111110100001101101;
assign LUT_2[26553] = 32'b11111111111111111011011010000110;
assign LUT_2[26554] = 32'b00000000000000000101011010101001;
assign LUT_2[26555] = 32'b00000000000000000010010011000010;
assign LUT_2[26556] = 32'b11111111111111111010111111010101;
assign LUT_2[26557] = 32'b11111111111111110111110111101110;
assign LUT_2[26558] = 32'b00000000000000000001111000010001;
assign LUT_2[26559] = 32'b11111111111111111110110000101010;
assign LUT_2[26560] = 32'b00000000000000000000111001000000;
assign LUT_2[26561] = 32'b11111111111111111101110001011001;
assign LUT_2[26562] = 32'b00000000000000000111110001111100;
assign LUT_2[26563] = 32'b00000000000000000100101010010101;
assign LUT_2[26564] = 32'b11111111111111111101010110101000;
assign LUT_2[26565] = 32'b11111111111111111010001111000001;
assign LUT_2[26566] = 32'b00000000000000000100001111100100;
assign LUT_2[26567] = 32'b00000000000000000001000111111101;
assign LUT_2[26568] = 32'b11111111111111111011101010011101;
assign LUT_2[26569] = 32'b11111111111111111000100010110110;
assign LUT_2[26570] = 32'b00000000000000000010100011011001;
assign LUT_2[26571] = 32'b11111111111111111111011011110010;
assign LUT_2[26572] = 32'b11111111111111111000001000000101;
assign LUT_2[26573] = 32'b11111111111111110101000000011110;
assign LUT_2[26574] = 32'b11111111111111111111000001000001;
assign LUT_2[26575] = 32'b11111111111111111011111001011010;
assign LUT_2[26576] = 32'b11111111111111111011011101001010;
assign LUT_2[26577] = 32'b11111111111111111000010101100011;
assign LUT_2[26578] = 32'b00000000000000000010010110000110;
assign LUT_2[26579] = 32'b11111111111111111111001110011111;
assign LUT_2[26580] = 32'b11111111111111110111111010110010;
assign LUT_2[26581] = 32'b11111111111111110100110011001011;
assign LUT_2[26582] = 32'b11111111111111111110110011101110;
assign LUT_2[26583] = 32'b11111111111111111011101100000111;
assign LUT_2[26584] = 32'b11111111111111110110001110100111;
assign LUT_2[26585] = 32'b11111111111111110011000111000000;
assign LUT_2[26586] = 32'b11111111111111111101000111100011;
assign LUT_2[26587] = 32'b11111111111111111001111111111100;
assign LUT_2[26588] = 32'b11111111111111110010101100001111;
assign LUT_2[26589] = 32'b11111111111111101111100100101000;
assign LUT_2[26590] = 32'b11111111111111111001100101001011;
assign LUT_2[26591] = 32'b11111111111111110110011101100100;
assign LUT_2[26592] = 32'b00000000000000000001010100101001;
assign LUT_2[26593] = 32'b11111111111111111110001101000010;
assign LUT_2[26594] = 32'b00000000000000001000001101100101;
assign LUT_2[26595] = 32'b00000000000000000101000101111110;
assign LUT_2[26596] = 32'b11111111111111111101110010010001;
assign LUT_2[26597] = 32'b11111111111111111010101010101010;
assign LUT_2[26598] = 32'b00000000000000000100101011001101;
assign LUT_2[26599] = 32'b00000000000000000001100011100110;
assign LUT_2[26600] = 32'b11111111111111111100000110000110;
assign LUT_2[26601] = 32'b11111111111111111000111110011111;
assign LUT_2[26602] = 32'b00000000000000000010111111000010;
assign LUT_2[26603] = 32'b11111111111111111111110111011011;
assign LUT_2[26604] = 32'b11111111111111111000100011101110;
assign LUT_2[26605] = 32'b11111111111111110101011100000111;
assign LUT_2[26606] = 32'b11111111111111111111011100101010;
assign LUT_2[26607] = 32'b11111111111111111100010101000011;
assign LUT_2[26608] = 32'b11111111111111111011111000110011;
assign LUT_2[26609] = 32'b11111111111111111000110001001100;
assign LUT_2[26610] = 32'b00000000000000000010110001101111;
assign LUT_2[26611] = 32'b11111111111111111111101010001000;
assign LUT_2[26612] = 32'b11111111111111111000010110011011;
assign LUT_2[26613] = 32'b11111111111111110101001110110100;
assign LUT_2[26614] = 32'b11111111111111111111001111010111;
assign LUT_2[26615] = 32'b11111111111111111100000111110000;
assign LUT_2[26616] = 32'b11111111111111110110101010010000;
assign LUT_2[26617] = 32'b11111111111111110011100010101001;
assign LUT_2[26618] = 32'b11111111111111111101100011001100;
assign LUT_2[26619] = 32'b11111111111111111010011011100101;
assign LUT_2[26620] = 32'b11111111111111110011000111111000;
assign LUT_2[26621] = 32'b11111111111111110000000000010001;
assign LUT_2[26622] = 32'b11111111111111111010000000110100;
assign LUT_2[26623] = 32'b11111111111111110110111001001101;
assign LUT_2[26624] = 32'b11111111111111110000110101101101;
assign LUT_2[26625] = 32'b11111111111111101101101110000110;
assign LUT_2[26626] = 32'b11111111111111110111101110101001;
assign LUT_2[26627] = 32'b11111111111111110100100111000010;
assign LUT_2[26628] = 32'b11111111111111101101010011010101;
assign LUT_2[26629] = 32'b11111111111111101010001011101110;
assign LUT_2[26630] = 32'b11111111111111110100001100010001;
assign LUT_2[26631] = 32'b11111111111111110001000100101010;
assign LUT_2[26632] = 32'b11111111111111101011100111001010;
assign LUT_2[26633] = 32'b11111111111111101000011111100011;
assign LUT_2[26634] = 32'b11111111111111110010100000000110;
assign LUT_2[26635] = 32'b11111111111111101111011000011111;
assign LUT_2[26636] = 32'b11111111111111101000000100110010;
assign LUT_2[26637] = 32'b11111111111111100100111101001011;
assign LUT_2[26638] = 32'b11111111111111101110111101101110;
assign LUT_2[26639] = 32'b11111111111111101011110110000111;
assign LUT_2[26640] = 32'b11111111111111101011011001110111;
assign LUT_2[26641] = 32'b11111111111111101000010010010000;
assign LUT_2[26642] = 32'b11111111111111110010010010110011;
assign LUT_2[26643] = 32'b11111111111111101111001011001100;
assign LUT_2[26644] = 32'b11111111111111100111110111011111;
assign LUT_2[26645] = 32'b11111111111111100100101111111000;
assign LUT_2[26646] = 32'b11111111111111101110110000011011;
assign LUT_2[26647] = 32'b11111111111111101011101000110100;
assign LUT_2[26648] = 32'b11111111111111100110001011010100;
assign LUT_2[26649] = 32'b11111111111111100011000011101101;
assign LUT_2[26650] = 32'b11111111111111101101000100010000;
assign LUT_2[26651] = 32'b11111111111111101001111100101001;
assign LUT_2[26652] = 32'b11111111111111100010101000111100;
assign LUT_2[26653] = 32'b11111111111111011111100001010101;
assign LUT_2[26654] = 32'b11111111111111101001100001111000;
assign LUT_2[26655] = 32'b11111111111111100110011010010001;
assign LUT_2[26656] = 32'b11111111111111110001010001010110;
assign LUT_2[26657] = 32'b11111111111111101110001001101111;
assign LUT_2[26658] = 32'b11111111111111111000001010010010;
assign LUT_2[26659] = 32'b11111111111111110101000010101011;
assign LUT_2[26660] = 32'b11111111111111101101101110111110;
assign LUT_2[26661] = 32'b11111111111111101010100111010111;
assign LUT_2[26662] = 32'b11111111111111110100100111111010;
assign LUT_2[26663] = 32'b11111111111111110001100000010011;
assign LUT_2[26664] = 32'b11111111111111101100000010110011;
assign LUT_2[26665] = 32'b11111111111111101000111011001100;
assign LUT_2[26666] = 32'b11111111111111110010111011101111;
assign LUT_2[26667] = 32'b11111111111111101111110100001000;
assign LUT_2[26668] = 32'b11111111111111101000100000011011;
assign LUT_2[26669] = 32'b11111111111111100101011000110100;
assign LUT_2[26670] = 32'b11111111111111101111011001010111;
assign LUT_2[26671] = 32'b11111111111111101100010001110000;
assign LUT_2[26672] = 32'b11111111111111101011110101100000;
assign LUT_2[26673] = 32'b11111111111111101000101101111001;
assign LUT_2[26674] = 32'b11111111111111110010101110011100;
assign LUT_2[26675] = 32'b11111111111111101111100110110101;
assign LUT_2[26676] = 32'b11111111111111101000010011001000;
assign LUT_2[26677] = 32'b11111111111111100101001011100001;
assign LUT_2[26678] = 32'b11111111111111101111001100000100;
assign LUT_2[26679] = 32'b11111111111111101100000100011101;
assign LUT_2[26680] = 32'b11111111111111100110100110111101;
assign LUT_2[26681] = 32'b11111111111111100011011111010110;
assign LUT_2[26682] = 32'b11111111111111101101011111111001;
assign LUT_2[26683] = 32'b11111111111111101010011000010010;
assign LUT_2[26684] = 32'b11111111111111100011000100100101;
assign LUT_2[26685] = 32'b11111111111111011111111100111110;
assign LUT_2[26686] = 32'b11111111111111101001111101100001;
assign LUT_2[26687] = 32'b11111111111111100110110101111010;
assign LUT_2[26688] = 32'b11111111111111101000111110010000;
assign LUT_2[26689] = 32'b11111111111111100101110110101001;
assign LUT_2[26690] = 32'b11111111111111101111110111001100;
assign LUT_2[26691] = 32'b11111111111111101100101111100101;
assign LUT_2[26692] = 32'b11111111111111100101011011111000;
assign LUT_2[26693] = 32'b11111111111111100010010100010001;
assign LUT_2[26694] = 32'b11111111111111101100010100110100;
assign LUT_2[26695] = 32'b11111111111111101001001101001101;
assign LUT_2[26696] = 32'b11111111111111100011101111101101;
assign LUT_2[26697] = 32'b11111111111111100000101000000110;
assign LUT_2[26698] = 32'b11111111111111101010101000101001;
assign LUT_2[26699] = 32'b11111111111111100111100001000010;
assign LUT_2[26700] = 32'b11111111111111100000001101010101;
assign LUT_2[26701] = 32'b11111111111111011101000101101110;
assign LUT_2[26702] = 32'b11111111111111100111000110010001;
assign LUT_2[26703] = 32'b11111111111111100011111110101010;
assign LUT_2[26704] = 32'b11111111111111100011100010011010;
assign LUT_2[26705] = 32'b11111111111111100000011010110011;
assign LUT_2[26706] = 32'b11111111111111101010011011010110;
assign LUT_2[26707] = 32'b11111111111111100111010011101111;
assign LUT_2[26708] = 32'b11111111111111100000000000000010;
assign LUT_2[26709] = 32'b11111111111111011100111000011011;
assign LUT_2[26710] = 32'b11111111111111100110111000111110;
assign LUT_2[26711] = 32'b11111111111111100011110001010111;
assign LUT_2[26712] = 32'b11111111111111011110010011110111;
assign LUT_2[26713] = 32'b11111111111111011011001100010000;
assign LUT_2[26714] = 32'b11111111111111100101001100110011;
assign LUT_2[26715] = 32'b11111111111111100010000101001100;
assign LUT_2[26716] = 32'b11111111111111011010110001011111;
assign LUT_2[26717] = 32'b11111111111111010111101001111000;
assign LUT_2[26718] = 32'b11111111111111100001101010011011;
assign LUT_2[26719] = 32'b11111111111111011110100010110100;
assign LUT_2[26720] = 32'b11111111111111101001011001111001;
assign LUT_2[26721] = 32'b11111111111111100110010010010010;
assign LUT_2[26722] = 32'b11111111111111110000010010110101;
assign LUT_2[26723] = 32'b11111111111111101101001011001110;
assign LUT_2[26724] = 32'b11111111111111100101110111100001;
assign LUT_2[26725] = 32'b11111111111111100010101111111010;
assign LUT_2[26726] = 32'b11111111111111101100110000011101;
assign LUT_2[26727] = 32'b11111111111111101001101000110110;
assign LUT_2[26728] = 32'b11111111111111100100001011010110;
assign LUT_2[26729] = 32'b11111111111111100001000011101111;
assign LUT_2[26730] = 32'b11111111111111101011000100010010;
assign LUT_2[26731] = 32'b11111111111111100111111100101011;
assign LUT_2[26732] = 32'b11111111111111100000101000111110;
assign LUT_2[26733] = 32'b11111111111111011101100001010111;
assign LUT_2[26734] = 32'b11111111111111100111100001111010;
assign LUT_2[26735] = 32'b11111111111111100100011010010011;
assign LUT_2[26736] = 32'b11111111111111100011111110000011;
assign LUT_2[26737] = 32'b11111111111111100000110110011100;
assign LUT_2[26738] = 32'b11111111111111101010110110111111;
assign LUT_2[26739] = 32'b11111111111111100111101111011000;
assign LUT_2[26740] = 32'b11111111111111100000011011101011;
assign LUT_2[26741] = 32'b11111111111111011101010100000100;
assign LUT_2[26742] = 32'b11111111111111100111010100100111;
assign LUT_2[26743] = 32'b11111111111111100100001101000000;
assign LUT_2[26744] = 32'b11111111111111011110101111100000;
assign LUT_2[26745] = 32'b11111111111111011011100111111001;
assign LUT_2[26746] = 32'b11111111111111100101101000011100;
assign LUT_2[26747] = 32'b11111111111111100010100000110101;
assign LUT_2[26748] = 32'b11111111111111011011001101001000;
assign LUT_2[26749] = 32'b11111111111111011000000101100001;
assign LUT_2[26750] = 32'b11111111111111100010000110000100;
assign LUT_2[26751] = 32'b11111111111111011110111110011101;
assign LUT_2[26752] = 32'b11111111111111110101001001111100;
assign LUT_2[26753] = 32'b11111111111111110010000010010101;
assign LUT_2[26754] = 32'b11111111111111111100000010111000;
assign LUT_2[26755] = 32'b11111111111111111000111011010001;
assign LUT_2[26756] = 32'b11111111111111110001100111100100;
assign LUT_2[26757] = 32'b11111111111111101110011111111101;
assign LUT_2[26758] = 32'b11111111111111111000100000100000;
assign LUT_2[26759] = 32'b11111111111111110101011000111001;
assign LUT_2[26760] = 32'b11111111111111101111111011011001;
assign LUT_2[26761] = 32'b11111111111111101100110011110010;
assign LUT_2[26762] = 32'b11111111111111110110110100010101;
assign LUT_2[26763] = 32'b11111111111111110011101100101110;
assign LUT_2[26764] = 32'b11111111111111101100011001000001;
assign LUT_2[26765] = 32'b11111111111111101001010001011010;
assign LUT_2[26766] = 32'b11111111111111110011010001111101;
assign LUT_2[26767] = 32'b11111111111111110000001010010110;
assign LUT_2[26768] = 32'b11111111111111101111101110000110;
assign LUT_2[26769] = 32'b11111111111111101100100110011111;
assign LUT_2[26770] = 32'b11111111111111110110100111000010;
assign LUT_2[26771] = 32'b11111111111111110011011111011011;
assign LUT_2[26772] = 32'b11111111111111101100001011101110;
assign LUT_2[26773] = 32'b11111111111111101001000100000111;
assign LUT_2[26774] = 32'b11111111111111110011000100101010;
assign LUT_2[26775] = 32'b11111111111111101111111101000011;
assign LUT_2[26776] = 32'b11111111111111101010011111100011;
assign LUT_2[26777] = 32'b11111111111111100111010111111100;
assign LUT_2[26778] = 32'b11111111111111110001011000011111;
assign LUT_2[26779] = 32'b11111111111111101110010000111000;
assign LUT_2[26780] = 32'b11111111111111100110111101001011;
assign LUT_2[26781] = 32'b11111111111111100011110101100100;
assign LUT_2[26782] = 32'b11111111111111101101110110000111;
assign LUT_2[26783] = 32'b11111111111111101010101110100000;
assign LUT_2[26784] = 32'b11111111111111110101100101100101;
assign LUT_2[26785] = 32'b11111111111111110010011101111110;
assign LUT_2[26786] = 32'b11111111111111111100011110100001;
assign LUT_2[26787] = 32'b11111111111111111001010110111010;
assign LUT_2[26788] = 32'b11111111111111110010000011001101;
assign LUT_2[26789] = 32'b11111111111111101110111011100110;
assign LUT_2[26790] = 32'b11111111111111111000111100001001;
assign LUT_2[26791] = 32'b11111111111111110101110100100010;
assign LUT_2[26792] = 32'b11111111111111110000010111000010;
assign LUT_2[26793] = 32'b11111111111111101101001111011011;
assign LUT_2[26794] = 32'b11111111111111110111001111111110;
assign LUT_2[26795] = 32'b11111111111111110100001000010111;
assign LUT_2[26796] = 32'b11111111111111101100110100101010;
assign LUT_2[26797] = 32'b11111111111111101001101101000011;
assign LUT_2[26798] = 32'b11111111111111110011101101100110;
assign LUT_2[26799] = 32'b11111111111111110000100101111111;
assign LUT_2[26800] = 32'b11111111111111110000001001101111;
assign LUT_2[26801] = 32'b11111111111111101101000010001000;
assign LUT_2[26802] = 32'b11111111111111110111000010101011;
assign LUT_2[26803] = 32'b11111111111111110011111011000100;
assign LUT_2[26804] = 32'b11111111111111101100100111010111;
assign LUT_2[26805] = 32'b11111111111111101001011111110000;
assign LUT_2[26806] = 32'b11111111111111110011100000010011;
assign LUT_2[26807] = 32'b11111111111111110000011000101100;
assign LUT_2[26808] = 32'b11111111111111101010111011001100;
assign LUT_2[26809] = 32'b11111111111111100111110011100101;
assign LUT_2[26810] = 32'b11111111111111110001110100001000;
assign LUT_2[26811] = 32'b11111111111111101110101100100001;
assign LUT_2[26812] = 32'b11111111111111100111011000110100;
assign LUT_2[26813] = 32'b11111111111111100100010001001101;
assign LUT_2[26814] = 32'b11111111111111101110010001110000;
assign LUT_2[26815] = 32'b11111111111111101011001010001001;
assign LUT_2[26816] = 32'b11111111111111101101010010011111;
assign LUT_2[26817] = 32'b11111111111111101010001010111000;
assign LUT_2[26818] = 32'b11111111111111110100001011011011;
assign LUT_2[26819] = 32'b11111111111111110001000011110100;
assign LUT_2[26820] = 32'b11111111111111101001110000000111;
assign LUT_2[26821] = 32'b11111111111111100110101000100000;
assign LUT_2[26822] = 32'b11111111111111110000101001000011;
assign LUT_2[26823] = 32'b11111111111111101101100001011100;
assign LUT_2[26824] = 32'b11111111111111101000000011111100;
assign LUT_2[26825] = 32'b11111111111111100100111100010101;
assign LUT_2[26826] = 32'b11111111111111101110111100111000;
assign LUT_2[26827] = 32'b11111111111111101011110101010001;
assign LUT_2[26828] = 32'b11111111111111100100100001100100;
assign LUT_2[26829] = 32'b11111111111111100001011001111101;
assign LUT_2[26830] = 32'b11111111111111101011011010100000;
assign LUT_2[26831] = 32'b11111111111111101000010010111001;
assign LUT_2[26832] = 32'b11111111111111100111110110101001;
assign LUT_2[26833] = 32'b11111111111111100100101111000010;
assign LUT_2[26834] = 32'b11111111111111101110101111100101;
assign LUT_2[26835] = 32'b11111111111111101011100111111110;
assign LUT_2[26836] = 32'b11111111111111100100010100010001;
assign LUT_2[26837] = 32'b11111111111111100001001100101010;
assign LUT_2[26838] = 32'b11111111111111101011001101001101;
assign LUT_2[26839] = 32'b11111111111111101000000101100110;
assign LUT_2[26840] = 32'b11111111111111100010101000000110;
assign LUT_2[26841] = 32'b11111111111111011111100000011111;
assign LUT_2[26842] = 32'b11111111111111101001100001000010;
assign LUT_2[26843] = 32'b11111111111111100110011001011011;
assign LUT_2[26844] = 32'b11111111111111011111000101101110;
assign LUT_2[26845] = 32'b11111111111111011011111110000111;
assign LUT_2[26846] = 32'b11111111111111100101111110101010;
assign LUT_2[26847] = 32'b11111111111111100010110111000011;
assign LUT_2[26848] = 32'b11111111111111101101101110001000;
assign LUT_2[26849] = 32'b11111111111111101010100110100001;
assign LUT_2[26850] = 32'b11111111111111110100100111000100;
assign LUT_2[26851] = 32'b11111111111111110001011111011101;
assign LUT_2[26852] = 32'b11111111111111101010001011110000;
assign LUT_2[26853] = 32'b11111111111111100111000100001001;
assign LUT_2[26854] = 32'b11111111111111110001000100101100;
assign LUT_2[26855] = 32'b11111111111111101101111101000101;
assign LUT_2[26856] = 32'b11111111111111101000011111100101;
assign LUT_2[26857] = 32'b11111111111111100101010111111110;
assign LUT_2[26858] = 32'b11111111111111101111011000100001;
assign LUT_2[26859] = 32'b11111111111111101100010000111010;
assign LUT_2[26860] = 32'b11111111111111100100111101001101;
assign LUT_2[26861] = 32'b11111111111111100001110101100110;
assign LUT_2[26862] = 32'b11111111111111101011110110001001;
assign LUT_2[26863] = 32'b11111111111111101000101110100010;
assign LUT_2[26864] = 32'b11111111111111101000010010010010;
assign LUT_2[26865] = 32'b11111111111111100101001010101011;
assign LUT_2[26866] = 32'b11111111111111101111001011001110;
assign LUT_2[26867] = 32'b11111111111111101100000011100111;
assign LUT_2[26868] = 32'b11111111111111100100101111111010;
assign LUT_2[26869] = 32'b11111111111111100001101000010011;
assign LUT_2[26870] = 32'b11111111111111101011101000110110;
assign LUT_2[26871] = 32'b11111111111111101000100001001111;
assign LUT_2[26872] = 32'b11111111111111100011000011101111;
assign LUT_2[26873] = 32'b11111111111111011111111100001000;
assign LUT_2[26874] = 32'b11111111111111101001111100101011;
assign LUT_2[26875] = 32'b11111111111111100110110101000100;
assign LUT_2[26876] = 32'b11111111111111011111100001010111;
assign LUT_2[26877] = 32'b11111111111111011100011001110000;
assign LUT_2[26878] = 32'b11111111111111100110011010010011;
assign LUT_2[26879] = 32'b11111111111111100011010010101100;
assign LUT_2[26880] = 32'b11111111111111110100110100010011;
assign LUT_2[26881] = 32'b11111111111111110001101100101100;
assign LUT_2[26882] = 32'b11111111111111111011101101001111;
assign LUT_2[26883] = 32'b11111111111111111000100101101000;
assign LUT_2[26884] = 32'b11111111111111110001010001111011;
assign LUT_2[26885] = 32'b11111111111111101110001010010100;
assign LUT_2[26886] = 32'b11111111111111111000001010110111;
assign LUT_2[26887] = 32'b11111111111111110101000011010000;
assign LUT_2[26888] = 32'b11111111111111101111100101110000;
assign LUT_2[26889] = 32'b11111111111111101100011110001001;
assign LUT_2[26890] = 32'b11111111111111110110011110101100;
assign LUT_2[26891] = 32'b11111111111111110011010111000101;
assign LUT_2[26892] = 32'b11111111111111101100000011011000;
assign LUT_2[26893] = 32'b11111111111111101000111011110001;
assign LUT_2[26894] = 32'b11111111111111110010111100010100;
assign LUT_2[26895] = 32'b11111111111111101111110100101101;
assign LUT_2[26896] = 32'b11111111111111101111011000011101;
assign LUT_2[26897] = 32'b11111111111111101100010000110110;
assign LUT_2[26898] = 32'b11111111111111110110010001011001;
assign LUT_2[26899] = 32'b11111111111111110011001001110010;
assign LUT_2[26900] = 32'b11111111111111101011110110000101;
assign LUT_2[26901] = 32'b11111111111111101000101110011110;
assign LUT_2[26902] = 32'b11111111111111110010101111000001;
assign LUT_2[26903] = 32'b11111111111111101111100111011010;
assign LUT_2[26904] = 32'b11111111111111101010001001111010;
assign LUT_2[26905] = 32'b11111111111111100111000010010011;
assign LUT_2[26906] = 32'b11111111111111110001000010110110;
assign LUT_2[26907] = 32'b11111111111111101101111011001111;
assign LUT_2[26908] = 32'b11111111111111100110100111100010;
assign LUT_2[26909] = 32'b11111111111111100011011111111011;
assign LUT_2[26910] = 32'b11111111111111101101100000011110;
assign LUT_2[26911] = 32'b11111111111111101010011000110111;
assign LUT_2[26912] = 32'b11111111111111110101001111111100;
assign LUT_2[26913] = 32'b11111111111111110010001000010101;
assign LUT_2[26914] = 32'b11111111111111111100001000111000;
assign LUT_2[26915] = 32'b11111111111111111001000001010001;
assign LUT_2[26916] = 32'b11111111111111110001101101100100;
assign LUT_2[26917] = 32'b11111111111111101110100101111101;
assign LUT_2[26918] = 32'b11111111111111111000100110100000;
assign LUT_2[26919] = 32'b11111111111111110101011110111001;
assign LUT_2[26920] = 32'b11111111111111110000000001011001;
assign LUT_2[26921] = 32'b11111111111111101100111001110010;
assign LUT_2[26922] = 32'b11111111111111110110111010010101;
assign LUT_2[26923] = 32'b11111111111111110011110010101110;
assign LUT_2[26924] = 32'b11111111111111101100011111000001;
assign LUT_2[26925] = 32'b11111111111111101001010111011010;
assign LUT_2[26926] = 32'b11111111111111110011010111111101;
assign LUT_2[26927] = 32'b11111111111111110000010000010110;
assign LUT_2[26928] = 32'b11111111111111101111110100000110;
assign LUT_2[26929] = 32'b11111111111111101100101100011111;
assign LUT_2[26930] = 32'b11111111111111110110101101000010;
assign LUT_2[26931] = 32'b11111111111111110011100101011011;
assign LUT_2[26932] = 32'b11111111111111101100010001101110;
assign LUT_2[26933] = 32'b11111111111111101001001010000111;
assign LUT_2[26934] = 32'b11111111111111110011001010101010;
assign LUT_2[26935] = 32'b11111111111111110000000011000011;
assign LUT_2[26936] = 32'b11111111111111101010100101100011;
assign LUT_2[26937] = 32'b11111111111111100111011101111100;
assign LUT_2[26938] = 32'b11111111111111110001011110011111;
assign LUT_2[26939] = 32'b11111111111111101110010110111000;
assign LUT_2[26940] = 32'b11111111111111100111000011001011;
assign LUT_2[26941] = 32'b11111111111111100011111011100100;
assign LUT_2[26942] = 32'b11111111111111101101111100000111;
assign LUT_2[26943] = 32'b11111111111111101010110100100000;
assign LUT_2[26944] = 32'b11111111111111101100111100110110;
assign LUT_2[26945] = 32'b11111111111111101001110101001111;
assign LUT_2[26946] = 32'b11111111111111110011110101110010;
assign LUT_2[26947] = 32'b11111111111111110000101110001011;
assign LUT_2[26948] = 32'b11111111111111101001011010011110;
assign LUT_2[26949] = 32'b11111111111111100110010010110111;
assign LUT_2[26950] = 32'b11111111111111110000010011011010;
assign LUT_2[26951] = 32'b11111111111111101101001011110011;
assign LUT_2[26952] = 32'b11111111111111100111101110010011;
assign LUT_2[26953] = 32'b11111111111111100100100110101100;
assign LUT_2[26954] = 32'b11111111111111101110100111001111;
assign LUT_2[26955] = 32'b11111111111111101011011111101000;
assign LUT_2[26956] = 32'b11111111111111100100001011111011;
assign LUT_2[26957] = 32'b11111111111111100001000100010100;
assign LUT_2[26958] = 32'b11111111111111101011000100110111;
assign LUT_2[26959] = 32'b11111111111111100111111101010000;
assign LUT_2[26960] = 32'b11111111111111100111100001000000;
assign LUT_2[26961] = 32'b11111111111111100100011001011001;
assign LUT_2[26962] = 32'b11111111111111101110011001111100;
assign LUT_2[26963] = 32'b11111111111111101011010010010101;
assign LUT_2[26964] = 32'b11111111111111100011111110101000;
assign LUT_2[26965] = 32'b11111111111111100000110111000001;
assign LUT_2[26966] = 32'b11111111111111101010110111100100;
assign LUT_2[26967] = 32'b11111111111111100111101111111101;
assign LUT_2[26968] = 32'b11111111111111100010010010011101;
assign LUT_2[26969] = 32'b11111111111111011111001010110110;
assign LUT_2[26970] = 32'b11111111111111101001001011011001;
assign LUT_2[26971] = 32'b11111111111111100110000011110010;
assign LUT_2[26972] = 32'b11111111111111011110110000000101;
assign LUT_2[26973] = 32'b11111111111111011011101000011110;
assign LUT_2[26974] = 32'b11111111111111100101101001000001;
assign LUT_2[26975] = 32'b11111111111111100010100001011010;
assign LUT_2[26976] = 32'b11111111111111101101011000011111;
assign LUT_2[26977] = 32'b11111111111111101010010000111000;
assign LUT_2[26978] = 32'b11111111111111110100010001011011;
assign LUT_2[26979] = 32'b11111111111111110001001001110100;
assign LUT_2[26980] = 32'b11111111111111101001110110000111;
assign LUT_2[26981] = 32'b11111111111111100110101110100000;
assign LUT_2[26982] = 32'b11111111111111110000101111000011;
assign LUT_2[26983] = 32'b11111111111111101101100111011100;
assign LUT_2[26984] = 32'b11111111111111101000001001111100;
assign LUT_2[26985] = 32'b11111111111111100101000010010101;
assign LUT_2[26986] = 32'b11111111111111101111000010111000;
assign LUT_2[26987] = 32'b11111111111111101011111011010001;
assign LUT_2[26988] = 32'b11111111111111100100100111100100;
assign LUT_2[26989] = 32'b11111111111111100001011111111101;
assign LUT_2[26990] = 32'b11111111111111101011100000100000;
assign LUT_2[26991] = 32'b11111111111111101000011000111001;
assign LUT_2[26992] = 32'b11111111111111100111111100101001;
assign LUT_2[26993] = 32'b11111111111111100100110101000010;
assign LUT_2[26994] = 32'b11111111111111101110110101100101;
assign LUT_2[26995] = 32'b11111111111111101011101101111110;
assign LUT_2[26996] = 32'b11111111111111100100011010010001;
assign LUT_2[26997] = 32'b11111111111111100001010010101010;
assign LUT_2[26998] = 32'b11111111111111101011010011001101;
assign LUT_2[26999] = 32'b11111111111111101000001011100110;
assign LUT_2[27000] = 32'b11111111111111100010101110000110;
assign LUT_2[27001] = 32'b11111111111111011111100110011111;
assign LUT_2[27002] = 32'b11111111111111101001100111000010;
assign LUT_2[27003] = 32'b11111111111111100110011111011011;
assign LUT_2[27004] = 32'b11111111111111011111001011101110;
assign LUT_2[27005] = 32'b11111111111111011100000100000111;
assign LUT_2[27006] = 32'b11111111111111100110000100101010;
assign LUT_2[27007] = 32'b11111111111111100010111101000011;
assign LUT_2[27008] = 32'b11111111111111111001001000100010;
assign LUT_2[27009] = 32'b11111111111111110110000000111011;
assign LUT_2[27010] = 32'b00000000000000000000000001011110;
assign LUT_2[27011] = 32'b11111111111111111100111001110111;
assign LUT_2[27012] = 32'b11111111111111110101100110001010;
assign LUT_2[27013] = 32'b11111111111111110010011110100011;
assign LUT_2[27014] = 32'b11111111111111111100011111000110;
assign LUT_2[27015] = 32'b11111111111111111001010111011111;
assign LUT_2[27016] = 32'b11111111111111110011111001111111;
assign LUT_2[27017] = 32'b11111111111111110000110010011000;
assign LUT_2[27018] = 32'b11111111111111111010110010111011;
assign LUT_2[27019] = 32'b11111111111111110111101011010100;
assign LUT_2[27020] = 32'b11111111111111110000010111100111;
assign LUT_2[27021] = 32'b11111111111111101101010000000000;
assign LUT_2[27022] = 32'b11111111111111110111010000100011;
assign LUT_2[27023] = 32'b11111111111111110100001000111100;
assign LUT_2[27024] = 32'b11111111111111110011101100101100;
assign LUT_2[27025] = 32'b11111111111111110000100101000101;
assign LUT_2[27026] = 32'b11111111111111111010100101101000;
assign LUT_2[27027] = 32'b11111111111111110111011110000001;
assign LUT_2[27028] = 32'b11111111111111110000001010010100;
assign LUT_2[27029] = 32'b11111111111111101101000010101101;
assign LUT_2[27030] = 32'b11111111111111110111000011010000;
assign LUT_2[27031] = 32'b11111111111111110011111011101001;
assign LUT_2[27032] = 32'b11111111111111101110011110001001;
assign LUT_2[27033] = 32'b11111111111111101011010110100010;
assign LUT_2[27034] = 32'b11111111111111110101010111000101;
assign LUT_2[27035] = 32'b11111111111111110010001111011110;
assign LUT_2[27036] = 32'b11111111111111101010111011110001;
assign LUT_2[27037] = 32'b11111111111111100111110100001010;
assign LUT_2[27038] = 32'b11111111111111110001110100101101;
assign LUT_2[27039] = 32'b11111111111111101110101101000110;
assign LUT_2[27040] = 32'b11111111111111111001100100001011;
assign LUT_2[27041] = 32'b11111111111111110110011100100100;
assign LUT_2[27042] = 32'b00000000000000000000011101000111;
assign LUT_2[27043] = 32'b11111111111111111101010101100000;
assign LUT_2[27044] = 32'b11111111111111110110000001110011;
assign LUT_2[27045] = 32'b11111111111111110010111010001100;
assign LUT_2[27046] = 32'b11111111111111111100111010101111;
assign LUT_2[27047] = 32'b11111111111111111001110011001000;
assign LUT_2[27048] = 32'b11111111111111110100010101101000;
assign LUT_2[27049] = 32'b11111111111111110001001110000001;
assign LUT_2[27050] = 32'b11111111111111111011001110100100;
assign LUT_2[27051] = 32'b11111111111111111000000110111101;
assign LUT_2[27052] = 32'b11111111111111110000110011010000;
assign LUT_2[27053] = 32'b11111111111111101101101011101001;
assign LUT_2[27054] = 32'b11111111111111110111101100001100;
assign LUT_2[27055] = 32'b11111111111111110100100100100101;
assign LUT_2[27056] = 32'b11111111111111110100001000010101;
assign LUT_2[27057] = 32'b11111111111111110001000000101110;
assign LUT_2[27058] = 32'b11111111111111111011000001010001;
assign LUT_2[27059] = 32'b11111111111111110111111001101010;
assign LUT_2[27060] = 32'b11111111111111110000100101111101;
assign LUT_2[27061] = 32'b11111111111111101101011110010110;
assign LUT_2[27062] = 32'b11111111111111110111011110111001;
assign LUT_2[27063] = 32'b11111111111111110100010111010010;
assign LUT_2[27064] = 32'b11111111111111101110111001110010;
assign LUT_2[27065] = 32'b11111111111111101011110010001011;
assign LUT_2[27066] = 32'b11111111111111110101110010101110;
assign LUT_2[27067] = 32'b11111111111111110010101011000111;
assign LUT_2[27068] = 32'b11111111111111101011010111011010;
assign LUT_2[27069] = 32'b11111111111111101000001111110011;
assign LUT_2[27070] = 32'b11111111111111110010010000010110;
assign LUT_2[27071] = 32'b11111111111111101111001000101111;
assign LUT_2[27072] = 32'b11111111111111110001010001000101;
assign LUT_2[27073] = 32'b11111111111111101110001001011110;
assign LUT_2[27074] = 32'b11111111111111111000001010000001;
assign LUT_2[27075] = 32'b11111111111111110101000010011010;
assign LUT_2[27076] = 32'b11111111111111101101101110101101;
assign LUT_2[27077] = 32'b11111111111111101010100111000110;
assign LUT_2[27078] = 32'b11111111111111110100100111101001;
assign LUT_2[27079] = 32'b11111111111111110001100000000010;
assign LUT_2[27080] = 32'b11111111111111101100000010100010;
assign LUT_2[27081] = 32'b11111111111111101000111010111011;
assign LUT_2[27082] = 32'b11111111111111110010111011011110;
assign LUT_2[27083] = 32'b11111111111111101111110011110111;
assign LUT_2[27084] = 32'b11111111111111101000100000001010;
assign LUT_2[27085] = 32'b11111111111111100101011000100011;
assign LUT_2[27086] = 32'b11111111111111101111011001000110;
assign LUT_2[27087] = 32'b11111111111111101100010001011111;
assign LUT_2[27088] = 32'b11111111111111101011110101001111;
assign LUT_2[27089] = 32'b11111111111111101000101101101000;
assign LUT_2[27090] = 32'b11111111111111110010101110001011;
assign LUT_2[27091] = 32'b11111111111111101111100110100100;
assign LUT_2[27092] = 32'b11111111111111101000010010110111;
assign LUT_2[27093] = 32'b11111111111111100101001011010000;
assign LUT_2[27094] = 32'b11111111111111101111001011110011;
assign LUT_2[27095] = 32'b11111111111111101100000100001100;
assign LUT_2[27096] = 32'b11111111111111100110100110101100;
assign LUT_2[27097] = 32'b11111111111111100011011111000101;
assign LUT_2[27098] = 32'b11111111111111101101011111101000;
assign LUT_2[27099] = 32'b11111111111111101010011000000001;
assign LUT_2[27100] = 32'b11111111111111100011000100010100;
assign LUT_2[27101] = 32'b11111111111111011111111100101101;
assign LUT_2[27102] = 32'b11111111111111101001111101010000;
assign LUT_2[27103] = 32'b11111111111111100110110101101001;
assign LUT_2[27104] = 32'b11111111111111110001101100101110;
assign LUT_2[27105] = 32'b11111111111111101110100101000111;
assign LUT_2[27106] = 32'b11111111111111111000100101101010;
assign LUT_2[27107] = 32'b11111111111111110101011110000011;
assign LUT_2[27108] = 32'b11111111111111101110001010010110;
assign LUT_2[27109] = 32'b11111111111111101011000010101111;
assign LUT_2[27110] = 32'b11111111111111110101000011010010;
assign LUT_2[27111] = 32'b11111111111111110001111011101011;
assign LUT_2[27112] = 32'b11111111111111101100011110001011;
assign LUT_2[27113] = 32'b11111111111111101001010110100100;
assign LUT_2[27114] = 32'b11111111111111110011010111000111;
assign LUT_2[27115] = 32'b11111111111111110000001111100000;
assign LUT_2[27116] = 32'b11111111111111101000111011110011;
assign LUT_2[27117] = 32'b11111111111111100101110100001100;
assign LUT_2[27118] = 32'b11111111111111101111110100101111;
assign LUT_2[27119] = 32'b11111111111111101100101101001000;
assign LUT_2[27120] = 32'b11111111111111101100010000111000;
assign LUT_2[27121] = 32'b11111111111111101001001001010001;
assign LUT_2[27122] = 32'b11111111111111110011001001110100;
assign LUT_2[27123] = 32'b11111111111111110000000010001101;
assign LUT_2[27124] = 32'b11111111111111101000101110100000;
assign LUT_2[27125] = 32'b11111111111111100101100110111001;
assign LUT_2[27126] = 32'b11111111111111101111100111011100;
assign LUT_2[27127] = 32'b11111111111111101100011111110101;
assign LUT_2[27128] = 32'b11111111111111100111000010010101;
assign LUT_2[27129] = 32'b11111111111111100011111010101110;
assign LUT_2[27130] = 32'b11111111111111101101111011010001;
assign LUT_2[27131] = 32'b11111111111111101010110011101010;
assign LUT_2[27132] = 32'b11111111111111100011011111111101;
assign LUT_2[27133] = 32'b11111111111111100000011000010110;
assign LUT_2[27134] = 32'b11111111111111101010011000111001;
assign LUT_2[27135] = 32'b11111111111111100111010001010010;
assign LUT_2[27136] = 32'b11111111111111110101100111011111;
assign LUT_2[27137] = 32'b11111111111111110010011111111000;
assign LUT_2[27138] = 32'b11111111111111111100100000011011;
assign LUT_2[27139] = 32'b11111111111111111001011000110100;
assign LUT_2[27140] = 32'b11111111111111110010000101000111;
assign LUT_2[27141] = 32'b11111111111111101110111101100000;
assign LUT_2[27142] = 32'b11111111111111111000111110000011;
assign LUT_2[27143] = 32'b11111111111111110101110110011100;
assign LUT_2[27144] = 32'b11111111111111110000011000111100;
assign LUT_2[27145] = 32'b11111111111111101101010001010101;
assign LUT_2[27146] = 32'b11111111111111110111010001111000;
assign LUT_2[27147] = 32'b11111111111111110100001010010001;
assign LUT_2[27148] = 32'b11111111111111101100110110100100;
assign LUT_2[27149] = 32'b11111111111111101001101110111101;
assign LUT_2[27150] = 32'b11111111111111110011101111100000;
assign LUT_2[27151] = 32'b11111111111111110000100111111001;
assign LUT_2[27152] = 32'b11111111111111110000001011101001;
assign LUT_2[27153] = 32'b11111111111111101101000100000010;
assign LUT_2[27154] = 32'b11111111111111110111000100100101;
assign LUT_2[27155] = 32'b11111111111111110011111100111110;
assign LUT_2[27156] = 32'b11111111111111101100101001010001;
assign LUT_2[27157] = 32'b11111111111111101001100001101010;
assign LUT_2[27158] = 32'b11111111111111110011100010001101;
assign LUT_2[27159] = 32'b11111111111111110000011010100110;
assign LUT_2[27160] = 32'b11111111111111101010111101000110;
assign LUT_2[27161] = 32'b11111111111111100111110101011111;
assign LUT_2[27162] = 32'b11111111111111110001110110000010;
assign LUT_2[27163] = 32'b11111111111111101110101110011011;
assign LUT_2[27164] = 32'b11111111111111100111011010101110;
assign LUT_2[27165] = 32'b11111111111111100100010011000111;
assign LUT_2[27166] = 32'b11111111111111101110010011101010;
assign LUT_2[27167] = 32'b11111111111111101011001100000011;
assign LUT_2[27168] = 32'b11111111111111110110000011001000;
assign LUT_2[27169] = 32'b11111111111111110010111011100001;
assign LUT_2[27170] = 32'b11111111111111111100111100000100;
assign LUT_2[27171] = 32'b11111111111111111001110100011101;
assign LUT_2[27172] = 32'b11111111111111110010100000110000;
assign LUT_2[27173] = 32'b11111111111111101111011001001001;
assign LUT_2[27174] = 32'b11111111111111111001011001101100;
assign LUT_2[27175] = 32'b11111111111111110110010010000101;
assign LUT_2[27176] = 32'b11111111111111110000110100100101;
assign LUT_2[27177] = 32'b11111111111111101101101100111110;
assign LUT_2[27178] = 32'b11111111111111110111101101100001;
assign LUT_2[27179] = 32'b11111111111111110100100101111010;
assign LUT_2[27180] = 32'b11111111111111101101010010001101;
assign LUT_2[27181] = 32'b11111111111111101010001010100110;
assign LUT_2[27182] = 32'b11111111111111110100001011001001;
assign LUT_2[27183] = 32'b11111111111111110001000011100010;
assign LUT_2[27184] = 32'b11111111111111110000100111010010;
assign LUT_2[27185] = 32'b11111111111111101101011111101011;
assign LUT_2[27186] = 32'b11111111111111110111100000001110;
assign LUT_2[27187] = 32'b11111111111111110100011000100111;
assign LUT_2[27188] = 32'b11111111111111101101000100111010;
assign LUT_2[27189] = 32'b11111111111111101001111101010011;
assign LUT_2[27190] = 32'b11111111111111110011111101110110;
assign LUT_2[27191] = 32'b11111111111111110000110110001111;
assign LUT_2[27192] = 32'b11111111111111101011011000101111;
assign LUT_2[27193] = 32'b11111111111111101000010001001000;
assign LUT_2[27194] = 32'b11111111111111110010010001101011;
assign LUT_2[27195] = 32'b11111111111111101111001010000100;
assign LUT_2[27196] = 32'b11111111111111100111110110010111;
assign LUT_2[27197] = 32'b11111111111111100100101110110000;
assign LUT_2[27198] = 32'b11111111111111101110101111010011;
assign LUT_2[27199] = 32'b11111111111111101011100111101100;
assign LUT_2[27200] = 32'b11111111111111101101110000000010;
assign LUT_2[27201] = 32'b11111111111111101010101000011011;
assign LUT_2[27202] = 32'b11111111111111110100101000111110;
assign LUT_2[27203] = 32'b11111111111111110001100001010111;
assign LUT_2[27204] = 32'b11111111111111101010001101101010;
assign LUT_2[27205] = 32'b11111111111111100111000110000011;
assign LUT_2[27206] = 32'b11111111111111110001000110100110;
assign LUT_2[27207] = 32'b11111111111111101101111110111111;
assign LUT_2[27208] = 32'b11111111111111101000100001011111;
assign LUT_2[27209] = 32'b11111111111111100101011001111000;
assign LUT_2[27210] = 32'b11111111111111101111011010011011;
assign LUT_2[27211] = 32'b11111111111111101100010010110100;
assign LUT_2[27212] = 32'b11111111111111100100111111000111;
assign LUT_2[27213] = 32'b11111111111111100001110111100000;
assign LUT_2[27214] = 32'b11111111111111101011111000000011;
assign LUT_2[27215] = 32'b11111111111111101000110000011100;
assign LUT_2[27216] = 32'b11111111111111101000010100001100;
assign LUT_2[27217] = 32'b11111111111111100101001100100101;
assign LUT_2[27218] = 32'b11111111111111101111001101001000;
assign LUT_2[27219] = 32'b11111111111111101100000101100001;
assign LUT_2[27220] = 32'b11111111111111100100110001110100;
assign LUT_2[27221] = 32'b11111111111111100001101010001101;
assign LUT_2[27222] = 32'b11111111111111101011101010110000;
assign LUT_2[27223] = 32'b11111111111111101000100011001001;
assign LUT_2[27224] = 32'b11111111111111100011000101101001;
assign LUT_2[27225] = 32'b11111111111111011111111110000010;
assign LUT_2[27226] = 32'b11111111111111101001111110100101;
assign LUT_2[27227] = 32'b11111111111111100110110110111110;
assign LUT_2[27228] = 32'b11111111111111011111100011010001;
assign LUT_2[27229] = 32'b11111111111111011100011011101010;
assign LUT_2[27230] = 32'b11111111111111100110011100001101;
assign LUT_2[27231] = 32'b11111111111111100011010100100110;
assign LUT_2[27232] = 32'b11111111111111101110001011101011;
assign LUT_2[27233] = 32'b11111111111111101011000100000100;
assign LUT_2[27234] = 32'b11111111111111110101000100100111;
assign LUT_2[27235] = 32'b11111111111111110001111101000000;
assign LUT_2[27236] = 32'b11111111111111101010101001010011;
assign LUT_2[27237] = 32'b11111111111111100111100001101100;
assign LUT_2[27238] = 32'b11111111111111110001100010001111;
assign LUT_2[27239] = 32'b11111111111111101110011010101000;
assign LUT_2[27240] = 32'b11111111111111101000111101001000;
assign LUT_2[27241] = 32'b11111111111111100101110101100001;
assign LUT_2[27242] = 32'b11111111111111101111110110000100;
assign LUT_2[27243] = 32'b11111111111111101100101110011101;
assign LUT_2[27244] = 32'b11111111111111100101011010110000;
assign LUT_2[27245] = 32'b11111111111111100010010011001001;
assign LUT_2[27246] = 32'b11111111111111101100010011101100;
assign LUT_2[27247] = 32'b11111111111111101001001100000101;
assign LUT_2[27248] = 32'b11111111111111101000101111110101;
assign LUT_2[27249] = 32'b11111111111111100101101000001110;
assign LUT_2[27250] = 32'b11111111111111101111101000110001;
assign LUT_2[27251] = 32'b11111111111111101100100001001010;
assign LUT_2[27252] = 32'b11111111111111100101001101011101;
assign LUT_2[27253] = 32'b11111111111111100010000101110110;
assign LUT_2[27254] = 32'b11111111111111101100000110011001;
assign LUT_2[27255] = 32'b11111111111111101000111110110010;
assign LUT_2[27256] = 32'b11111111111111100011100001010010;
assign LUT_2[27257] = 32'b11111111111111100000011001101011;
assign LUT_2[27258] = 32'b11111111111111101010011010001110;
assign LUT_2[27259] = 32'b11111111111111100111010010100111;
assign LUT_2[27260] = 32'b11111111111111011111111110111010;
assign LUT_2[27261] = 32'b11111111111111011100110111010011;
assign LUT_2[27262] = 32'b11111111111111100110110111110110;
assign LUT_2[27263] = 32'b11111111111111100011110000001111;
assign LUT_2[27264] = 32'b11111111111111111001111011101110;
assign LUT_2[27265] = 32'b11111111111111110110110100000111;
assign LUT_2[27266] = 32'b00000000000000000000110100101010;
assign LUT_2[27267] = 32'b11111111111111111101101101000011;
assign LUT_2[27268] = 32'b11111111111111110110011001010110;
assign LUT_2[27269] = 32'b11111111111111110011010001101111;
assign LUT_2[27270] = 32'b11111111111111111101010010010010;
assign LUT_2[27271] = 32'b11111111111111111010001010101011;
assign LUT_2[27272] = 32'b11111111111111110100101101001011;
assign LUT_2[27273] = 32'b11111111111111110001100101100100;
assign LUT_2[27274] = 32'b11111111111111111011100110000111;
assign LUT_2[27275] = 32'b11111111111111111000011110100000;
assign LUT_2[27276] = 32'b11111111111111110001001010110011;
assign LUT_2[27277] = 32'b11111111111111101110000011001100;
assign LUT_2[27278] = 32'b11111111111111111000000011101111;
assign LUT_2[27279] = 32'b11111111111111110100111100001000;
assign LUT_2[27280] = 32'b11111111111111110100011111111000;
assign LUT_2[27281] = 32'b11111111111111110001011000010001;
assign LUT_2[27282] = 32'b11111111111111111011011000110100;
assign LUT_2[27283] = 32'b11111111111111111000010001001101;
assign LUT_2[27284] = 32'b11111111111111110000111101100000;
assign LUT_2[27285] = 32'b11111111111111101101110101111001;
assign LUT_2[27286] = 32'b11111111111111110111110110011100;
assign LUT_2[27287] = 32'b11111111111111110100101110110101;
assign LUT_2[27288] = 32'b11111111111111101111010001010101;
assign LUT_2[27289] = 32'b11111111111111101100001001101110;
assign LUT_2[27290] = 32'b11111111111111110110001010010001;
assign LUT_2[27291] = 32'b11111111111111110011000010101010;
assign LUT_2[27292] = 32'b11111111111111101011101110111101;
assign LUT_2[27293] = 32'b11111111111111101000100111010110;
assign LUT_2[27294] = 32'b11111111111111110010100111111001;
assign LUT_2[27295] = 32'b11111111111111101111100000010010;
assign LUT_2[27296] = 32'b11111111111111111010010111010111;
assign LUT_2[27297] = 32'b11111111111111110111001111110000;
assign LUT_2[27298] = 32'b00000000000000000001010000010011;
assign LUT_2[27299] = 32'b11111111111111111110001000101100;
assign LUT_2[27300] = 32'b11111111111111110110110100111111;
assign LUT_2[27301] = 32'b11111111111111110011101101011000;
assign LUT_2[27302] = 32'b11111111111111111101101101111011;
assign LUT_2[27303] = 32'b11111111111111111010100110010100;
assign LUT_2[27304] = 32'b11111111111111110101001000110100;
assign LUT_2[27305] = 32'b11111111111111110010000001001101;
assign LUT_2[27306] = 32'b11111111111111111100000001110000;
assign LUT_2[27307] = 32'b11111111111111111000111010001001;
assign LUT_2[27308] = 32'b11111111111111110001100110011100;
assign LUT_2[27309] = 32'b11111111111111101110011110110101;
assign LUT_2[27310] = 32'b11111111111111111000011111011000;
assign LUT_2[27311] = 32'b11111111111111110101010111110001;
assign LUT_2[27312] = 32'b11111111111111110100111011100001;
assign LUT_2[27313] = 32'b11111111111111110001110011111010;
assign LUT_2[27314] = 32'b11111111111111111011110100011101;
assign LUT_2[27315] = 32'b11111111111111111000101100110110;
assign LUT_2[27316] = 32'b11111111111111110001011001001001;
assign LUT_2[27317] = 32'b11111111111111101110010001100010;
assign LUT_2[27318] = 32'b11111111111111111000010010000101;
assign LUT_2[27319] = 32'b11111111111111110101001010011110;
assign LUT_2[27320] = 32'b11111111111111101111101100111110;
assign LUT_2[27321] = 32'b11111111111111101100100101010111;
assign LUT_2[27322] = 32'b11111111111111110110100101111010;
assign LUT_2[27323] = 32'b11111111111111110011011110010011;
assign LUT_2[27324] = 32'b11111111111111101100001010100110;
assign LUT_2[27325] = 32'b11111111111111101001000010111111;
assign LUT_2[27326] = 32'b11111111111111110011000011100010;
assign LUT_2[27327] = 32'b11111111111111101111111011111011;
assign LUT_2[27328] = 32'b11111111111111110010000100010001;
assign LUT_2[27329] = 32'b11111111111111101110111100101010;
assign LUT_2[27330] = 32'b11111111111111111000111101001101;
assign LUT_2[27331] = 32'b11111111111111110101110101100110;
assign LUT_2[27332] = 32'b11111111111111101110100001111001;
assign LUT_2[27333] = 32'b11111111111111101011011010010010;
assign LUT_2[27334] = 32'b11111111111111110101011010110101;
assign LUT_2[27335] = 32'b11111111111111110010010011001110;
assign LUT_2[27336] = 32'b11111111111111101100110101101110;
assign LUT_2[27337] = 32'b11111111111111101001101110000111;
assign LUT_2[27338] = 32'b11111111111111110011101110101010;
assign LUT_2[27339] = 32'b11111111111111110000100111000011;
assign LUT_2[27340] = 32'b11111111111111101001010011010110;
assign LUT_2[27341] = 32'b11111111111111100110001011101111;
assign LUT_2[27342] = 32'b11111111111111110000001100010010;
assign LUT_2[27343] = 32'b11111111111111101101000100101011;
assign LUT_2[27344] = 32'b11111111111111101100101000011011;
assign LUT_2[27345] = 32'b11111111111111101001100000110100;
assign LUT_2[27346] = 32'b11111111111111110011100001010111;
assign LUT_2[27347] = 32'b11111111111111110000011001110000;
assign LUT_2[27348] = 32'b11111111111111101001000110000011;
assign LUT_2[27349] = 32'b11111111111111100101111110011100;
assign LUT_2[27350] = 32'b11111111111111101111111110111111;
assign LUT_2[27351] = 32'b11111111111111101100110111011000;
assign LUT_2[27352] = 32'b11111111111111100111011001111000;
assign LUT_2[27353] = 32'b11111111111111100100010010010001;
assign LUT_2[27354] = 32'b11111111111111101110010010110100;
assign LUT_2[27355] = 32'b11111111111111101011001011001101;
assign LUT_2[27356] = 32'b11111111111111100011110111100000;
assign LUT_2[27357] = 32'b11111111111111100000101111111001;
assign LUT_2[27358] = 32'b11111111111111101010110000011100;
assign LUT_2[27359] = 32'b11111111111111100111101000110101;
assign LUT_2[27360] = 32'b11111111111111110010011111111010;
assign LUT_2[27361] = 32'b11111111111111101111011000010011;
assign LUT_2[27362] = 32'b11111111111111111001011000110110;
assign LUT_2[27363] = 32'b11111111111111110110010001001111;
assign LUT_2[27364] = 32'b11111111111111101110111101100010;
assign LUT_2[27365] = 32'b11111111111111101011110101111011;
assign LUT_2[27366] = 32'b11111111111111110101110110011110;
assign LUT_2[27367] = 32'b11111111111111110010101110110111;
assign LUT_2[27368] = 32'b11111111111111101101010001010111;
assign LUT_2[27369] = 32'b11111111111111101010001001110000;
assign LUT_2[27370] = 32'b11111111111111110100001010010011;
assign LUT_2[27371] = 32'b11111111111111110001000010101100;
assign LUT_2[27372] = 32'b11111111111111101001101110111111;
assign LUT_2[27373] = 32'b11111111111111100110100111011000;
assign LUT_2[27374] = 32'b11111111111111110000100111111011;
assign LUT_2[27375] = 32'b11111111111111101101100000010100;
assign LUT_2[27376] = 32'b11111111111111101101000100000100;
assign LUT_2[27377] = 32'b11111111111111101001111100011101;
assign LUT_2[27378] = 32'b11111111111111110011111101000000;
assign LUT_2[27379] = 32'b11111111111111110000110101011001;
assign LUT_2[27380] = 32'b11111111111111101001100001101100;
assign LUT_2[27381] = 32'b11111111111111100110011010000101;
assign LUT_2[27382] = 32'b11111111111111110000011010101000;
assign LUT_2[27383] = 32'b11111111111111101101010011000001;
assign LUT_2[27384] = 32'b11111111111111100111110101100001;
assign LUT_2[27385] = 32'b11111111111111100100101101111010;
assign LUT_2[27386] = 32'b11111111111111101110101110011101;
assign LUT_2[27387] = 32'b11111111111111101011100110110110;
assign LUT_2[27388] = 32'b11111111111111100100010011001001;
assign LUT_2[27389] = 32'b11111111111111100001001011100010;
assign LUT_2[27390] = 32'b11111111111111101011001100000101;
assign LUT_2[27391] = 32'b11111111111111101000000100011110;
assign LUT_2[27392] = 32'b11111111111111111001100110000101;
assign LUT_2[27393] = 32'b11111111111111110110011110011110;
assign LUT_2[27394] = 32'b00000000000000000000011111000001;
assign LUT_2[27395] = 32'b11111111111111111101010111011010;
assign LUT_2[27396] = 32'b11111111111111110110000011101101;
assign LUT_2[27397] = 32'b11111111111111110010111100000110;
assign LUT_2[27398] = 32'b11111111111111111100111100101001;
assign LUT_2[27399] = 32'b11111111111111111001110101000010;
assign LUT_2[27400] = 32'b11111111111111110100010111100010;
assign LUT_2[27401] = 32'b11111111111111110001001111111011;
assign LUT_2[27402] = 32'b11111111111111111011010000011110;
assign LUT_2[27403] = 32'b11111111111111111000001000110111;
assign LUT_2[27404] = 32'b11111111111111110000110101001010;
assign LUT_2[27405] = 32'b11111111111111101101101101100011;
assign LUT_2[27406] = 32'b11111111111111110111101110000110;
assign LUT_2[27407] = 32'b11111111111111110100100110011111;
assign LUT_2[27408] = 32'b11111111111111110100001010001111;
assign LUT_2[27409] = 32'b11111111111111110001000010101000;
assign LUT_2[27410] = 32'b11111111111111111011000011001011;
assign LUT_2[27411] = 32'b11111111111111110111111011100100;
assign LUT_2[27412] = 32'b11111111111111110000100111110111;
assign LUT_2[27413] = 32'b11111111111111101101100000010000;
assign LUT_2[27414] = 32'b11111111111111110111100000110011;
assign LUT_2[27415] = 32'b11111111111111110100011001001100;
assign LUT_2[27416] = 32'b11111111111111101110111011101100;
assign LUT_2[27417] = 32'b11111111111111101011110100000101;
assign LUT_2[27418] = 32'b11111111111111110101110100101000;
assign LUT_2[27419] = 32'b11111111111111110010101101000001;
assign LUT_2[27420] = 32'b11111111111111101011011001010100;
assign LUT_2[27421] = 32'b11111111111111101000010001101101;
assign LUT_2[27422] = 32'b11111111111111110010010010010000;
assign LUT_2[27423] = 32'b11111111111111101111001010101001;
assign LUT_2[27424] = 32'b11111111111111111010000001101110;
assign LUT_2[27425] = 32'b11111111111111110110111010000111;
assign LUT_2[27426] = 32'b00000000000000000000111010101010;
assign LUT_2[27427] = 32'b11111111111111111101110011000011;
assign LUT_2[27428] = 32'b11111111111111110110011111010110;
assign LUT_2[27429] = 32'b11111111111111110011010111101111;
assign LUT_2[27430] = 32'b11111111111111111101011000010010;
assign LUT_2[27431] = 32'b11111111111111111010010000101011;
assign LUT_2[27432] = 32'b11111111111111110100110011001011;
assign LUT_2[27433] = 32'b11111111111111110001101011100100;
assign LUT_2[27434] = 32'b11111111111111111011101100000111;
assign LUT_2[27435] = 32'b11111111111111111000100100100000;
assign LUT_2[27436] = 32'b11111111111111110001010000110011;
assign LUT_2[27437] = 32'b11111111111111101110001001001100;
assign LUT_2[27438] = 32'b11111111111111111000001001101111;
assign LUT_2[27439] = 32'b11111111111111110101000010001000;
assign LUT_2[27440] = 32'b11111111111111110100100101111000;
assign LUT_2[27441] = 32'b11111111111111110001011110010001;
assign LUT_2[27442] = 32'b11111111111111111011011110110100;
assign LUT_2[27443] = 32'b11111111111111111000010111001101;
assign LUT_2[27444] = 32'b11111111111111110001000011100000;
assign LUT_2[27445] = 32'b11111111111111101101111011111001;
assign LUT_2[27446] = 32'b11111111111111110111111100011100;
assign LUT_2[27447] = 32'b11111111111111110100110100110101;
assign LUT_2[27448] = 32'b11111111111111101111010111010101;
assign LUT_2[27449] = 32'b11111111111111101100001111101110;
assign LUT_2[27450] = 32'b11111111111111110110010000010001;
assign LUT_2[27451] = 32'b11111111111111110011001000101010;
assign LUT_2[27452] = 32'b11111111111111101011110100111101;
assign LUT_2[27453] = 32'b11111111111111101000101101010110;
assign LUT_2[27454] = 32'b11111111111111110010101101111001;
assign LUT_2[27455] = 32'b11111111111111101111100110010010;
assign LUT_2[27456] = 32'b11111111111111110001101110101000;
assign LUT_2[27457] = 32'b11111111111111101110100111000001;
assign LUT_2[27458] = 32'b11111111111111111000100111100100;
assign LUT_2[27459] = 32'b11111111111111110101011111111101;
assign LUT_2[27460] = 32'b11111111111111101110001100010000;
assign LUT_2[27461] = 32'b11111111111111101011000100101001;
assign LUT_2[27462] = 32'b11111111111111110101000101001100;
assign LUT_2[27463] = 32'b11111111111111110001111101100101;
assign LUT_2[27464] = 32'b11111111111111101100100000000101;
assign LUT_2[27465] = 32'b11111111111111101001011000011110;
assign LUT_2[27466] = 32'b11111111111111110011011001000001;
assign LUT_2[27467] = 32'b11111111111111110000010001011010;
assign LUT_2[27468] = 32'b11111111111111101000111101101101;
assign LUT_2[27469] = 32'b11111111111111100101110110000110;
assign LUT_2[27470] = 32'b11111111111111101111110110101001;
assign LUT_2[27471] = 32'b11111111111111101100101111000010;
assign LUT_2[27472] = 32'b11111111111111101100010010110010;
assign LUT_2[27473] = 32'b11111111111111101001001011001011;
assign LUT_2[27474] = 32'b11111111111111110011001011101110;
assign LUT_2[27475] = 32'b11111111111111110000000100000111;
assign LUT_2[27476] = 32'b11111111111111101000110000011010;
assign LUT_2[27477] = 32'b11111111111111100101101000110011;
assign LUT_2[27478] = 32'b11111111111111101111101001010110;
assign LUT_2[27479] = 32'b11111111111111101100100001101111;
assign LUT_2[27480] = 32'b11111111111111100111000100001111;
assign LUT_2[27481] = 32'b11111111111111100011111100101000;
assign LUT_2[27482] = 32'b11111111111111101101111101001011;
assign LUT_2[27483] = 32'b11111111111111101010110101100100;
assign LUT_2[27484] = 32'b11111111111111100011100001110111;
assign LUT_2[27485] = 32'b11111111111111100000011010010000;
assign LUT_2[27486] = 32'b11111111111111101010011010110011;
assign LUT_2[27487] = 32'b11111111111111100111010011001100;
assign LUT_2[27488] = 32'b11111111111111110010001010010001;
assign LUT_2[27489] = 32'b11111111111111101111000010101010;
assign LUT_2[27490] = 32'b11111111111111111001000011001101;
assign LUT_2[27491] = 32'b11111111111111110101111011100110;
assign LUT_2[27492] = 32'b11111111111111101110100111111001;
assign LUT_2[27493] = 32'b11111111111111101011100000010010;
assign LUT_2[27494] = 32'b11111111111111110101100000110101;
assign LUT_2[27495] = 32'b11111111111111110010011001001110;
assign LUT_2[27496] = 32'b11111111111111101100111011101110;
assign LUT_2[27497] = 32'b11111111111111101001110100000111;
assign LUT_2[27498] = 32'b11111111111111110011110100101010;
assign LUT_2[27499] = 32'b11111111111111110000101101000011;
assign LUT_2[27500] = 32'b11111111111111101001011001010110;
assign LUT_2[27501] = 32'b11111111111111100110010001101111;
assign LUT_2[27502] = 32'b11111111111111110000010010010010;
assign LUT_2[27503] = 32'b11111111111111101101001010101011;
assign LUT_2[27504] = 32'b11111111111111101100101110011011;
assign LUT_2[27505] = 32'b11111111111111101001100110110100;
assign LUT_2[27506] = 32'b11111111111111110011100111010111;
assign LUT_2[27507] = 32'b11111111111111110000011111110000;
assign LUT_2[27508] = 32'b11111111111111101001001100000011;
assign LUT_2[27509] = 32'b11111111111111100110000100011100;
assign LUT_2[27510] = 32'b11111111111111110000000100111111;
assign LUT_2[27511] = 32'b11111111111111101100111101011000;
assign LUT_2[27512] = 32'b11111111111111100111011111111000;
assign LUT_2[27513] = 32'b11111111111111100100011000010001;
assign LUT_2[27514] = 32'b11111111111111101110011000110100;
assign LUT_2[27515] = 32'b11111111111111101011010001001101;
assign LUT_2[27516] = 32'b11111111111111100011111101100000;
assign LUT_2[27517] = 32'b11111111111111100000110101111001;
assign LUT_2[27518] = 32'b11111111111111101010110110011100;
assign LUT_2[27519] = 32'b11111111111111100111101110110101;
assign LUT_2[27520] = 32'b11111111111111111101111010010100;
assign LUT_2[27521] = 32'b11111111111111111010110010101101;
assign LUT_2[27522] = 32'b00000000000000000100110011010000;
assign LUT_2[27523] = 32'b00000000000000000001101011101001;
assign LUT_2[27524] = 32'b11111111111111111010010111111100;
assign LUT_2[27525] = 32'b11111111111111110111010000010101;
assign LUT_2[27526] = 32'b00000000000000000001010000111000;
assign LUT_2[27527] = 32'b11111111111111111110001001010001;
assign LUT_2[27528] = 32'b11111111111111111000101011110001;
assign LUT_2[27529] = 32'b11111111111111110101100100001010;
assign LUT_2[27530] = 32'b11111111111111111111100100101101;
assign LUT_2[27531] = 32'b11111111111111111100011101000110;
assign LUT_2[27532] = 32'b11111111111111110101001001011001;
assign LUT_2[27533] = 32'b11111111111111110010000001110010;
assign LUT_2[27534] = 32'b11111111111111111100000010010101;
assign LUT_2[27535] = 32'b11111111111111111000111010101110;
assign LUT_2[27536] = 32'b11111111111111111000011110011110;
assign LUT_2[27537] = 32'b11111111111111110101010110110111;
assign LUT_2[27538] = 32'b11111111111111111111010111011010;
assign LUT_2[27539] = 32'b11111111111111111100001111110011;
assign LUT_2[27540] = 32'b11111111111111110100111100000110;
assign LUT_2[27541] = 32'b11111111111111110001110100011111;
assign LUT_2[27542] = 32'b11111111111111111011110101000010;
assign LUT_2[27543] = 32'b11111111111111111000101101011011;
assign LUT_2[27544] = 32'b11111111111111110011001111111011;
assign LUT_2[27545] = 32'b11111111111111110000001000010100;
assign LUT_2[27546] = 32'b11111111111111111010001000110111;
assign LUT_2[27547] = 32'b11111111111111110111000001010000;
assign LUT_2[27548] = 32'b11111111111111101111101101100011;
assign LUT_2[27549] = 32'b11111111111111101100100101111100;
assign LUT_2[27550] = 32'b11111111111111110110100110011111;
assign LUT_2[27551] = 32'b11111111111111110011011110111000;
assign LUT_2[27552] = 32'b11111111111111111110010101111101;
assign LUT_2[27553] = 32'b11111111111111111011001110010110;
assign LUT_2[27554] = 32'b00000000000000000101001110111001;
assign LUT_2[27555] = 32'b00000000000000000010000111010010;
assign LUT_2[27556] = 32'b11111111111111111010110011100101;
assign LUT_2[27557] = 32'b11111111111111110111101011111110;
assign LUT_2[27558] = 32'b00000000000000000001101100100001;
assign LUT_2[27559] = 32'b11111111111111111110100100111010;
assign LUT_2[27560] = 32'b11111111111111111001000111011010;
assign LUT_2[27561] = 32'b11111111111111110101111111110011;
assign LUT_2[27562] = 32'b00000000000000000000000000010110;
assign LUT_2[27563] = 32'b11111111111111111100111000101111;
assign LUT_2[27564] = 32'b11111111111111110101100101000010;
assign LUT_2[27565] = 32'b11111111111111110010011101011011;
assign LUT_2[27566] = 32'b11111111111111111100011101111110;
assign LUT_2[27567] = 32'b11111111111111111001010110010111;
assign LUT_2[27568] = 32'b11111111111111111000111010000111;
assign LUT_2[27569] = 32'b11111111111111110101110010100000;
assign LUT_2[27570] = 32'b11111111111111111111110011000011;
assign LUT_2[27571] = 32'b11111111111111111100101011011100;
assign LUT_2[27572] = 32'b11111111111111110101010111101111;
assign LUT_2[27573] = 32'b11111111111111110010010000001000;
assign LUT_2[27574] = 32'b11111111111111111100010000101011;
assign LUT_2[27575] = 32'b11111111111111111001001001000100;
assign LUT_2[27576] = 32'b11111111111111110011101011100100;
assign LUT_2[27577] = 32'b11111111111111110000100011111101;
assign LUT_2[27578] = 32'b11111111111111111010100100100000;
assign LUT_2[27579] = 32'b11111111111111110111011100111001;
assign LUT_2[27580] = 32'b11111111111111110000001001001100;
assign LUT_2[27581] = 32'b11111111111111101101000001100101;
assign LUT_2[27582] = 32'b11111111111111110111000010001000;
assign LUT_2[27583] = 32'b11111111111111110011111010100001;
assign LUT_2[27584] = 32'b11111111111111110110000010110111;
assign LUT_2[27585] = 32'b11111111111111110010111011010000;
assign LUT_2[27586] = 32'b11111111111111111100111011110011;
assign LUT_2[27587] = 32'b11111111111111111001110100001100;
assign LUT_2[27588] = 32'b11111111111111110010100000011111;
assign LUT_2[27589] = 32'b11111111111111101111011000111000;
assign LUT_2[27590] = 32'b11111111111111111001011001011011;
assign LUT_2[27591] = 32'b11111111111111110110010001110100;
assign LUT_2[27592] = 32'b11111111111111110000110100010100;
assign LUT_2[27593] = 32'b11111111111111101101101100101101;
assign LUT_2[27594] = 32'b11111111111111110111101101010000;
assign LUT_2[27595] = 32'b11111111111111110100100101101001;
assign LUT_2[27596] = 32'b11111111111111101101010001111100;
assign LUT_2[27597] = 32'b11111111111111101010001010010101;
assign LUT_2[27598] = 32'b11111111111111110100001010111000;
assign LUT_2[27599] = 32'b11111111111111110001000011010001;
assign LUT_2[27600] = 32'b11111111111111110000100111000001;
assign LUT_2[27601] = 32'b11111111111111101101011111011010;
assign LUT_2[27602] = 32'b11111111111111110111011111111101;
assign LUT_2[27603] = 32'b11111111111111110100011000010110;
assign LUT_2[27604] = 32'b11111111111111101101000100101001;
assign LUT_2[27605] = 32'b11111111111111101001111101000010;
assign LUT_2[27606] = 32'b11111111111111110011111101100101;
assign LUT_2[27607] = 32'b11111111111111110000110101111110;
assign LUT_2[27608] = 32'b11111111111111101011011000011110;
assign LUT_2[27609] = 32'b11111111111111101000010000110111;
assign LUT_2[27610] = 32'b11111111111111110010010001011010;
assign LUT_2[27611] = 32'b11111111111111101111001001110011;
assign LUT_2[27612] = 32'b11111111111111100111110110000110;
assign LUT_2[27613] = 32'b11111111111111100100101110011111;
assign LUT_2[27614] = 32'b11111111111111101110101111000010;
assign LUT_2[27615] = 32'b11111111111111101011100111011011;
assign LUT_2[27616] = 32'b11111111111111110110011110100000;
assign LUT_2[27617] = 32'b11111111111111110011010110111001;
assign LUT_2[27618] = 32'b11111111111111111101010111011100;
assign LUT_2[27619] = 32'b11111111111111111010001111110101;
assign LUT_2[27620] = 32'b11111111111111110010111100001000;
assign LUT_2[27621] = 32'b11111111111111101111110100100001;
assign LUT_2[27622] = 32'b11111111111111111001110101000100;
assign LUT_2[27623] = 32'b11111111111111110110101101011101;
assign LUT_2[27624] = 32'b11111111111111110001001111111101;
assign LUT_2[27625] = 32'b11111111111111101110001000010110;
assign LUT_2[27626] = 32'b11111111111111111000001000111001;
assign LUT_2[27627] = 32'b11111111111111110101000001010010;
assign LUT_2[27628] = 32'b11111111111111101101101101100101;
assign LUT_2[27629] = 32'b11111111111111101010100101111110;
assign LUT_2[27630] = 32'b11111111111111110100100110100001;
assign LUT_2[27631] = 32'b11111111111111110001011110111010;
assign LUT_2[27632] = 32'b11111111111111110001000010101010;
assign LUT_2[27633] = 32'b11111111111111101101111011000011;
assign LUT_2[27634] = 32'b11111111111111110111111011100110;
assign LUT_2[27635] = 32'b11111111111111110100110011111111;
assign LUT_2[27636] = 32'b11111111111111101101100000010010;
assign LUT_2[27637] = 32'b11111111111111101010011000101011;
assign LUT_2[27638] = 32'b11111111111111110100011001001110;
assign LUT_2[27639] = 32'b11111111111111110001010001100111;
assign LUT_2[27640] = 32'b11111111111111101011110100000111;
assign LUT_2[27641] = 32'b11111111111111101000101100100000;
assign LUT_2[27642] = 32'b11111111111111110010101101000011;
assign LUT_2[27643] = 32'b11111111111111101111100101011100;
assign LUT_2[27644] = 32'b11111111111111101000010001101111;
assign LUT_2[27645] = 32'b11111111111111100101001010001000;
assign LUT_2[27646] = 32'b11111111111111101111001010101011;
assign LUT_2[27647] = 32'b11111111111111101100000011000100;
assign LUT_2[27648] = 32'b11111111111111110111100001110010;
assign LUT_2[27649] = 32'b11111111111111110100011010001011;
assign LUT_2[27650] = 32'b11111111111111111110011010101110;
assign LUT_2[27651] = 32'b11111111111111111011010011000111;
assign LUT_2[27652] = 32'b11111111111111110011111111011010;
assign LUT_2[27653] = 32'b11111111111111110000110111110011;
assign LUT_2[27654] = 32'b11111111111111111010111000010110;
assign LUT_2[27655] = 32'b11111111111111110111110000101111;
assign LUT_2[27656] = 32'b11111111111111110010010011001111;
assign LUT_2[27657] = 32'b11111111111111101111001011101000;
assign LUT_2[27658] = 32'b11111111111111111001001100001011;
assign LUT_2[27659] = 32'b11111111111111110110000100100100;
assign LUT_2[27660] = 32'b11111111111111101110110000110111;
assign LUT_2[27661] = 32'b11111111111111101011101001010000;
assign LUT_2[27662] = 32'b11111111111111110101101001110011;
assign LUT_2[27663] = 32'b11111111111111110010100010001100;
assign LUT_2[27664] = 32'b11111111111111110010000101111100;
assign LUT_2[27665] = 32'b11111111111111101110111110010101;
assign LUT_2[27666] = 32'b11111111111111111000111110111000;
assign LUT_2[27667] = 32'b11111111111111110101110111010001;
assign LUT_2[27668] = 32'b11111111111111101110100011100100;
assign LUT_2[27669] = 32'b11111111111111101011011011111101;
assign LUT_2[27670] = 32'b11111111111111110101011100100000;
assign LUT_2[27671] = 32'b11111111111111110010010100111001;
assign LUT_2[27672] = 32'b11111111111111101100110111011001;
assign LUT_2[27673] = 32'b11111111111111101001101111110010;
assign LUT_2[27674] = 32'b11111111111111110011110000010101;
assign LUT_2[27675] = 32'b11111111111111110000101000101110;
assign LUT_2[27676] = 32'b11111111111111101001010101000001;
assign LUT_2[27677] = 32'b11111111111111100110001101011010;
assign LUT_2[27678] = 32'b11111111111111110000001101111101;
assign LUT_2[27679] = 32'b11111111111111101101000110010110;
assign LUT_2[27680] = 32'b11111111111111110111111101011011;
assign LUT_2[27681] = 32'b11111111111111110100110101110100;
assign LUT_2[27682] = 32'b11111111111111111110110110010111;
assign LUT_2[27683] = 32'b11111111111111111011101110110000;
assign LUT_2[27684] = 32'b11111111111111110100011011000011;
assign LUT_2[27685] = 32'b11111111111111110001010011011100;
assign LUT_2[27686] = 32'b11111111111111111011010011111111;
assign LUT_2[27687] = 32'b11111111111111111000001100011000;
assign LUT_2[27688] = 32'b11111111111111110010101110111000;
assign LUT_2[27689] = 32'b11111111111111101111100111010001;
assign LUT_2[27690] = 32'b11111111111111111001100111110100;
assign LUT_2[27691] = 32'b11111111111111110110100000001101;
assign LUT_2[27692] = 32'b11111111111111101111001100100000;
assign LUT_2[27693] = 32'b11111111111111101100000100111001;
assign LUT_2[27694] = 32'b11111111111111110110000101011100;
assign LUT_2[27695] = 32'b11111111111111110010111101110101;
assign LUT_2[27696] = 32'b11111111111111110010100001100101;
assign LUT_2[27697] = 32'b11111111111111101111011001111110;
assign LUT_2[27698] = 32'b11111111111111111001011010100001;
assign LUT_2[27699] = 32'b11111111111111110110010010111010;
assign LUT_2[27700] = 32'b11111111111111101110111111001101;
assign LUT_2[27701] = 32'b11111111111111101011110111100110;
assign LUT_2[27702] = 32'b11111111111111110101111000001001;
assign LUT_2[27703] = 32'b11111111111111110010110000100010;
assign LUT_2[27704] = 32'b11111111111111101101010011000010;
assign LUT_2[27705] = 32'b11111111111111101010001011011011;
assign LUT_2[27706] = 32'b11111111111111110100001011111110;
assign LUT_2[27707] = 32'b11111111111111110001000100010111;
assign LUT_2[27708] = 32'b11111111111111101001110000101010;
assign LUT_2[27709] = 32'b11111111111111100110101001000011;
assign LUT_2[27710] = 32'b11111111111111110000101001100110;
assign LUT_2[27711] = 32'b11111111111111101101100001111111;
assign LUT_2[27712] = 32'b11111111111111101111101010010101;
assign LUT_2[27713] = 32'b11111111111111101100100010101110;
assign LUT_2[27714] = 32'b11111111111111110110100011010001;
assign LUT_2[27715] = 32'b11111111111111110011011011101010;
assign LUT_2[27716] = 32'b11111111111111101100000111111101;
assign LUT_2[27717] = 32'b11111111111111101001000000010110;
assign LUT_2[27718] = 32'b11111111111111110011000000111001;
assign LUT_2[27719] = 32'b11111111111111101111111001010010;
assign LUT_2[27720] = 32'b11111111111111101010011011110010;
assign LUT_2[27721] = 32'b11111111111111100111010100001011;
assign LUT_2[27722] = 32'b11111111111111110001010100101110;
assign LUT_2[27723] = 32'b11111111111111101110001101000111;
assign LUT_2[27724] = 32'b11111111111111100110111001011010;
assign LUT_2[27725] = 32'b11111111111111100011110001110011;
assign LUT_2[27726] = 32'b11111111111111101101110010010110;
assign LUT_2[27727] = 32'b11111111111111101010101010101111;
assign LUT_2[27728] = 32'b11111111111111101010001110011111;
assign LUT_2[27729] = 32'b11111111111111100111000110111000;
assign LUT_2[27730] = 32'b11111111111111110001000111011011;
assign LUT_2[27731] = 32'b11111111111111101101111111110100;
assign LUT_2[27732] = 32'b11111111111111100110101100000111;
assign LUT_2[27733] = 32'b11111111111111100011100100100000;
assign LUT_2[27734] = 32'b11111111111111101101100101000011;
assign LUT_2[27735] = 32'b11111111111111101010011101011100;
assign LUT_2[27736] = 32'b11111111111111100100111111111100;
assign LUT_2[27737] = 32'b11111111111111100001111000010101;
assign LUT_2[27738] = 32'b11111111111111101011111000111000;
assign LUT_2[27739] = 32'b11111111111111101000110001010001;
assign LUT_2[27740] = 32'b11111111111111100001011101100100;
assign LUT_2[27741] = 32'b11111111111111011110010101111101;
assign LUT_2[27742] = 32'b11111111111111101000010110100000;
assign LUT_2[27743] = 32'b11111111111111100101001110111001;
assign LUT_2[27744] = 32'b11111111111111110000000101111110;
assign LUT_2[27745] = 32'b11111111111111101100111110010111;
assign LUT_2[27746] = 32'b11111111111111110110111110111010;
assign LUT_2[27747] = 32'b11111111111111110011110111010011;
assign LUT_2[27748] = 32'b11111111111111101100100011100110;
assign LUT_2[27749] = 32'b11111111111111101001011011111111;
assign LUT_2[27750] = 32'b11111111111111110011011100100010;
assign LUT_2[27751] = 32'b11111111111111110000010100111011;
assign LUT_2[27752] = 32'b11111111111111101010110111011011;
assign LUT_2[27753] = 32'b11111111111111100111101111110100;
assign LUT_2[27754] = 32'b11111111111111110001110000010111;
assign LUT_2[27755] = 32'b11111111111111101110101000110000;
assign LUT_2[27756] = 32'b11111111111111100111010101000011;
assign LUT_2[27757] = 32'b11111111111111100100001101011100;
assign LUT_2[27758] = 32'b11111111111111101110001101111111;
assign LUT_2[27759] = 32'b11111111111111101011000110011000;
assign LUT_2[27760] = 32'b11111111111111101010101010001000;
assign LUT_2[27761] = 32'b11111111111111100111100010100001;
assign LUT_2[27762] = 32'b11111111111111110001100011000100;
assign LUT_2[27763] = 32'b11111111111111101110011011011101;
assign LUT_2[27764] = 32'b11111111111111100111000111110000;
assign LUT_2[27765] = 32'b11111111111111100100000000001001;
assign LUT_2[27766] = 32'b11111111111111101110000000101100;
assign LUT_2[27767] = 32'b11111111111111101010111001000101;
assign LUT_2[27768] = 32'b11111111111111100101011011100101;
assign LUT_2[27769] = 32'b11111111111111100010010011111110;
assign LUT_2[27770] = 32'b11111111111111101100010100100001;
assign LUT_2[27771] = 32'b11111111111111101001001100111010;
assign LUT_2[27772] = 32'b11111111111111100001111001001101;
assign LUT_2[27773] = 32'b11111111111111011110110001100110;
assign LUT_2[27774] = 32'b11111111111111101000110010001001;
assign LUT_2[27775] = 32'b11111111111111100101101010100010;
assign LUT_2[27776] = 32'b11111111111111111011110110000001;
assign LUT_2[27777] = 32'b11111111111111111000101110011010;
assign LUT_2[27778] = 32'b00000000000000000010101110111101;
assign LUT_2[27779] = 32'b11111111111111111111100111010110;
assign LUT_2[27780] = 32'b11111111111111111000010011101001;
assign LUT_2[27781] = 32'b11111111111111110101001100000010;
assign LUT_2[27782] = 32'b11111111111111111111001100100101;
assign LUT_2[27783] = 32'b11111111111111111100000100111110;
assign LUT_2[27784] = 32'b11111111111111110110100111011110;
assign LUT_2[27785] = 32'b11111111111111110011011111110111;
assign LUT_2[27786] = 32'b11111111111111111101100000011010;
assign LUT_2[27787] = 32'b11111111111111111010011000110011;
assign LUT_2[27788] = 32'b11111111111111110011000101000110;
assign LUT_2[27789] = 32'b11111111111111101111111101011111;
assign LUT_2[27790] = 32'b11111111111111111001111110000010;
assign LUT_2[27791] = 32'b11111111111111110110110110011011;
assign LUT_2[27792] = 32'b11111111111111110110011010001011;
assign LUT_2[27793] = 32'b11111111111111110011010010100100;
assign LUT_2[27794] = 32'b11111111111111111101010011000111;
assign LUT_2[27795] = 32'b11111111111111111010001011100000;
assign LUT_2[27796] = 32'b11111111111111110010110111110011;
assign LUT_2[27797] = 32'b11111111111111101111110000001100;
assign LUT_2[27798] = 32'b11111111111111111001110000101111;
assign LUT_2[27799] = 32'b11111111111111110110101001001000;
assign LUT_2[27800] = 32'b11111111111111110001001011101000;
assign LUT_2[27801] = 32'b11111111111111101110000100000001;
assign LUT_2[27802] = 32'b11111111111111111000000100100100;
assign LUT_2[27803] = 32'b11111111111111110100111100111101;
assign LUT_2[27804] = 32'b11111111111111101101101001010000;
assign LUT_2[27805] = 32'b11111111111111101010100001101001;
assign LUT_2[27806] = 32'b11111111111111110100100010001100;
assign LUT_2[27807] = 32'b11111111111111110001011010100101;
assign LUT_2[27808] = 32'b11111111111111111100010001101010;
assign LUT_2[27809] = 32'b11111111111111111001001010000011;
assign LUT_2[27810] = 32'b00000000000000000011001010100110;
assign LUT_2[27811] = 32'b00000000000000000000000010111111;
assign LUT_2[27812] = 32'b11111111111111111000101111010010;
assign LUT_2[27813] = 32'b11111111111111110101100111101011;
assign LUT_2[27814] = 32'b11111111111111111111101000001110;
assign LUT_2[27815] = 32'b11111111111111111100100000100111;
assign LUT_2[27816] = 32'b11111111111111110111000011000111;
assign LUT_2[27817] = 32'b11111111111111110011111011100000;
assign LUT_2[27818] = 32'b11111111111111111101111100000011;
assign LUT_2[27819] = 32'b11111111111111111010110100011100;
assign LUT_2[27820] = 32'b11111111111111110011100000101111;
assign LUT_2[27821] = 32'b11111111111111110000011001001000;
assign LUT_2[27822] = 32'b11111111111111111010011001101011;
assign LUT_2[27823] = 32'b11111111111111110111010010000100;
assign LUT_2[27824] = 32'b11111111111111110110110101110100;
assign LUT_2[27825] = 32'b11111111111111110011101110001101;
assign LUT_2[27826] = 32'b11111111111111111101101110110000;
assign LUT_2[27827] = 32'b11111111111111111010100111001001;
assign LUT_2[27828] = 32'b11111111111111110011010011011100;
assign LUT_2[27829] = 32'b11111111111111110000001011110101;
assign LUT_2[27830] = 32'b11111111111111111010001100011000;
assign LUT_2[27831] = 32'b11111111111111110111000100110001;
assign LUT_2[27832] = 32'b11111111111111110001100111010001;
assign LUT_2[27833] = 32'b11111111111111101110011111101010;
assign LUT_2[27834] = 32'b11111111111111111000100000001101;
assign LUT_2[27835] = 32'b11111111111111110101011000100110;
assign LUT_2[27836] = 32'b11111111111111101110000100111001;
assign LUT_2[27837] = 32'b11111111111111101010111101010010;
assign LUT_2[27838] = 32'b11111111111111110100111101110101;
assign LUT_2[27839] = 32'b11111111111111110001110110001110;
assign LUT_2[27840] = 32'b11111111111111110011111110100100;
assign LUT_2[27841] = 32'b11111111111111110000110110111101;
assign LUT_2[27842] = 32'b11111111111111111010110111100000;
assign LUT_2[27843] = 32'b11111111111111110111101111111001;
assign LUT_2[27844] = 32'b11111111111111110000011100001100;
assign LUT_2[27845] = 32'b11111111111111101101010100100101;
assign LUT_2[27846] = 32'b11111111111111110111010101001000;
assign LUT_2[27847] = 32'b11111111111111110100001101100001;
assign LUT_2[27848] = 32'b11111111111111101110110000000001;
assign LUT_2[27849] = 32'b11111111111111101011101000011010;
assign LUT_2[27850] = 32'b11111111111111110101101000111101;
assign LUT_2[27851] = 32'b11111111111111110010100001010110;
assign LUT_2[27852] = 32'b11111111111111101011001101101001;
assign LUT_2[27853] = 32'b11111111111111101000000110000010;
assign LUT_2[27854] = 32'b11111111111111110010000110100101;
assign LUT_2[27855] = 32'b11111111111111101110111110111110;
assign LUT_2[27856] = 32'b11111111111111101110100010101110;
assign LUT_2[27857] = 32'b11111111111111101011011011000111;
assign LUT_2[27858] = 32'b11111111111111110101011011101010;
assign LUT_2[27859] = 32'b11111111111111110010010100000011;
assign LUT_2[27860] = 32'b11111111111111101011000000010110;
assign LUT_2[27861] = 32'b11111111111111100111111000101111;
assign LUT_2[27862] = 32'b11111111111111110001111001010010;
assign LUT_2[27863] = 32'b11111111111111101110110001101011;
assign LUT_2[27864] = 32'b11111111111111101001010100001011;
assign LUT_2[27865] = 32'b11111111111111100110001100100100;
assign LUT_2[27866] = 32'b11111111111111110000001101000111;
assign LUT_2[27867] = 32'b11111111111111101101000101100000;
assign LUT_2[27868] = 32'b11111111111111100101110001110011;
assign LUT_2[27869] = 32'b11111111111111100010101010001100;
assign LUT_2[27870] = 32'b11111111111111101100101010101111;
assign LUT_2[27871] = 32'b11111111111111101001100011001000;
assign LUT_2[27872] = 32'b11111111111111110100011010001101;
assign LUT_2[27873] = 32'b11111111111111110001010010100110;
assign LUT_2[27874] = 32'b11111111111111111011010011001001;
assign LUT_2[27875] = 32'b11111111111111111000001011100010;
assign LUT_2[27876] = 32'b11111111111111110000110111110101;
assign LUT_2[27877] = 32'b11111111111111101101110000001110;
assign LUT_2[27878] = 32'b11111111111111110111110000110001;
assign LUT_2[27879] = 32'b11111111111111110100101001001010;
assign LUT_2[27880] = 32'b11111111111111101111001011101010;
assign LUT_2[27881] = 32'b11111111111111101100000100000011;
assign LUT_2[27882] = 32'b11111111111111110110000100100110;
assign LUT_2[27883] = 32'b11111111111111110010111100111111;
assign LUT_2[27884] = 32'b11111111111111101011101001010010;
assign LUT_2[27885] = 32'b11111111111111101000100001101011;
assign LUT_2[27886] = 32'b11111111111111110010100010001110;
assign LUT_2[27887] = 32'b11111111111111101111011010100111;
assign LUT_2[27888] = 32'b11111111111111101110111110010111;
assign LUT_2[27889] = 32'b11111111111111101011110110110000;
assign LUT_2[27890] = 32'b11111111111111110101110111010011;
assign LUT_2[27891] = 32'b11111111111111110010101111101100;
assign LUT_2[27892] = 32'b11111111111111101011011011111111;
assign LUT_2[27893] = 32'b11111111111111101000010100011000;
assign LUT_2[27894] = 32'b11111111111111110010010100111011;
assign LUT_2[27895] = 32'b11111111111111101111001101010100;
assign LUT_2[27896] = 32'b11111111111111101001101111110100;
assign LUT_2[27897] = 32'b11111111111111100110101000001101;
assign LUT_2[27898] = 32'b11111111111111110000101000110000;
assign LUT_2[27899] = 32'b11111111111111101101100001001001;
assign LUT_2[27900] = 32'b11111111111111100110001101011100;
assign LUT_2[27901] = 32'b11111111111111100011000101110101;
assign LUT_2[27902] = 32'b11111111111111101101000110011000;
assign LUT_2[27903] = 32'b11111111111111101001111110110001;
assign LUT_2[27904] = 32'b11111111111111111011100000011000;
assign LUT_2[27905] = 32'b11111111111111111000011000110001;
assign LUT_2[27906] = 32'b00000000000000000010011001010100;
assign LUT_2[27907] = 32'b11111111111111111111010001101101;
assign LUT_2[27908] = 32'b11111111111111110111111110000000;
assign LUT_2[27909] = 32'b11111111111111110100110110011001;
assign LUT_2[27910] = 32'b11111111111111111110110110111100;
assign LUT_2[27911] = 32'b11111111111111111011101111010101;
assign LUT_2[27912] = 32'b11111111111111110110010001110101;
assign LUT_2[27913] = 32'b11111111111111110011001010001110;
assign LUT_2[27914] = 32'b11111111111111111101001010110001;
assign LUT_2[27915] = 32'b11111111111111111010000011001010;
assign LUT_2[27916] = 32'b11111111111111110010101111011101;
assign LUT_2[27917] = 32'b11111111111111101111100111110110;
assign LUT_2[27918] = 32'b11111111111111111001101000011001;
assign LUT_2[27919] = 32'b11111111111111110110100000110010;
assign LUT_2[27920] = 32'b11111111111111110110000100100010;
assign LUT_2[27921] = 32'b11111111111111110010111100111011;
assign LUT_2[27922] = 32'b11111111111111111100111101011110;
assign LUT_2[27923] = 32'b11111111111111111001110101110111;
assign LUT_2[27924] = 32'b11111111111111110010100010001010;
assign LUT_2[27925] = 32'b11111111111111101111011010100011;
assign LUT_2[27926] = 32'b11111111111111111001011011000110;
assign LUT_2[27927] = 32'b11111111111111110110010011011111;
assign LUT_2[27928] = 32'b11111111111111110000110101111111;
assign LUT_2[27929] = 32'b11111111111111101101101110011000;
assign LUT_2[27930] = 32'b11111111111111110111101110111011;
assign LUT_2[27931] = 32'b11111111111111110100100111010100;
assign LUT_2[27932] = 32'b11111111111111101101010011100111;
assign LUT_2[27933] = 32'b11111111111111101010001100000000;
assign LUT_2[27934] = 32'b11111111111111110100001100100011;
assign LUT_2[27935] = 32'b11111111111111110001000100111100;
assign LUT_2[27936] = 32'b11111111111111111011111100000001;
assign LUT_2[27937] = 32'b11111111111111111000110100011010;
assign LUT_2[27938] = 32'b00000000000000000010110100111101;
assign LUT_2[27939] = 32'b11111111111111111111101101010110;
assign LUT_2[27940] = 32'b11111111111111111000011001101001;
assign LUT_2[27941] = 32'b11111111111111110101010010000010;
assign LUT_2[27942] = 32'b11111111111111111111010010100101;
assign LUT_2[27943] = 32'b11111111111111111100001010111110;
assign LUT_2[27944] = 32'b11111111111111110110101101011110;
assign LUT_2[27945] = 32'b11111111111111110011100101110111;
assign LUT_2[27946] = 32'b11111111111111111101100110011010;
assign LUT_2[27947] = 32'b11111111111111111010011110110011;
assign LUT_2[27948] = 32'b11111111111111110011001011000110;
assign LUT_2[27949] = 32'b11111111111111110000000011011111;
assign LUT_2[27950] = 32'b11111111111111111010000100000010;
assign LUT_2[27951] = 32'b11111111111111110110111100011011;
assign LUT_2[27952] = 32'b11111111111111110110100000001011;
assign LUT_2[27953] = 32'b11111111111111110011011000100100;
assign LUT_2[27954] = 32'b11111111111111111101011001000111;
assign LUT_2[27955] = 32'b11111111111111111010010001100000;
assign LUT_2[27956] = 32'b11111111111111110010111101110011;
assign LUT_2[27957] = 32'b11111111111111101111110110001100;
assign LUT_2[27958] = 32'b11111111111111111001110110101111;
assign LUT_2[27959] = 32'b11111111111111110110101111001000;
assign LUT_2[27960] = 32'b11111111111111110001010001101000;
assign LUT_2[27961] = 32'b11111111111111101110001010000001;
assign LUT_2[27962] = 32'b11111111111111111000001010100100;
assign LUT_2[27963] = 32'b11111111111111110101000010111101;
assign LUT_2[27964] = 32'b11111111111111101101101111010000;
assign LUT_2[27965] = 32'b11111111111111101010100111101001;
assign LUT_2[27966] = 32'b11111111111111110100101000001100;
assign LUT_2[27967] = 32'b11111111111111110001100000100101;
assign LUT_2[27968] = 32'b11111111111111110011101000111011;
assign LUT_2[27969] = 32'b11111111111111110000100001010100;
assign LUT_2[27970] = 32'b11111111111111111010100001110111;
assign LUT_2[27971] = 32'b11111111111111110111011010010000;
assign LUT_2[27972] = 32'b11111111111111110000000110100011;
assign LUT_2[27973] = 32'b11111111111111101100111110111100;
assign LUT_2[27974] = 32'b11111111111111110110111111011111;
assign LUT_2[27975] = 32'b11111111111111110011110111111000;
assign LUT_2[27976] = 32'b11111111111111101110011010011000;
assign LUT_2[27977] = 32'b11111111111111101011010010110001;
assign LUT_2[27978] = 32'b11111111111111110101010011010100;
assign LUT_2[27979] = 32'b11111111111111110010001011101101;
assign LUT_2[27980] = 32'b11111111111111101010111000000000;
assign LUT_2[27981] = 32'b11111111111111100111110000011001;
assign LUT_2[27982] = 32'b11111111111111110001110000111100;
assign LUT_2[27983] = 32'b11111111111111101110101001010101;
assign LUT_2[27984] = 32'b11111111111111101110001101000101;
assign LUT_2[27985] = 32'b11111111111111101011000101011110;
assign LUT_2[27986] = 32'b11111111111111110101000110000001;
assign LUT_2[27987] = 32'b11111111111111110001111110011010;
assign LUT_2[27988] = 32'b11111111111111101010101010101101;
assign LUT_2[27989] = 32'b11111111111111100111100011000110;
assign LUT_2[27990] = 32'b11111111111111110001100011101001;
assign LUT_2[27991] = 32'b11111111111111101110011100000010;
assign LUT_2[27992] = 32'b11111111111111101000111110100010;
assign LUT_2[27993] = 32'b11111111111111100101110110111011;
assign LUT_2[27994] = 32'b11111111111111101111110111011110;
assign LUT_2[27995] = 32'b11111111111111101100101111110111;
assign LUT_2[27996] = 32'b11111111111111100101011100001010;
assign LUT_2[27997] = 32'b11111111111111100010010100100011;
assign LUT_2[27998] = 32'b11111111111111101100010101000110;
assign LUT_2[27999] = 32'b11111111111111101001001101011111;
assign LUT_2[28000] = 32'b11111111111111110100000100100100;
assign LUT_2[28001] = 32'b11111111111111110000111100111101;
assign LUT_2[28002] = 32'b11111111111111111010111101100000;
assign LUT_2[28003] = 32'b11111111111111110111110101111001;
assign LUT_2[28004] = 32'b11111111111111110000100010001100;
assign LUT_2[28005] = 32'b11111111111111101101011010100101;
assign LUT_2[28006] = 32'b11111111111111110111011011001000;
assign LUT_2[28007] = 32'b11111111111111110100010011100001;
assign LUT_2[28008] = 32'b11111111111111101110110110000001;
assign LUT_2[28009] = 32'b11111111111111101011101110011010;
assign LUT_2[28010] = 32'b11111111111111110101101110111101;
assign LUT_2[28011] = 32'b11111111111111110010100111010110;
assign LUT_2[28012] = 32'b11111111111111101011010011101001;
assign LUT_2[28013] = 32'b11111111111111101000001100000010;
assign LUT_2[28014] = 32'b11111111111111110010001100100101;
assign LUT_2[28015] = 32'b11111111111111101111000100111110;
assign LUT_2[28016] = 32'b11111111111111101110101000101110;
assign LUT_2[28017] = 32'b11111111111111101011100001000111;
assign LUT_2[28018] = 32'b11111111111111110101100001101010;
assign LUT_2[28019] = 32'b11111111111111110010011010000011;
assign LUT_2[28020] = 32'b11111111111111101011000110010110;
assign LUT_2[28021] = 32'b11111111111111100111111110101111;
assign LUT_2[28022] = 32'b11111111111111110001111111010010;
assign LUT_2[28023] = 32'b11111111111111101110110111101011;
assign LUT_2[28024] = 32'b11111111111111101001011010001011;
assign LUT_2[28025] = 32'b11111111111111100110010010100100;
assign LUT_2[28026] = 32'b11111111111111110000010011000111;
assign LUT_2[28027] = 32'b11111111111111101101001011100000;
assign LUT_2[28028] = 32'b11111111111111100101110111110011;
assign LUT_2[28029] = 32'b11111111111111100010110000001100;
assign LUT_2[28030] = 32'b11111111111111101100110000101111;
assign LUT_2[28031] = 32'b11111111111111101001101001001000;
assign LUT_2[28032] = 32'b11111111111111111111110100100111;
assign LUT_2[28033] = 32'b11111111111111111100101101000000;
assign LUT_2[28034] = 32'b00000000000000000110101101100011;
assign LUT_2[28035] = 32'b00000000000000000011100101111100;
assign LUT_2[28036] = 32'b11111111111111111100010010001111;
assign LUT_2[28037] = 32'b11111111111111111001001010101000;
assign LUT_2[28038] = 32'b00000000000000000011001011001011;
assign LUT_2[28039] = 32'b00000000000000000000000011100100;
assign LUT_2[28040] = 32'b11111111111111111010100110000100;
assign LUT_2[28041] = 32'b11111111111111110111011110011101;
assign LUT_2[28042] = 32'b00000000000000000001011111000000;
assign LUT_2[28043] = 32'b11111111111111111110010111011001;
assign LUT_2[28044] = 32'b11111111111111110111000011101100;
assign LUT_2[28045] = 32'b11111111111111110011111100000101;
assign LUT_2[28046] = 32'b11111111111111111101111100101000;
assign LUT_2[28047] = 32'b11111111111111111010110101000001;
assign LUT_2[28048] = 32'b11111111111111111010011000110001;
assign LUT_2[28049] = 32'b11111111111111110111010001001010;
assign LUT_2[28050] = 32'b00000000000000000001010001101101;
assign LUT_2[28051] = 32'b11111111111111111110001010000110;
assign LUT_2[28052] = 32'b11111111111111110110110110011001;
assign LUT_2[28053] = 32'b11111111111111110011101110110010;
assign LUT_2[28054] = 32'b11111111111111111101101111010101;
assign LUT_2[28055] = 32'b11111111111111111010100111101110;
assign LUT_2[28056] = 32'b11111111111111110101001010001110;
assign LUT_2[28057] = 32'b11111111111111110010000010100111;
assign LUT_2[28058] = 32'b11111111111111111100000011001010;
assign LUT_2[28059] = 32'b11111111111111111000111011100011;
assign LUT_2[28060] = 32'b11111111111111110001100111110110;
assign LUT_2[28061] = 32'b11111111111111101110100000001111;
assign LUT_2[28062] = 32'b11111111111111111000100000110010;
assign LUT_2[28063] = 32'b11111111111111110101011001001011;
assign LUT_2[28064] = 32'b00000000000000000000010000010000;
assign LUT_2[28065] = 32'b11111111111111111101001000101001;
assign LUT_2[28066] = 32'b00000000000000000111001001001100;
assign LUT_2[28067] = 32'b00000000000000000100000001100101;
assign LUT_2[28068] = 32'b11111111111111111100101101111000;
assign LUT_2[28069] = 32'b11111111111111111001100110010001;
assign LUT_2[28070] = 32'b00000000000000000011100110110100;
assign LUT_2[28071] = 32'b00000000000000000000011111001101;
assign LUT_2[28072] = 32'b11111111111111111011000001101101;
assign LUT_2[28073] = 32'b11111111111111110111111010000110;
assign LUT_2[28074] = 32'b00000000000000000001111010101001;
assign LUT_2[28075] = 32'b11111111111111111110110011000010;
assign LUT_2[28076] = 32'b11111111111111110111011111010101;
assign LUT_2[28077] = 32'b11111111111111110100010111101110;
assign LUT_2[28078] = 32'b11111111111111111110011000010001;
assign LUT_2[28079] = 32'b11111111111111111011010000101010;
assign LUT_2[28080] = 32'b11111111111111111010110100011010;
assign LUT_2[28081] = 32'b11111111111111110111101100110011;
assign LUT_2[28082] = 32'b00000000000000000001101101010110;
assign LUT_2[28083] = 32'b11111111111111111110100101101111;
assign LUT_2[28084] = 32'b11111111111111110111010010000010;
assign LUT_2[28085] = 32'b11111111111111110100001010011011;
assign LUT_2[28086] = 32'b11111111111111111110001010111110;
assign LUT_2[28087] = 32'b11111111111111111011000011010111;
assign LUT_2[28088] = 32'b11111111111111110101100101110111;
assign LUT_2[28089] = 32'b11111111111111110010011110010000;
assign LUT_2[28090] = 32'b11111111111111111100011110110011;
assign LUT_2[28091] = 32'b11111111111111111001010111001100;
assign LUT_2[28092] = 32'b11111111111111110010000011011111;
assign LUT_2[28093] = 32'b11111111111111101110111011111000;
assign LUT_2[28094] = 32'b11111111111111111000111100011011;
assign LUT_2[28095] = 32'b11111111111111110101110100110100;
assign LUT_2[28096] = 32'b11111111111111110111111101001010;
assign LUT_2[28097] = 32'b11111111111111110100110101100011;
assign LUT_2[28098] = 32'b11111111111111111110110110000110;
assign LUT_2[28099] = 32'b11111111111111111011101110011111;
assign LUT_2[28100] = 32'b11111111111111110100011010110010;
assign LUT_2[28101] = 32'b11111111111111110001010011001011;
assign LUT_2[28102] = 32'b11111111111111111011010011101110;
assign LUT_2[28103] = 32'b11111111111111111000001100000111;
assign LUT_2[28104] = 32'b11111111111111110010101110100111;
assign LUT_2[28105] = 32'b11111111111111101111100111000000;
assign LUT_2[28106] = 32'b11111111111111111001100111100011;
assign LUT_2[28107] = 32'b11111111111111110110011111111100;
assign LUT_2[28108] = 32'b11111111111111101111001100001111;
assign LUT_2[28109] = 32'b11111111111111101100000100101000;
assign LUT_2[28110] = 32'b11111111111111110110000101001011;
assign LUT_2[28111] = 32'b11111111111111110010111101100100;
assign LUT_2[28112] = 32'b11111111111111110010100001010100;
assign LUT_2[28113] = 32'b11111111111111101111011001101101;
assign LUT_2[28114] = 32'b11111111111111111001011010010000;
assign LUT_2[28115] = 32'b11111111111111110110010010101001;
assign LUT_2[28116] = 32'b11111111111111101110111110111100;
assign LUT_2[28117] = 32'b11111111111111101011110111010101;
assign LUT_2[28118] = 32'b11111111111111110101110111111000;
assign LUT_2[28119] = 32'b11111111111111110010110000010001;
assign LUT_2[28120] = 32'b11111111111111101101010010110001;
assign LUT_2[28121] = 32'b11111111111111101010001011001010;
assign LUT_2[28122] = 32'b11111111111111110100001011101101;
assign LUT_2[28123] = 32'b11111111111111110001000100000110;
assign LUT_2[28124] = 32'b11111111111111101001110000011001;
assign LUT_2[28125] = 32'b11111111111111100110101000110010;
assign LUT_2[28126] = 32'b11111111111111110000101001010101;
assign LUT_2[28127] = 32'b11111111111111101101100001101110;
assign LUT_2[28128] = 32'b11111111111111111000011000110011;
assign LUT_2[28129] = 32'b11111111111111110101010001001100;
assign LUT_2[28130] = 32'b11111111111111111111010001101111;
assign LUT_2[28131] = 32'b11111111111111111100001010001000;
assign LUT_2[28132] = 32'b11111111111111110100110110011011;
assign LUT_2[28133] = 32'b11111111111111110001101110110100;
assign LUT_2[28134] = 32'b11111111111111111011101111010111;
assign LUT_2[28135] = 32'b11111111111111111000100111110000;
assign LUT_2[28136] = 32'b11111111111111110011001010010000;
assign LUT_2[28137] = 32'b11111111111111110000000010101001;
assign LUT_2[28138] = 32'b11111111111111111010000011001100;
assign LUT_2[28139] = 32'b11111111111111110110111011100101;
assign LUT_2[28140] = 32'b11111111111111101111100111111000;
assign LUT_2[28141] = 32'b11111111111111101100100000010001;
assign LUT_2[28142] = 32'b11111111111111110110100000110100;
assign LUT_2[28143] = 32'b11111111111111110011011001001101;
assign LUT_2[28144] = 32'b11111111111111110010111100111101;
assign LUT_2[28145] = 32'b11111111111111101111110101010110;
assign LUT_2[28146] = 32'b11111111111111111001110101111001;
assign LUT_2[28147] = 32'b11111111111111110110101110010010;
assign LUT_2[28148] = 32'b11111111111111101111011010100101;
assign LUT_2[28149] = 32'b11111111111111101100010010111110;
assign LUT_2[28150] = 32'b11111111111111110110010011100001;
assign LUT_2[28151] = 32'b11111111111111110011001011111010;
assign LUT_2[28152] = 32'b11111111111111101101101110011010;
assign LUT_2[28153] = 32'b11111111111111101010100110110011;
assign LUT_2[28154] = 32'b11111111111111110100100111010110;
assign LUT_2[28155] = 32'b11111111111111110001011111101111;
assign LUT_2[28156] = 32'b11111111111111101010001100000010;
assign LUT_2[28157] = 32'b11111111111111100111000100011011;
assign LUT_2[28158] = 32'b11111111111111110001000100111110;
assign LUT_2[28159] = 32'b11111111111111101101111101010111;
assign LUT_2[28160] = 32'b11111111111111111100010011100100;
assign LUT_2[28161] = 32'b11111111111111111001001011111101;
assign LUT_2[28162] = 32'b00000000000000000011001100100000;
assign LUT_2[28163] = 32'b00000000000000000000000100111001;
assign LUT_2[28164] = 32'b11111111111111111000110001001100;
assign LUT_2[28165] = 32'b11111111111111110101101001100101;
assign LUT_2[28166] = 32'b11111111111111111111101010001000;
assign LUT_2[28167] = 32'b11111111111111111100100010100001;
assign LUT_2[28168] = 32'b11111111111111110111000101000001;
assign LUT_2[28169] = 32'b11111111111111110011111101011010;
assign LUT_2[28170] = 32'b11111111111111111101111101111101;
assign LUT_2[28171] = 32'b11111111111111111010110110010110;
assign LUT_2[28172] = 32'b11111111111111110011100010101001;
assign LUT_2[28173] = 32'b11111111111111110000011011000010;
assign LUT_2[28174] = 32'b11111111111111111010011011100101;
assign LUT_2[28175] = 32'b11111111111111110111010011111110;
assign LUT_2[28176] = 32'b11111111111111110110110111101110;
assign LUT_2[28177] = 32'b11111111111111110011110000000111;
assign LUT_2[28178] = 32'b11111111111111111101110000101010;
assign LUT_2[28179] = 32'b11111111111111111010101001000011;
assign LUT_2[28180] = 32'b11111111111111110011010101010110;
assign LUT_2[28181] = 32'b11111111111111110000001101101111;
assign LUT_2[28182] = 32'b11111111111111111010001110010010;
assign LUT_2[28183] = 32'b11111111111111110111000110101011;
assign LUT_2[28184] = 32'b11111111111111110001101001001011;
assign LUT_2[28185] = 32'b11111111111111101110100001100100;
assign LUT_2[28186] = 32'b11111111111111111000100010000111;
assign LUT_2[28187] = 32'b11111111111111110101011010100000;
assign LUT_2[28188] = 32'b11111111111111101110000110110011;
assign LUT_2[28189] = 32'b11111111111111101010111111001100;
assign LUT_2[28190] = 32'b11111111111111110100111111101111;
assign LUT_2[28191] = 32'b11111111111111110001111000001000;
assign LUT_2[28192] = 32'b11111111111111111100101111001101;
assign LUT_2[28193] = 32'b11111111111111111001100111100110;
assign LUT_2[28194] = 32'b00000000000000000011101000001001;
assign LUT_2[28195] = 32'b00000000000000000000100000100010;
assign LUT_2[28196] = 32'b11111111111111111001001100110101;
assign LUT_2[28197] = 32'b11111111111111110110000101001110;
assign LUT_2[28198] = 32'b00000000000000000000000101110001;
assign LUT_2[28199] = 32'b11111111111111111100111110001010;
assign LUT_2[28200] = 32'b11111111111111110111100000101010;
assign LUT_2[28201] = 32'b11111111111111110100011001000011;
assign LUT_2[28202] = 32'b11111111111111111110011001100110;
assign LUT_2[28203] = 32'b11111111111111111011010001111111;
assign LUT_2[28204] = 32'b11111111111111110011111110010010;
assign LUT_2[28205] = 32'b11111111111111110000110110101011;
assign LUT_2[28206] = 32'b11111111111111111010110111001110;
assign LUT_2[28207] = 32'b11111111111111110111101111100111;
assign LUT_2[28208] = 32'b11111111111111110111010011010111;
assign LUT_2[28209] = 32'b11111111111111110100001011110000;
assign LUT_2[28210] = 32'b11111111111111111110001100010011;
assign LUT_2[28211] = 32'b11111111111111111011000100101100;
assign LUT_2[28212] = 32'b11111111111111110011110000111111;
assign LUT_2[28213] = 32'b11111111111111110000101001011000;
assign LUT_2[28214] = 32'b11111111111111111010101001111011;
assign LUT_2[28215] = 32'b11111111111111110111100010010100;
assign LUT_2[28216] = 32'b11111111111111110010000100110100;
assign LUT_2[28217] = 32'b11111111111111101110111101001101;
assign LUT_2[28218] = 32'b11111111111111111000111101110000;
assign LUT_2[28219] = 32'b11111111111111110101110110001001;
assign LUT_2[28220] = 32'b11111111111111101110100010011100;
assign LUT_2[28221] = 32'b11111111111111101011011010110101;
assign LUT_2[28222] = 32'b11111111111111110101011011011000;
assign LUT_2[28223] = 32'b11111111111111110010010011110001;
assign LUT_2[28224] = 32'b11111111111111110100011100000111;
assign LUT_2[28225] = 32'b11111111111111110001010100100000;
assign LUT_2[28226] = 32'b11111111111111111011010101000011;
assign LUT_2[28227] = 32'b11111111111111111000001101011100;
assign LUT_2[28228] = 32'b11111111111111110000111001101111;
assign LUT_2[28229] = 32'b11111111111111101101110010001000;
assign LUT_2[28230] = 32'b11111111111111110111110010101011;
assign LUT_2[28231] = 32'b11111111111111110100101011000100;
assign LUT_2[28232] = 32'b11111111111111101111001101100100;
assign LUT_2[28233] = 32'b11111111111111101100000101111101;
assign LUT_2[28234] = 32'b11111111111111110110000110100000;
assign LUT_2[28235] = 32'b11111111111111110010111110111001;
assign LUT_2[28236] = 32'b11111111111111101011101011001100;
assign LUT_2[28237] = 32'b11111111111111101000100011100101;
assign LUT_2[28238] = 32'b11111111111111110010100100001000;
assign LUT_2[28239] = 32'b11111111111111101111011100100001;
assign LUT_2[28240] = 32'b11111111111111101111000000010001;
assign LUT_2[28241] = 32'b11111111111111101011111000101010;
assign LUT_2[28242] = 32'b11111111111111110101111001001101;
assign LUT_2[28243] = 32'b11111111111111110010110001100110;
assign LUT_2[28244] = 32'b11111111111111101011011101111001;
assign LUT_2[28245] = 32'b11111111111111101000010110010010;
assign LUT_2[28246] = 32'b11111111111111110010010110110101;
assign LUT_2[28247] = 32'b11111111111111101111001111001110;
assign LUT_2[28248] = 32'b11111111111111101001110001101110;
assign LUT_2[28249] = 32'b11111111111111100110101010000111;
assign LUT_2[28250] = 32'b11111111111111110000101010101010;
assign LUT_2[28251] = 32'b11111111111111101101100011000011;
assign LUT_2[28252] = 32'b11111111111111100110001111010110;
assign LUT_2[28253] = 32'b11111111111111100011000111101111;
assign LUT_2[28254] = 32'b11111111111111101101001000010010;
assign LUT_2[28255] = 32'b11111111111111101010000000101011;
assign LUT_2[28256] = 32'b11111111111111110100110111110000;
assign LUT_2[28257] = 32'b11111111111111110001110000001001;
assign LUT_2[28258] = 32'b11111111111111111011110000101100;
assign LUT_2[28259] = 32'b11111111111111111000101001000101;
assign LUT_2[28260] = 32'b11111111111111110001010101011000;
assign LUT_2[28261] = 32'b11111111111111101110001101110001;
assign LUT_2[28262] = 32'b11111111111111111000001110010100;
assign LUT_2[28263] = 32'b11111111111111110101000110101101;
assign LUT_2[28264] = 32'b11111111111111101111101001001101;
assign LUT_2[28265] = 32'b11111111111111101100100001100110;
assign LUT_2[28266] = 32'b11111111111111110110100010001001;
assign LUT_2[28267] = 32'b11111111111111110011011010100010;
assign LUT_2[28268] = 32'b11111111111111101100000110110101;
assign LUT_2[28269] = 32'b11111111111111101000111111001110;
assign LUT_2[28270] = 32'b11111111111111110010111111110001;
assign LUT_2[28271] = 32'b11111111111111101111111000001010;
assign LUT_2[28272] = 32'b11111111111111101111011011111010;
assign LUT_2[28273] = 32'b11111111111111101100010100010011;
assign LUT_2[28274] = 32'b11111111111111110110010100110110;
assign LUT_2[28275] = 32'b11111111111111110011001101001111;
assign LUT_2[28276] = 32'b11111111111111101011111001100010;
assign LUT_2[28277] = 32'b11111111111111101000110001111011;
assign LUT_2[28278] = 32'b11111111111111110010110010011110;
assign LUT_2[28279] = 32'b11111111111111101111101010110111;
assign LUT_2[28280] = 32'b11111111111111101010001101010111;
assign LUT_2[28281] = 32'b11111111111111100111000101110000;
assign LUT_2[28282] = 32'b11111111111111110001000110010011;
assign LUT_2[28283] = 32'b11111111111111101101111110101100;
assign LUT_2[28284] = 32'b11111111111111100110101010111111;
assign LUT_2[28285] = 32'b11111111111111100011100011011000;
assign LUT_2[28286] = 32'b11111111111111101101100011111011;
assign LUT_2[28287] = 32'b11111111111111101010011100010100;
assign LUT_2[28288] = 32'b00000000000000000000100111110011;
assign LUT_2[28289] = 32'b11111111111111111101100000001100;
assign LUT_2[28290] = 32'b00000000000000000111100000101111;
assign LUT_2[28291] = 32'b00000000000000000100011001001000;
assign LUT_2[28292] = 32'b11111111111111111101000101011011;
assign LUT_2[28293] = 32'b11111111111111111001111101110100;
assign LUT_2[28294] = 32'b00000000000000000011111110010111;
assign LUT_2[28295] = 32'b00000000000000000000110110110000;
assign LUT_2[28296] = 32'b11111111111111111011011001010000;
assign LUT_2[28297] = 32'b11111111111111111000010001101001;
assign LUT_2[28298] = 32'b00000000000000000010010010001100;
assign LUT_2[28299] = 32'b11111111111111111111001010100101;
assign LUT_2[28300] = 32'b11111111111111110111110110111000;
assign LUT_2[28301] = 32'b11111111111111110100101111010001;
assign LUT_2[28302] = 32'b11111111111111111110101111110100;
assign LUT_2[28303] = 32'b11111111111111111011101000001101;
assign LUT_2[28304] = 32'b11111111111111111011001011111101;
assign LUT_2[28305] = 32'b11111111111111111000000100010110;
assign LUT_2[28306] = 32'b00000000000000000010000100111001;
assign LUT_2[28307] = 32'b11111111111111111110111101010010;
assign LUT_2[28308] = 32'b11111111111111110111101001100101;
assign LUT_2[28309] = 32'b11111111111111110100100001111110;
assign LUT_2[28310] = 32'b11111111111111111110100010100001;
assign LUT_2[28311] = 32'b11111111111111111011011010111010;
assign LUT_2[28312] = 32'b11111111111111110101111101011010;
assign LUT_2[28313] = 32'b11111111111111110010110101110011;
assign LUT_2[28314] = 32'b11111111111111111100110110010110;
assign LUT_2[28315] = 32'b11111111111111111001101110101111;
assign LUT_2[28316] = 32'b11111111111111110010011011000010;
assign LUT_2[28317] = 32'b11111111111111101111010011011011;
assign LUT_2[28318] = 32'b11111111111111111001010011111110;
assign LUT_2[28319] = 32'b11111111111111110110001100010111;
assign LUT_2[28320] = 32'b00000000000000000001000011011100;
assign LUT_2[28321] = 32'b11111111111111111101111011110101;
assign LUT_2[28322] = 32'b00000000000000000111111100011000;
assign LUT_2[28323] = 32'b00000000000000000100110100110001;
assign LUT_2[28324] = 32'b11111111111111111101100001000100;
assign LUT_2[28325] = 32'b11111111111111111010011001011101;
assign LUT_2[28326] = 32'b00000000000000000100011010000000;
assign LUT_2[28327] = 32'b00000000000000000001010010011001;
assign LUT_2[28328] = 32'b11111111111111111011110100111001;
assign LUT_2[28329] = 32'b11111111111111111000101101010010;
assign LUT_2[28330] = 32'b00000000000000000010101101110101;
assign LUT_2[28331] = 32'b11111111111111111111100110001110;
assign LUT_2[28332] = 32'b11111111111111111000010010100001;
assign LUT_2[28333] = 32'b11111111111111110101001010111010;
assign LUT_2[28334] = 32'b11111111111111111111001011011101;
assign LUT_2[28335] = 32'b11111111111111111100000011110110;
assign LUT_2[28336] = 32'b11111111111111111011100111100110;
assign LUT_2[28337] = 32'b11111111111111111000011111111111;
assign LUT_2[28338] = 32'b00000000000000000010100000100010;
assign LUT_2[28339] = 32'b11111111111111111111011000111011;
assign LUT_2[28340] = 32'b11111111111111111000000101001110;
assign LUT_2[28341] = 32'b11111111111111110100111101100111;
assign LUT_2[28342] = 32'b11111111111111111110111110001010;
assign LUT_2[28343] = 32'b11111111111111111011110110100011;
assign LUT_2[28344] = 32'b11111111111111110110011001000011;
assign LUT_2[28345] = 32'b11111111111111110011010001011100;
assign LUT_2[28346] = 32'b11111111111111111101010001111111;
assign LUT_2[28347] = 32'b11111111111111111010001010011000;
assign LUT_2[28348] = 32'b11111111111111110010110110101011;
assign LUT_2[28349] = 32'b11111111111111101111101111000100;
assign LUT_2[28350] = 32'b11111111111111111001101111100111;
assign LUT_2[28351] = 32'b11111111111111110110101000000000;
assign LUT_2[28352] = 32'b11111111111111111000110000010110;
assign LUT_2[28353] = 32'b11111111111111110101101000101111;
assign LUT_2[28354] = 32'b11111111111111111111101001010010;
assign LUT_2[28355] = 32'b11111111111111111100100001101011;
assign LUT_2[28356] = 32'b11111111111111110101001101111110;
assign LUT_2[28357] = 32'b11111111111111110010000110010111;
assign LUT_2[28358] = 32'b11111111111111111100000110111010;
assign LUT_2[28359] = 32'b11111111111111111000111111010011;
assign LUT_2[28360] = 32'b11111111111111110011100001110011;
assign LUT_2[28361] = 32'b11111111111111110000011010001100;
assign LUT_2[28362] = 32'b11111111111111111010011010101111;
assign LUT_2[28363] = 32'b11111111111111110111010011001000;
assign LUT_2[28364] = 32'b11111111111111101111111111011011;
assign LUT_2[28365] = 32'b11111111111111101100110111110100;
assign LUT_2[28366] = 32'b11111111111111110110111000010111;
assign LUT_2[28367] = 32'b11111111111111110011110000110000;
assign LUT_2[28368] = 32'b11111111111111110011010100100000;
assign LUT_2[28369] = 32'b11111111111111110000001100111001;
assign LUT_2[28370] = 32'b11111111111111111010001101011100;
assign LUT_2[28371] = 32'b11111111111111110111000101110101;
assign LUT_2[28372] = 32'b11111111111111101111110010001000;
assign LUT_2[28373] = 32'b11111111111111101100101010100001;
assign LUT_2[28374] = 32'b11111111111111110110101011000100;
assign LUT_2[28375] = 32'b11111111111111110011100011011101;
assign LUT_2[28376] = 32'b11111111111111101110000101111101;
assign LUT_2[28377] = 32'b11111111111111101010111110010110;
assign LUT_2[28378] = 32'b11111111111111110100111110111001;
assign LUT_2[28379] = 32'b11111111111111110001110111010010;
assign LUT_2[28380] = 32'b11111111111111101010100011100101;
assign LUT_2[28381] = 32'b11111111111111100111011011111110;
assign LUT_2[28382] = 32'b11111111111111110001011100100001;
assign LUT_2[28383] = 32'b11111111111111101110010100111010;
assign LUT_2[28384] = 32'b11111111111111111001001011111111;
assign LUT_2[28385] = 32'b11111111111111110110000100011000;
assign LUT_2[28386] = 32'b00000000000000000000000100111011;
assign LUT_2[28387] = 32'b11111111111111111100111101010100;
assign LUT_2[28388] = 32'b11111111111111110101101001100111;
assign LUT_2[28389] = 32'b11111111111111110010100010000000;
assign LUT_2[28390] = 32'b11111111111111111100100010100011;
assign LUT_2[28391] = 32'b11111111111111111001011010111100;
assign LUT_2[28392] = 32'b11111111111111110011111101011100;
assign LUT_2[28393] = 32'b11111111111111110000110101110101;
assign LUT_2[28394] = 32'b11111111111111111010110110011000;
assign LUT_2[28395] = 32'b11111111111111110111101110110001;
assign LUT_2[28396] = 32'b11111111111111110000011011000100;
assign LUT_2[28397] = 32'b11111111111111101101010011011101;
assign LUT_2[28398] = 32'b11111111111111110111010100000000;
assign LUT_2[28399] = 32'b11111111111111110100001100011001;
assign LUT_2[28400] = 32'b11111111111111110011110000001001;
assign LUT_2[28401] = 32'b11111111111111110000101000100010;
assign LUT_2[28402] = 32'b11111111111111111010101001000101;
assign LUT_2[28403] = 32'b11111111111111110111100001011110;
assign LUT_2[28404] = 32'b11111111111111110000001101110001;
assign LUT_2[28405] = 32'b11111111111111101101000110001010;
assign LUT_2[28406] = 32'b11111111111111110111000110101101;
assign LUT_2[28407] = 32'b11111111111111110011111111000110;
assign LUT_2[28408] = 32'b11111111111111101110100001100110;
assign LUT_2[28409] = 32'b11111111111111101011011001111111;
assign LUT_2[28410] = 32'b11111111111111110101011010100010;
assign LUT_2[28411] = 32'b11111111111111110010010010111011;
assign LUT_2[28412] = 32'b11111111111111101010111111001110;
assign LUT_2[28413] = 32'b11111111111111100111110111100111;
assign LUT_2[28414] = 32'b11111111111111110001111000001010;
assign LUT_2[28415] = 32'b11111111111111101110110000100011;
assign LUT_2[28416] = 32'b00000000000000000000010010001010;
assign LUT_2[28417] = 32'b11111111111111111101001010100011;
assign LUT_2[28418] = 32'b00000000000000000111001011000110;
assign LUT_2[28419] = 32'b00000000000000000100000011011111;
assign LUT_2[28420] = 32'b11111111111111111100101111110010;
assign LUT_2[28421] = 32'b11111111111111111001101000001011;
assign LUT_2[28422] = 32'b00000000000000000011101000101110;
assign LUT_2[28423] = 32'b00000000000000000000100001000111;
assign LUT_2[28424] = 32'b11111111111111111011000011100111;
assign LUT_2[28425] = 32'b11111111111111110111111100000000;
assign LUT_2[28426] = 32'b00000000000000000001111100100011;
assign LUT_2[28427] = 32'b11111111111111111110110100111100;
assign LUT_2[28428] = 32'b11111111111111110111100001001111;
assign LUT_2[28429] = 32'b11111111111111110100011001101000;
assign LUT_2[28430] = 32'b11111111111111111110011010001011;
assign LUT_2[28431] = 32'b11111111111111111011010010100100;
assign LUT_2[28432] = 32'b11111111111111111010110110010100;
assign LUT_2[28433] = 32'b11111111111111110111101110101101;
assign LUT_2[28434] = 32'b00000000000000000001101111010000;
assign LUT_2[28435] = 32'b11111111111111111110100111101001;
assign LUT_2[28436] = 32'b11111111111111110111010011111100;
assign LUT_2[28437] = 32'b11111111111111110100001100010101;
assign LUT_2[28438] = 32'b11111111111111111110001100111000;
assign LUT_2[28439] = 32'b11111111111111111011000101010001;
assign LUT_2[28440] = 32'b11111111111111110101100111110001;
assign LUT_2[28441] = 32'b11111111111111110010100000001010;
assign LUT_2[28442] = 32'b11111111111111111100100000101101;
assign LUT_2[28443] = 32'b11111111111111111001011001000110;
assign LUT_2[28444] = 32'b11111111111111110010000101011001;
assign LUT_2[28445] = 32'b11111111111111101110111101110010;
assign LUT_2[28446] = 32'b11111111111111111000111110010101;
assign LUT_2[28447] = 32'b11111111111111110101110110101110;
assign LUT_2[28448] = 32'b00000000000000000000101101110011;
assign LUT_2[28449] = 32'b11111111111111111101100110001100;
assign LUT_2[28450] = 32'b00000000000000000111100110101111;
assign LUT_2[28451] = 32'b00000000000000000100011111001000;
assign LUT_2[28452] = 32'b11111111111111111101001011011011;
assign LUT_2[28453] = 32'b11111111111111111010000011110100;
assign LUT_2[28454] = 32'b00000000000000000100000100010111;
assign LUT_2[28455] = 32'b00000000000000000000111100110000;
assign LUT_2[28456] = 32'b11111111111111111011011111010000;
assign LUT_2[28457] = 32'b11111111111111111000010111101001;
assign LUT_2[28458] = 32'b00000000000000000010011000001100;
assign LUT_2[28459] = 32'b11111111111111111111010000100101;
assign LUT_2[28460] = 32'b11111111111111110111111100111000;
assign LUT_2[28461] = 32'b11111111111111110100110101010001;
assign LUT_2[28462] = 32'b11111111111111111110110101110100;
assign LUT_2[28463] = 32'b11111111111111111011101110001101;
assign LUT_2[28464] = 32'b11111111111111111011010001111101;
assign LUT_2[28465] = 32'b11111111111111111000001010010110;
assign LUT_2[28466] = 32'b00000000000000000010001010111001;
assign LUT_2[28467] = 32'b11111111111111111111000011010010;
assign LUT_2[28468] = 32'b11111111111111110111101111100101;
assign LUT_2[28469] = 32'b11111111111111110100100111111110;
assign LUT_2[28470] = 32'b11111111111111111110101000100001;
assign LUT_2[28471] = 32'b11111111111111111011100000111010;
assign LUT_2[28472] = 32'b11111111111111110110000011011010;
assign LUT_2[28473] = 32'b11111111111111110010111011110011;
assign LUT_2[28474] = 32'b11111111111111111100111100010110;
assign LUT_2[28475] = 32'b11111111111111111001110100101111;
assign LUT_2[28476] = 32'b11111111111111110010100001000010;
assign LUT_2[28477] = 32'b11111111111111101111011001011011;
assign LUT_2[28478] = 32'b11111111111111111001011001111110;
assign LUT_2[28479] = 32'b11111111111111110110010010010111;
assign LUT_2[28480] = 32'b11111111111111111000011010101101;
assign LUT_2[28481] = 32'b11111111111111110101010011000110;
assign LUT_2[28482] = 32'b11111111111111111111010011101001;
assign LUT_2[28483] = 32'b11111111111111111100001100000010;
assign LUT_2[28484] = 32'b11111111111111110100111000010101;
assign LUT_2[28485] = 32'b11111111111111110001110000101110;
assign LUT_2[28486] = 32'b11111111111111111011110001010001;
assign LUT_2[28487] = 32'b11111111111111111000101001101010;
assign LUT_2[28488] = 32'b11111111111111110011001100001010;
assign LUT_2[28489] = 32'b11111111111111110000000100100011;
assign LUT_2[28490] = 32'b11111111111111111010000101000110;
assign LUT_2[28491] = 32'b11111111111111110110111101011111;
assign LUT_2[28492] = 32'b11111111111111101111101001110010;
assign LUT_2[28493] = 32'b11111111111111101100100010001011;
assign LUT_2[28494] = 32'b11111111111111110110100010101110;
assign LUT_2[28495] = 32'b11111111111111110011011011000111;
assign LUT_2[28496] = 32'b11111111111111110010111110110111;
assign LUT_2[28497] = 32'b11111111111111101111110111010000;
assign LUT_2[28498] = 32'b11111111111111111001110111110011;
assign LUT_2[28499] = 32'b11111111111111110110110000001100;
assign LUT_2[28500] = 32'b11111111111111101111011100011111;
assign LUT_2[28501] = 32'b11111111111111101100010100111000;
assign LUT_2[28502] = 32'b11111111111111110110010101011011;
assign LUT_2[28503] = 32'b11111111111111110011001101110100;
assign LUT_2[28504] = 32'b11111111111111101101110000010100;
assign LUT_2[28505] = 32'b11111111111111101010101000101101;
assign LUT_2[28506] = 32'b11111111111111110100101001010000;
assign LUT_2[28507] = 32'b11111111111111110001100001101001;
assign LUT_2[28508] = 32'b11111111111111101010001101111100;
assign LUT_2[28509] = 32'b11111111111111100111000110010101;
assign LUT_2[28510] = 32'b11111111111111110001000110111000;
assign LUT_2[28511] = 32'b11111111111111101101111111010001;
assign LUT_2[28512] = 32'b11111111111111111000110110010110;
assign LUT_2[28513] = 32'b11111111111111110101101110101111;
assign LUT_2[28514] = 32'b11111111111111111111101111010010;
assign LUT_2[28515] = 32'b11111111111111111100100111101011;
assign LUT_2[28516] = 32'b11111111111111110101010011111110;
assign LUT_2[28517] = 32'b11111111111111110010001100010111;
assign LUT_2[28518] = 32'b11111111111111111100001100111010;
assign LUT_2[28519] = 32'b11111111111111111001000101010011;
assign LUT_2[28520] = 32'b11111111111111110011100111110011;
assign LUT_2[28521] = 32'b11111111111111110000100000001100;
assign LUT_2[28522] = 32'b11111111111111111010100000101111;
assign LUT_2[28523] = 32'b11111111111111110111011001001000;
assign LUT_2[28524] = 32'b11111111111111110000000101011011;
assign LUT_2[28525] = 32'b11111111111111101100111101110100;
assign LUT_2[28526] = 32'b11111111111111110110111110010111;
assign LUT_2[28527] = 32'b11111111111111110011110110110000;
assign LUT_2[28528] = 32'b11111111111111110011011010100000;
assign LUT_2[28529] = 32'b11111111111111110000010010111001;
assign LUT_2[28530] = 32'b11111111111111111010010011011100;
assign LUT_2[28531] = 32'b11111111111111110111001011110101;
assign LUT_2[28532] = 32'b11111111111111101111111000001000;
assign LUT_2[28533] = 32'b11111111111111101100110000100001;
assign LUT_2[28534] = 32'b11111111111111110110110001000100;
assign LUT_2[28535] = 32'b11111111111111110011101001011101;
assign LUT_2[28536] = 32'b11111111111111101110001011111101;
assign LUT_2[28537] = 32'b11111111111111101011000100010110;
assign LUT_2[28538] = 32'b11111111111111110101000100111001;
assign LUT_2[28539] = 32'b11111111111111110001111101010010;
assign LUT_2[28540] = 32'b11111111111111101010101001100101;
assign LUT_2[28541] = 32'b11111111111111100111100001111110;
assign LUT_2[28542] = 32'b11111111111111110001100010100001;
assign LUT_2[28543] = 32'b11111111111111101110011010111010;
assign LUT_2[28544] = 32'b00000000000000000100100110011001;
assign LUT_2[28545] = 32'b00000000000000000001011110110010;
assign LUT_2[28546] = 32'b00000000000000001011011111010101;
assign LUT_2[28547] = 32'b00000000000000001000010111101110;
assign LUT_2[28548] = 32'b00000000000000000001000100000001;
assign LUT_2[28549] = 32'b11111111111111111101111100011010;
assign LUT_2[28550] = 32'b00000000000000000111111100111101;
assign LUT_2[28551] = 32'b00000000000000000100110101010110;
assign LUT_2[28552] = 32'b11111111111111111111010111110110;
assign LUT_2[28553] = 32'b11111111111111111100010000001111;
assign LUT_2[28554] = 32'b00000000000000000110010000110010;
assign LUT_2[28555] = 32'b00000000000000000011001001001011;
assign LUT_2[28556] = 32'b11111111111111111011110101011110;
assign LUT_2[28557] = 32'b11111111111111111000101101110111;
assign LUT_2[28558] = 32'b00000000000000000010101110011010;
assign LUT_2[28559] = 32'b11111111111111111111100110110011;
assign LUT_2[28560] = 32'b11111111111111111111001010100011;
assign LUT_2[28561] = 32'b11111111111111111100000010111100;
assign LUT_2[28562] = 32'b00000000000000000110000011011111;
assign LUT_2[28563] = 32'b00000000000000000010111011111000;
assign LUT_2[28564] = 32'b11111111111111111011101000001011;
assign LUT_2[28565] = 32'b11111111111111111000100000100100;
assign LUT_2[28566] = 32'b00000000000000000010100001000111;
assign LUT_2[28567] = 32'b11111111111111111111011001100000;
assign LUT_2[28568] = 32'b11111111111111111001111100000000;
assign LUT_2[28569] = 32'b11111111111111110110110100011001;
assign LUT_2[28570] = 32'b00000000000000000000110100111100;
assign LUT_2[28571] = 32'b11111111111111111101101101010101;
assign LUT_2[28572] = 32'b11111111111111110110011001101000;
assign LUT_2[28573] = 32'b11111111111111110011010010000001;
assign LUT_2[28574] = 32'b11111111111111111101010010100100;
assign LUT_2[28575] = 32'b11111111111111111010001010111101;
assign LUT_2[28576] = 32'b00000000000000000101000010000010;
assign LUT_2[28577] = 32'b00000000000000000001111010011011;
assign LUT_2[28578] = 32'b00000000000000001011111010111110;
assign LUT_2[28579] = 32'b00000000000000001000110011010111;
assign LUT_2[28580] = 32'b00000000000000000001011111101010;
assign LUT_2[28581] = 32'b11111111111111111110011000000011;
assign LUT_2[28582] = 32'b00000000000000001000011000100110;
assign LUT_2[28583] = 32'b00000000000000000101010000111111;
assign LUT_2[28584] = 32'b11111111111111111111110011011111;
assign LUT_2[28585] = 32'b11111111111111111100101011111000;
assign LUT_2[28586] = 32'b00000000000000000110101100011011;
assign LUT_2[28587] = 32'b00000000000000000011100100110100;
assign LUT_2[28588] = 32'b11111111111111111100010001000111;
assign LUT_2[28589] = 32'b11111111111111111001001001100000;
assign LUT_2[28590] = 32'b00000000000000000011001010000011;
assign LUT_2[28591] = 32'b00000000000000000000000010011100;
assign LUT_2[28592] = 32'b11111111111111111111100110001100;
assign LUT_2[28593] = 32'b11111111111111111100011110100101;
assign LUT_2[28594] = 32'b00000000000000000110011111001000;
assign LUT_2[28595] = 32'b00000000000000000011010111100001;
assign LUT_2[28596] = 32'b11111111111111111100000011110100;
assign LUT_2[28597] = 32'b11111111111111111000111100001101;
assign LUT_2[28598] = 32'b00000000000000000010111100110000;
assign LUT_2[28599] = 32'b11111111111111111111110101001001;
assign LUT_2[28600] = 32'b11111111111111111010010111101001;
assign LUT_2[28601] = 32'b11111111111111110111010000000010;
assign LUT_2[28602] = 32'b00000000000000000001010000100101;
assign LUT_2[28603] = 32'b11111111111111111110001000111110;
assign LUT_2[28604] = 32'b11111111111111110110110101010001;
assign LUT_2[28605] = 32'b11111111111111110011101101101010;
assign LUT_2[28606] = 32'b11111111111111111101101110001101;
assign LUT_2[28607] = 32'b11111111111111111010100110100110;
assign LUT_2[28608] = 32'b11111111111111111100101110111100;
assign LUT_2[28609] = 32'b11111111111111111001100111010101;
assign LUT_2[28610] = 32'b00000000000000000011100111111000;
assign LUT_2[28611] = 32'b00000000000000000000100000010001;
assign LUT_2[28612] = 32'b11111111111111111001001100100100;
assign LUT_2[28613] = 32'b11111111111111110110000100111101;
assign LUT_2[28614] = 32'b00000000000000000000000101100000;
assign LUT_2[28615] = 32'b11111111111111111100111101111001;
assign LUT_2[28616] = 32'b11111111111111110111100000011001;
assign LUT_2[28617] = 32'b11111111111111110100011000110010;
assign LUT_2[28618] = 32'b11111111111111111110011001010101;
assign LUT_2[28619] = 32'b11111111111111111011010001101110;
assign LUT_2[28620] = 32'b11111111111111110011111110000001;
assign LUT_2[28621] = 32'b11111111111111110000110110011010;
assign LUT_2[28622] = 32'b11111111111111111010110110111101;
assign LUT_2[28623] = 32'b11111111111111110111101111010110;
assign LUT_2[28624] = 32'b11111111111111110111010011000110;
assign LUT_2[28625] = 32'b11111111111111110100001011011111;
assign LUT_2[28626] = 32'b11111111111111111110001100000010;
assign LUT_2[28627] = 32'b11111111111111111011000100011011;
assign LUT_2[28628] = 32'b11111111111111110011110000101110;
assign LUT_2[28629] = 32'b11111111111111110000101001000111;
assign LUT_2[28630] = 32'b11111111111111111010101001101010;
assign LUT_2[28631] = 32'b11111111111111110111100010000011;
assign LUT_2[28632] = 32'b11111111111111110010000100100011;
assign LUT_2[28633] = 32'b11111111111111101110111100111100;
assign LUT_2[28634] = 32'b11111111111111111000111101011111;
assign LUT_2[28635] = 32'b11111111111111110101110101111000;
assign LUT_2[28636] = 32'b11111111111111101110100010001011;
assign LUT_2[28637] = 32'b11111111111111101011011010100100;
assign LUT_2[28638] = 32'b11111111111111110101011011000111;
assign LUT_2[28639] = 32'b11111111111111110010010011100000;
assign LUT_2[28640] = 32'b11111111111111111101001010100101;
assign LUT_2[28641] = 32'b11111111111111111010000010111110;
assign LUT_2[28642] = 32'b00000000000000000100000011100001;
assign LUT_2[28643] = 32'b00000000000000000000111011111010;
assign LUT_2[28644] = 32'b11111111111111111001101000001101;
assign LUT_2[28645] = 32'b11111111111111110110100000100110;
assign LUT_2[28646] = 32'b00000000000000000000100001001001;
assign LUT_2[28647] = 32'b11111111111111111101011001100010;
assign LUT_2[28648] = 32'b11111111111111110111111100000010;
assign LUT_2[28649] = 32'b11111111111111110100110100011011;
assign LUT_2[28650] = 32'b11111111111111111110110100111110;
assign LUT_2[28651] = 32'b11111111111111111011101101010111;
assign LUT_2[28652] = 32'b11111111111111110100011001101010;
assign LUT_2[28653] = 32'b11111111111111110001010010000011;
assign LUT_2[28654] = 32'b11111111111111111011010010100110;
assign LUT_2[28655] = 32'b11111111111111111000001010111111;
assign LUT_2[28656] = 32'b11111111111111110111101110101111;
assign LUT_2[28657] = 32'b11111111111111110100100111001000;
assign LUT_2[28658] = 32'b11111111111111111110100111101011;
assign LUT_2[28659] = 32'b11111111111111111011100000000100;
assign LUT_2[28660] = 32'b11111111111111110100001100010111;
assign LUT_2[28661] = 32'b11111111111111110001000100110000;
assign LUT_2[28662] = 32'b11111111111111111011000101010011;
assign LUT_2[28663] = 32'b11111111111111110111111101101100;
assign LUT_2[28664] = 32'b11111111111111110010100000001100;
assign LUT_2[28665] = 32'b11111111111111101111011000100101;
assign LUT_2[28666] = 32'b11111111111111111001011001001000;
assign LUT_2[28667] = 32'b11111111111111110110010001100001;
assign LUT_2[28668] = 32'b11111111111111101110111101110100;
assign LUT_2[28669] = 32'b11111111111111101011110110001101;
assign LUT_2[28670] = 32'b11111111111111110101110110110000;
assign LUT_2[28671] = 32'b11111111111111110010101111001001;
assign LUT_2[28672] = 32'b11111111111111110100000011111100;
assign LUT_2[28673] = 32'b11111111111111110000111100010101;
assign LUT_2[28674] = 32'b11111111111111111010111100111000;
assign LUT_2[28675] = 32'b11111111111111110111110101010001;
assign LUT_2[28676] = 32'b11111111111111110000100001100100;
assign LUT_2[28677] = 32'b11111111111111101101011001111101;
assign LUT_2[28678] = 32'b11111111111111110111011010100000;
assign LUT_2[28679] = 32'b11111111111111110100010010111001;
assign LUT_2[28680] = 32'b11111111111111101110110101011001;
assign LUT_2[28681] = 32'b11111111111111101011101101110010;
assign LUT_2[28682] = 32'b11111111111111110101101110010101;
assign LUT_2[28683] = 32'b11111111111111110010100110101110;
assign LUT_2[28684] = 32'b11111111111111101011010011000001;
assign LUT_2[28685] = 32'b11111111111111101000001011011010;
assign LUT_2[28686] = 32'b11111111111111110010001011111101;
assign LUT_2[28687] = 32'b11111111111111101111000100010110;
assign LUT_2[28688] = 32'b11111111111111101110101000000110;
assign LUT_2[28689] = 32'b11111111111111101011100000011111;
assign LUT_2[28690] = 32'b11111111111111110101100001000010;
assign LUT_2[28691] = 32'b11111111111111110010011001011011;
assign LUT_2[28692] = 32'b11111111111111101011000101101110;
assign LUT_2[28693] = 32'b11111111111111100111111110000111;
assign LUT_2[28694] = 32'b11111111111111110001111110101010;
assign LUT_2[28695] = 32'b11111111111111101110110111000011;
assign LUT_2[28696] = 32'b11111111111111101001011001100011;
assign LUT_2[28697] = 32'b11111111111111100110010001111100;
assign LUT_2[28698] = 32'b11111111111111110000010010011111;
assign LUT_2[28699] = 32'b11111111111111101101001010111000;
assign LUT_2[28700] = 32'b11111111111111100101110111001011;
assign LUT_2[28701] = 32'b11111111111111100010101111100100;
assign LUT_2[28702] = 32'b11111111111111101100110000000111;
assign LUT_2[28703] = 32'b11111111111111101001101000100000;
assign LUT_2[28704] = 32'b11111111111111110100011111100101;
assign LUT_2[28705] = 32'b11111111111111110001010111111110;
assign LUT_2[28706] = 32'b11111111111111111011011000100001;
assign LUT_2[28707] = 32'b11111111111111111000010000111010;
assign LUT_2[28708] = 32'b11111111111111110000111101001101;
assign LUT_2[28709] = 32'b11111111111111101101110101100110;
assign LUT_2[28710] = 32'b11111111111111110111110110001001;
assign LUT_2[28711] = 32'b11111111111111110100101110100010;
assign LUT_2[28712] = 32'b11111111111111101111010001000010;
assign LUT_2[28713] = 32'b11111111111111101100001001011011;
assign LUT_2[28714] = 32'b11111111111111110110001001111110;
assign LUT_2[28715] = 32'b11111111111111110011000010010111;
assign LUT_2[28716] = 32'b11111111111111101011101110101010;
assign LUT_2[28717] = 32'b11111111111111101000100111000011;
assign LUT_2[28718] = 32'b11111111111111110010100111100110;
assign LUT_2[28719] = 32'b11111111111111101111011111111111;
assign LUT_2[28720] = 32'b11111111111111101111000011101111;
assign LUT_2[28721] = 32'b11111111111111101011111100001000;
assign LUT_2[28722] = 32'b11111111111111110101111100101011;
assign LUT_2[28723] = 32'b11111111111111110010110101000100;
assign LUT_2[28724] = 32'b11111111111111101011100001010111;
assign LUT_2[28725] = 32'b11111111111111101000011001110000;
assign LUT_2[28726] = 32'b11111111111111110010011010010011;
assign LUT_2[28727] = 32'b11111111111111101111010010101100;
assign LUT_2[28728] = 32'b11111111111111101001110101001100;
assign LUT_2[28729] = 32'b11111111111111100110101101100101;
assign LUT_2[28730] = 32'b11111111111111110000101110001000;
assign LUT_2[28731] = 32'b11111111111111101101100110100001;
assign LUT_2[28732] = 32'b11111111111111100110010010110100;
assign LUT_2[28733] = 32'b11111111111111100011001011001101;
assign LUT_2[28734] = 32'b11111111111111101101001011110000;
assign LUT_2[28735] = 32'b11111111111111101010000100001001;
assign LUT_2[28736] = 32'b11111111111111101100001100011111;
assign LUT_2[28737] = 32'b11111111111111101001000100111000;
assign LUT_2[28738] = 32'b11111111111111110011000101011011;
assign LUT_2[28739] = 32'b11111111111111101111111101110100;
assign LUT_2[28740] = 32'b11111111111111101000101010000111;
assign LUT_2[28741] = 32'b11111111111111100101100010100000;
assign LUT_2[28742] = 32'b11111111111111101111100011000011;
assign LUT_2[28743] = 32'b11111111111111101100011011011100;
assign LUT_2[28744] = 32'b11111111111111100110111101111100;
assign LUT_2[28745] = 32'b11111111111111100011110110010101;
assign LUT_2[28746] = 32'b11111111111111101101110110111000;
assign LUT_2[28747] = 32'b11111111111111101010101111010001;
assign LUT_2[28748] = 32'b11111111111111100011011011100100;
assign LUT_2[28749] = 32'b11111111111111100000010011111101;
assign LUT_2[28750] = 32'b11111111111111101010010100100000;
assign LUT_2[28751] = 32'b11111111111111100111001100111001;
assign LUT_2[28752] = 32'b11111111111111100110110000101001;
assign LUT_2[28753] = 32'b11111111111111100011101001000010;
assign LUT_2[28754] = 32'b11111111111111101101101001100101;
assign LUT_2[28755] = 32'b11111111111111101010100001111110;
assign LUT_2[28756] = 32'b11111111111111100011001110010001;
assign LUT_2[28757] = 32'b11111111111111100000000110101010;
assign LUT_2[28758] = 32'b11111111111111101010000111001101;
assign LUT_2[28759] = 32'b11111111111111100110111111100110;
assign LUT_2[28760] = 32'b11111111111111100001100010000110;
assign LUT_2[28761] = 32'b11111111111111011110011010011111;
assign LUT_2[28762] = 32'b11111111111111101000011011000010;
assign LUT_2[28763] = 32'b11111111111111100101010011011011;
assign LUT_2[28764] = 32'b11111111111111011101111111101110;
assign LUT_2[28765] = 32'b11111111111111011010111000000111;
assign LUT_2[28766] = 32'b11111111111111100100111000101010;
assign LUT_2[28767] = 32'b11111111111111100001110001000011;
assign LUT_2[28768] = 32'b11111111111111101100101000001000;
assign LUT_2[28769] = 32'b11111111111111101001100000100001;
assign LUT_2[28770] = 32'b11111111111111110011100001000100;
assign LUT_2[28771] = 32'b11111111111111110000011001011101;
assign LUT_2[28772] = 32'b11111111111111101001000101110000;
assign LUT_2[28773] = 32'b11111111111111100101111110001001;
assign LUT_2[28774] = 32'b11111111111111101111111110101100;
assign LUT_2[28775] = 32'b11111111111111101100110111000101;
assign LUT_2[28776] = 32'b11111111111111100111011001100101;
assign LUT_2[28777] = 32'b11111111111111100100010001111110;
assign LUT_2[28778] = 32'b11111111111111101110010010100001;
assign LUT_2[28779] = 32'b11111111111111101011001010111010;
assign LUT_2[28780] = 32'b11111111111111100011110111001101;
assign LUT_2[28781] = 32'b11111111111111100000101111100110;
assign LUT_2[28782] = 32'b11111111111111101010110000001001;
assign LUT_2[28783] = 32'b11111111111111100111101000100010;
assign LUT_2[28784] = 32'b11111111111111100111001100010010;
assign LUT_2[28785] = 32'b11111111111111100100000100101011;
assign LUT_2[28786] = 32'b11111111111111101110000101001110;
assign LUT_2[28787] = 32'b11111111111111101010111101100111;
assign LUT_2[28788] = 32'b11111111111111100011101001111010;
assign LUT_2[28789] = 32'b11111111111111100000100010010011;
assign LUT_2[28790] = 32'b11111111111111101010100010110110;
assign LUT_2[28791] = 32'b11111111111111100111011011001111;
assign LUT_2[28792] = 32'b11111111111111100001111101101111;
assign LUT_2[28793] = 32'b11111111111111011110110110001000;
assign LUT_2[28794] = 32'b11111111111111101000110110101011;
assign LUT_2[28795] = 32'b11111111111111100101101111000100;
assign LUT_2[28796] = 32'b11111111111111011110011011010111;
assign LUT_2[28797] = 32'b11111111111111011011010011110000;
assign LUT_2[28798] = 32'b11111111111111100101010100010011;
assign LUT_2[28799] = 32'b11111111111111100010001100101100;
assign LUT_2[28800] = 32'b11111111111111111000011000001011;
assign LUT_2[28801] = 32'b11111111111111110101010000100100;
assign LUT_2[28802] = 32'b11111111111111111111010001000111;
assign LUT_2[28803] = 32'b11111111111111111100001001100000;
assign LUT_2[28804] = 32'b11111111111111110100110101110011;
assign LUT_2[28805] = 32'b11111111111111110001101110001100;
assign LUT_2[28806] = 32'b11111111111111111011101110101111;
assign LUT_2[28807] = 32'b11111111111111111000100111001000;
assign LUT_2[28808] = 32'b11111111111111110011001001101000;
assign LUT_2[28809] = 32'b11111111111111110000000010000001;
assign LUT_2[28810] = 32'b11111111111111111010000010100100;
assign LUT_2[28811] = 32'b11111111111111110110111010111101;
assign LUT_2[28812] = 32'b11111111111111101111100111010000;
assign LUT_2[28813] = 32'b11111111111111101100011111101001;
assign LUT_2[28814] = 32'b11111111111111110110100000001100;
assign LUT_2[28815] = 32'b11111111111111110011011000100101;
assign LUT_2[28816] = 32'b11111111111111110010111100010101;
assign LUT_2[28817] = 32'b11111111111111101111110100101110;
assign LUT_2[28818] = 32'b11111111111111111001110101010001;
assign LUT_2[28819] = 32'b11111111111111110110101101101010;
assign LUT_2[28820] = 32'b11111111111111101111011001111101;
assign LUT_2[28821] = 32'b11111111111111101100010010010110;
assign LUT_2[28822] = 32'b11111111111111110110010010111001;
assign LUT_2[28823] = 32'b11111111111111110011001011010010;
assign LUT_2[28824] = 32'b11111111111111101101101101110010;
assign LUT_2[28825] = 32'b11111111111111101010100110001011;
assign LUT_2[28826] = 32'b11111111111111110100100110101110;
assign LUT_2[28827] = 32'b11111111111111110001011111000111;
assign LUT_2[28828] = 32'b11111111111111101010001011011010;
assign LUT_2[28829] = 32'b11111111111111100111000011110011;
assign LUT_2[28830] = 32'b11111111111111110001000100010110;
assign LUT_2[28831] = 32'b11111111111111101101111100101111;
assign LUT_2[28832] = 32'b11111111111111111000110011110100;
assign LUT_2[28833] = 32'b11111111111111110101101100001101;
assign LUT_2[28834] = 32'b11111111111111111111101100110000;
assign LUT_2[28835] = 32'b11111111111111111100100101001001;
assign LUT_2[28836] = 32'b11111111111111110101010001011100;
assign LUT_2[28837] = 32'b11111111111111110010001001110101;
assign LUT_2[28838] = 32'b11111111111111111100001010011000;
assign LUT_2[28839] = 32'b11111111111111111001000010110001;
assign LUT_2[28840] = 32'b11111111111111110011100101010001;
assign LUT_2[28841] = 32'b11111111111111110000011101101010;
assign LUT_2[28842] = 32'b11111111111111111010011110001101;
assign LUT_2[28843] = 32'b11111111111111110111010110100110;
assign LUT_2[28844] = 32'b11111111111111110000000010111001;
assign LUT_2[28845] = 32'b11111111111111101100111011010010;
assign LUT_2[28846] = 32'b11111111111111110110111011110101;
assign LUT_2[28847] = 32'b11111111111111110011110100001110;
assign LUT_2[28848] = 32'b11111111111111110011010111111110;
assign LUT_2[28849] = 32'b11111111111111110000010000010111;
assign LUT_2[28850] = 32'b11111111111111111010010000111010;
assign LUT_2[28851] = 32'b11111111111111110111001001010011;
assign LUT_2[28852] = 32'b11111111111111101111110101100110;
assign LUT_2[28853] = 32'b11111111111111101100101101111111;
assign LUT_2[28854] = 32'b11111111111111110110101110100010;
assign LUT_2[28855] = 32'b11111111111111110011100110111011;
assign LUT_2[28856] = 32'b11111111111111101110001001011011;
assign LUT_2[28857] = 32'b11111111111111101011000001110100;
assign LUT_2[28858] = 32'b11111111111111110101000010010111;
assign LUT_2[28859] = 32'b11111111111111110001111010110000;
assign LUT_2[28860] = 32'b11111111111111101010100111000011;
assign LUT_2[28861] = 32'b11111111111111100111011111011100;
assign LUT_2[28862] = 32'b11111111111111110001011111111111;
assign LUT_2[28863] = 32'b11111111111111101110011000011000;
assign LUT_2[28864] = 32'b11111111111111110000100000101110;
assign LUT_2[28865] = 32'b11111111111111101101011001000111;
assign LUT_2[28866] = 32'b11111111111111110111011001101010;
assign LUT_2[28867] = 32'b11111111111111110100010010000011;
assign LUT_2[28868] = 32'b11111111111111101100111110010110;
assign LUT_2[28869] = 32'b11111111111111101001110110101111;
assign LUT_2[28870] = 32'b11111111111111110011110111010010;
assign LUT_2[28871] = 32'b11111111111111110000101111101011;
assign LUT_2[28872] = 32'b11111111111111101011010010001011;
assign LUT_2[28873] = 32'b11111111111111101000001010100100;
assign LUT_2[28874] = 32'b11111111111111110010001011000111;
assign LUT_2[28875] = 32'b11111111111111101111000011100000;
assign LUT_2[28876] = 32'b11111111111111100111101111110011;
assign LUT_2[28877] = 32'b11111111111111100100101000001100;
assign LUT_2[28878] = 32'b11111111111111101110101000101111;
assign LUT_2[28879] = 32'b11111111111111101011100001001000;
assign LUT_2[28880] = 32'b11111111111111101011000100111000;
assign LUT_2[28881] = 32'b11111111111111100111111101010001;
assign LUT_2[28882] = 32'b11111111111111110001111101110100;
assign LUT_2[28883] = 32'b11111111111111101110110110001101;
assign LUT_2[28884] = 32'b11111111111111100111100010100000;
assign LUT_2[28885] = 32'b11111111111111100100011010111001;
assign LUT_2[28886] = 32'b11111111111111101110011011011100;
assign LUT_2[28887] = 32'b11111111111111101011010011110101;
assign LUT_2[28888] = 32'b11111111111111100101110110010101;
assign LUT_2[28889] = 32'b11111111111111100010101110101110;
assign LUT_2[28890] = 32'b11111111111111101100101111010001;
assign LUT_2[28891] = 32'b11111111111111101001100111101010;
assign LUT_2[28892] = 32'b11111111111111100010010011111101;
assign LUT_2[28893] = 32'b11111111111111011111001100010110;
assign LUT_2[28894] = 32'b11111111111111101001001100111001;
assign LUT_2[28895] = 32'b11111111111111100110000101010010;
assign LUT_2[28896] = 32'b11111111111111110000111100010111;
assign LUT_2[28897] = 32'b11111111111111101101110100110000;
assign LUT_2[28898] = 32'b11111111111111110111110101010011;
assign LUT_2[28899] = 32'b11111111111111110100101101101100;
assign LUT_2[28900] = 32'b11111111111111101101011001111111;
assign LUT_2[28901] = 32'b11111111111111101010010010011000;
assign LUT_2[28902] = 32'b11111111111111110100010010111011;
assign LUT_2[28903] = 32'b11111111111111110001001011010100;
assign LUT_2[28904] = 32'b11111111111111101011101101110100;
assign LUT_2[28905] = 32'b11111111111111101000100110001101;
assign LUT_2[28906] = 32'b11111111111111110010100110110000;
assign LUT_2[28907] = 32'b11111111111111101111011111001001;
assign LUT_2[28908] = 32'b11111111111111101000001011011100;
assign LUT_2[28909] = 32'b11111111111111100101000011110101;
assign LUT_2[28910] = 32'b11111111111111101111000100011000;
assign LUT_2[28911] = 32'b11111111111111101011111100110001;
assign LUT_2[28912] = 32'b11111111111111101011100000100001;
assign LUT_2[28913] = 32'b11111111111111101000011000111010;
assign LUT_2[28914] = 32'b11111111111111110010011001011101;
assign LUT_2[28915] = 32'b11111111111111101111010001110110;
assign LUT_2[28916] = 32'b11111111111111100111111110001001;
assign LUT_2[28917] = 32'b11111111111111100100110110100010;
assign LUT_2[28918] = 32'b11111111111111101110110111000101;
assign LUT_2[28919] = 32'b11111111111111101011101111011110;
assign LUT_2[28920] = 32'b11111111111111100110010001111110;
assign LUT_2[28921] = 32'b11111111111111100011001010010111;
assign LUT_2[28922] = 32'b11111111111111101101001010111010;
assign LUT_2[28923] = 32'b11111111111111101010000011010011;
assign LUT_2[28924] = 32'b11111111111111100010101111100110;
assign LUT_2[28925] = 32'b11111111111111011111100111111111;
assign LUT_2[28926] = 32'b11111111111111101001101000100010;
assign LUT_2[28927] = 32'b11111111111111100110100000111011;
assign LUT_2[28928] = 32'b11111111111111111000000010100010;
assign LUT_2[28929] = 32'b11111111111111110100111010111011;
assign LUT_2[28930] = 32'b11111111111111111110111011011110;
assign LUT_2[28931] = 32'b11111111111111111011110011110111;
assign LUT_2[28932] = 32'b11111111111111110100100000001010;
assign LUT_2[28933] = 32'b11111111111111110001011000100011;
assign LUT_2[28934] = 32'b11111111111111111011011001000110;
assign LUT_2[28935] = 32'b11111111111111111000010001011111;
assign LUT_2[28936] = 32'b11111111111111110010110011111111;
assign LUT_2[28937] = 32'b11111111111111101111101100011000;
assign LUT_2[28938] = 32'b11111111111111111001101100111011;
assign LUT_2[28939] = 32'b11111111111111110110100101010100;
assign LUT_2[28940] = 32'b11111111111111101111010001100111;
assign LUT_2[28941] = 32'b11111111111111101100001010000000;
assign LUT_2[28942] = 32'b11111111111111110110001010100011;
assign LUT_2[28943] = 32'b11111111111111110011000010111100;
assign LUT_2[28944] = 32'b11111111111111110010100110101100;
assign LUT_2[28945] = 32'b11111111111111101111011111000101;
assign LUT_2[28946] = 32'b11111111111111111001011111101000;
assign LUT_2[28947] = 32'b11111111111111110110011000000001;
assign LUT_2[28948] = 32'b11111111111111101111000100010100;
assign LUT_2[28949] = 32'b11111111111111101011111100101101;
assign LUT_2[28950] = 32'b11111111111111110101111101010000;
assign LUT_2[28951] = 32'b11111111111111110010110101101001;
assign LUT_2[28952] = 32'b11111111111111101101011000001001;
assign LUT_2[28953] = 32'b11111111111111101010010000100010;
assign LUT_2[28954] = 32'b11111111111111110100010001000101;
assign LUT_2[28955] = 32'b11111111111111110001001001011110;
assign LUT_2[28956] = 32'b11111111111111101001110101110001;
assign LUT_2[28957] = 32'b11111111111111100110101110001010;
assign LUT_2[28958] = 32'b11111111111111110000101110101101;
assign LUT_2[28959] = 32'b11111111111111101101100111000110;
assign LUT_2[28960] = 32'b11111111111111111000011110001011;
assign LUT_2[28961] = 32'b11111111111111110101010110100100;
assign LUT_2[28962] = 32'b11111111111111111111010111000111;
assign LUT_2[28963] = 32'b11111111111111111100001111100000;
assign LUT_2[28964] = 32'b11111111111111110100111011110011;
assign LUT_2[28965] = 32'b11111111111111110001110100001100;
assign LUT_2[28966] = 32'b11111111111111111011110100101111;
assign LUT_2[28967] = 32'b11111111111111111000101101001000;
assign LUT_2[28968] = 32'b11111111111111110011001111101000;
assign LUT_2[28969] = 32'b11111111111111110000001000000001;
assign LUT_2[28970] = 32'b11111111111111111010001000100100;
assign LUT_2[28971] = 32'b11111111111111110111000000111101;
assign LUT_2[28972] = 32'b11111111111111101111101101010000;
assign LUT_2[28973] = 32'b11111111111111101100100101101001;
assign LUT_2[28974] = 32'b11111111111111110110100110001100;
assign LUT_2[28975] = 32'b11111111111111110011011110100101;
assign LUT_2[28976] = 32'b11111111111111110011000010010101;
assign LUT_2[28977] = 32'b11111111111111101111111010101110;
assign LUT_2[28978] = 32'b11111111111111111001111011010001;
assign LUT_2[28979] = 32'b11111111111111110110110011101010;
assign LUT_2[28980] = 32'b11111111111111101111011111111101;
assign LUT_2[28981] = 32'b11111111111111101100011000010110;
assign LUT_2[28982] = 32'b11111111111111110110011000111001;
assign LUT_2[28983] = 32'b11111111111111110011010001010010;
assign LUT_2[28984] = 32'b11111111111111101101110011110010;
assign LUT_2[28985] = 32'b11111111111111101010101100001011;
assign LUT_2[28986] = 32'b11111111111111110100101100101110;
assign LUT_2[28987] = 32'b11111111111111110001100101000111;
assign LUT_2[28988] = 32'b11111111111111101010010001011010;
assign LUT_2[28989] = 32'b11111111111111100111001001110011;
assign LUT_2[28990] = 32'b11111111111111110001001010010110;
assign LUT_2[28991] = 32'b11111111111111101110000010101111;
assign LUT_2[28992] = 32'b11111111111111110000001011000101;
assign LUT_2[28993] = 32'b11111111111111101101000011011110;
assign LUT_2[28994] = 32'b11111111111111110111000100000001;
assign LUT_2[28995] = 32'b11111111111111110011111100011010;
assign LUT_2[28996] = 32'b11111111111111101100101000101101;
assign LUT_2[28997] = 32'b11111111111111101001100001000110;
assign LUT_2[28998] = 32'b11111111111111110011100001101001;
assign LUT_2[28999] = 32'b11111111111111110000011010000010;
assign LUT_2[29000] = 32'b11111111111111101010111100100010;
assign LUT_2[29001] = 32'b11111111111111100111110100111011;
assign LUT_2[29002] = 32'b11111111111111110001110101011110;
assign LUT_2[29003] = 32'b11111111111111101110101101110111;
assign LUT_2[29004] = 32'b11111111111111100111011010001010;
assign LUT_2[29005] = 32'b11111111111111100100010010100011;
assign LUT_2[29006] = 32'b11111111111111101110010011000110;
assign LUT_2[29007] = 32'b11111111111111101011001011011111;
assign LUT_2[29008] = 32'b11111111111111101010101111001111;
assign LUT_2[29009] = 32'b11111111111111100111100111101000;
assign LUT_2[29010] = 32'b11111111111111110001101000001011;
assign LUT_2[29011] = 32'b11111111111111101110100000100100;
assign LUT_2[29012] = 32'b11111111111111100111001100110111;
assign LUT_2[29013] = 32'b11111111111111100100000101010000;
assign LUT_2[29014] = 32'b11111111111111101110000101110011;
assign LUT_2[29015] = 32'b11111111111111101010111110001100;
assign LUT_2[29016] = 32'b11111111111111100101100000101100;
assign LUT_2[29017] = 32'b11111111111111100010011001000101;
assign LUT_2[29018] = 32'b11111111111111101100011001101000;
assign LUT_2[29019] = 32'b11111111111111101001010010000001;
assign LUT_2[29020] = 32'b11111111111111100001111110010100;
assign LUT_2[29021] = 32'b11111111111111011110110110101101;
assign LUT_2[29022] = 32'b11111111111111101000110111010000;
assign LUT_2[29023] = 32'b11111111111111100101101111101001;
assign LUT_2[29024] = 32'b11111111111111110000100110101110;
assign LUT_2[29025] = 32'b11111111111111101101011111000111;
assign LUT_2[29026] = 32'b11111111111111110111011111101010;
assign LUT_2[29027] = 32'b11111111111111110100011000000011;
assign LUT_2[29028] = 32'b11111111111111101101000100010110;
assign LUT_2[29029] = 32'b11111111111111101001111100101111;
assign LUT_2[29030] = 32'b11111111111111110011111101010010;
assign LUT_2[29031] = 32'b11111111111111110000110101101011;
assign LUT_2[29032] = 32'b11111111111111101011011000001011;
assign LUT_2[29033] = 32'b11111111111111101000010000100100;
assign LUT_2[29034] = 32'b11111111111111110010010001000111;
assign LUT_2[29035] = 32'b11111111111111101111001001100000;
assign LUT_2[29036] = 32'b11111111111111100111110101110011;
assign LUT_2[29037] = 32'b11111111111111100100101110001100;
assign LUT_2[29038] = 32'b11111111111111101110101110101111;
assign LUT_2[29039] = 32'b11111111111111101011100111001000;
assign LUT_2[29040] = 32'b11111111111111101011001010111000;
assign LUT_2[29041] = 32'b11111111111111101000000011010001;
assign LUT_2[29042] = 32'b11111111111111110010000011110100;
assign LUT_2[29043] = 32'b11111111111111101110111100001101;
assign LUT_2[29044] = 32'b11111111111111100111101000100000;
assign LUT_2[29045] = 32'b11111111111111100100100000111001;
assign LUT_2[29046] = 32'b11111111111111101110100001011100;
assign LUT_2[29047] = 32'b11111111111111101011011001110101;
assign LUT_2[29048] = 32'b11111111111111100101111100010101;
assign LUT_2[29049] = 32'b11111111111111100010110100101110;
assign LUT_2[29050] = 32'b11111111111111101100110101010001;
assign LUT_2[29051] = 32'b11111111111111101001101101101010;
assign LUT_2[29052] = 32'b11111111111111100010011001111101;
assign LUT_2[29053] = 32'b11111111111111011111010010010110;
assign LUT_2[29054] = 32'b11111111111111101001010010111001;
assign LUT_2[29055] = 32'b11111111111111100110001011010010;
assign LUT_2[29056] = 32'b11111111111111111100010110110001;
assign LUT_2[29057] = 32'b11111111111111111001001111001010;
assign LUT_2[29058] = 32'b00000000000000000011001111101101;
assign LUT_2[29059] = 32'b00000000000000000000001000000110;
assign LUT_2[29060] = 32'b11111111111111111000110100011001;
assign LUT_2[29061] = 32'b11111111111111110101101100110010;
assign LUT_2[29062] = 32'b11111111111111111111101101010101;
assign LUT_2[29063] = 32'b11111111111111111100100101101110;
assign LUT_2[29064] = 32'b11111111111111110111001000001110;
assign LUT_2[29065] = 32'b11111111111111110100000000100111;
assign LUT_2[29066] = 32'b11111111111111111110000001001010;
assign LUT_2[29067] = 32'b11111111111111111010111001100011;
assign LUT_2[29068] = 32'b11111111111111110011100101110110;
assign LUT_2[29069] = 32'b11111111111111110000011110001111;
assign LUT_2[29070] = 32'b11111111111111111010011110110010;
assign LUT_2[29071] = 32'b11111111111111110111010111001011;
assign LUT_2[29072] = 32'b11111111111111110110111010111011;
assign LUT_2[29073] = 32'b11111111111111110011110011010100;
assign LUT_2[29074] = 32'b11111111111111111101110011110111;
assign LUT_2[29075] = 32'b11111111111111111010101100010000;
assign LUT_2[29076] = 32'b11111111111111110011011000100011;
assign LUT_2[29077] = 32'b11111111111111110000010000111100;
assign LUT_2[29078] = 32'b11111111111111111010010001011111;
assign LUT_2[29079] = 32'b11111111111111110111001001111000;
assign LUT_2[29080] = 32'b11111111111111110001101100011000;
assign LUT_2[29081] = 32'b11111111111111101110100100110001;
assign LUT_2[29082] = 32'b11111111111111111000100101010100;
assign LUT_2[29083] = 32'b11111111111111110101011101101101;
assign LUT_2[29084] = 32'b11111111111111101110001010000000;
assign LUT_2[29085] = 32'b11111111111111101011000010011001;
assign LUT_2[29086] = 32'b11111111111111110101000010111100;
assign LUT_2[29087] = 32'b11111111111111110001111011010101;
assign LUT_2[29088] = 32'b11111111111111111100110010011010;
assign LUT_2[29089] = 32'b11111111111111111001101010110011;
assign LUT_2[29090] = 32'b00000000000000000011101011010110;
assign LUT_2[29091] = 32'b00000000000000000000100011101111;
assign LUT_2[29092] = 32'b11111111111111111001010000000010;
assign LUT_2[29093] = 32'b11111111111111110110001000011011;
assign LUT_2[29094] = 32'b00000000000000000000001000111110;
assign LUT_2[29095] = 32'b11111111111111111101000001010111;
assign LUT_2[29096] = 32'b11111111111111110111100011110111;
assign LUT_2[29097] = 32'b11111111111111110100011100010000;
assign LUT_2[29098] = 32'b11111111111111111110011100110011;
assign LUT_2[29099] = 32'b11111111111111111011010101001100;
assign LUT_2[29100] = 32'b11111111111111110100000001011111;
assign LUT_2[29101] = 32'b11111111111111110000111001111000;
assign LUT_2[29102] = 32'b11111111111111111010111010011011;
assign LUT_2[29103] = 32'b11111111111111110111110010110100;
assign LUT_2[29104] = 32'b11111111111111110111010110100100;
assign LUT_2[29105] = 32'b11111111111111110100001110111101;
assign LUT_2[29106] = 32'b11111111111111111110001111100000;
assign LUT_2[29107] = 32'b11111111111111111011000111111001;
assign LUT_2[29108] = 32'b11111111111111110011110100001100;
assign LUT_2[29109] = 32'b11111111111111110000101100100101;
assign LUT_2[29110] = 32'b11111111111111111010101101001000;
assign LUT_2[29111] = 32'b11111111111111110111100101100001;
assign LUT_2[29112] = 32'b11111111111111110010001000000001;
assign LUT_2[29113] = 32'b11111111111111101111000000011010;
assign LUT_2[29114] = 32'b11111111111111111001000000111101;
assign LUT_2[29115] = 32'b11111111111111110101111001010110;
assign LUT_2[29116] = 32'b11111111111111101110100101101001;
assign LUT_2[29117] = 32'b11111111111111101011011110000010;
assign LUT_2[29118] = 32'b11111111111111110101011110100101;
assign LUT_2[29119] = 32'b11111111111111110010010110111110;
assign LUT_2[29120] = 32'b11111111111111110100011111010100;
assign LUT_2[29121] = 32'b11111111111111110001010111101101;
assign LUT_2[29122] = 32'b11111111111111111011011000010000;
assign LUT_2[29123] = 32'b11111111111111111000010000101001;
assign LUT_2[29124] = 32'b11111111111111110000111100111100;
assign LUT_2[29125] = 32'b11111111111111101101110101010101;
assign LUT_2[29126] = 32'b11111111111111110111110101111000;
assign LUT_2[29127] = 32'b11111111111111110100101110010001;
assign LUT_2[29128] = 32'b11111111111111101111010000110001;
assign LUT_2[29129] = 32'b11111111111111101100001001001010;
assign LUT_2[29130] = 32'b11111111111111110110001001101101;
assign LUT_2[29131] = 32'b11111111111111110011000010000110;
assign LUT_2[29132] = 32'b11111111111111101011101110011001;
assign LUT_2[29133] = 32'b11111111111111101000100110110010;
assign LUT_2[29134] = 32'b11111111111111110010100111010101;
assign LUT_2[29135] = 32'b11111111111111101111011111101110;
assign LUT_2[29136] = 32'b11111111111111101111000011011110;
assign LUT_2[29137] = 32'b11111111111111101011111011110111;
assign LUT_2[29138] = 32'b11111111111111110101111100011010;
assign LUT_2[29139] = 32'b11111111111111110010110100110011;
assign LUT_2[29140] = 32'b11111111111111101011100001000110;
assign LUT_2[29141] = 32'b11111111111111101000011001011111;
assign LUT_2[29142] = 32'b11111111111111110010011010000010;
assign LUT_2[29143] = 32'b11111111111111101111010010011011;
assign LUT_2[29144] = 32'b11111111111111101001110100111011;
assign LUT_2[29145] = 32'b11111111111111100110101101010100;
assign LUT_2[29146] = 32'b11111111111111110000101101110111;
assign LUT_2[29147] = 32'b11111111111111101101100110010000;
assign LUT_2[29148] = 32'b11111111111111100110010010100011;
assign LUT_2[29149] = 32'b11111111111111100011001010111100;
assign LUT_2[29150] = 32'b11111111111111101101001011011111;
assign LUT_2[29151] = 32'b11111111111111101010000011111000;
assign LUT_2[29152] = 32'b11111111111111110100111010111101;
assign LUT_2[29153] = 32'b11111111111111110001110011010110;
assign LUT_2[29154] = 32'b11111111111111111011110011111001;
assign LUT_2[29155] = 32'b11111111111111111000101100010010;
assign LUT_2[29156] = 32'b11111111111111110001011000100101;
assign LUT_2[29157] = 32'b11111111111111101110010000111110;
assign LUT_2[29158] = 32'b11111111111111111000010001100001;
assign LUT_2[29159] = 32'b11111111111111110101001001111010;
assign LUT_2[29160] = 32'b11111111111111101111101100011010;
assign LUT_2[29161] = 32'b11111111111111101100100100110011;
assign LUT_2[29162] = 32'b11111111111111110110100101010110;
assign LUT_2[29163] = 32'b11111111111111110011011101101111;
assign LUT_2[29164] = 32'b11111111111111101100001010000010;
assign LUT_2[29165] = 32'b11111111111111101001000010011011;
assign LUT_2[29166] = 32'b11111111111111110011000010111110;
assign LUT_2[29167] = 32'b11111111111111101111111011010111;
assign LUT_2[29168] = 32'b11111111111111101111011111000111;
assign LUT_2[29169] = 32'b11111111111111101100010111100000;
assign LUT_2[29170] = 32'b11111111111111110110011000000011;
assign LUT_2[29171] = 32'b11111111111111110011010000011100;
assign LUT_2[29172] = 32'b11111111111111101011111100101111;
assign LUT_2[29173] = 32'b11111111111111101000110101001000;
assign LUT_2[29174] = 32'b11111111111111110010110101101011;
assign LUT_2[29175] = 32'b11111111111111101111101110000100;
assign LUT_2[29176] = 32'b11111111111111101010010000100100;
assign LUT_2[29177] = 32'b11111111111111100111001000111101;
assign LUT_2[29178] = 32'b11111111111111110001001001100000;
assign LUT_2[29179] = 32'b11111111111111101110000001111001;
assign LUT_2[29180] = 32'b11111111111111100110101110001100;
assign LUT_2[29181] = 32'b11111111111111100011100110100101;
assign LUT_2[29182] = 32'b11111111111111101101100111001000;
assign LUT_2[29183] = 32'b11111111111111101010011111100001;
assign LUT_2[29184] = 32'b11111111111111111000110101101110;
assign LUT_2[29185] = 32'b11111111111111110101101110000111;
assign LUT_2[29186] = 32'b11111111111111111111101110101010;
assign LUT_2[29187] = 32'b11111111111111111100100111000011;
assign LUT_2[29188] = 32'b11111111111111110101010011010110;
assign LUT_2[29189] = 32'b11111111111111110010001011101111;
assign LUT_2[29190] = 32'b11111111111111111100001100010010;
assign LUT_2[29191] = 32'b11111111111111111001000100101011;
assign LUT_2[29192] = 32'b11111111111111110011100111001011;
assign LUT_2[29193] = 32'b11111111111111110000011111100100;
assign LUT_2[29194] = 32'b11111111111111111010100000000111;
assign LUT_2[29195] = 32'b11111111111111110111011000100000;
assign LUT_2[29196] = 32'b11111111111111110000000100110011;
assign LUT_2[29197] = 32'b11111111111111101100111101001100;
assign LUT_2[29198] = 32'b11111111111111110110111101101111;
assign LUT_2[29199] = 32'b11111111111111110011110110001000;
assign LUT_2[29200] = 32'b11111111111111110011011001111000;
assign LUT_2[29201] = 32'b11111111111111110000010010010001;
assign LUT_2[29202] = 32'b11111111111111111010010010110100;
assign LUT_2[29203] = 32'b11111111111111110111001011001101;
assign LUT_2[29204] = 32'b11111111111111101111110111100000;
assign LUT_2[29205] = 32'b11111111111111101100101111111001;
assign LUT_2[29206] = 32'b11111111111111110110110000011100;
assign LUT_2[29207] = 32'b11111111111111110011101000110101;
assign LUT_2[29208] = 32'b11111111111111101110001011010101;
assign LUT_2[29209] = 32'b11111111111111101011000011101110;
assign LUT_2[29210] = 32'b11111111111111110101000100010001;
assign LUT_2[29211] = 32'b11111111111111110001111100101010;
assign LUT_2[29212] = 32'b11111111111111101010101000111101;
assign LUT_2[29213] = 32'b11111111111111100111100001010110;
assign LUT_2[29214] = 32'b11111111111111110001100001111001;
assign LUT_2[29215] = 32'b11111111111111101110011010010010;
assign LUT_2[29216] = 32'b11111111111111111001010001010111;
assign LUT_2[29217] = 32'b11111111111111110110001001110000;
assign LUT_2[29218] = 32'b00000000000000000000001010010011;
assign LUT_2[29219] = 32'b11111111111111111101000010101100;
assign LUT_2[29220] = 32'b11111111111111110101101110111111;
assign LUT_2[29221] = 32'b11111111111111110010100111011000;
assign LUT_2[29222] = 32'b11111111111111111100100111111011;
assign LUT_2[29223] = 32'b11111111111111111001100000010100;
assign LUT_2[29224] = 32'b11111111111111110100000010110100;
assign LUT_2[29225] = 32'b11111111111111110000111011001101;
assign LUT_2[29226] = 32'b11111111111111111010111011110000;
assign LUT_2[29227] = 32'b11111111111111110111110100001001;
assign LUT_2[29228] = 32'b11111111111111110000100000011100;
assign LUT_2[29229] = 32'b11111111111111101101011000110101;
assign LUT_2[29230] = 32'b11111111111111110111011001011000;
assign LUT_2[29231] = 32'b11111111111111110100010001110001;
assign LUT_2[29232] = 32'b11111111111111110011110101100001;
assign LUT_2[29233] = 32'b11111111111111110000101101111010;
assign LUT_2[29234] = 32'b11111111111111111010101110011101;
assign LUT_2[29235] = 32'b11111111111111110111100110110110;
assign LUT_2[29236] = 32'b11111111111111110000010011001001;
assign LUT_2[29237] = 32'b11111111111111101101001011100010;
assign LUT_2[29238] = 32'b11111111111111110111001100000101;
assign LUT_2[29239] = 32'b11111111111111110100000100011110;
assign LUT_2[29240] = 32'b11111111111111101110100110111110;
assign LUT_2[29241] = 32'b11111111111111101011011111010111;
assign LUT_2[29242] = 32'b11111111111111110101011111111010;
assign LUT_2[29243] = 32'b11111111111111110010011000010011;
assign LUT_2[29244] = 32'b11111111111111101011000100100110;
assign LUT_2[29245] = 32'b11111111111111100111111100111111;
assign LUT_2[29246] = 32'b11111111111111110001111101100010;
assign LUT_2[29247] = 32'b11111111111111101110110101111011;
assign LUT_2[29248] = 32'b11111111111111110000111110010001;
assign LUT_2[29249] = 32'b11111111111111101101110110101010;
assign LUT_2[29250] = 32'b11111111111111110111110111001101;
assign LUT_2[29251] = 32'b11111111111111110100101111100110;
assign LUT_2[29252] = 32'b11111111111111101101011011111001;
assign LUT_2[29253] = 32'b11111111111111101010010100010010;
assign LUT_2[29254] = 32'b11111111111111110100010100110101;
assign LUT_2[29255] = 32'b11111111111111110001001101001110;
assign LUT_2[29256] = 32'b11111111111111101011101111101110;
assign LUT_2[29257] = 32'b11111111111111101000101000000111;
assign LUT_2[29258] = 32'b11111111111111110010101000101010;
assign LUT_2[29259] = 32'b11111111111111101111100001000011;
assign LUT_2[29260] = 32'b11111111111111101000001101010110;
assign LUT_2[29261] = 32'b11111111111111100101000101101111;
assign LUT_2[29262] = 32'b11111111111111101111000110010010;
assign LUT_2[29263] = 32'b11111111111111101011111110101011;
assign LUT_2[29264] = 32'b11111111111111101011100010011011;
assign LUT_2[29265] = 32'b11111111111111101000011010110100;
assign LUT_2[29266] = 32'b11111111111111110010011011010111;
assign LUT_2[29267] = 32'b11111111111111101111010011110000;
assign LUT_2[29268] = 32'b11111111111111101000000000000011;
assign LUT_2[29269] = 32'b11111111111111100100111000011100;
assign LUT_2[29270] = 32'b11111111111111101110111000111111;
assign LUT_2[29271] = 32'b11111111111111101011110001011000;
assign LUT_2[29272] = 32'b11111111111111100110010011111000;
assign LUT_2[29273] = 32'b11111111111111100011001100010001;
assign LUT_2[29274] = 32'b11111111111111101101001100110100;
assign LUT_2[29275] = 32'b11111111111111101010000101001101;
assign LUT_2[29276] = 32'b11111111111111100010110001100000;
assign LUT_2[29277] = 32'b11111111111111011111101001111001;
assign LUT_2[29278] = 32'b11111111111111101001101010011100;
assign LUT_2[29279] = 32'b11111111111111100110100010110101;
assign LUT_2[29280] = 32'b11111111111111110001011001111010;
assign LUT_2[29281] = 32'b11111111111111101110010010010011;
assign LUT_2[29282] = 32'b11111111111111111000010010110110;
assign LUT_2[29283] = 32'b11111111111111110101001011001111;
assign LUT_2[29284] = 32'b11111111111111101101110111100010;
assign LUT_2[29285] = 32'b11111111111111101010101111111011;
assign LUT_2[29286] = 32'b11111111111111110100110000011110;
assign LUT_2[29287] = 32'b11111111111111110001101000110111;
assign LUT_2[29288] = 32'b11111111111111101100001011010111;
assign LUT_2[29289] = 32'b11111111111111101001000011110000;
assign LUT_2[29290] = 32'b11111111111111110011000100010011;
assign LUT_2[29291] = 32'b11111111111111101111111100101100;
assign LUT_2[29292] = 32'b11111111111111101000101000111111;
assign LUT_2[29293] = 32'b11111111111111100101100001011000;
assign LUT_2[29294] = 32'b11111111111111101111100001111011;
assign LUT_2[29295] = 32'b11111111111111101100011010010100;
assign LUT_2[29296] = 32'b11111111111111101011111110000100;
assign LUT_2[29297] = 32'b11111111111111101000110110011101;
assign LUT_2[29298] = 32'b11111111111111110010110111000000;
assign LUT_2[29299] = 32'b11111111111111101111101111011001;
assign LUT_2[29300] = 32'b11111111111111101000011011101100;
assign LUT_2[29301] = 32'b11111111111111100101010100000101;
assign LUT_2[29302] = 32'b11111111111111101111010100101000;
assign LUT_2[29303] = 32'b11111111111111101100001101000001;
assign LUT_2[29304] = 32'b11111111111111100110101111100001;
assign LUT_2[29305] = 32'b11111111111111100011100111111010;
assign LUT_2[29306] = 32'b11111111111111101101101000011101;
assign LUT_2[29307] = 32'b11111111111111101010100000110110;
assign LUT_2[29308] = 32'b11111111111111100011001101001001;
assign LUT_2[29309] = 32'b11111111111111100000000101100010;
assign LUT_2[29310] = 32'b11111111111111101010000110000101;
assign LUT_2[29311] = 32'b11111111111111100110111110011110;
assign LUT_2[29312] = 32'b11111111111111111101001001111101;
assign LUT_2[29313] = 32'b11111111111111111010000010010110;
assign LUT_2[29314] = 32'b00000000000000000100000010111001;
assign LUT_2[29315] = 32'b00000000000000000000111011010010;
assign LUT_2[29316] = 32'b11111111111111111001100111100101;
assign LUT_2[29317] = 32'b11111111111111110110011111111110;
assign LUT_2[29318] = 32'b00000000000000000000100000100001;
assign LUT_2[29319] = 32'b11111111111111111101011000111010;
assign LUT_2[29320] = 32'b11111111111111110111111011011010;
assign LUT_2[29321] = 32'b11111111111111110100110011110011;
assign LUT_2[29322] = 32'b11111111111111111110110100010110;
assign LUT_2[29323] = 32'b11111111111111111011101100101111;
assign LUT_2[29324] = 32'b11111111111111110100011001000010;
assign LUT_2[29325] = 32'b11111111111111110001010001011011;
assign LUT_2[29326] = 32'b11111111111111111011010001111110;
assign LUT_2[29327] = 32'b11111111111111111000001010010111;
assign LUT_2[29328] = 32'b11111111111111110111101110000111;
assign LUT_2[29329] = 32'b11111111111111110100100110100000;
assign LUT_2[29330] = 32'b11111111111111111110100111000011;
assign LUT_2[29331] = 32'b11111111111111111011011111011100;
assign LUT_2[29332] = 32'b11111111111111110100001011101111;
assign LUT_2[29333] = 32'b11111111111111110001000100001000;
assign LUT_2[29334] = 32'b11111111111111111011000100101011;
assign LUT_2[29335] = 32'b11111111111111110111111101000100;
assign LUT_2[29336] = 32'b11111111111111110010011111100100;
assign LUT_2[29337] = 32'b11111111111111101111010111111101;
assign LUT_2[29338] = 32'b11111111111111111001011000100000;
assign LUT_2[29339] = 32'b11111111111111110110010000111001;
assign LUT_2[29340] = 32'b11111111111111101110111101001100;
assign LUT_2[29341] = 32'b11111111111111101011110101100101;
assign LUT_2[29342] = 32'b11111111111111110101110110001000;
assign LUT_2[29343] = 32'b11111111111111110010101110100001;
assign LUT_2[29344] = 32'b11111111111111111101100101100110;
assign LUT_2[29345] = 32'b11111111111111111010011101111111;
assign LUT_2[29346] = 32'b00000000000000000100011110100010;
assign LUT_2[29347] = 32'b00000000000000000001010110111011;
assign LUT_2[29348] = 32'b11111111111111111010000011001110;
assign LUT_2[29349] = 32'b11111111111111110110111011100111;
assign LUT_2[29350] = 32'b00000000000000000000111100001010;
assign LUT_2[29351] = 32'b11111111111111111101110100100011;
assign LUT_2[29352] = 32'b11111111111111111000010111000011;
assign LUT_2[29353] = 32'b11111111111111110101001111011100;
assign LUT_2[29354] = 32'b11111111111111111111001111111111;
assign LUT_2[29355] = 32'b11111111111111111100001000011000;
assign LUT_2[29356] = 32'b11111111111111110100110100101011;
assign LUT_2[29357] = 32'b11111111111111110001101101000100;
assign LUT_2[29358] = 32'b11111111111111111011101101100111;
assign LUT_2[29359] = 32'b11111111111111111000100110000000;
assign LUT_2[29360] = 32'b11111111111111111000001001110000;
assign LUT_2[29361] = 32'b11111111111111110101000010001001;
assign LUT_2[29362] = 32'b11111111111111111111000010101100;
assign LUT_2[29363] = 32'b11111111111111111011111011000101;
assign LUT_2[29364] = 32'b11111111111111110100100111011000;
assign LUT_2[29365] = 32'b11111111111111110001011111110001;
assign LUT_2[29366] = 32'b11111111111111111011100000010100;
assign LUT_2[29367] = 32'b11111111111111111000011000101101;
assign LUT_2[29368] = 32'b11111111111111110010111011001101;
assign LUT_2[29369] = 32'b11111111111111101111110011100110;
assign LUT_2[29370] = 32'b11111111111111111001110100001001;
assign LUT_2[29371] = 32'b11111111111111110110101100100010;
assign LUT_2[29372] = 32'b11111111111111101111011000110101;
assign LUT_2[29373] = 32'b11111111111111101100010001001110;
assign LUT_2[29374] = 32'b11111111111111110110010001110001;
assign LUT_2[29375] = 32'b11111111111111110011001010001010;
assign LUT_2[29376] = 32'b11111111111111110101010010100000;
assign LUT_2[29377] = 32'b11111111111111110010001010111001;
assign LUT_2[29378] = 32'b11111111111111111100001011011100;
assign LUT_2[29379] = 32'b11111111111111111001000011110101;
assign LUT_2[29380] = 32'b11111111111111110001110000001000;
assign LUT_2[29381] = 32'b11111111111111101110101000100001;
assign LUT_2[29382] = 32'b11111111111111111000101001000100;
assign LUT_2[29383] = 32'b11111111111111110101100001011101;
assign LUT_2[29384] = 32'b11111111111111110000000011111101;
assign LUT_2[29385] = 32'b11111111111111101100111100010110;
assign LUT_2[29386] = 32'b11111111111111110110111100111001;
assign LUT_2[29387] = 32'b11111111111111110011110101010010;
assign LUT_2[29388] = 32'b11111111111111101100100001100101;
assign LUT_2[29389] = 32'b11111111111111101001011001111110;
assign LUT_2[29390] = 32'b11111111111111110011011010100001;
assign LUT_2[29391] = 32'b11111111111111110000010010111010;
assign LUT_2[29392] = 32'b11111111111111101111110110101010;
assign LUT_2[29393] = 32'b11111111111111101100101111000011;
assign LUT_2[29394] = 32'b11111111111111110110101111100110;
assign LUT_2[29395] = 32'b11111111111111110011100111111111;
assign LUT_2[29396] = 32'b11111111111111101100010100010010;
assign LUT_2[29397] = 32'b11111111111111101001001100101011;
assign LUT_2[29398] = 32'b11111111111111110011001101001110;
assign LUT_2[29399] = 32'b11111111111111110000000101100111;
assign LUT_2[29400] = 32'b11111111111111101010101000000111;
assign LUT_2[29401] = 32'b11111111111111100111100000100000;
assign LUT_2[29402] = 32'b11111111111111110001100001000011;
assign LUT_2[29403] = 32'b11111111111111101110011001011100;
assign LUT_2[29404] = 32'b11111111111111100111000101101111;
assign LUT_2[29405] = 32'b11111111111111100011111110001000;
assign LUT_2[29406] = 32'b11111111111111101101111110101011;
assign LUT_2[29407] = 32'b11111111111111101010110111000100;
assign LUT_2[29408] = 32'b11111111111111110101101110001001;
assign LUT_2[29409] = 32'b11111111111111110010100110100010;
assign LUT_2[29410] = 32'b11111111111111111100100111000101;
assign LUT_2[29411] = 32'b11111111111111111001011111011110;
assign LUT_2[29412] = 32'b11111111111111110010001011110001;
assign LUT_2[29413] = 32'b11111111111111101111000100001010;
assign LUT_2[29414] = 32'b11111111111111111001000100101101;
assign LUT_2[29415] = 32'b11111111111111110101111101000110;
assign LUT_2[29416] = 32'b11111111111111110000011111100110;
assign LUT_2[29417] = 32'b11111111111111101101010111111111;
assign LUT_2[29418] = 32'b11111111111111110111011000100010;
assign LUT_2[29419] = 32'b11111111111111110100010000111011;
assign LUT_2[29420] = 32'b11111111111111101100111101001110;
assign LUT_2[29421] = 32'b11111111111111101001110101100111;
assign LUT_2[29422] = 32'b11111111111111110011110110001010;
assign LUT_2[29423] = 32'b11111111111111110000101110100011;
assign LUT_2[29424] = 32'b11111111111111110000010010010011;
assign LUT_2[29425] = 32'b11111111111111101101001010101100;
assign LUT_2[29426] = 32'b11111111111111110111001011001111;
assign LUT_2[29427] = 32'b11111111111111110100000011101000;
assign LUT_2[29428] = 32'b11111111111111101100101111111011;
assign LUT_2[29429] = 32'b11111111111111101001101000010100;
assign LUT_2[29430] = 32'b11111111111111110011101000110111;
assign LUT_2[29431] = 32'b11111111111111110000100001010000;
assign LUT_2[29432] = 32'b11111111111111101011000011110000;
assign LUT_2[29433] = 32'b11111111111111100111111100001001;
assign LUT_2[29434] = 32'b11111111111111110001111100101100;
assign LUT_2[29435] = 32'b11111111111111101110110101000101;
assign LUT_2[29436] = 32'b11111111111111100111100001011000;
assign LUT_2[29437] = 32'b11111111111111100100011001110001;
assign LUT_2[29438] = 32'b11111111111111101110011010010100;
assign LUT_2[29439] = 32'b11111111111111101011010010101101;
assign LUT_2[29440] = 32'b11111111111111111100110100010100;
assign LUT_2[29441] = 32'b11111111111111111001101100101101;
assign LUT_2[29442] = 32'b00000000000000000011101101010000;
assign LUT_2[29443] = 32'b00000000000000000000100101101001;
assign LUT_2[29444] = 32'b11111111111111111001010001111100;
assign LUT_2[29445] = 32'b11111111111111110110001010010101;
assign LUT_2[29446] = 32'b00000000000000000000001010111000;
assign LUT_2[29447] = 32'b11111111111111111101000011010001;
assign LUT_2[29448] = 32'b11111111111111110111100101110001;
assign LUT_2[29449] = 32'b11111111111111110100011110001010;
assign LUT_2[29450] = 32'b11111111111111111110011110101101;
assign LUT_2[29451] = 32'b11111111111111111011010111000110;
assign LUT_2[29452] = 32'b11111111111111110100000011011001;
assign LUT_2[29453] = 32'b11111111111111110000111011110010;
assign LUT_2[29454] = 32'b11111111111111111010111100010101;
assign LUT_2[29455] = 32'b11111111111111110111110100101110;
assign LUT_2[29456] = 32'b11111111111111110111011000011110;
assign LUT_2[29457] = 32'b11111111111111110100010000110111;
assign LUT_2[29458] = 32'b11111111111111111110010001011010;
assign LUT_2[29459] = 32'b11111111111111111011001001110011;
assign LUT_2[29460] = 32'b11111111111111110011110110000110;
assign LUT_2[29461] = 32'b11111111111111110000101110011111;
assign LUT_2[29462] = 32'b11111111111111111010101111000010;
assign LUT_2[29463] = 32'b11111111111111110111100111011011;
assign LUT_2[29464] = 32'b11111111111111110010001001111011;
assign LUT_2[29465] = 32'b11111111111111101111000010010100;
assign LUT_2[29466] = 32'b11111111111111111001000010110111;
assign LUT_2[29467] = 32'b11111111111111110101111011010000;
assign LUT_2[29468] = 32'b11111111111111101110100111100011;
assign LUT_2[29469] = 32'b11111111111111101011011111111100;
assign LUT_2[29470] = 32'b11111111111111110101100000011111;
assign LUT_2[29471] = 32'b11111111111111110010011000111000;
assign LUT_2[29472] = 32'b11111111111111111101001111111101;
assign LUT_2[29473] = 32'b11111111111111111010001000010110;
assign LUT_2[29474] = 32'b00000000000000000100001000111001;
assign LUT_2[29475] = 32'b00000000000000000001000001010010;
assign LUT_2[29476] = 32'b11111111111111111001101101100101;
assign LUT_2[29477] = 32'b11111111111111110110100101111110;
assign LUT_2[29478] = 32'b00000000000000000000100110100001;
assign LUT_2[29479] = 32'b11111111111111111101011110111010;
assign LUT_2[29480] = 32'b11111111111111111000000001011010;
assign LUT_2[29481] = 32'b11111111111111110100111001110011;
assign LUT_2[29482] = 32'b11111111111111111110111010010110;
assign LUT_2[29483] = 32'b11111111111111111011110010101111;
assign LUT_2[29484] = 32'b11111111111111110100011111000010;
assign LUT_2[29485] = 32'b11111111111111110001010111011011;
assign LUT_2[29486] = 32'b11111111111111111011010111111110;
assign LUT_2[29487] = 32'b11111111111111111000010000010111;
assign LUT_2[29488] = 32'b11111111111111110111110100000111;
assign LUT_2[29489] = 32'b11111111111111110100101100100000;
assign LUT_2[29490] = 32'b11111111111111111110101101000011;
assign LUT_2[29491] = 32'b11111111111111111011100101011100;
assign LUT_2[29492] = 32'b11111111111111110100010001101111;
assign LUT_2[29493] = 32'b11111111111111110001001010001000;
assign LUT_2[29494] = 32'b11111111111111111011001010101011;
assign LUT_2[29495] = 32'b11111111111111111000000011000100;
assign LUT_2[29496] = 32'b11111111111111110010100101100100;
assign LUT_2[29497] = 32'b11111111111111101111011101111101;
assign LUT_2[29498] = 32'b11111111111111111001011110100000;
assign LUT_2[29499] = 32'b11111111111111110110010110111001;
assign LUT_2[29500] = 32'b11111111111111101111000011001100;
assign LUT_2[29501] = 32'b11111111111111101011111011100101;
assign LUT_2[29502] = 32'b11111111111111110101111100001000;
assign LUT_2[29503] = 32'b11111111111111110010110100100001;
assign LUT_2[29504] = 32'b11111111111111110100111100110111;
assign LUT_2[29505] = 32'b11111111111111110001110101010000;
assign LUT_2[29506] = 32'b11111111111111111011110101110011;
assign LUT_2[29507] = 32'b11111111111111111000101110001100;
assign LUT_2[29508] = 32'b11111111111111110001011010011111;
assign LUT_2[29509] = 32'b11111111111111101110010010111000;
assign LUT_2[29510] = 32'b11111111111111111000010011011011;
assign LUT_2[29511] = 32'b11111111111111110101001011110100;
assign LUT_2[29512] = 32'b11111111111111101111101110010100;
assign LUT_2[29513] = 32'b11111111111111101100100110101101;
assign LUT_2[29514] = 32'b11111111111111110110100111010000;
assign LUT_2[29515] = 32'b11111111111111110011011111101001;
assign LUT_2[29516] = 32'b11111111111111101100001011111100;
assign LUT_2[29517] = 32'b11111111111111101001000100010101;
assign LUT_2[29518] = 32'b11111111111111110011000100111000;
assign LUT_2[29519] = 32'b11111111111111101111111101010001;
assign LUT_2[29520] = 32'b11111111111111101111100001000001;
assign LUT_2[29521] = 32'b11111111111111101100011001011010;
assign LUT_2[29522] = 32'b11111111111111110110011001111101;
assign LUT_2[29523] = 32'b11111111111111110011010010010110;
assign LUT_2[29524] = 32'b11111111111111101011111110101001;
assign LUT_2[29525] = 32'b11111111111111101000110111000010;
assign LUT_2[29526] = 32'b11111111111111110010110111100101;
assign LUT_2[29527] = 32'b11111111111111101111101111111110;
assign LUT_2[29528] = 32'b11111111111111101010010010011110;
assign LUT_2[29529] = 32'b11111111111111100111001010110111;
assign LUT_2[29530] = 32'b11111111111111110001001011011010;
assign LUT_2[29531] = 32'b11111111111111101110000011110011;
assign LUT_2[29532] = 32'b11111111111111100110110000000110;
assign LUT_2[29533] = 32'b11111111111111100011101000011111;
assign LUT_2[29534] = 32'b11111111111111101101101001000010;
assign LUT_2[29535] = 32'b11111111111111101010100001011011;
assign LUT_2[29536] = 32'b11111111111111110101011000100000;
assign LUT_2[29537] = 32'b11111111111111110010010000111001;
assign LUT_2[29538] = 32'b11111111111111111100010001011100;
assign LUT_2[29539] = 32'b11111111111111111001001001110101;
assign LUT_2[29540] = 32'b11111111111111110001110110001000;
assign LUT_2[29541] = 32'b11111111111111101110101110100001;
assign LUT_2[29542] = 32'b11111111111111111000101111000100;
assign LUT_2[29543] = 32'b11111111111111110101100111011101;
assign LUT_2[29544] = 32'b11111111111111110000001001111101;
assign LUT_2[29545] = 32'b11111111111111101101000010010110;
assign LUT_2[29546] = 32'b11111111111111110111000010111001;
assign LUT_2[29547] = 32'b11111111111111110011111011010010;
assign LUT_2[29548] = 32'b11111111111111101100100111100101;
assign LUT_2[29549] = 32'b11111111111111101001011111111110;
assign LUT_2[29550] = 32'b11111111111111110011100000100001;
assign LUT_2[29551] = 32'b11111111111111110000011000111010;
assign LUT_2[29552] = 32'b11111111111111101111111100101010;
assign LUT_2[29553] = 32'b11111111111111101100110101000011;
assign LUT_2[29554] = 32'b11111111111111110110110101100110;
assign LUT_2[29555] = 32'b11111111111111110011101101111111;
assign LUT_2[29556] = 32'b11111111111111101100011010010010;
assign LUT_2[29557] = 32'b11111111111111101001010010101011;
assign LUT_2[29558] = 32'b11111111111111110011010011001110;
assign LUT_2[29559] = 32'b11111111111111110000001011100111;
assign LUT_2[29560] = 32'b11111111111111101010101110000111;
assign LUT_2[29561] = 32'b11111111111111100111100110100000;
assign LUT_2[29562] = 32'b11111111111111110001100111000011;
assign LUT_2[29563] = 32'b11111111111111101110011111011100;
assign LUT_2[29564] = 32'b11111111111111100111001011101111;
assign LUT_2[29565] = 32'b11111111111111100100000100001000;
assign LUT_2[29566] = 32'b11111111111111101110000100101011;
assign LUT_2[29567] = 32'b11111111111111101010111101000100;
assign LUT_2[29568] = 32'b00000000000000000001001000100011;
assign LUT_2[29569] = 32'b11111111111111111110000000111100;
assign LUT_2[29570] = 32'b00000000000000001000000001011111;
assign LUT_2[29571] = 32'b00000000000000000100111001111000;
assign LUT_2[29572] = 32'b11111111111111111101100110001011;
assign LUT_2[29573] = 32'b11111111111111111010011110100100;
assign LUT_2[29574] = 32'b00000000000000000100011111000111;
assign LUT_2[29575] = 32'b00000000000000000001010111100000;
assign LUT_2[29576] = 32'b11111111111111111011111010000000;
assign LUT_2[29577] = 32'b11111111111111111000110010011001;
assign LUT_2[29578] = 32'b00000000000000000010110010111100;
assign LUT_2[29579] = 32'b11111111111111111111101011010101;
assign LUT_2[29580] = 32'b11111111111111111000010111101000;
assign LUT_2[29581] = 32'b11111111111111110101010000000001;
assign LUT_2[29582] = 32'b11111111111111111111010000100100;
assign LUT_2[29583] = 32'b11111111111111111100001000111101;
assign LUT_2[29584] = 32'b11111111111111111011101100101101;
assign LUT_2[29585] = 32'b11111111111111111000100101000110;
assign LUT_2[29586] = 32'b00000000000000000010100101101001;
assign LUT_2[29587] = 32'b11111111111111111111011110000010;
assign LUT_2[29588] = 32'b11111111111111111000001010010101;
assign LUT_2[29589] = 32'b11111111111111110101000010101110;
assign LUT_2[29590] = 32'b11111111111111111111000011010001;
assign LUT_2[29591] = 32'b11111111111111111011111011101010;
assign LUT_2[29592] = 32'b11111111111111110110011110001010;
assign LUT_2[29593] = 32'b11111111111111110011010110100011;
assign LUT_2[29594] = 32'b11111111111111111101010111000110;
assign LUT_2[29595] = 32'b11111111111111111010001111011111;
assign LUT_2[29596] = 32'b11111111111111110010111011110010;
assign LUT_2[29597] = 32'b11111111111111101111110100001011;
assign LUT_2[29598] = 32'b11111111111111111001110100101110;
assign LUT_2[29599] = 32'b11111111111111110110101101000111;
assign LUT_2[29600] = 32'b00000000000000000001100100001100;
assign LUT_2[29601] = 32'b11111111111111111110011100100101;
assign LUT_2[29602] = 32'b00000000000000001000011101001000;
assign LUT_2[29603] = 32'b00000000000000000101010101100001;
assign LUT_2[29604] = 32'b11111111111111111110000001110100;
assign LUT_2[29605] = 32'b11111111111111111010111010001101;
assign LUT_2[29606] = 32'b00000000000000000100111010110000;
assign LUT_2[29607] = 32'b00000000000000000001110011001001;
assign LUT_2[29608] = 32'b11111111111111111100010101101001;
assign LUT_2[29609] = 32'b11111111111111111001001110000010;
assign LUT_2[29610] = 32'b00000000000000000011001110100101;
assign LUT_2[29611] = 32'b00000000000000000000000110111110;
assign LUT_2[29612] = 32'b11111111111111111000110011010001;
assign LUT_2[29613] = 32'b11111111111111110101101011101010;
assign LUT_2[29614] = 32'b11111111111111111111101100001101;
assign LUT_2[29615] = 32'b11111111111111111100100100100110;
assign LUT_2[29616] = 32'b11111111111111111100001000010110;
assign LUT_2[29617] = 32'b11111111111111111001000000101111;
assign LUT_2[29618] = 32'b00000000000000000011000001010010;
assign LUT_2[29619] = 32'b11111111111111111111111001101011;
assign LUT_2[29620] = 32'b11111111111111111000100101111110;
assign LUT_2[29621] = 32'b11111111111111110101011110010111;
assign LUT_2[29622] = 32'b11111111111111111111011110111010;
assign LUT_2[29623] = 32'b11111111111111111100010111010011;
assign LUT_2[29624] = 32'b11111111111111110110111001110011;
assign LUT_2[29625] = 32'b11111111111111110011110010001100;
assign LUT_2[29626] = 32'b11111111111111111101110010101111;
assign LUT_2[29627] = 32'b11111111111111111010101011001000;
assign LUT_2[29628] = 32'b11111111111111110011010111011011;
assign LUT_2[29629] = 32'b11111111111111110000001111110100;
assign LUT_2[29630] = 32'b11111111111111111010010000010111;
assign LUT_2[29631] = 32'b11111111111111110111001000110000;
assign LUT_2[29632] = 32'b11111111111111111001010001000110;
assign LUT_2[29633] = 32'b11111111111111110110001001011111;
assign LUT_2[29634] = 32'b00000000000000000000001010000010;
assign LUT_2[29635] = 32'b11111111111111111101000010011011;
assign LUT_2[29636] = 32'b11111111111111110101101110101110;
assign LUT_2[29637] = 32'b11111111111111110010100111000111;
assign LUT_2[29638] = 32'b11111111111111111100100111101010;
assign LUT_2[29639] = 32'b11111111111111111001100000000011;
assign LUT_2[29640] = 32'b11111111111111110100000010100011;
assign LUT_2[29641] = 32'b11111111111111110000111010111100;
assign LUT_2[29642] = 32'b11111111111111111010111011011111;
assign LUT_2[29643] = 32'b11111111111111110111110011111000;
assign LUT_2[29644] = 32'b11111111111111110000100000001011;
assign LUT_2[29645] = 32'b11111111111111101101011000100100;
assign LUT_2[29646] = 32'b11111111111111110111011001000111;
assign LUT_2[29647] = 32'b11111111111111110100010001100000;
assign LUT_2[29648] = 32'b11111111111111110011110101010000;
assign LUT_2[29649] = 32'b11111111111111110000101101101001;
assign LUT_2[29650] = 32'b11111111111111111010101110001100;
assign LUT_2[29651] = 32'b11111111111111110111100110100101;
assign LUT_2[29652] = 32'b11111111111111110000010010111000;
assign LUT_2[29653] = 32'b11111111111111101101001011010001;
assign LUT_2[29654] = 32'b11111111111111110111001011110100;
assign LUT_2[29655] = 32'b11111111111111110100000100001101;
assign LUT_2[29656] = 32'b11111111111111101110100110101101;
assign LUT_2[29657] = 32'b11111111111111101011011111000110;
assign LUT_2[29658] = 32'b11111111111111110101011111101001;
assign LUT_2[29659] = 32'b11111111111111110010011000000010;
assign LUT_2[29660] = 32'b11111111111111101011000100010101;
assign LUT_2[29661] = 32'b11111111111111100111111100101110;
assign LUT_2[29662] = 32'b11111111111111110001111101010001;
assign LUT_2[29663] = 32'b11111111111111101110110101101010;
assign LUT_2[29664] = 32'b11111111111111111001101100101111;
assign LUT_2[29665] = 32'b11111111111111110110100101001000;
assign LUT_2[29666] = 32'b00000000000000000000100101101011;
assign LUT_2[29667] = 32'b11111111111111111101011110000100;
assign LUT_2[29668] = 32'b11111111111111110110001010010111;
assign LUT_2[29669] = 32'b11111111111111110011000010110000;
assign LUT_2[29670] = 32'b11111111111111111101000011010011;
assign LUT_2[29671] = 32'b11111111111111111001111011101100;
assign LUT_2[29672] = 32'b11111111111111110100011110001100;
assign LUT_2[29673] = 32'b11111111111111110001010110100101;
assign LUT_2[29674] = 32'b11111111111111111011010111001000;
assign LUT_2[29675] = 32'b11111111111111111000001111100001;
assign LUT_2[29676] = 32'b11111111111111110000111011110100;
assign LUT_2[29677] = 32'b11111111111111101101110100001101;
assign LUT_2[29678] = 32'b11111111111111110111110100110000;
assign LUT_2[29679] = 32'b11111111111111110100101101001001;
assign LUT_2[29680] = 32'b11111111111111110100010000111001;
assign LUT_2[29681] = 32'b11111111111111110001001001010010;
assign LUT_2[29682] = 32'b11111111111111111011001001110101;
assign LUT_2[29683] = 32'b11111111111111111000000010001110;
assign LUT_2[29684] = 32'b11111111111111110000101110100001;
assign LUT_2[29685] = 32'b11111111111111101101100110111010;
assign LUT_2[29686] = 32'b11111111111111110111100111011101;
assign LUT_2[29687] = 32'b11111111111111110100011111110110;
assign LUT_2[29688] = 32'b11111111111111101111000010010110;
assign LUT_2[29689] = 32'b11111111111111101011111010101111;
assign LUT_2[29690] = 32'b11111111111111110101111011010010;
assign LUT_2[29691] = 32'b11111111111111110010110011101011;
assign LUT_2[29692] = 32'b11111111111111101011011111111110;
assign LUT_2[29693] = 32'b11111111111111101000011000010111;
assign LUT_2[29694] = 32'b11111111111111110010011000111010;
assign LUT_2[29695] = 32'b11111111111111101111010001010011;
assign LUT_2[29696] = 32'b11111111111111111010110000000001;
assign LUT_2[29697] = 32'b11111111111111110111101000011010;
assign LUT_2[29698] = 32'b00000000000000000001101000111101;
assign LUT_2[29699] = 32'b11111111111111111110100001010110;
assign LUT_2[29700] = 32'b11111111111111110111001101101001;
assign LUT_2[29701] = 32'b11111111111111110100000110000010;
assign LUT_2[29702] = 32'b11111111111111111110000110100101;
assign LUT_2[29703] = 32'b11111111111111111010111110111110;
assign LUT_2[29704] = 32'b11111111111111110101100001011110;
assign LUT_2[29705] = 32'b11111111111111110010011001110111;
assign LUT_2[29706] = 32'b11111111111111111100011010011010;
assign LUT_2[29707] = 32'b11111111111111111001010010110011;
assign LUT_2[29708] = 32'b11111111111111110001111111000110;
assign LUT_2[29709] = 32'b11111111111111101110110111011111;
assign LUT_2[29710] = 32'b11111111111111111000111000000010;
assign LUT_2[29711] = 32'b11111111111111110101110000011011;
assign LUT_2[29712] = 32'b11111111111111110101010100001011;
assign LUT_2[29713] = 32'b11111111111111110010001100100100;
assign LUT_2[29714] = 32'b11111111111111111100001101000111;
assign LUT_2[29715] = 32'b11111111111111111001000101100000;
assign LUT_2[29716] = 32'b11111111111111110001110001110011;
assign LUT_2[29717] = 32'b11111111111111101110101010001100;
assign LUT_2[29718] = 32'b11111111111111111000101010101111;
assign LUT_2[29719] = 32'b11111111111111110101100011001000;
assign LUT_2[29720] = 32'b11111111111111110000000101101000;
assign LUT_2[29721] = 32'b11111111111111101100111110000001;
assign LUT_2[29722] = 32'b11111111111111110110111110100100;
assign LUT_2[29723] = 32'b11111111111111110011110110111101;
assign LUT_2[29724] = 32'b11111111111111101100100011010000;
assign LUT_2[29725] = 32'b11111111111111101001011011101001;
assign LUT_2[29726] = 32'b11111111111111110011011100001100;
assign LUT_2[29727] = 32'b11111111111111110000010100100101;
assign LUT_2[29728] = 32'b11111111111111111011001011101010;
assign LUT_2[29729] = 32'b11111111111111111000000100000011;
assign LUT_2[29730] = 32'b00000000000000000010000100100110;
assign LUT_2[29731] = 32'b11111111111111111110111100111111;
assign LUT_2[29732] = 32'b11111111111111110111101001010010;
assign LUT_2[29733] = 32'b11111111111111110100100001101011;
assign LUT_2[29734] = 32'b11111111111111111110100010001110;
assign LUT_2[29735] = 32'b11111111111111111011011010100111;
assign LUT_2[29736] = 32'b11111111111111110101111101000111;
assign LUT_2[29737] = 32'b11111111111111110010110101100000;
assign LUT_2[29738] = 32'b11111111111111111100110110000011;
assign LUT_2[29739] = 32'b11111111111111111001101110011100;
assign LUT_2[29740] = 32'b11111111111111110010011010101111;
assign LUT_2[29741] = 32'b11111111111111101111010011001000;
assign LUT_2[29742] = 32'b11111111111111111001010011101011;
assign LUT_2[29743] = 32'b11111111111111110110001100000100;
assign LUT_2[29744] = 32'b11111111111111110101101111110100;
assign LUT_2[29745] = 32'b11111111111111110010101000001101;
assign LUT_2[29746] = 32'b11111111111111111100101000110000;
assign LUT_2[29747] = 32'b11111111111111111001100001001001;
assign LUT_2[29748] = 32'b11111111111111110010001101011100;
assign LUT_2[29749] = 32'b11111111111111101111000101110101;
assign LUT_2[29750] = 32'b11111111111111111001000110011000;
assign LUT_2[29751] = 32'b11111111111111110101111110110001;
assign LUT_2[29752] = 32'b11111111111111110000100001010001;
assign LUT_2[29753] = 32'b11111111111111101101011001101010;
assign LUT_2[29754] = 32'b11111111111111110111011010001101;
assign LUT_2[29755] = 32'b11111111111111110100010010100110;
assign LUT_2[29756] = 32'b11111111111111101100111110111001;
assign LUT_2[29757] = 32'b11111111111111101001110111010010;
assign LUT_2[29758] = 32'b11111111111111110011110111110101;
assign LUT_2[29759] = 32'b11111111111111110000110000001110;
assign LUT_2[29760] = 32'b11111111111111110010111000100100;
assign LUT_2[29761] = 32'b11111111111111101111110000111101;
assign LUT_2[29762] = 32'b11111111111111111001110001100000;
assign LUT_2[29763] = 32'b11111111111111110110101001111001;
assign LUT_2[29764] = 32'b11111111111111101111010110001100;
assign LUT_2[29765] = 32'b11111111111111101100001110100101;
assign LUT_2[29766] = 32'b11111111111111110110001111001000;
assign LUT_2[29767] = 32'b11111111111111110011000111100001;
assign LUT_2[29768] = 32'b11111111111111101101101010000001;
assign LUT_2[29769] = 32'b11111111111111101010100010011010;
assign LUT_2[29770] = 32'b11111111111111110100100010111101;
assign LUT_2[29771] = 32'b11111111111111110001011011010110;
assign LUT_2[29772] = 32'b11111111111111101010000111101001;
assign LUT_2[29773] = 32'b11111111111111100111000000000010;
assign LUT_2[29774] = 32'b11111111111111110001000000100101;
assign LUT_2[29775] = 32'b11111111111111101101111000111110;
assign LUT_2[29776] = 32'b11111111111111101101011100101110;
assign LUT_2[29777] = 32'b11111111111111101010010101000111;
assign LUT_2[29778] = 32'b11111111111111110100010101101010;
assign LUT_2[29779] = 32'b11111111111111110001001110000011;
assign LUT_2[29780] = 32'b11111111111111101001111010010110;
assign LUT_2[29781] = 32'b11111111111111100110110010101111;
assign LUT_2[29782] = 32'b11111111111111110000110011010010;
assign LUT_2[29783] = 32'b11111111111111101101101011101011;
assign LUT_2[29784] = 32'b11111111111111101000001110001011;
assign LUT_2[29785] = 32'b11111111111111100101000110100100;
assign LUT_2[29786] = 32'b11111111111111101111000111000111;
assign LUT_2[29787] = 32'b11111111111111101011111111100000;
assign LUT_2[29788] = 32'b11111111111111100100101011110011;
assign LUT_2[29789] = 32'b11111111111111100001100100001100;
assign LUT_2[29790] = 32'b11111111111111101011100100101111;
assign LUT_2[29791] = 32'b11111111111111101000011101001000;
assign LUT_2[29792] = 32'b11111111111111110011010100001101;
assign LUT_2[29793] = 32'b11111111111111110000001100100110;
assign LUT_2[29794] = 32'b11111111111111111010001101001001;
assign LUT_2[29795] = 32'b11111111111111110111000101100010;
assign LUT_2[29796] = 32'b11111111111111101111110001110101;
assign LUT_2[29797] = 32'b11111111111111101100101010001110;
assign LUT_2[29798] = 32'b11111111111111110110101010110001;
assign LUT_2[29799] = 32'b11111111111111110011100011001010;
assign LUT_2[29800] = 32'b11111111111111101110000101101010;
assign LUT_2[29801] = 32'b11111111111111101010111110000011;
assign LUT_2[29802] = 32'b11111111111111110100111110100110;
assign LUT_2[29803] = 32'b11111111111111110001110110111111;
assign LUT_2[29804] = 32'b11111111111111101010100011010010;
assign LUT_2[29805] = 32'b11111111111111100111011011101011;
assign LUT_2[29806] = 32'b11111111111111110001011100001110;
assign LUT_2[29807] = 32'b11111111111111101110010100100111;
assign LUT_2[29808] = 32'b11111111111111101101111000010111;
assign LUT_2[29809] = 32'b11111111111111101010110000110000;
assign LUT_2[29810] = 32'b11111111111111110100110001010011;
assign LUT_2[29811] = 32'b11111111111111110001101001101100;
assign LUT_2[29812] = 32'b11111111111111101010010101111111;
assign LUT_2[29813] = 32'b11111111111111100111001110011000;
assign LUT_2[29814] = 32'b11111111111111110001001110111011;
assign LUT_2[29815] = 32'b11111111111111101110000111010100;
assign LUT_2[29816] = 32'b11111111111111101000101001110100;
assign LUT_2[29817] = 32'b11111111111111100101100010001101;
assign LUT_2[29818] = 32'b11111111111111101111100010110000;
assign LUT_2[29819] = 32'b11111111111111101100011011001001;
assign LUT_2[29820] = 32'b11111111111111100101000111011100;
assign LUT_2[29821] = 32'b11111111111111100001111111110101;
assign LUT_2[29822] = 32'b11111111111111101100000000011000;
assign LUT_2[29823] = 32'b11111111111111101000111000110001;
assign LUT_2[29824] = 32'b11111111111111111111000100010000;
assign LUT_2[29825] = 32'b11111111111111111011111100101001;
assign LUT_2[29826] = 32'b00000000000000000101111101001100;
assign LUT_2[29827] = 32'b00000000000000000010110101100101;
assign LUT_2[29828] = 32'b11111111111111111011100001111000;
assign LUT_2[29829] = 32'b11111111111111111000011010010001;
assign LUT_2[29830] = 32'b00000000000000000010011010110100;
assign LUT_2[29831] = 32'b11111111111111111111010011001101;
assign LUT_2[29832] = 32'b11111111111111111001110101101101;
assign LUT_2[29833] = 32'b11111111111111110110101110000110;
assign LUT_2[29834] = 32'b00000000000000000000101110101001;
assign LUT_2[29835] = 32'b11111111111111111101100111000010;
assign LUT_2[29836] = 32'b11111111111111110110010011010101;
assign LUT_2[29837] = 32'b11111111111111110011001011101110;
assign LUT_2[29838] = 32'b11111111111111111101001100010001;
assign LUT_2[29839] = 32'b11111111111111111010000100101010;
assign LUT_2[29840] = 32'b11111111111111111001101000011010;
assign LUT_2[29841] = 32'b11111111111111110110100000110011;
assign LUT_2[29842] = 32'b00000000000000000000100001010110;
assign LUT_2[29843] = 32'b11111111111111111101011001101111;
assign LUT_2[29844] = 32'b11111111111111110110000110000010;
assign LUT_2[29845] = 32'b11111111111111110010111110011011;
assign LUT_2[29846] = 32'b11111111111111111100111110111110;
assign LUT_2[29847] = 32'b11111111111111111001110111010111;
assign LUT_2[29848] = 32'b11111111111111110100011001110111;
assign LUT_2[29849] = 32'b11111111111111110001010010010000;
assign LUT_2[29850] = 32'b11111111111111111011010010110011;
assign LUT_2[29851] = 32'b11111111111111111000001011001100;
assign LUT_2[29852] = 32'b11111111111111110000110111011111;
assign LUT_2[29853] = 32'b11111111111111101101101111111000;
assign LUT_2[29854] = 32'b11111111111111110111110000011011;
assign LUT_2[29855] = 32'b11111111111111110100101000110100;
assign LUT_2[29856] = 32'b11111111111111111111011111111001;
assign LUT_2[29857] = 32'b11111111111111111100011000010010;
assign LUT_2[29858] = 32'b00000000000000000110011000110101;
assign LUT_2[29859] = 32'b00000000000000000011010001001110;
assign LUT_2[29860] = 32'b11111111111111111011111101100001;
assign LUT_2[29861] = 32'b11111111111111111000110101111010;
assign LUT_2[29862] = 32'b00000000000000000010110110011101;
assign LUT_2[29863] = 32'b11111111111111111111101110110110;
assign LUT_2[29864] = 32'b11111111111111111010010001010110;
assign LUT_2[29865] = 32'b11111111111111110111001001101111;
assign LUT_2[29866] = 32'b00000000000000000001001010010010;
assign LUT_2[29867] = 32'b11111111111111111110000010101011;
assign LUT_2[29868] = 32'b11111111111111110110101110111110;
assign LUT_2[29869] = 32'b11111111111111110011100111010111;
assign LUT_2[29870] = 32'b11111111111111111101100111111010;
assign LUT_2[29871] = 32'b11111111111111111010100000010011;
assign LUT_2[29872] = 32'b11111111111111111010000100000011;
assign LUT_2[29873] = 32'b11111111111111110110111100011100;
assign LUT_2[29874] = 32'b00000000000000000000111100111111;
assign LUT_2[29875] = 32'b11111111111111111101110101011000;
assign LUT_2[29876] = 32'b11111111111111110110100001101011;
assign LUT_2[29877] = 32'b11111111111111110011011010000100;
assign LUT_2[29878] = 32'b11111111111111111101011010100111;
assign LUT_2[29879] = 32'b11111111111111111010010011000000;
assign LUT_2[29880] = 32'b11111111111111110100110101100000;
assign LUT_2[29881] = 32'b11111111111111110001101101111001;
assign LUT_2[29882] = 32'b11111111111111111011101110011100;
assign LUT_2[29883] = 32'b11111111111111111000100110110101;
assign LUT_2[29884] = 32'b11111111111111110001010011001000;
assign LUT_2[29885] = 32'b11111111111111101110001011100001;
assign LUT_2[29886] = 32'b11111111111111111000001100000100;
assign LUT_2[29887] = 32'b11111111111111110101000100011101;
assign LUT_2[29888] = 32'b11111111111111110111001100110011;
assign LUT_2[29889] = 32'b11111111111111110100000101001100;
assign LUT_2[29890] = 32'b11111111111111111110000101101111;
assign LUT_2[29891] = 32'b11111111111111111010111110001000;
assign LUT_2[29892] = 32'b11111111111111110011101010011011;
assign LUT_2[29893] = 32'b11111111111111110000100010110100;
assign LUT_2[29894] = 32'b11111111111111111010100011010111;
assign LUT_2[29895] = 32'b11111111111111110111011011110000;
assign LUT_2[29896] = 32'b11111111111111110001111110010000;
assign LUT_2[29897] = 32'b11111111111111101110110110101001;
assign LUT_2[29898] = 32'b11111111111111111000110111001100;
assign LUT_2[29899] = 32'b11111111111111110101101111100101;
assign LUT_2[29900] = 32'b11111111111111101110011011111000;
assign LUT_2[29901] = 32'b11111111111111101011010100010001;
assign LUT_2[29902] = 32'b11111111111111110101010100110100;
assign LUT_2[29903] = 32'b11111111111111110010001101001101;
assign LUT_2[29904] = 32'b11111111111111110001110000111101;
assign LUT_2[29905] = 32'b11111111111111101110101001010110;
assign LUT_2[29906] = 32'b11111111111111111000101001111001;
assign LUT_2[29907] = 32'b11111111111111110101100010010010;
assign LUT_2[29908] = 32'b11111111111111101110001110100101;
assign LUT_2[29909] = 32'b11111111111111101011000110111110;
assign LUT_2[29910] = 32'b11111111111111110101000111100001;
assign LUT_2[29911] = 32'b11111111111111110001111111111010;
assign LUT_2[29912] = 32'b11111111111111101100100010011010;
assign LUT_2[29913] = 32'b11111111111111101001011010110011;
assign LUT_2[29914] = 32'b11111111111111110011011011010110;
assign LUT_2[29915] = 32'b11111111111111110000010011101111;
assign LUT_2[29916] = 32'b11111111111111101001000000000010;
assign LUT_2[29917] = 32'b11111111111111100101111000011011;
assign LUT_2[29918] = 32'b11111111111111101111111000111110;
assign LUT_2[29919] = 32'b11111111111111101100110001010111;
assign LUT_2[29920] = 32'b11111111111111110111101000011100;
assign LUT_2[29921] = 32'b11111111111111110100100000110101;
assign LUT_2[29922] = 32'b11111111111111111110100001011000;
assign LUT_2[29923] = 32'b11111111111111111011011001110001;
assign LUT_2[29924] = 32'b11111111111111110100000110000100;
assign LUT_2[29925] = 32'b11111111111111110000111110011101;
assign LUT_2[29926] = 32'b11111111111111111010111111000000;
assign LUT_2[29927] = 32'b11111111111111110111110111011001;
assign LUT_2[29928] = 32'b11111111111111110010011001111001;
assign LUT_2[29929] = 32'b11111111111111101111010010010010;
assign LUT_2[29930] = 32'b11111111111111111001010010110101;
assign LUT_2[29931] = 32'b11111111111111110110001011001110;
assign LUT_2[29932] = 32'b11111111111111101110110111100001;
assign LUT_2[29933] = 32'b11111111111111101011101111111010;
assign LUT_2[29934] = 32'b11111111111111110101110000011101;
assign LUT_2[29935] = 32'b11111111111111110010101000110110;
assign LUT_2[29936] = 32'b11111111111111110010001100100110;
assign LUT_2[29937] = 32'b11111111111111101111000100111111;
assign LUT_2[29938] = 32'b11111111111111111001000101100010;
assign LUT_2[29939] = 32'b11111111111111110101111101111011;
assign LUT_2[29940] = 32'b11111111111111101110101010001110;
assign LUT_2[29941] = 32'b11111111111111101011100010100111;
assign LUT_2[29942] = 32'b11111111111111110101100011001010;
assign LUT_2[29943] = 32'b11111111111111110010011011100011;
assign LUT_2[29944] = 32'b11111111111111101100111110000011;
assign LUT_2[29945] = 32'b11111111111111101001110110011100;
assign LUT_2[29946] = 32'b11111111111111110011110110111111;
assign LUT_2[29947] = 32'b11111111111111110000101111011000;
assign LUT_2[29948] = 32'b11111111111111101001011011101011;
assign LUT_2[29949] = 32'b11111111111111100110010100000100;
assign LUT_2[29950] = 32'b11111111111111110000010100100111;
assign LUT_2[29951] = 32'b11111111111111101101001101000000;
assign LUT_2[29952] = 32'b11111111111111111110101110100111;
assign LUT_2[29953] = 32'b11111111111111111011100111000000;
assign LUT_2[29954] = 32'b00000000000000000101100111100011;
assign LUT_2[29955] = 32'b00000000000000000010011111111100;
assign LUT_2[29956] = 32'b11111111111111111011001100001111;
assign LUT_2[29957] = 32'b11111111111111111000000100101000;
assign LUT_2[29958] = 32'b00000000000000000010000101001011;
assign LUT_2[29959] = 32'b11111111111111111110111101100100;
assign LUT_2[29960] = 32'b11111111111111111001100000000100;
assign LUT_2[29961] = 32'b11111111111111110110011000011101;
assign LUT_2[29962] = 32'b00000000000000000000011001000000;
assign LUT_2[29963] = 32'b11111111111111111101010001011001;
assign LUT_2[29964] = 32'b11111111111111110101111101101100;
assign LUT_2[29965] = 32'b11111111111111110010110110000101;
assign LUT_2[29966] = 32'b11111111111111111100110110101000;
assign LUT_2[29967] = 32'b11111111111111111001101111000001;
assign LUT_2[29968] = 32'b11111111111111111001010010110001;
assign LUT_2[29969] = 32'b11111111111111110110001011001010;
assign LUT_2[29970] = 32'b00000000000000000000001011101101;
assign LUT_2[29971] = 32'b11111111111111111101000100000110;
assign LUT_2[29972] = 32'b11111111111111110101110000011001;
assign LUT_2[29973] = 32'b11111111111111110010101000110010;
assign LUT_2[29974] = 32'b11111111111111111100101001010101;
assign LUT_2[29975] = 32'b11111111111111111001100001101110;
assign LUT_2[29976] = 32'b11111111111111110100000100001110;
assign LUT_2[29977] = 32'b11111111111111110000111100100111;
assign LUT_2[29978] = 32'b11111111111111111010111101001010;
assign LUT_2[29979] = 32'b11111111111111110111110101100011;
assign LUT_2[29980] = 32'b11111111111111110000100001110110;
assign LUT_2[29981] = 32'b11111111111111101101011010001111;
assign LUT_2[29982] = 32'b11111111111111110111011010110010;
assign LUT_2[29983] = 32'b11111111111111110100010011001011;
assign LUT_2[29984] = 32'b11111111111111111111001010010000;
assign LUT_2[29985] = 32'b11111111111111111100000010101001;
assign LUT_2[29986] = 32'b00000000000000000110000011001100;
assign LUT_2[29987] = 32'b00000000000000000010111011100101;
assign LUT_2[29988] = 32'b11111111111111111011100111111000;
assign LUT_2[29989] = 32'b11111111111111111000100000010001;
assign LUT_2[29990] = 32'b00000000000000000010100000110100;
assign LUT_2[29991] = 32'b11111111111111111111011001001101;
assign LUT_2[29992] = 32'b11111111111111111001111011101101;
assign LUT_2[29993] = 32'b11111111111111110110110100000110;
assign LUT_2[29994] = 32'b00000000000000000000110100101001;
assign LUT_2[29995] = 32'b11111111111111111101101101000010;
assign LUT_2[29996] = 32'b11111111111111110110011001010101;
assign LUT_2[29997] = 32'b11111111111111110011010001101110;
assign LUT_2[29998] = 32'b11111111111111111101010010010001;
assign LUT_2[29999] = 32'b11111111111111111010001010101010;
assign LUT_2[30000] = 32'b11111111111111111001101110011010;
assign LUT_2[30001] = 32'b11111111111111110110100110110011;
assign LUT_2[30002] = 32'b00000000000000000000100111010110;
assign LUT_2[30003] = 32'b11111111111111111101011111101111;
assign LUT_2[30004] = 32'b11111111111111110110001100000010;
assign LUT_2[30005] = 32'b11111111111111110011000100011011;
assign LUT_2[30006] = 32'b11111111111111111101000100111110;
assign LUT_2[30007] = 32'b11111111111111111001111101010111;
assign LUT_2[30008] = 32'b11111111111111110100011111110111;
assign LUT_2[30009] = 32'b11111111111111110001011000010000;
assign LUT_2[30010] = 32'b11111111111111111011011000110011;
assign LUT_2[30011] = 32'b11111111111111111000010001001100;
assign LUT_2[30012] = 32'b11111111111111110000111101011111;
assign LUT_2[30013] = 32'b11111111111111101101110101111000;
assign LUT_2[30014] = 32'b11111111111111110111110110011011;
assign LUT_2[30015] = 32'b11111111111111110100101110110100;
assign LUT_2[30016] = 32'b11111111111111110110110111001010;
assign LUT_2[30017] = 32'b11111111111111110011101111100011;
assign LUT_2[30018] = 32'b11111111111111111101110000000110;
assign LUT_2[30019] = 32'b11111111111111111010101000011111;
assign LUT_2[30020] = 32'b11111111111111110011010100110010;
assign LUT_2[30021] = 32'b11111111111111110000001101001011;
assign LUT_2[30022] = 32'b11111111111111111010001101101110;
assign LUT_2[30023] = 32'b11111111111111110111000110000111;
assign LUT_2[30024] = 32'b11111111111111110001101000100111;
assign LUT_2[30025] = 32'b11111111111111101110100001000000;
assign LUT_2[30026] = 32'b11111111111111111000100001100011;
assign LUT_2[30027] = 32'b11111111111111110101011001111100;
assign LUT_2[30028] = 32'b11111111111111101110000110001111;
assign LUT_2[30029] = 32'b11111111111111101010111110101000;
assign LUT_2[30030] = 32'b11111111111111110100111111001011;
assign LUT_2[30031] = 32'b11111111111111110001110111100100;
assign LUT_2[30032] = 32'b11111111111111110001011011010100;
assign LUT_2[30033] = 32'b11111111111111101110010011101101;
assign LUT_2[30034] = 32'b11111111111111111000010100010000;
assign LUT_2[30035] = 32'b11111111111111110101001100101001;
assign LUT_2[30036] = 32'b11111111111111101101111000111100;
assign LUT_2[30037] = 32'b11111111111111101010110001010101;
assign LUT_2[30038] = 32'b11111111111111110100110001111000;
assign LUT_2[30039] = 32'b11111111111111110001101010010001;
assign LUT_2[30040] = 32'b11111111111111101100001100110001;
assign LUT_2[30041] = 32'b11111111111111101001000101001010;
assign LUT_2[30042] = 32'b11111111111111110011000101101101;
assign LUT_2[30043] = 32'b11111111111111101111111110000110;
assign LUT_2[30044] = 32'b11111111111111101000101010011001;
assign LUT_2[30045] = 32'b11111111111111100101100010110010;
assign LUT_2[30046] = 32'b11111111111111101111100011010101;
assign LUT_2[30047] = 32'b11111111111111101100011011101110;
assign LUT_2[30048] = 32'b11111111111111110111010010110011;
assign LUT_2[30049] = 32'b11111111111111110100001011001100;
assign LUT_2[30050] = 32'b11111111111111111110001011101111;
assign LUT_2[30051] = 32'b11111111111111111011000100001000;
assign LUT_2[30052] = 32'b11111111111111110011110000011011;
assign LUT_2[30053] = 32'b11111111111111110000101000110100;
assign LUT_2[30054] = 32'b11111111111111111010101001010111;
assign LUT_2[30055] = 32'b11111111111111110111100001110000;
assign LUT_2[30056] = 32'b11111111111111110010000100010000;
assign LUT_2[30057] = 32'b11111111111111101110111100101001;
assign LUT_2[30058] = 32'b11111111111111111000111101001100;
assign LUT_2[30059] = 32'b11111111111111110101110101100101;
assign LUT_2[30060] = 32'b11111111111111101110100001111000;
assign LUT_2[30061] = 32'b11111111111111101011011010010001;
assign LUT_2[30062] = 32'b11111111111111110101011010110100;
assign LUT_2[30063] = 32'b11111111111111110010010011001101;
assign LUT_2[30064] = 32'b11111111111111110001110110111101;
assign LUT_2[30065] = 32'b11111111111111101110101111010110;
assign LUT_2[30066] = 32'b11111111111111111000101111111001;
assign LUT_2[30067] = 32'b11111111111111110101101000010010;
assign LUT_2[30068] = 32'b11111111111111101110010100100101;
assign LUT_2[30069] = 32'b11111111111111101011001100111110;
assign LUT_2[30070] = 32'b11111111111111110101001101100001;
assign LUT_2[30071] = 32'b11111111111111110010000101111010;
assign LUT_2[30072] = 32'b11111111111111101100101000011010;
assign LUT_2[30073] = 32'b11111111111111101001100000110011;
assign LUT_2[30074] = 32'b11111111111111110011100001010110;
assign LUT_2[30075] = 32'b11111111111111110000011001101111;
assign LUT_2[30076] = 32'b11111111111111101001000110000010;
assign LUT_2[30077] = 32'b11111111111111100101111110011011;
assign LUT_2[30078] = 32'b11111111111111101111111110111110;
assign LUT_2[30079] = 32'b11111111111111101100110111010111;
assign LUT_2[30080] = 32'b00000000000000000011000010110110;
assign LUT_2[30081] = 32'b11111111111111111111111011001111;
assign LUT_2[30082] = 32'b00000000000000001001111011110010;
assign LUT_2[30083] = 32'b00000000000000000110110100001011;
assign LUT_2[30084] = 32'b11111111111111111111100000011110;
assign LUT_2[30085] = 32'b11111111111111111100011000110111;
assign LUT_2[30086] = 32'b00000000000000000110011001011010;
assign LUT_2[30087] = 32'b00000000000000000011010001110011;
assign LUT_2[30088] = 32'b11111111111111111101110100010011;
assign LUT_2[30089] = 32'b11111111111111111010101100101100;
assign LUT_2[30090] = 32'b00000000000000000100101101001111;
assign LUT_2[30091] = 32'b00000000000000000001100101101000;
assign LUT_2[30092] = 32'b11111111111111111010010001111011;
assign LUT_2[30093] = 32'b11111111111111110111001010010100;
assign LUT_2[30094] = 32'b00000000000000000001001010110111;
assign LUT_2[30095] = 32'b11111111111111111110000011010000;
assign LUT_2[30096] = 32'b11111111111111111101100111000000;
assign LUT_2[30097] = 32'b11111111111111111010011111011001;
assign LUT_2[30098] = 32'b00000000000000000100011111111100;
assign LUT_2[30099] = 32'b00000000000000000001011000010101;
assign LUT_2[30100] = 32'b11111111111111111010000100101000;
assign LUT_2[30101] = 32'b11111111111111110110111101000001;
assign LUT_2[30102] = 32'b00000000000000000000111101100100;
assign LUT_2[30103] = 32'b11111111111111111101110101111101;
assign LUT_2[30104] = 32'b11111111111111111000011000011101;
assign LUT_2[30105] = 32'b11111111111111110101010000110110;
assign LUT_2[30106] = 32'b11111111111111111111010001011001;
assign LUT_2[30107] = 32'b11111111111111111100001001110010;
assign LUT_2[30108] = 32'b11111111111111110100110110000101;
assign LUT_2[30109] = 32'b11111111111111110001101110011110;
assign LUT_2[30110] = 32'b11111111111111111011101111000001;
assign LUT_2[30111] = 32'b11111111111111111000100111011010;
assign LUT_2[30112] = 32'b00000000000000000011011110011111;
assign LUT_2[30113] = 32'b00000000000000000000010110111000;
assign LUT_2[30114] = 32'b00000000000000001010010111011011;
assign LUT_2[30115] = 32'b00000000000000000111001111110100;
assign LUT_2[30116] = 32'b11111111111111111111111100000111;
assign LUT_2[30117] = 32'b11111111111111111100110100100000;
assign LUT_2[30118] = 32'b00000000000000000110110101000011;
assign LUT_2[30119] = 32'b00000000000000000011101101011100;
assign LUT_2[30120] = 32'b11111111111111111110001111111100;
assign LUT_2[30121] = 32'b11111111111111111011001000010101;
assign LUT_2[30122] = 32'b00000000000000000101001000111000;
assign LUT_2[30123] = 32'b00000000000000000010000001010001;
assign LUT_2[30124] = 32'b11111111111111111010101101100100;
assign LUT_2[30125] = 32'b11111111111111110111100101111101;
assign LUT_2[30126] = 32'b00000000000000000001100110100000;
assign LUT_2[30127] = 32'b11111111111111111110011110111001;
assign LUT_2[30128] = 32'b11111111111111111110000010101001;
assign LUT_2[30129] = 32'b11111111111111111010111011000010;
assign LUT_2[30130] = 32'b00000000000000000100111011100101;
assign LUT_2[30131] = 32'b00000000000000000001110011111110;
assign LUT_2[30132] = 32'b11111111111111111010100000010001;
assign LUT_2[30133] = 32'b11111111111111110111011000101010;
assign LUT_2[30134] = 32'b00000000000000000001011001001101;
assign LUT_2[30135] = 32'b11111111111111111110010001100110;
assign LUT_2[30136] = 32'b11111111111111111000110100000110;
assign LUT_2[30137] = 32'b11111111111111110101101100011111;
assign LUT_2[30138] = 32'b11111111111111111111101101000010;
assign LUT_2[30139] = 32'b11111111111111111100100101011011;
assign LUT_2[30140] = 32'b11111111111111110101010001101110;
assign LUT_2[30141] = 32'b11111111111111110010001010000111;
assign LUT_2[30142] = 32'b11111111111111111100001010101010;
assign LUT_2[30143] = 32'b11111111111111111001000011000011;
assign LUT_2[30144] = 32'b11111111111111111011001011011001;
assign LUT_2[30145] = 32'b11111111111111111000000011110010;
assign LUT_2[30146] = 32'b00000000000000000010000100010101;
assign LUT_2[30147] = 32'b11111111111111111110111100101110;
assign LUT_2[30148] = 32'b11111111111111110111101001000001;
assign LUT_2[30149] = 32'b11111111111111110100100001011010;
assign LUT_2[30150] = 32'b11111111111111111110100001111101;
assign LUT_2[30151] = 32'b11111111111111111011011010010110;
assign LUT_2[30152] = 32'b11111111111111110101111100110110;
assign LUT_2[30153] = 32'b11111111111111110010110101001111;
assign LUT_2[30154] = 32'b11111111111111111100110101110010;
assign LUT_2[30155] = 32'b11111111111111111001101110001011;
assign LUT_2[30156] = 32'b11111111111111110010011010011110;
assign LUT_2[30157] = 32'b11111111111111101111010010110111;
assign LUT_2[30158] = 32'b11111111111111111001010011011010;
assign LUT_2[30159] = 32'b11111111111111110110001011110011;
assign LUT_2[30160] = 32'b11111111111111110101101111100011;
assign LUT_2[30161] = 32'b11111111111111110010100111111100;
assign LUT_2[30162] = 32'b11111111111111111100101000011111;
assign LUT_2[30163] = 32'b11111111111111111001100000111000;
assign LUT_2[30164] = 32'b11111111111111110010001101001011;
assign LUT_2[30165] = 32'b11111111111111101111000101100100;
assign LUT_2[30166] = 32'b11111111111111111001000110000111;
assign LUT_2[30167] = 32'b11111111111111110101111110100000;
assign LUT_2[30168] = 32'b11111111111111110000100001000000;
assign LUT_2[30169] = 32'b11111111111111101101011001011001;
assign LUT_2[30170] = 32'b11111111111111110111011001111100;
assign LUT_2[30171] = 32'b11111111111111110100010010010101;
assign LUT_2[30172] = 32'b11111111111111101100111110101000;
assign LUT_2[30173] = 32'b11111111111111101001110111000001;
assign LUT_2[30174] = 32'b11111111111111110011110111100100;
assign LUT_2[30175] = 32'b11111111111111110000101111111101;
assign LUT_2[30176] = 32'b11111111111111111011100111000010;
assign LUT_2[30177] = 32'b11111111111111111000011111011011;
assign LUT_2[30178] = 32'b00000000000000000010011111111110;
assign LUT_2[30179] = 32'b11111111111111111111011000010111;
assign LUT_2[30180] = 32'b11111111111111111000000100101010;
assign LUT_2[30181] = 32'b11111111111111110100111101000011;
assign LUT_2[30182] = 32'b11111111111111111110111101100110;
assign LUT_2[30183] = 32'b11111111111111111011110101111111;
assign LUT_2[30184] = 32'b11111111111111110110011000011111;
assign LUT_2[30185] = 32'b11111111111111110011010000111000;
assign LUT_2[30186] = 32'b11111111111111111101010001011011;
assign LUT_2[30187] = 32'b11111111111111111010001001110100;
assign LUT_2[30188] = 32'b11111111111111110010110110000111;
assign LUT_2[30189] = 32'b11111111111111101111101110100000;
assign LUT_2[30190] = 32'b11111111111111111001101111000011;
assign LUT_2[30191] = 32'b11111111111111110110100111011100;
assign LUT_2[30192] = 32'b11111111111111110110001011001100;
assign LUT_2[30193] = 32'b11111111111111110011000011100101;
assign LUT_2[30194] = 32'b11111111111111111101000100001000;
assign LUT_2[30195] = 32'b11111111111111111001111100100001;
assign LUT_2[30196] = 32'b11111111111111110010101000110100;
assign LUT_2[30197] = 32'b11111111111111101111100001001101;
assign LUT_2[30198] = 32'b11111111111111111001100001110000;
assign LUT_2[30199] = 32'b11111111111111110110011010001001;
assign LUT_2[30200] = 32'b11111111111111110000111100101001;
assign LUT_2[30201] = 32'b11111111111111101101110101000010;
assign LUT_2[30202] = 32'b11111111111111110111110101100101;
assign LUT_2[30203] = 32'b11111111111111110100101101111110;
assign LUT_2[30204] = 32'b11111111111111101101011010010001;
assign LUT_2[30205] = 32'b11111111111111101010010010101010;
assign LUT_2[30206] = 32'b11111111111111110100010011001101;
assign LUT_2[30207] = 32'b11111111111111110001001011100110;
assign LUT_2[30208] = 32'b11111111111111111111100001110011;
assign LUT_2[30209] = 32'b11111111111111111100011010001100;
assign LUT_2[30210] = 32'b00000000000000000110011010101111;
assign LUT_2[30211] = 32'b00000000000000000011010011001000;
assign LUT_2[30212] = 32'b11111111111111111011111111011011;
assign LUT_2[30213] = 32'b11111111111111111000110111110100;
assign LUT_2[30214] = 32'b00000000000000000010111000010111;
assign LUT_2[30215] = 32'b11111111111111111111110000110000;
assign LUT_2[30216] = 32'b11111111111111111010010011010000;
assign LUT_2[30217] = 32'b11111111111111110111001011101001;
assign LUT_2[30218] = 32'b00000000000000000001001100001100;
assign LUT_2[30219] = 32'b11111111111111111110000100100101;
assign LUT_2[30220] = 32'b11111111111111110110110000111000;
assign LUT_2[30221] = 32'b11111111111111110011101001010001;
assign LUT_2[30222] = 32'b11111111111111111101101001110100;
assign LUT_2[30223] = 32'b11111111111111111010100010001101;
assign LUT_2[30224] = 32'b11111111111111111010000101111101;
assign LUT_2[30225] = 32'b11111111111111110110111110010110;
assign LUT_2[30226] = 32'b00000000000000000000111110111001;
assign LUT_2[30227] = 32'b11111111111111111101110111010010;
assign LUT_2[30228] = 32'b11111111111111110110100011100101;
assign LUT_2[30229] = 32'b11111111111111110011011011111110;
assign LUT_2[30230] = 32'b11111111111111111101011100100001;
assign LUT_2[30231] = 32'b11111111111111111010010100111010;
assign LUT_2[30232] = 32'b11111111111111110100110111011010;
assign LUT_2[30233] = 32'b11111111111111110001101111110011;
assign LUT_2[30234] = 32'b11111111111111111011110000010110;
assign LUT_2[30235] = 32'b11111111111111111000101000101111;
assign LUT_2[30236] = 32'b11111111111111110001010101000010;
assign LUT_2[30237] = 32'b11111111111111101110001101011011;
assign LUT_2[30238] = 32'b11111111111111111000001101111110;
assign LUT_2[30239] = 32'b11111111111111110101000110010111;
assign LUT_2[30240] = 32'b11111111111111111111111101011100;
assign LUT_2[30241] = 32'b11111111111111111100110101110101;
assign LUT_2[30242] = 32'b00000000000000000110110110011000;
assign LUT_2[30243] = 32'b00000000000000000011101110110001;
assign LUT_2[30244] = 32'b11111111111111111100011011000100;
assign LUT_2[30245] = 32'b11111111111111111001010011011101;
assign LUT_2[30246] = 32'b00000000000000000011010100000000;
assign LUT_2[30247] = 32'b00000000000000000000001100011001;
assign LUT_2[30248] = 32'b11111111111111111010101110111001;
assign LUT_2[30249] = 32'b11111111111111110111100111010010;
assign LUT_2[30250] = 32'b00000000000000000001100111110101;
assign LUT_2[30251] = 32'b11111111111111111110100000001110;
assign LUT_2[30252] = 32'b11111111111111110111001100100001;
assign LUT_2[30253] = 32'b11111111111111110100000100111010;
assign LUT_2[30254] = 32'b11111111111111111110000101011101;
assign LUT_2[30255] = 32'b11111111111111111010111101110110;
assign LUT_2[30256] = 32'b11111111111111111010100001100110;
assign LUT_2[30257] = 32'b11111111111111110111011001111111;
assign LUT_2[30258] = 32'b00000000000000000001011010100010;
assign LUT_2[30259] = 32'b11111111111111111110010010111011;
assign LUT_2[30260] = 32'b11111111111111110110111111001110;
assign LUT_2[30261] = 32'b11111111111111110011110111100111;
assign LUT_2[30262] = 32'b11111111111111111101111000001010;
assign LUT_2[30263] = 32'b11111111111111111010110000100011;
assign LUT_2[30264] = 32'b11111111111111110101010011000011;
assign LUT_2[30265] = 32'b11111111111111110010001011011100;
assign LUT_2[30266] = 32'b11111111111111111100001011111111;
assign LUT_2[30267] = 32'b11111111111111111001000100011000;
assign LUT_2[30268] = 32'b11111111111111110001110000101011;
assign LUT_2[30269] = 32'b11111111111111101110101001000100;
assign LUT_2[30270] = 32'b11111111111111111000101001100111;
assign LUT_2[30271] = 32'b11111111111111110101100010000000;
assign LUT_2[30272] = 32'b11111111111111110111101010010110;
assign LUT_2[30273] = 32'b11111111111111110100100010101111;
assign LUT_2[30274] = 32'b11111111111111111110100011010010;
assign LUT_2[30275] = 32'b11111111111111111011011011101011;
assign LUT_2[30276] = 32'b11111111111111110100000111111110;
assign LUT_2[30277] = 32'b11111111111111110001000000010111;
assign LUT_2[30278] = 32'b11111111111111111011000000111010;
assign LUT_2[30279] = 32'b11111111111111110111111001010011;
assign LUT_2[30280] = 32'b11111111111111110010011011110011;
assign LUT_2[30281] = 32'b11111111111111101111010100001100;
assign LUT_2[30282] = 32'b11111111111111111001010100101111;
assign LUT_2[30283] = 32'b11111111111111110110001101001000;
assign LUT_2[30284] = 32'b11111111111111101110111001011011;
assign LUT_2[30285] = 32'b11111111111111101011110001110100;
assign LUT_2[30286] = 32'b11111111111111110101110010010111;
assign LUT_2[30287] = 32'b11111111111111110010101010110000;
assign LUT_2[30288] = 32'b11111111111111110010001110100000;
assign LUT_2[30289] = 32'b11111111111111101111000110111001;
assign LUT_2[30290] = 32'b11111111111111111001000111011100;
assign LUT_2[30291] = 32'b11111111111111110101111111110101;
assign LUT_2[30292] = 32'b11111111111111101110101100001000;
assign LUT_2[30293] = 32'b11111111111111101011100100100001;
assign LUT_2[30294] = 32'b11111111111111110101100101000100;
assign LUT_2[30295] = 32'b11111111111111110010011101011101;
assign LUT_2[30296] = 32'b11111111111111101100111111111101;
assign LUT_2[30297] = 32'b11111111111111101001111000010110;
assign LUT_2[30298] = 32'b11111111111111110011111000111001;
assign LUT_2[30299] = 32'b11111111111111110000110001010010;
assign LUT_2[30300] = 32'b11111111111111101001011101100101;
assign LUT_2[30301] = 32'b11111111111111100110010101111110;
assign LUT_2[30302] = 32'b11111111111111110000010110100001;
assign LUT_2[30303] = 32'b11111111111111101101001110111010;
assign LUT_2[30304] = 32'b11111111111111111000000101111111;
assign LUT_2[30305] = 32'b11111111111111110100111110011000;
assign LUT_2[30306] = 32'b11111111111111111110111110111011;
assign LUT_2[30307] = 32'b11111111111111111011110111010100;
assign LUT_2[30308] = 32'b11111111111111110100100011100111;
assign LUT_2[30309] = 32'b11111111111111110001011100000000;
assign LUT_2[30310] = 32'b11111111111111111011011100100011;
assign LUT_2[30311] = 32'b11111111111111111000010100111100;
assign LUT_2[30312] = 32'b11111111111111110010110111011100;
assign LUT_2[30313] = 32'b11111111111111101111101111110101;
assign LUT_2[30314] = 32'b11111111111111111001110000011000;
assign LUT_2[30315] = 32'b11111111111111110110101000110001;
assign LUT_2[30316] = 32'b11111111111111101111010101000100;
assign LUT_2[30317] = 32'b11111111111111101100001101011101;
assign LUT_2[30318] = 32'b11111111111111110110001110000000;
assign LUT_2[30319] = 32'b11111111111111110011000110011001;
assign LUT_2[30320] = 32'b11111111111111110010101010001001;
assign LUT_2[30321] = 32'b11111111111111101111100010100010;
assign LUT_2[30322] = 32'b11111111111111111001100011000101;
assign LUT_2[30323] = 32'b11111111111111110110011011011110;
assign LUT_2[30324] = 32'b11111111111111101111000111110001;
assign LUT_2[30325] = 32'b11111111111111101100000000001010;
assign LUT_2[30326] = 32'b11111111111111110110000000101101;
assign LUT_2[30327] = 32'b11111111111111110010111001000110;
assign LUT_2[30328] = 32'b11111111111111101101011011100110;
assign LUT_2[30329] = 32'b11111111111111101010010011111111;
assign LUT_2[30330] = 32'b11111111111111110100010100100010;
assign LUT_2[30331] = 32'b11111111111111110001001100111011;
assign LUT_2[30332] = 32'b11111111111111101001111001001110;
assign LUT_2[30333] = 32'b11111111111111100110110001100111;
assign LUT_2[30334] = 32'b11111111111111110000110010001010;
assign LUT_2[30335] = 32'b11111111111111101101101010100011;
assign LUT_2[30336] = 32'b00000000000000000011110110000010;
assign LUT_2[30337] = 32'b00000000000000000000101110011011;
assign LUT_2[30338] = 32'b00000000000000001010101110111110;
assign LUT_2[30339] = 32'b00000000000000000111100111010111;
assign LUT_2[30340] = 32'b00000000000000000000010011101010;
assign LUT_2[30341] = 32'b11111111111111111101001100000011;
assign LUT_2[30342] = 32'b00000000000000000111001100100110;
assign LUT_2[30343] = 32'b00000000000000000100000100111111;
assign LUT_2[30344] = 32'b11111111111111111110100111011111;
assign LUT_2[30345] = 32'b11111111111111111011011111111000;
assign LUT_2[30346] = 32'b00000000000000000101100000011011;
assign LUT_2[30347] = 32'b00000000000000000010011000110100;
assign LUT_2[30348] = 32'b11111111111111111011000101000111;
assign LUT_2[30349] = 32'b11111111111111110111111101100000;
assign LUT_2[30350] = 32'b00000000000000000001111110000011;
assign LUT_2[30351] = 32'b11111111111111111110110110011100;
assign LUT_2[30352] = 32'b11111111111111111110011010001100;
assign LUT_2[30353] = 32'b11111111111111111011010010100101;
assign LUT_2[30354] = 32'b00000000000000000101010011001000;
assign LUT_2[30355] = 32'b00000000000000000010001011100001;
assign LUT_2[30356] = 32'b11111111111111111010110111110100;
assign LUT_2[30357] = 32'b11111111111111110111110000001101;
assign LUT_2[30358] = 32'b00000000000000000001110000110000;
assign LUT_2[30359] = 32'b11111111111111111110101001001001;
assign LUT_2[30360] = 32'b11111111111111111001001011101001;
assign LUT_2[30361] = 32'b11111111111111110110000100000010;
assign LUT_2[30362] = 32'b00000000000000000000000100100101;
assign LUT_2[30363] = 32'b11111111111111111100111100111110;
assign LUT_2[30364] = 32'b11111111111111110101101001010001;
assign LUT_2[30365] = 32'b11111111111111110010100001101010;
assign LUT_2[30366] = 32'b11111111111111111100100010001101;
assign LUT_2[30367] = 32'b11111111111111111001011010100110;
assign LUT_2[30368] = 32'b00000000000000000100010001101011;
assign LUT_2[30369] = 32'b00000000000000000001001010000100;
assign LUT_2[30370] = 32'b00000000000000001011001010100111;
assign LUT_2[30371] = 32'b00000000000000001000000011000000;
assign LUT_2[30372] = 32'b00000000000000000000101111010011;
assign LUT_2[30373] = 32'b11111111111111111101100111101100;
assign LUT_2[30374] = 32'b00000000000000000111101000001111;
assign LUT_2[30375] = 32'b00000000000000000100100000101000;
assign LUT_2[30376] = 32'b11111111111111111111000011001000;
assign LUT_2[30377] = 32'b11111111111111111011111011100001;
assign LUT_2[30378] = 32'b00000000000000000101111100000100;
assign LUT_2[30379] = 32'b00000000000000000010110100011101;
assign LUT_2[30380] = 32'b11111111111111111011100000110000;
assign LUT_2[30381] = 32'b11111111111111111000011001001001;
assign LUT_2[30382] = 32'b00000000000000000010011001101100;
assign LUT_2[30383] = 32'b11111111111111111111010010000101;
assign LUT_2[30384] = 32'b11111111111111111110110101110101;
assign LUT_2[30385] = 32'b11111111111111111011101110001110;
assign LUT_2[30386] = 32'b00000000000000000101101110110001;
assign LUT_2[30387] = 32'b00000000000000000010100111001010;
assign LUT_2[30388] = 32'b11111111111111111011010011011101;
assign LUT_2[30389] = 32'b11111111111111111000001011110110;
assign LUT_2[30390] = 32'b00000000000000000010001100011001;
assign LUT_2[30391] = 32'b11111111111111111111000100110010;
assign LUT_2[30392] = 32'b11111111111111111001100111010010;
assign LUT_2[30393] = 32'b11111111111111110110011111101011;
assign LUT_2[30394] = 32'b00000000000000000000100000001110;
assign LUT_2[30395] = 32'b11111111111111111101011000100111;
assign LUT_2[30396] = 32'b11111111111111110110000100111010;
assign LUT_2[30397] = 32'b11111111111111110010111101010011;
assign LUT_2[30398] = 32'b11111111111111111100111101110110;
assign LUT_2[30399] = 32'b11111111111111111001110110001111;
assign LUT_2[30400] = 32'b11111111111111111011111110100101;
assign LUT_2[30401] = 32'b11111111111111111000110110111110;
assign LUT_2[30402] = 32'b00000000000000000010110111100001;
assign LUT_2[30403] = 32'b11111111111111111111101111111010;
assign LUT_2[30404] = 32'b11111111111111111000011100001101;
assign LUT_2[30405] = 32'b11111111111111110101010100100110;
assign LUT_2[30406] = 32'b11111111111111111111010101001001;
assign LUT_2[30407] = 32'b11111111111111111100001101100010;
assign LUT_2[30408] = 32'b11111111111111110110110000000010;
assign LUT_2[30409] = 32'b11111111111111110011101000011011;
assign LUT_2[30410] = 32'b11111111111111111101101000111110;
assign LUT_2[30411] = 32'b11111111111111111010100001010111;
assign LUT_2[30412] = 32'b11111111111111110011001101101010;
assign LUT_2[30413] = 32'b11111111111111110000000110000011;
assign LUT_2[30414] = 32'b11111111111111111010000110100110;
assign LUT_2[30415] = 32'b11111111111111110110111110111111;
assign LUT_2[30416] = 32'b11111111111111110110100010101111;
assign LUT_2[30417] = 32'b11111111111111110011011011001000;
assign LUT_2[30418] = 32'b11111111111111111101011011101011;
assign LUT_2[30419] = 32'b11111111111111111010010100000100;
assign LUT_2[30420] = 32'b11111111111111110011000000010111;
assign LUT_2[30421] = 32'b11111111111111101111111000110000;
assign LUT_2[30422] = 32'b11111111111111111001111001010011;
assign LUT_2[30423] = 32'b11111111111111110110110001101100;
assign LUT_2[30424] = 32'b11111111111111110001010100001100;
assign LUT_2[30425] = 32'b11111111111111101110001100100101;
assign LUT_2[30426] = 32'b11111111111111111000001101001000;
assign LUT_2[30427] = 32'b11111111111111110101000101100001;
assign LUT_2[30428] = 32'b11111111111111101101110001110100;
assign LUT_2[30429] = 32'b11111111111111101010101010001101;
assign LUT_2[30430] = 32'b11111111111111110100101010110000;
assign LUT_2[30431] = 32'b11111111111111110001100011001001;
assign LUT_2[30432] = 32'b11111111111111111100011010001110;
assign LUT_2[30433] = 32'b11111111111111111001010010100111;
assign LUT_2[30434] = 32'b00000000000000000011010011001010;
assign LUT_2[30435] = 32'b00000000000000000000001011100011;
assign LUT_2[30436] = 32'b11111111111111111000110111110110;
assign LUT_2[30437] = 32'b11111111111111110101110000001111;
assign LUT_2[30438] = 32'b11111111111111111111110000110010;
assign LUT_2[30439] = 32'b11111111111111111100101001001011;
assign LUT_2[30440] = 32'b11111111111111110111001011101011;
assign LUT_2[30441] = 32'b11111111111111110100000100000100;
assign LUT_2[30442] = 32'b11111111111111111110000100100111;
assign LUT_2[30443] = 32'b11111111111111111010111101000000;
assign LUT_2[30444] = 32'b11111111111111110011101001010011;
assign LUT_2[30445] = 32'b11111111111111110000100001101100;
assign LUT_2[30446] = 32'b11111111111111111010100010001111;
assign LUT_2[30447] = 32'b11111111111111110111011010101000;
assign LUT_2[30448] = 32'b11111111111111110110111110011000;
assign LUT_2[30449] = 32'b11111111111111110011110110110001;
assign LUT_2[30450] = 32'b11111111111111111101110111010100;
assign LUT_2[30451] = 32'b11111111111111111010101111101101;
assign LUT_2[30452] = 32'b11111111111111110011011100000000;
assign LUT_2[30453] = 32'b11111111111111110000010100011001;
assign LUT_2[30454] = 32'b11111111111111111010010100111100;
assign LUT_2[30455] = 32'b11111111111111110111001101010101;
assign LUT_2[30456] = 32'b11111111111111110001101111110101;
assign LUT_2[30457] = 32'b11111111111111101110101000001110;
assign LUT_2[30458] = 32'b11111111111111111000101000110001;
assign LUT_2[30459] = 32'b11111111111111110101100001001010;
assign LUT_2[30460] = 32'b11111111111111101110001101011101;
assign LUT_2[30461] = 32'b11111111111111101011000101110110;
assign LUT_2[30462] = 32'b11111111111111110101000110011001;
assign LUT_2[30463] = 32'b11111111111111110001111110110010;
assign LUT_2[30464] = 32'b00000000000000000011100000011001;
assign LUT_2[30465] = 32'b00000000000000000000011000110010;
assign LUT_2[30466] = 32'b00000000000000001010011001010101;
assign LUT_2[30467] = 32'b00000000000000000111010001101110;
assign LUT_2[30468] = 32'b11111111111111111111111110000001;
assign LUT_2[30469] = 32'b11111111111111111100110110011010;
assign LUT_2[30470] = 32'b00000000000000000110110110111101;
assign LUT_2[30471] = 32'b00000000000000000011101111010110;
assign LUT_2[30472] = 32'b11111111111111111110010001110110;
assign LUT_2[30473] = 32'b11111111111111111011001010001111;
assign LUT_2[30474] = 32'b00000000000000000101001010110010;
assign LUT_2[30475] = 32'b00000000000000000010000011001011;
assign LUT_2[30476] = 32'b11111111111111111010101111011110;
assign LUT_2[30477] = 32'b11111111111111110111100111110111;
assign LUT_2[30478] = 32'b00000000000000000001101000011010;
assign LUT_2[30479] = 32'b11111111111111111110100000110011;
assign LUT_2[30480] = 32'b11111111111111111110000100100011;
assign LUT_2[30481] = 32'b11111111111111111010111100111100;
assign LUT_2[30482] = 32'b00000000000000000100111101011111;
assign LUT_2[30483] = 32'b00000000000000000001110101111000;
assign LUT_2[30484] = 32'b11111111111111111010100010001011;
assign LUT_2[30485] = 32'b11111111111111110111011010100100;
assign LUT_2[30486] = 32'b00000000000000000001011011000111;
assign LUT_2[30487] = 32'b11111111111111111110010011100000;
assign LUT_2[30488] = 32'b11111111111111111000110110000000;
assign LUT_2[30489] = 32'b11111111111111110101101110011001;
assign LUT_2[30490] = 32'b11111111111111111111101110111100;
assign LUT_2[30491] = 32'b11111111111111111100100111010101;
assign LUT_2[30492] = 32'b11111111111111110101010011101000;
assign LUT_2[30493] = 32'b11111111111111110010001100000001;
assign LUT_2[30494] = 32'b11111111111111111100001100100100;
assign LUT_2[30495] = 32'b11111111111111111001000100111101;
assign LUT_2[30496] = 32'b00000000000000000011111100000010;
assign LUT_2[30497] = 32'b00000000000000000000110100011011;
assign LUT_2[30498] = 32'b00000000000000001010110100111110;
assign LUT_2[30499] = 32'b00000000000000000111101101010111;
assign LUT_2[30500] = 32'b00000000000000000000011001101010;
assign LUT_2[30501] = 32'b11111111111111111101010010000011;
assign LUT_2[30502] = 32'b00000000000000000111010010100110;
assign LUT_2[30503] = 32'b00000000000000000100001010111111;
assign LUT_2[30504] = 32'b11111111111111111110101101011111;
assign LUT_2[30505] = 32'b11111111111111111011100101111000;
assign LUT_2[30506] = 32'b00000000000000000101100110011011;
assign LUT_2[30507] = 32'b00000000000000000010011110110100;
assign LUT_2[30508] = 32'b11111111111111111011001011000111;
assign LUT_2[30509] = 32'b11111111111111111000000011100000;
assign LUT_2[30510] = 32'b00000000000000000010000100000011;
assign LUT_2[30511] = 32'b11111111111111111110111100011100;
assign LUT_2[30512] = 32'b11111111111111111110100000001100;
assign LUT_2[30513] = 32'b11111111111111111011011000100101;
assign LUT_2[30514] = 32'b00000000000000000101011001001000;
assign LUT_2[30515] = 32'b00000000000000000010010001100001;
assign LUT_2[30516] = 32'b11111111111111111010111101110100;
assign LUT_2[30517] = 32'b11111111111111110111110110001101;
assign LUT_2[30518] = 32'b00000000000000000001110110110000;
assign LUT_2[30519] = 32'b11111111111111111110101111001001;
assign LUT_2[30520] = 32'b11111111111111111001010001101001;
assign LUT_2[30521] = 32'b11111111111111110110001010000010;
assign LUT_2[30522] = 32'b00000000000000000000001010100101;
assign LUT_2[30523] = 32'b11111111111111111101000010111110;
assign LUT_2[30524] = 32'b11111111111111110101101111010001;
assign LUT_2[30525] = 32'b11111111111111110010100111101010;
assign LUT_2[30526] = 32'b11111111111111111100101000001101;
assign LUT_2[30527] = 32'b11111111111111111001100000100110;
assign LUT_2[30528] = 32'b11111111111111111011101000111100;
assign LUT_2[30529] = 32'b11111111111111111000100001010101;
assign LUT_2[30530] = 32'b00000000000000000010100001111000;
assign LUT_2[30531] = 32'b11111111111111111111011010010001;
assign LUT_2[30532] = 32'b11111111111111111000000110100100;
assign LUT_2[30533] = 32'b11111111111111110100111110111101;
assign LUT_2[30534] = 32'b11111111111111111110111111100000;
assign LUT_2[30535] = 32'b11111111111111111011110111111001;
assign LUT_2[30536] = 32'b11111111111111110110011010011001;
assign LUT_2[30537] = 32'b11111111111111110011010010110010;
assign LUT_2[30538] = 32'b11111111111111111101010011010101;
assign LUT_2[30539] = 32'b11111111111111111010001011101110;
assign LUT_2[30540] = 32'b11111111111111110010111000000001;
assign LUT_2[30541] = 32'b11111111111111101111110000011010;
assign LUT_2[30542] = 32'b11111111111111111001110000111101;
assign LUT_2[30543] = 32'b11111111111111110110101001010110;
assign LUT_2[30544] = 32'b11111111111111110110001101000110;
assign LUT_2[30545] = 32'b11111111111111110011000101011111;
assign LUT_2[30546] = 32'b11111111111111111101000110000010;
assign LUT_2[30547] = 32'b11111111111111111001111110011011;
assign LUT_2[30548] = 32'b11111111111111110010101010101110;
assign LUT_2[30549] = 32'b11111111111111101111100011000111;
assign LUT_2[30550] = 32'b11111111111111111001100011101010;
assign LUT_2[30551] = 32'b11111111111111110110011100000011;
assign LUT_2[30552] = 32'b11111111111111110000111110100011;
assign LUT_2[30553] = 32'b11111111111111101101110110111100;
assign LUT_2[30554] = 32'b11111111111111110111110111011111;
assign LUT_2[30555] = 32'b11111111111111110100101111111000;
assign LUT_2[30556] = 32'b11111111111111101101011100001011;
assign LUT_2[30557] = 32'b11111111111111101010010100100100;
assign LUT_2[30558] = 32'b11111111111111110100010101000111;
assign LUT_2[30559] = 32'b11111111111111110001001101100000;
assign LUT_2[30560] = 32'b11111111111111111100000100100101;
assign LUT_2[30561] = 32'b11111111111111111000111100111110;
assign LUT_2[30562] = 32'b00000000000000000010111101100001;
assign LUT_2[30563] = 32'b11111111111111111111110101111010;
assign LUT_2[30564] = 32'b11111111111111111000100010001101;
assign LUT_2[30565] = 32'b11111111111111110101011010100110;
assign LUT_2[30566] = 32'b11111111111111111111011011001001;
assign LUT_2[30567] = 32'b11111111111111111100010011100010;
assign LUT_2[30568] = 32'b11111111111111110110110110000010;
assign LUT_2[30569] = 32'b11111111111111110011101110011011;
assign LUT_2[30570] = 32'b11111111111111111101101110111110;
assign LUT_2[30571] = 32'b11111111111111111010100111010111;
assign LUT_2[30572] = 32'b11111111111111110011010011101010;
assign LUT_2[30573] = 32'b11111111111111110000001100000011;
assign LUT_2[30574] = 32'b11111111111111111010001100100110;
assign LUT_2[30575] = 32'b11111111111111110111000100111111;
assign LUT_2[30576] = 32'b11111111111111110110101000101111;
assign LUT_2[30577] = 32'b11111111111111110011100001001000;
assign LUT_2[30578] = 32'b11111111111111111101100001101011;
assign LUT_2[30579] = 32'b11111111111111111010011010000100;
assign LUT_2[30580] = 32'b11111111111111110011000110010111;
assign LUT_2[30581] = 32'b11111111111111101111111110110000;
assign LUT_2[30582] = 32'b11111111111111111001111111010011;
assign LUT_2[30583] = 32'b11111111111111110110110111101100;
assign LUT_2[30584] = 32'b11111111111111110001011010001100;
assign LUT_2[30585] = 32'b11111111111111101110010010100101;
assign LUT_2[30586] = 32'b11111111111111111000010011001000;
assign LUT_2[30587] = 32'b11111111111111110101001011100001;
assign LUT_2[30588] = 32'b11111111111111101101110111110100;
assign LUT_2[30589] = 32'b11111111111111101010110000001101;
assign LUT_2[30590] = 32'b11111111111111110100110000110000;
assign LUT_2[30591] = 32'b11111111111111110001101001001001;
assign LUT_2[30592] = 32'b00000000000000000111110100101000;
assign LUT_2[30593] = 32'b00000000000000000100101101000001;
assign LUT_2[30594] = 32'b00000000000000001110101101100100;
assign LUT_2[30595] = 32'b00000000000000001011100101111101;
assign LUT_2[30596] = 32'b00000000000000000100010010010000;
assign LUT_2[30597] = 32'b00000000000000000001001010101001;
assign LUT_2[30598] = 32'b00000000000000001011001011001100;
assign LUT_2[30599] = 32'b00000000000000001000000011100101;
assign LUT_2[30600] = 32'b00000000000000000010100110000101;
assign LUT_2[30601] = 32'b11111111111111111111011110011110;
assign LUT_2[30602] = 32'b00000000000000001001011111000001;
assign LUT_2[30603] = 32'b00000000000000000110010111011010;
assign LUT_2[30604] = 32'b11111111111111111111000011101101;
assign LUT_2[30605] = 32'b11111111111111111011111100000110;
assign LUT_2[30606] = 32'b00000000000000000101111100101001;
assign LUT_2[30607] = 32'b00000000000000000010110101000010;
assign LUT_2[30608] = 32'b00000000000000000010011000110010;
assign LUT_2[30609] = 32'b11111111111111111111010001001011;
assign LUT_2[30610] = 32'b00000000000000001001010001101110;
assign LUT_2[30611] = 32'b00000000000000000110001010000111;
assign LUT_2[30612] = 32'b11111111111111111110110110011010;
assign LUT_2[30613] = 32'b11111111111111111011101110110011;
assign LUT_2[30614] = 32'b00000000000000000101101111010110;
assign LUT_2[30615] = 32'b00000000000000000010100111101111;
assign LUT_2[30616] = 32'b11111111111111111101001010001111;
assign LUT_2[30617] = 32'b11111111111111111010000010101000;
assign LUT_2[30618] = 32'b00000000000000000100000011001011;
assign LUT_2[30619] = 32'b00000000000000000000111011100100;
assign LUT_2[30620] = 32'b11111111111111111001100111110111;
assign LUT_2[30621] = 32'b11111111111111110110100000010000;
assign LUT_2[30622] = 32'b00000000000000000000100000110011;
assign LUT_2[30623] = 32'b11111111111111111101011001001100;
assign LUT_2[30624] = 32'b00000000000000001000010000010001;
assign LUT_2[30625] = 32'b00000000000000000101001000101010;
assign LUT_2[30626] = 32'b00000000000000001111001001001101;
assign LUT_2[30627] = 32'b00000000000000001100000001100110;
assign LUT_2[30628] = 32'b00000000000000000100101101111001;
assign LUT_2[30629] = 32'b00000000000000000001100110010010;
assign LUT_2[30630] = 32'b00000000000000001011100110110101;
assign LUT_2[30631] = 32'b00000000000000001000011111001110;
assign LUT_2[30632] = 32'b00000000000000000011000001101110;
assign LUT_2[30633] = 32'b11111111111111111111111010000111;
assign LUT_2[30634] = 32'b00000000000000001001111010101010;
assign LUT_2[30635] = 32'b00000000000000000110110011000011;
assign LUT_2[30636] = 32'b11111111111111111111011111010110;
assign LUT_2[30637] = 32'b11111111111111111100010111101111;
assign LUT_2[30638] = 32'b00000000000000000110011000010010;
assign LUT_2[30639] = 32'b00000000000000000011010000101011;
assign LUT_2[30640] = 32'b00000000000000000010110100011011;
assign LUT_2[30641] = 32'b11111111111111111111101100110100;
assign LUT_2[30642] = 32'b00000000000000001001101101010111;
assign LUT_2[30643] = 32'b00000000000000000110100101110000;
assign LUT_2[30644] = 32'b11111111111111111111010010000011;
assign LUT_2[30645] = 32'b11111111111111111100001010011100;
assign LUT_2[30646] = 32'b00000000000000000110001010111111;
assign LUT_2[30647] = 32'b00000000000000000011000011011000;
assign LUT_2[30648] = 32'b11111111111111111101100101111000;
assign LUT_2[30649] = 32'b11111111111111111010011110010001;
assign LUT_2[30650] = 32'b00000000000000000100011110110100;
assign LUT_2[30651] = 32'b00000000000000000001010111001101;
assign LUT_2[30652] = 32'b11111111111111111010000011100000;
assign LUT_2[30653] = 32'b11111111111111110110111011111001;
assign LUT_2[30654] = 32'b00000000000000000000111100011100;
assign LUT_2[30655] = 32'b11111111111111111101110100110101;
assign LUT_2[30656] = 32'b11111111111111111111111101001011;
assign LUT_2[30657] = 32'b11111111111111111100110101100100;
assign LUT_2[30658] = 32'b00000000000000000110110110000111;
assign LUT_2[30659] = 32'b00000000000000000011101110100000;
assign LUT_2[30660] = 32'b11111111111111111100011010110011;
assign LUT_2[30661] = 32'b11111111111111111001010011001100;
assign LUT_2[30662] = 32'b00000000000000000011010011101111;
assign LUT_2[30663] = 32'b00000000000000000000001100001000;
assign LUT_2[30664] = 32'b11111111111111111010101110101000;
assign LUT_2[30665] = 32'b11111111111111110111100111000001;
assign LUT_2[30666] = 32'b00000000000000000001100111100100;
assign LUT_2[30667] = 32'b11111111111111111110011111111101;
assign LUT_2[30668] = 32'b11111111111111110111001100010000;
assign LUT_2[30669] = 32'b11111111111111110100000100101001;
assign LUT_2[30670] = 32'b11111111111111111110000101001100;
assign LUT_2[30671] = 32'b11111111111111111010111101100101;
assign LUT_2[30672] = 32'b11111111111111111010100001010101;
assign LUT_2[30673] = 32'b11111111111111110111011001101110;
assign LUT_2[30674] = 32'b00000000000000000001011010010001;
assign LUT_2[30675] = 32'b11111111111111111110010010101010;
assign LUT_2[30676] = 32'b11111111111111110110111110111101;
assign LUT_2[30677] = 32'b11111111111111110011110111010110;
assign LUT_2[30678] = 32'b11111111111111111101110111111001;
assign LUT_2[30679] = 32'b11111111111111111010110000010010;
assign LUT_2[30680] = 32'b11111111111111110101010010110010;
assign LUT_2[30681] = 32'b11111111111111110010001011001011;
assign LUT_2[30682] = 32'b11111111111111111100001011101110;
assign LUT_2[30683] = 32'b11111111111111111001000100000111;
assign LUT_2[30684] = 32'b11111111111111110001110000011010;
assign LUT_2[30685] = 32'b11111111111111101110101000110011;
assign LUT_2[30686] = 32'b11111111111111111000101001010110;
assign LUT_2[30687] = 32'b11111111111111110101100001101111;
assign LUT_2[30688] = 32'b00000000000000000000011000110100;
assign LUT_2[30689] = 32'b11111111111111111101010001001101;
assign LUT_2[30690] = 32'b00000000000000000111010001110000;
assign LUT_2[30691] = 32'b00000000000000000100001010001001;
assign LUT_2[30692] = 32'b11111111111111111100110110011100;
assign LUT_2[30693] = 32'b11111111111111111001101110110101;
assign LUT_2[30694] = 32'b00000000000000000011101111011000;
assign LUT_2[30695] = 32'b00000000000000000000100111110001;
assign LUT_2[30696] = 32'b11111111111111111011001010010001;
assign LUT_2[30697] = 32'b11111111111111111000000010101010;
assign LUT_2[30698] = 32'b00000000000000000010000011001101;
assign LUT_2[30699] = 32'b11111111111111111110111011100110;
assign LUT_2[30700] = 32'b11111111111111110111100111111001;
assign LUT_2[30701] = 32'b11111111111111110100100000010010;
assign LUT_2[30702] = 32'b11111111111111111110100000110101;
assign LUT_2[30703] = 32'b11111111111111111011011001001110;
assign LUT_2[30704] = 32'b11111111111111111010111100111110;
assign LUT_2[30705] = 32'b11111111111111110111110101010111;
assign LUT_2[30706] = 32'b00000000000000000001110101111010;
assign LUT_2[30707] = 32'b11111111111111111110101110010011;
assign LUT_2[30708] = 32'b11111111111111110111011010100110;
assign LUT_2[30709] = 32'b11111111111111110100010010111111;
assign LUT_2[30710] = 32'b11111111111111111110010011100010;
assign LUT_2[30711] = 32'b11111111111111111011001011111011;
assign LUT_2[30712] = 32'b11111111111111110101101110011011;
assign LUT_2[30713] = 32'b11111111111111110010100110110100;
assign LUT_2[30714] = 32'b11111111111111111100100111010111;
assign LUT_2[30715] = 32'b11111111111111111001011111110000;
assign LUT_2[30716] = 32'b11111111111111110010001100000011;
assign LUT_2[30717] = 32'b11111111111111101111000100011100;
assign LUT_2[30718] = 32'b11111111111111111001000100111111;
assign LUT_2[30719] = 32'b11111111111111110101111101011000;
assign LUT_2[30720] = 32'b11111111111111101111111001111000;
assign LUT_2[30721] = 32'b11111111111111101100110010010001;
assign LUT_2[30722] = 32'b11111111111111110110110010110100;
assign LUT_2[30723] = 32'b11111111111111110011101011001101;
assign LUT_2[30724] = 32'b11111111111111101100010111100000;
assign LUT_2[30725] = 32'b11111111111111101001001111111001;
assign LUT_2[30726] = 32'b11111111111111110011010000011100;
assign LUT_2[30727] = 32'b11111111111111110000001000110101;
assign LUT_2[30728] = 32'b11111111111111101010101011010101;
assign LUT_2[30729] = 32'b11111111111111100111100011101110;
assign LUT_2[30730] = 32'b11111111111111110001100100010001;
assign LUT_2[30731] = 32'b11111111111111101110011100101010;
assign LUT_2[30732] = 32'b11111111111111100111001000111101;
assign LUT_2[30733] = 32'b11111111111111100100000001010110;
assign LUT_2[30734] = 32'b11111111111111101110000001111001;
assign LUT_2[30735] = 32'b11111111111111101010111010010010;
assign LUT_2[30736] = 32'b11111111111111101010011110000010;
assign LUT_2[30737] = 32'b11111111111111100111010110011011;
assign LUT_2[30738] = 32'b11111111111111110001010110111110;
assign LUT_2[30739] = 32'b11111111111111101110001111010111;
assign LUT_2[30740] = 32'b11111111111111100110111011101010;
assign LUT_2[30741] = 32'b11111111111111100011110100000011;
assign LUT_2[30742] = 32'b11111111111111101101110100100110;
assign LUT_2[30743] = 32'b11111111111111101010101100111111;
assign LUT_2[30744] = 32'b11111111111111100101001111011111;
assign LUT_2[30745] = 32'b11111111111111100010000111111000;
assign LUT_2[30746] = 32'b11111111111111101100001000011011;
assign LUT_2[30747] = 32'b11111111111111101001000000110100;
assign LUT_2[30748] = 32'b11111111111111100001101101000111;
assign LUT_2[30749] = 32'b11111111111111011110100101100000;
assign LUT_2[30750] = 32'b11111111111111101000100110000011;
assign LUT_2[30751] = 32'b11111111111111100101011110011100;
assign LUT_2[30752] = 32'b11111111111111110000010101100001;
assign LUT_2[30753] = 32'b11111111111111101101001101111010;
assign LUT_2[30754] = 32'b11111111111111110111001110011101;
assign LUT_2[30755] = 32'b11111111111111110100000110110110;
assign LUT_2[30756] = 32'b11111111111111101100110011001001;
assign LUT_2[30757] = 32'b11111111111111101001101011100010;
assign LUT_2[30758] = 32'b11111111111111110011101100000101;
assign LUT_2[30759] = 32'b11111111111111110000100100011110;
assign LUT_2[30760] = 32'b11111111111111101011000110111110;
assign LUT_2[30761] = 32'b11111111111111100111111111010111;
assign LUT_2[30762] = 32'b11111111111111110001111111111010;
assign LUT_2[30763] = 32'b11111111111111101110111000010011;
assign LUT_2[30764] = 32'b11111111111111100111100100100110;
assign LUT_2[30765] = 32'b11111111111111100100011100111111;
assign LUT_2[30766] = 32'b11111111111111101110011101100010;
assign LUT_2[30767] = 32'b11111111111111101011010101111011;
assign LUT_2[30768] = 32'b11111111111111101010111001101011;
assign LUT_2[30769] = 32'b11111111111111100111110010000100;
assign LUT_2[30770] = 32'b11111111111111110001110010100111;
assign LUT_2[30771] = 32'b11111111111111101110101011000000;
assign LUT_2[30772] = 32'b11111111111111100111010111010011;
assign LUT_2[30773] = 32'b11111111111111100100001111101100;
assign LUT_2[30774] = 32'b11111111111111101110010000001111;
assign LUT_2[30775] = 32'b11111111111111101011001000101000;
assign LUT_2[30776] = 32'b11111111111111100101101011001000;
assign LUT_2[30777] = 32'b11111111111111100010100011100001;
assign LUT_2[30778] = 32'b11111111111111101100100100000100;
assign LUT_2[30779] = 32'b11111111111111101001011100011101;
assign LUT_2[30780] = 32'b11111111111111100010001000110000;
assign LUT_2[30781] = 32'b11111111111111011111000001001001;
assign LUT_2[30782] = 32'b11111111111111101001000001101100;
assign LUT_2[30783] = 32'b11111111111111100101111010000101;
assign LUT_2[30784] = 32'b11111111111111101000000010011011;
assign LUT_2[30785] = 32'b11111111111111100100111010110100;
assign LUT_2[30786] = 32'b11111111111111101110111011010111;
assign LUT_2[30787] = 32'b11111111111111101011110011110000;
assign LUT_2[30788] = 32'b11111111111111100100100000000011;
assign LUT_2[30789] = 32'b11111111111111100001011000011100;
assign LUT_2[30790] = 32'b11111111111111101011011000111111;
assign LUT_2[30791] = 32'b11111111111111101000010001011000;
assign LUT_2[30792] = 32'b11111111111111100010110011111000;
assign LUT_2[30793] = 32'b11111111111111011111101100010001;
assign LUT_2[30794] = 32'b11111111111111101001101100110100;
assign LUT_2[30795] = 32'b11111111111111100110100101001101;
assign LUT_2[30796] = 32'b11111111111111011111010001100000;
assign LUT_2[30797] = 32'b11111111111111011100001001111001;
assign LUT_2[30798] = 32'b11111111111111100110001010011100;
assign LUT_2[30799] = 32'b11111111111111100011000010110101;
assign LUT_2[30800] = 32'b11111111111111100010100110100101;
assign LUT_2[30801] = 32'b11111111111111011111011110111110;
assign LUT_2[30802] = 32'b11111111111111101001011111100001;
assign LUT_2[30803] = 32'b11111111111111100110010111111010;
assign LUT_2[30804] = 32'b11111111111111011111000100001101;
assign LUT_2[30805] = 32'b11111111111111011011111100100110;
assign LUT_2[30806] = 32'b11111111111111100101111101001001;
assign LUT_2[30807] = 32'b11111111111111100010110101100010;
assign LUT_2[30808] = 32'b11111111111111011101011000000010;
assign LUT_2[30809] = 32'b11111111111111011010010000011011;
assign LUT_2[30810] = 32'b11111111111111100100010000111110;
assign LUT_2[30811] = 32'b11111111111111100001001001010111;
assign LUT_2[30812] = 32'b11111111111111011001110101101010;
assign LUT_2[30813] = 32'b11111111111111010110101110000011;
assign LUT_2[30814] = 32'b11111111111111100000101110100110;
assign LUT_2[30815] = 32'b11111111111111011101100110111111;
assign LUT_2[30816] = 32'b11111111111111101000011110000100;
assign LUT_2[30817] = 32'b11111111111111100101010110011101;
assign LUT_2[30818] = 32'b11111111111111101111010111000000;
assign LUT_2[30819] = 32'b11111111111111101100001111011001;
assign LUT_2[30820] = 32'b11111111111111100100111011101100;
assign LUT_2[30821] = 32'b11111111111111100001110100000101;
assign LUT_2[30822] = 32'b11111111111111101011110100101000;
assign LUT_2[30823] = 32'b11111111111111101000101101000001;
assign LUT_2[30824] = 32'b11111111111111100011001111100001;
assign LUT_2[30825] = 32'b11111111111111100000000111111010;
assign LUT_2[30826] = 32'b11111111111111101010001000011101;
assign LUT_2[30827] = 32'b11111111111111100111000000110110;
assign LUT_2[30828] = 32'b11111111111111011111101101001001;
assign LUT_2[30829] = 32'b11111111111111011100100101100010;
assign LUT_2[30830] = 32'b11111111111111100110100110000101;
assign LUT_2[30831] = 32'b11111111111111100011011110011110;
assign LUT_2[30832] = 32'b11111111111111100011000010001110;
assign LUT_2[30833] = 32'b11111111111111011111111010100111;
assign LUT_2[30834] = 32'b11111111111111101001111011001010;
assign LUT_2[30835] = 32'b11111111111111100110110011100011;
assign LUT_2[30836] = 32'b11111111111111011111011111110110;
assign LUT_2[30837] = 32'b11111111111111011100011000001111;
assign LUT_2[30838] = 32'b11111111111111100110011000110010;
assign LUT_2[30839] = 32'b11111111111111100011010001001011;
assign LUT_2[30840] = 32'b11111111111111011101110011101011;
assign LUT_2[30841] = 32'b11111111111111011010101100000100;
assign LUT_2[30842] = 32'b11111111111111100100101100100111;
assign LUT_2[30843] = 32'b11111111111111100001100101000000;
assign LUT_2[30844] = 32'b11111111111111011010010001010011;
assign LUT_2[30845] = 32'b11111111111111010111001001101100;
assign LUT_2[30846] = 32'b11111111111111100001001010001111;
assign LUT_2[30847] = 32'b11111111111111011110000010101000;
assign LUT_2[30848] = 32'b11111111111111110100001110000111;
assign LUT_2[30849] = 32'b11111111111111110001000110100000;
assign LUT_2[30850] = 32'b11111111111111111011000111000011;
assign LUT_2[30851] = 32'b11111111111111110111111111011100;
assign LUT_2[30852] = 32'b11111111111111110000101011101111;
assign LUT_2[30853] = 32'b11111111111111101101100100001000;
assign LUT_2[30854] = 32'b11111111111111110111100100101011;
assign LUT_2[30855] = 32'b11111111111111110100011101000100;
assign LUT_2[30856] = 32'b11111111111111101110111111100100;
assign LUT_2[30857] = 32'b11111111111111101011110111111101;
assign LUT_2[30858] = 32'b11111111111111110101111000100000;
assign LUT_2[30859] = 32'b11111111111111110010110000111001;
assign LUT_2[30860] = 32'b11111111111111101011011101001100;
assign LUT_2[30861] = 32'b11111111111111101000010101100101;
assign LUT_2[30862] = 32'b11111111111111110010010110001000;
assign LUT_2[30863] = 32'b11111111111111101111001110100001;
assign LUT_2[30864] = 32'b11111111111111101110110010010001;
assign LUT_2[30865] = 32'b11111111111111101011101010101010;
assign LUT_2[30866] = 32'b11111111111111110101101011001101;
assign LUT_2[30867] = 32'b11111111111111110010100011100110;
assign LUT_2[30868] = 32'b11111111111111101011001111111001;
assign LUT_2[30869] = 32'b11111111111111101000001000010010;
assign LUT_2[30870] = 32'b11111111111111110010001000110101;
assign LUT_2[30871] = 32'b11111111111111101111000001001110;
assign LUT_2[30872] = 32'b11111111111111101001100011101110;
assign LUT_2[30873] = 32'b11111111111111100110011100000111;
assign LUT_2[30874] = 32'b11111111111111110000011100101010;
assign LUT_2[30875] = 32'b11111111111111101101010101000011;
assign LUT_2[30876] = 32'b11111111111111100110000001010110;
assign LUT_2[30877] = 32'b11111111111111100010111001101111;
assign LUT_2[30878] = 32'b11111111111111101100111010010010;
assign LUT_2[30879] = 32'b11111111111111101001110010101011;
assign LUT_2[30880] = 32'b11111111111111110100101001110000;
assign LUT_2[30881] = 32'b11111111111111110001100010001001;
assign LUT_2[30882] = 32'b11111111111111111011100010101100;
assign LUT_2[30883] = 32'b11111111111111111000011011000101;
assign LUT_2[30884] = 32'b11111111111111110001000111011000;
assign LUT_2[30885] = 32'b11111111111111101101111111110001;
assign LUT_2[30886] = 32'b11111111111111111000000000010100;
assign LUT_2[30887] = 32'b11111111111111110100111000101101;
assign LUT_2[30888] = 32'b11111111111111101111011011001101;
assign LUT_2[30889] = 32'b11111111111111101100010011100110;
assign LUT_2[30890] = 32'b11111111111111110110010100001001;
assign LUT_2[30891] = 32'b11111111111111110011001100100010;
assign LUT_2[30892] = 32'b11111111111111101011111000110101;
assign LUT_2[30893] = 32'b11111111111111101000110001001110;
assign LUT_2[30894] = 32'b11111111111111110010110001110001;
assign LUT_2[30895] = 32'b11111111111111101111101010001010;
assign LUT_2[30896] = 32'b11111111111111101111001101111010;
assign LUT_2[30897] = 32'b11111111111111101100000110010011;
assign LUT_2[30898] = 32'b11111111111111110110000110110110;
assign LUT_2[30899] = 32'b11111111111111110010111111001111;
assign LUT_2[30900] = 32'b11111111111111101011101011100010;
assign LUT_2[30901] = 32'b11111111111111101000100011111011;
assign LUT_2[30902] = 32'b11111111111111110010100100011110;
assign LUT_2[30903] = 32'b11111111111111101111011100110111;
assign LUT_2[30904] = 32'b11111111111111101001111111010111;
assign LUT_2[30905] = 32'b11111111111111100110110111110000;
assign LUT_2[30906] = 32'b11111111111111110000111000010011;
assign LUT_2[30907] = 32'b11111111111111101101110000101100;
assign LUT_2[30908] = 32'b11111111111111100110011100111111;
assign LUT_2[30909] = 32'b11111111111111100011010101011000;
assign LUT_2[30910] = 32'b11111111111111101101010101111011;
assign LUT_2[30911] = 32'b11111111111111101010001110010100;
assign LUT_2[30912] = 32'b11111111111111101100010110101010;
assign LUT_2[30913] = 32'b11111111111111101001001111000011;
assign LUT_2[30914] = 32'b11111111111111110011001111100110;
assign LUT_2[30915] = 32'b11111111111111110000000111111111;
assign LUT_2[30916] = 32'b11111111111111101000110100010010;
assign LUT_2[30917] = 32'b11111111111111100101101100101011;
assign LUT_2[30918] = 32'b11111111111111101111101101001110;
assign LUT_2[30919] = 32'b11111111111111101100100101100111;
assign LUT_2[30920] = 32'b11111111111111100111001000000111;
assign LUT_2[30921] = 32'b11111111111111100100000000100000;
assign LUT_2[30922] = 32'b11111111111111101110000001000011;
assign LUT_2[30923] = 32'b11111111111111101010111001011100;
assign LUT_2[30924] = 32'b11111111111111100011100101101111;
assign LUT_2[30925] = 32'b11111111111111100000011110001000;
assign LUT_2[30926] = 32'b11111111111111101010011110101011;
assign LUT_2[30927] = 32'b11111111111111100111010111000100;
assign LUT_2[30928] = 32'b11111111111111100110111010110100;
assign LUT_2[30929] = 32'b11111111111111100011110011001101;
assign LUT_2[30930] = 32'b11111111111111101101110011110000;
assign LUT_2[30931] = 32'b11111111111111101010101100001001;
assign LUT_2[30932] = 32'b11111111111111100011011000011100;
assign LUT_2[30933] = 32'b11111111111111100000010000110101;
assign LUT_2[30934] = 32'b11111111111111101010010001011000;
assign LUT_2[30935] = 32'b11111111111111100111001001110001;
assign LUT_2[30936] = 32'b11111111111111100001101100010001;
assign LUT_2[30937] = 32'b11111111111111011110100100101010;
assign LUT_2[30938] = 32'b11111111111111101000100101001101;
assign LUT_2[30939] = 32'b11111111111111100101011101100110;
assign LUT_2[30940] = 32'b11111111111111011110001001111001;
assign LUT_2[30941] = 32'b11111111111111011011000010010010;
assign LUT_2[30942] = 32'b11111111111111100101000010110101;
assign LUT_2[30943] = 32'b11111111111111100001111011001110;
assign LUT_2[30944] = 32'b11111111111111101100110010010011;
assign LUT_2[30945] = 32'b11111111111111101001101010101100;
assign LUT_2[30946] = 32'b11111111111111110011101011001111;
assign LUT_2[30947] = 32'b11111111111111110000100011101000;
assign LUT_2[30948] = 32'b11111111111111101001001111111011;
assign LUT_2[30949] = 32'b11111111111111100110001000010100;
assign LUT_2[30950] = 32'b11111111111111110000001000110111;
assign LUT_2[30951] = 32'b11111111111111101101000001010000;
assign LUT_2[30952] = 32'b11111111111111100111100011110000;
assign LUT_2[30953] = 32'b11111111111111100100011100001001;
assign LUT_2[30954] = 32'b11111111111111101110011100101100;
assign LUT_2[30955] = 32'b11111111111111101011010101000101;
assign LUT_2[30956] = 32'b11111111111111100100000001011000;
assign LUT_2[30957] = 32'b11111111111111100000111001110001;
assign LUT_2[30958] = 32'b11111111111111101010111010010100;
assign LUT_2[30959] = 32'b11111111111111100111110010101101;
assign LUT_2[30960] = 32'b11111111111111100111010110011101;
assign LUT_2[30961] = 32'b11111111111111100100001110110110;
assign LUT_2[30962] = 32'b11111111111111101110001111011001;
assign LUT_2[30963] = 32'b11111111111111101011000111110010;
assign LUT_2[30964] = 32'b11111111111111100011110100000101;
assign LUT_2[30965] = 32'b11111111111111100000101100011110;
assign LUT_2[30966] = 32'b11111111111111101010101101000001;
assign LUT_2[30967] = 32'b11111111111111100111100101011010;
assign LUT_2[30968] = 32'b11111111111111100010000111111010;
assign LUT_2[30969] = 32'b11111111111111011111000000010011;
assign LUT_2[30970] = 32'b11111111111111101001000000110110;
assign LUT_2[30971] = 32'b11111111111111100101111001001111;
assign LUT_2[30972] = 32'b11111111111111011110100101100010;
assign LUT_2[30973] = 32'b11111111111111011011011101111011;
assign LUT_2[30974] = 32'b11111111111111100101011110011110;
assign LUT_2[30975] = 32'b11111111111111100010010110110111;
assign LUT_2[30976] = 32'b11111111111111110011111000011110;
assign LUT_2[30977] = 32'b11111111111111110000110000110111;
assign LUT_2[30978] = 32'b11111111111111111010110001011010;
assign LUT_2[30979] = 32'b11111111111111110111101001110011;
assign LUT_2[30980] = 32'b11111111111111110000010110000110;
assign LUT_2[30981] = 32'b11111111111111101101001110011111;
assign LUT_2[30982] = 32'b11111111111111110111001111000010;
assign LUT_2[30983] = 32'b11111111111111110100000111011011;
assign LUT_2[30984] = 32'b11111111111111101110101001111011;
assign LUT_2[30985] = 32'b11111111111111101011100010010100;
assign LUT_2[30986] = 32'b11111111111111110101100010110111;
assign LUT_2[30987] = 32'b11111111111111110010011011010000;
assign LUT_2[30988] = 32'b11111111111111101011000111100011;
assign LUT_2[30989] = 32'b11111111111111100111111111111100;
assign LUT_2[30990] = 32'b11111111111111110010000000011111;
assign LUT_2[30991] = 32'b11111111111111101110111000111000;
assign LUT_2[30992] = 32'b11111111111111101110011100101000;
assign LUT_2[30993] = 32'b11111111111111101011010101000001;
assign LUT_2[30994] = 32'b11111111111111110101010101100100;
assign LUT_2[30995] = 32'b11111111111111110010001101111101;
assign LUT_2[30996] = 32'b11111111111111101010111010010000;
assign LUT_2[30997] = 32'b11111111111111100111110010101001;
assign LUT_2[30998] = 32'b11111111111111110001110011001100;
assign LUT_2[30999] = 32'b11111111111111101110101011100101;
assign LUT_2[31000] = 32'b11111111111111101001001110000101;
assign LUT_2[31001] = 32'b11111111111111100110000110011110;
assign LUT_2[31002] = 32'b11111111111111110000000111000001;
assign LUT_2[31003] = 32'b11111111111111101100111111011010;
assign LUT_2[31004] = 32'b11111111111111100101101011101101;
assign LUT_2[31005] = 32'b11111111111111100010100100000110;
assign LUT_2[31006] = 32'b11111111111111101100100100101001;
assign LUT_2[31007] = 32'b11111111111111101001011101000010;
assign LUT_2[31008] = 32'b11111111111111110100010100000111;
assign LUT_2[31009] = 32'b11111111111111110001001100100000;
assign LUT_2[31010] = 32'b11111111111111111011001101000011;
assign LUT_2[31011] = 32'b11111111111111111000000101011100;
assign LUT_2[31012] = 32'b11111111111111110000110001101111;
assign LUT_2[31013] = 32'b11111111111111101101101010001000;
assign LUT_2[31014] = 32'b11111111111111110111101010101011;
assign LUT_2[31015] = 32'b11111111111111110100100011000100;
assign LUT_2[31016] = 32'b11111111111111101111000101100100;
assign LUT_2[31017] = 32'b11111111111111101011111101111101;
assign LUT_2[31018] = 32'b11111111111111110101111110100000;
assign LUT_2[31019] = 32'b11111111111111110010110110111001;
assign LUT_2[31020] = 32'b11111111111111101011100011001100;
assign LUT_2[31021] = 32'b11111111111111101000011011100101;
assign LUT_2[31022] = 32'b11111111111111110010011100001000;
assign LUT_2[31023] = 32'b11111111111111101111010100100001;
assign LUT_2[31024] = 32'b11111111111111101110111000010001;
assign LUT_2[31025] = 32'b11111111111111101011110000101010;
assign LUT_2[31026] = 32'b11111111111111110101110001001101;
assign LUT_2[31027] = 32'b11111111111111110010101001100110;
assign LUT_2[31028] = 32'b11111111111111101011010101111001;
assign LUT_2[31029] = 32'b11111111111111101000001110010010;
assign LUT_2[31030] = 32'b11111111111111110010001110110101;
assign LUT_2[31031] = 32'b11111111111111101111000111001110;
assign LUT_2[31032] = 32'b11111111111111101001101001101110;
assign LUT_2[31033] = 32'b11111111111111100110100010000111;
assign LUT_2[31034] = 32'b11111111111111110000100010101010;
assign LUT_2[31035] = 32'b11111111111111101101011011000011;
assign LUT_2[31036] = 32'b11111111111111100110000111010110;
assign LUT_2[31037] = 32'b11111111111111100010111111101111;
assign LUT_2[31038] = 32'b11111111111111101101000000010010;
assign LUT_2[31039] = 32'b11111111111111101001111000101011;
assign LUT_2[31040] = 32'b11111111111111101100000001000001;
assign LUT_2[31041] = 32'b11111111111111101000111001011010;
assign LUT_2[31042] = 32'b11111111111111110010111001111101;
assign LUT_2[31043] = 32'b11111111111111101111110010010110;
assign LUT_2[31044] = 32'b11111111111111101000011110101001;
assign LUT_2[31045] = 32'b11111111111111100101010111000010;
assign LUT_2[31046] = 32'b11111111111111101111010111100101;
assign LUT_2[31047] = 32'b11111111111111101100001111111110;
assign LUT_2[31048] = 32'b11111111111111100110110010011110;
assign LUT_2[31049] = 32'b11111111111111100011101010110111;
assign LUT_2[31050] = 32'b11111111111111101101101011011010;
assign LUT_2[31051] = 32'b11111111111111101010100011110011;
assign LUT_2[31052] = 32'b11111111111111100011010000000110;
assign LUT_2[31053] = 32'b11111111111111100000001000011111;
assign LUT_2[31054] = 32'b11111111111111101010001001000010;
assign LUT_2[31055] = 32'b11111111111111100111000001011011;
assign LUT_2[31056] = 32'b11111111111111100110100101001011;
assign LUT_2[31057] = 32'b11111111111111100011011101100100;
assign LUT_2[31058] = 32'b11111111111111101101011110000111;
assign LUT_2[31059] = 32'b11111111111111101010010110100000;
assign LUT_2[31060] = 32'b11111111111111100011000010110011;
assign LUT_2[31061] = 32'b11111111111111011111111011001100;
assign LUT_2[31062] = 32'b11111111111111101001111011101111;
assign LUT_2[31063] = 32'b11111111111111100110110100001000;
assign LUT_2[31064] = 32'b11111111111111100001010110101000;
assign LUT_2[31065] = 32'b11111111111111011110001111000001;
assign LUT_2[31066] = 32'b11111111111111101000001111100100;
assign LUT_2[31067] = 32'b11111111111111100101000111111101;
assign LUT_2[31068] = 32'b11111111111111011101110100010000;
assign LUT_2[31069] = 32'b11111111111111011010101100101001;
assign LUT_2[31070] = 32'b11111111111111100100101101001100;
assign LUT_2[31071] = 32'b11111111111111100001100101100101;
assign LUT_2[31072] = 32'b11111111111111101100011100101010;
assign LUT_2[31073] = 32'b11111111111111101001010101000011;
assign LUT_2[31074] = 32'b11111111111111110011010101100110;
assign LUT_2[31075] = 32'b11111111111111110000001101111111;
assign LUT_2[31076] = 32'b11111111111111101000111010010010;
assign LUT_2[31077] = 32'b11111111111111100101110010101011;
assign LUT_2[31078] = 32'b11111111111111101111110011001110;
assign LUT_2[31079] = 32'b11111111111111101100101011100111;
assign LUT_2[31080] = 32'b11111111111111100111001110000111;
assign LUT_2[31081] = 32'b11111111111111100100000110100000;
assign LUT_2[31082] = 32'b11111111111111101110000111000011;
assign LUT_2[31083] = 32'b11111111111111101010111111011100;
assign LUT_2[31084] = 32'b11111111111111100011101011101111;
assign LUT_2[31085] = 32'b11111111111111100000100100001000;
assign LUT_2[31086] = 32'b11111111111111101010100100101011;
assign LUT_2[31087] = 32'b11111111111111100111011101000100;
assign LUT_2[31088] = 32'b11111111111111100111000000110100;
assign LUT_2[31089] = 32'b11111111111111100011111001001101;
assign LUT_2[31090] = 32'b11111111111111101101111001110000;
assign LUT_2[31091] = 32'b11111111111111101010110010001001;
assign LUT_2[31092] = 32'b11111111111111100011011110011100;
assign LUT_2[31093] = 32'b11111111111111100000010110110101;
assign LUT_2[31094] = 32'b11111111111111101010010111011000;
assign LUT_2[31095] = 32'b11111111111111100111001111110001;
assign LUT_2[31096] = 32'b11111111111111100001110010010001;
assign LUT_2[31097] = 32'b11111111111111011110101010101010;
assign LUT_2[31098] = 32'b11111111111111101000101011001101;
assign LUT_2[31099] = 32'b11111111111111100101100011100110;
assign LUT_2[31100] = 32'b11111111111111011110001111111001;
assign LUT_2[31101] = 32'b11111111111111011011001000010010;
assign LUT_2[31102] = 32'b11111111111111100101001000110101;
assign LUT_2[31103] = 32'b11111111111111100010000001001110;
assign LUT_2[31104] = 32'b11111111111111111000001100101101;
assign LUT_2[31105] = 32'b11111111111111110101000101000110;
assign LUT_2[31106] = 32'b11111111111111111111000101101001;
assign LUT_2[31107] = 32'b11111111111111111011111110000010;
assign LUT_2[31108] = 32'b11111111111111110100101010010101;
assign LUT_2[31109] = 32'b11111111111111110001100010101110;
assign LUT_2[31110] = 32'b11111111111111111011100011010001;
assign LUT_2[31111] = 32'b11111111111111111000011011101010;
assign LUT_2[31112] = 32'b11111111111111110010111110001010;
assign LUT_2[31113] = 32'b11111111111111101111110110100011;
assign LUT_2[31114] = 32'b11111111111111111001110111000110;
assign LUT_2[31115] = 32'b11111111111111110110101111011111;
assign LUT_2[31116] = 32'b11111111111111101111011011110010;
assign LUT_2[31117] = 32'b11111111111111101100010100001011;
assign LUT_2[31118] = 32'b11111111111111110110010100101110;
assign LUT_2[31119] = 32'b11111111111111110011001101000111;
assign LUT_2[31120] = 32'b11111111111111110010110000110111;
assign LUT_2[31121] = 32'b11111111111111101111101001010000;
assign LUT_2[31122] = 32'b11111111111111111001101001110011;
assign LUT_2[31123] = 32'b11111111111111110110100010001100;
assign LUT_2[31124] = 32'b11111111111111101111001110011111;
assign LUT_2[31125] = 32'b11111111111111101100000110111000;
assign LUT_2[31126] = 32'b11111111111111110110000111011011;
assign LUT_2[31127] = 32'b11111111111111110010111111110100;
assign LUT_2[31128] = 32'b11111111111111101101100010010100;
assign LUT_2[31129] = 32'b11111111111111101010011010101101;
assign LUT_2[31130] = 32'b11111111111111110100011011010000;
assign LUT_2[31131] = 32'b11111111111111110001010011101001;
assign LUT_2[31132] = 32'b11111111111111101001111111111100;
assign LUT_2[31133] = 32'b11111111111111100110111000010101;
assign LUT_2[31134] = 32'b11111111111111110000111000111000;
assign LUT_2[31135] = 32'b11111111111111101101110001010001;
assign LUT_2[31136] = 32'b11111111111111111000101000010110;
assign LUT_2[31137] = 32'b11111111111111110101100000101111;
assign LUT_2[31138] = 32'b11111111111111111111100001010010;
assign LUT_2[31139] = 32'b11111111111111111100011001101011;
assign LUT_2[31140] = 32'b11111111111111110101000101111110;
assign LUT_2[31141] = 32'b11111111111111110001111110010111;
assign LUT_2[31142] = 32'b11111111111111111011111110111010;
assign LUT_2[31143] = 32'b11111111111111111000110111010011;
assign LUT_2[31144] = 32'b11111111111111110011011001110011;
assign LUT_2[31145] = 32'b11111111111111110000010010001100;
assign LUT_2[31146] = 32'b11111111111111111010010010101111;
assign LUT_2[31147] = 32'b11111111111111110111001011001000;
assign LUT_2[31148] = 32'b11111111111111101111110111011011;
assign LUT_2[31149] = 32'b11111111111111101100101111110100;
assign LUT_2[31150] = 32'b11111111111111110110110000010111;
assign LUT_2[31151] = 32'b11111111111111110011101000110000;
assign LUT_2[31152] = 32'b11111111111111110011001100100000;
assign LUT_2[31153] = 32'b11111111111111110000000100111001;
assign LUT_2[31154] = 32'b11111111111111111010000101011100;
assign LUT_2[31155] = 32'b11111111111111110110111101110101;
assign LUT_2[31156] = 32'b11111111111111101111101010001000;
assign LUT_2[31157] = 32'b11111111111111101100100010100001;
assign LUT_2[31158] = 32'b11111111111111110110100011000100;
assign LUT_2[31159] = 32'b11111111111111110011011011011101;
assign LUT_2[31160] = 32'b11111111111111101101111101111101;
assign LUT_2[31161] = 32'b11111111111111101010110110010110;
assign LUT_2[31162] = 32'b11111111111111110100110110111001;
assign LUT_2[31163] = 32'b11111111111111110001101111010010;
assign LUT_2[31164] = 32'b11111111111111101010011011100101;
assign LUT_2[31165] = 32'b11111111111111100111010011111110;
assign LUT_2[31166] = 32'b11111111111111110001010100100001;
assign LUT_2[31167] = 32'b11111111111111101110001100111010;
assign LUT_2[31168] = 32'b11111111111111110000010101010000;
assign LUT_2[31169] = 32'b11111111111111101101001101101001;
assign LUT_2[31170] = 32'b11111111111111110111001110001100;
assign LUT_2[31171] = 32'b11111111111111110100000110100101;
assign LUT_2[31172] = 32'b11111111111111101100110010111000;
assign LUT_2[31173] = 32'b11111111111111101001101011010001;
assign LUT_2[31174] = 32'b11111111111111110011101011110100;
assign LUT_2[31175] = 32'b11111111111111110000100100001101;
assign LUT_2[31176] = 32'b11111111111111101011000110101101;
assign LUT_2[31177] = 32'b11111111111111100111111111000110;
assign LUT_2[31178] = 32'b11111111111111110001111111101001;
assign LUT_2[31179] = 32'b11111111111111101110111000000010;
assign LUT_2[31180] = 32'b11111111111111100111100100010101;
assign LUT_2[31181] = 32'b11111111111111100100011100101110;
assign LUT_2[31182] = 32'b11111111111111101110011101010001;
assign LUT_2[31183] = 32'b11111111111111101011010101101010;
assign LUT_2[31184] = 32'b11111111111111101010111001011010;
assign LUT_2[31185] = 32'b11111111111111100111110001110011;
assign LUT_2[31186] = 32'b11111111111111110001110010010110;
assign LUT_2[31187] = 32'b11111111111111101110101010101111;
assign LUT_2[31188] = 32'b11111111111111100111010111000010;
assign LUT_2[31189] = 32'b11111111111111100100001111011011;
assign LUT_2[31190] = 32'b11111111111111101110001111111110;
assign LUT_2[31191] = 32'b11111111111111101011001000010111;
assign LUT_2[31192] = 32'b11111111111111100101101010110111;
assign LUT_2[31193] = 32'b11111111111111100010100011010000;
assign LUT_2[31194] = 32'b11111111111111101100100011110011;
assign LUT_2[31195] = 32'b11111111111111101001011100001100;
assign LUT_2[31196] = 32'b11111111111111100010001000011111;
assign LUT_2[31197] = 32'b11111111111111011111000000111000;
assign LUT_2[31198] = 32'b11111111111111101001000001011011;
assign LUT_2[31199] = 32'b11111111111111100101111001110100;
assign LUT_2[31200] = 32'b11111111111111110000110000111001;
assign LUT_2[31201] = 32'b11111111111111101101101001010010;
assign LUT_2[31202] = 32'b11111111111111110111101001110101;
assign LUT_2[31203] = 32'b11111111111111110100100010001110;
assign LUT_2[31204] = 32'b11111111111111101101001110100001;
assign LUT_2[31205] = 32'b11111111111111101010000110111010;
assign LUT_2[31206] = 32'b11111111111111110100000111011101;
assign LUT_2[31207] = 32'b11111111111111110000111111110110;
assign LUT_2[31208] = 32'b11111111111111101011100010010110;
assign LUT_2[31209] = 32'b11111111111111101000011010101111;
assign LUT_2[31210] = 32'b11111111111111110010011011010010;
assign LUT_2[31211] = 32'b11111111111111101111010011101011;
assign LUT_2[31212] = 32'b11111111111111100111111111111110;
assign LUT_2[31213] = 32'b11111111111111100100111000010111;
assign LUT_2[31214] = 32'b11111111111111101110111000111010;
assign LUT_2[31215] = 32'b11111111111111101011110001010011;
assign LUT_2[31216] = 32'b11111111111111101011010101000011;
assign LUT_2[31217] = 32'b11111111111111101000001101011100;
assign LUT_2[31218] = 32'b11111111111111110010001101111111;
assign LUT_2[31219] = 32'b11111111111111101111000110011000;
assign LUT_2[31220] = 32'b11111111111111100111110010101011;
assign LUT_2[31221] = 32'b11111111111111100100101011000100;
assign LUT_2[31222] = 32'b11111111111111101110101011100111;
assign LUT_2[31223] = 32'b11111111111111101011100100000000;
assign LUT_2[31224] = 32'b11111111111111100110000110100000;
assign LUT_2[31225] = 32'b11111111111111100010111110111001;
assign LUT_2[31226] = 32'b11111111111111101100111111011100;
assign LUT_2[31227] = 32'b11111111111111101001110111110101;
assign LUT_2[31228] = 32'b11111111111111100010100100001000;
assign LUT_2[31229] = 32'b11111111111111011111011100100001;
assign LUT_2[31230] = 32'b11111111111111101001011101000100;
assign LUT_2[31231] = 32'b11111111111111100110010101011101;
assign LUT_2[31232] = 32'b11111111111111110100101011101010;
assign LUT_2[31233] = 32'b11111111111111110001100100000011;
assign LUT_2[31234] = 32'b11111111111111111011100100100110;
assign LUT_2[31235] = 32'b11111111111111111000011100111111;
assign LUT_2[31236] = 32'b11111111111111110001001001010010;
assign LUT_2[31237] = 32'b11111111111111101110000001101011;
assign LUT_2[31238] = 32'b11111111111111111000000010001110;
assign LUT_2[31239] = 32'b11111111111111110100111010100111;
assign LUT_2[31240] = 32'b11111111111111101111011101000111;
assign LUT_2[31241] = 32'b11111111111111101100010101100000;
assign LUT_2[31242] = 32'b11111111111111110110010110000011;
assign LUT_2[31243] = 32'b11111111111111110011001110011100;
assign LUT_2[31244] = 32'b11111111111111101011111010101111;
assign LUT_2[31245] = 32'b11111111111111101000110011001000;
assign LUT_2[31246] = 32'b11111111111111110010110011101011;
assign LUT_2[31247] = 32'b11111111111111101111101100000100;
assign LUT_2[31248] = 32'b11111111111111101111001111110100;
assign LUT_2[31249] = 32'b11111111111111101100001000001101;
assign LUT_2[31250] = 32'b11111111111111110110001000110000;
assign LUT_2[31251] = 32'b11111111111111110011000001001001;
assign LUT_2[31252] = 32'b11111111111111101011101101011100;
assign LUT_2[31253] = 32'b11111111111111101000100101110101;
assign LUT_2[31254] = 32'b11111111111111110010100110011000;
assign LUT_2[31255] = 32'b11111111111111101111011110110001;
assign LUT_2[31256] = 32'b11111111111111101010000001010001;
assign LUT_2[31257] = 32'b11111111111111100110111001101010;
assign LUT_2[31258] = 32'b11111111111111110000111010001101;
assign LUT_2[31259] = 32'b11111111111111101101110010100110;
assign LUT_2[31260] = 32'b11111111111111100110011110111001;
assign LUT_2[31261] = 32'b11111111111111100011010111010010;
assign LUT_2[31262] = 32'b11111111111111101101010111110101;
assign LUT_2[31263] = 32'b11111111111111101010010000001110;
assign LUT_2[31264] = 32'b11111111111111110101000111010011;
assign LUT_2[31265] = 32'b11111111111111110001111111101100;
assign LUT_2[31266] = 32'b11111111111111111100000000001111;
assign LUT_2[31267] = 32'b11111111111111111000111000101000;
assign LUT_2[31268] = 32'b11111111111111110001100100111011;
assign LUT_2[31269] = 32'b11111111111111101110011101010100;
assign LUT_2[31270] = 32'b11111111111111111000011101110111;
assign LUT_2[31271] = 32'b11111111111111110101010110010000;
assign LUT_2[31272] = 32'b11111111111111101111111000110000;
assign LUT_2[31273] = 32'b11111111111111101100110001001001;
assign LUT_2[31274] = 32'b11111111111111110110110001101100;
assign LUT_2[31275] = 32'b11111111111111110011101010000101;
assign LUT_2[31276] = 32'b11111111111111101100010110011000;
assign LUT_2[31277] = 32'b11111111111111101001001110110001;
assign LUT_2[31278] = 32'b11111111111111110011001111010100;
assign LUT_2[31279] = 32'b11111111111111110000000111101101;
assign LUT_2[31280] = 32'b11111111111111101111101011011101;
assign LUT_2[31281] = 32'b11111111111111101100100011110110;
assign LUT_2[31282] = 32'b11111111111111110110100100011001;
assign LUT_2[31283] = 32'b11111111111111110011011100110010;
assign LUT_2[31284] = 32'b11111111111111101100001001000101;
assign LUT_2[31285] = 32'b11111111111111101001000001011110;
assign LUT_2[31286] = 32'b11111111111111110011000010000001;
assign LUT_2[31287] = 32'b11111111111111101111111010011010;
assign LUT_2[31288] = 32'b11111111111111101010011100111010;
assign LUT_2[31289] = 32'b11111111111111100111010101010011;
assign LUT_2[31290] = 32'b11111111111111110001010101110110;
assign LUT_2[31291] = 32'b11111111111111101110001110001111;
assign LUT_2[31292] = 32'b11111111111111100110111010100010;
assign LUT_2[31293] = 32'b11111111111111100011110010111011;
assign LUT_2[31294] = 32'b11111111111111101101110011011110;
assign LUT_2[31295] = 32'b11111111111111101010101011110111;
assign LUT_2[31296] = 32'b11111111111111101100110100001101;
assign LUT_2[31297] = 32'b11111111111111101001101100100110;
assign LUT_2[31298] = 32'b11111111111111110011101101001001;
assign LUT_2[31299] = 32'b11111111111111110000100101100010;
assign LUT_2[31300] = 32'b11111111111111101001010001110101;
assign LUT_2[31301] = 32'b11111111111111100110001010001110;
assign LUT_2[31302] = 32'b11111111111111110000001010110001;
assign LUT_2[31303] = 32'b11111111111111101101000011001010;
assign LUT_2[31304] = 32'b11111111111111100111100101101010;
assign LUT_2[31305] = 32'b11111111111111100100011110000011;
assign LUT_2[31306] = 32'b11111111111111101110011110100110;
assign LUT_2[31307] = 32'b11111111111111101011010110111111;
assign LUT_2[31308] = 32'b11111111111111100100000011010010;
assign LUT_2[31309] = 32'b11111111111111100000111011101011;
assign LUT_2[31310] = 32'b11111111111111101010111100001110;
assign LUT_2[31311] = 32'b11111111111111100111110100100111;
assign LUT_2[31312] = 32'b11111111111111100111011000010111;
assign LUT_2[31313] = 32'b11111111111111100100010000110000;
assign LUT_2[31314] = 32'b11111111111111101110010001010011;
assign LUT_2[31315] = 32'b11111111111111101011001001101100;
assign LUT_2[31316] = 32'b11111111111111100011110101111111;
assign LUT_2[31317] = 32'b11111111111111100000101110011000;
assign LUT_2[31318] = 32'b11111111111111101010101110111011;
assign LUT_2[31319] = 32'b11111111111111100111100111010100;
assign LUT_2[31320] = 32'b11111111111111100010001001110100;
assign LUT_2[31321] = 32'b11111111111111011111000010001101;
assign LUT_2[31322] = 32'b11111111111111101001000010110000;
assign LUT_2[31323] = 32'b11111111111111100101111011001001;
assign LUT_2[31324] = 32'b11111111111111011110100111011100;
assign LUT_2[31325] = 32'b11111111111111011011011111110101;
assign LUT_2[31326] = 32'b11111111111111100101100000011000;
assign LUT_2[31327] = 32'b11111111111111100010011000110001;
assign LUT_2[31328] = 32'b11111111111111101101001111110110;
assign LUT_2[31329] = 32'b11111111111111101010001000001111;
assign LUT_2[31330] = 32'b11111111111111110100001000110010;
assign LUT_2[31331] = 32'b11111111111111110001000001001011;
assign LUT_2[31332] = 32'b11111111111111101001101101011110;
assign LUT_2[31333] = 32'b11111111111111100110100101110111;
assign LUT_2[31334] = 32'b11111111111111110000100110011010;
assign LUT_2[31335] = 32'b11111111111111101101011110110011;
assign LUT_2[31336] = 32'b11111111111111101000000001010011;
assign LUT_2[31337] = 32'b11111111111111100100111001101100;
assign LUT_2[31338] = 32'b11111111111111101110111010001111;
assign LUT_2[31339] = 32'b11111111111111101011110010101000;
assign LUT_2[31340] = 32'b11111111111111100100011110111011;
assign LUT_2[31341] = 32'b11111111111111100001010111010100;
assign LUT_2[31342] = 32'b11111111111111101011010111110111;
assign LUT_2[31343] = 32'b11111111111111101000010000010000;
assign LUT_2[31344] = 32'b11111111111111100111110100000000;
assign LUT_2[31345] = 32'b11111111111111100100101100011001;
assign LUT_2[31346] = 32'b11111111111111101110101100111100;
assign LUT_2[31347] = 32'b11111111111111101011100101010101;
assign LUT_2[31348] = 32'b11111111111111100100010001101000;
assign LUT_2[31349] = 32'b11111111111111100001001010000001;
assign LUT_2[31350] = 32'b11111111111111101011001010100100;
assign LUT_2[31351] = 32'b11111111111111101000000010111101;
assign LUT_2[31352] = 32'b11111111111111100010100101011101;
assign LUT_2[31353] = 32'b11111111111111011111011101110110;
assign LUT_2[31354] = 32'b11111111111111101001011110011001;
assign LUT_2[31355] = 32'b11111111111111100110010110110010;
assign LUT_2[31356] = 32'b11111111111111011111000011000101;
assign LUT_2[31357] = 32'b11111111111111011011111011011110;
assign LUT_2[31358] = 32'b11111111111111100101111100000001;
assign LUT_2[31359] = 32'b11111111111111100010110100011010;
assign LUT_2[31360] = 32'b11111111111111111000111111111001;
assign LUT_2[31361] = 32'b11111111111111110101111000010010;
assign LUT_2[31362] = 32'b11111111111111111111111000110101;
assign LUT_2[31363] = 32'b11111111111111111100110001001110;
assign LUT_2[31364] = 32'b11111111111111110101011101100001;
assign LUT_2[31365] = 32'b11111111111111110010010101111010;
assign LUT_2[31366] = 32'b11111111111111111100010110011101;
assign LUT_2[31367] = 32'b11111111111111111001001110110110;
assign LUT_2[31368] = 32'b11111111111111110011110001010110;
assign LUT_2[31369] = 32'b11111111111111110000101001101111;
assign LUT_2[31370] = 32'b11111111111111111010101010010010;
assign LUT_2[31371] = 32'b11111111111111110111100010101011;
assign LUT_2[31372] = 32'b11111111111111110000001110111110;
assign LUT_2[31373] = 32'b11111111111111101101000111010111;
assign LUT_2[31374] = 32'b11111111111111110111000111111010;
assign LUT_2[31375] = 32'b11111111111111110100000000010011;
assign LUT_2[31376] = 32'b11111111111111110011100100000011;
assign LUT_2[31377] = 32'b11111111111111110000011100011100;
assign LUT_2[31378] = 32'b11111111111111111010011100111111;
assign LUT_2[31379] = 32'b11111111111111110111010101011000;
assign LUT_2[31380] = 32'b11111111111111110000000001101011;
assign LUT_2[31381] = 32'b11111111111111101100111010000100;
assign LUT_2[31382] = 32'b11111111111111110110111010100111;
assign LUT_2[31383] = 32'b11111111111111110011110011000000;
assign LUT_2[31384] = 32'b11111111111111101110010101100000;
assign LUT_2[31385] = 32'b11111111111111101011001101111001;
assign LUT_2[31386] = 32'b11111111111111110101001110011100;
assign LUT_2[31387] = 32'b11111111111111110010000110110101;
assign LUT_2[31388] = 32'b11111111111111101010110011001000;
assign LUT_2[31389] = 32'b11111111111111100111101011100001;
assign LUT_2[31390] = 32'b11111111111111110001101100000100;
assign LUT_2[31391] = 32'b11111111111111101110100100011101;
assign LUT_2[31392] = 32'b11111111111111111001011011100010;
assign LUT_2[31393] = 32'b11111111111111110110010011111011;
assign LUT_2[31394] = 32'b00000000000000000000010100011110;
assign LUT_2[31395] = 32'b11111111111111111101001100110111;
assign LUT_2[31396] = 32'b11111111111111110101111001001010;
assign LUT_2[31397] = 32'b11111111111111110010110001100011;
assign LUT_2[31398] = 32'b11111111111111111100110010000110;
assign LUT_2[31399] = 32'b11111111111111111001101010011111;
assign LUT_2[31400] = 32'b11111111111111110100001100111111;
assign LUT_2[31401] = 32'b11111111111111110001000101011000;
assign LUT_2[31402] = 32'b11111111111111111011000101111011;
assign LUT_2[31403] = 32'b11111111111111110111111110010100;
assign LUT_2[31404] = 32'b11111111111111110000101010100111;
assign LUT_2[31405] = 32'b11111111111111101101100011000000;
assign LUT_2[31406] = 32'b11111111111111110111100011100011;
assign LUT_2[31407] = 32'b11111111111111110100011011111100;
assign LUT_2[31408] = 32'b11111111111111110011111111101100;
assign LUT_2[31409] = 32'b11111111111111110000111000000101;
assign LUT_2[31410] = 32'b11111111111111111010111000101000;
assign LUT_2[31411] = 32'b11111111111111110111110001000001;
assign LUT_2[31412] = 32'b11111111111111110000011101010100;
assign LUT_2[31413] = 32'b11111111111111101101010101101101;
assign LUT_2[31414] = 32'b11111111111111110111010110010000;
assign LUT_2[31415] = 32'b11111111111111110100001110101001;
assign LUT_2[31416] = 32'b11111111111111101110110001001001;
assign LUT_2[31417] = 32'b11111111111111101011101001100010;
assign LUT_2[31418] = 32'b11111111111111110101101010000101;
assign LUT_2[31419] = 32'b11111111111111110010100010011110;
assign LUT_2[31420] = 32'b11111111111111101011001110110001;
assign LUT_2[31421] = 32'b11111111111111101000000111001010;
assign LUT_2[31422] = 32'b11111111111111110010000111101101;
assign LUT_2[31423] = 32'b11111111111111101111000000000110;
assign LUT_2[31424] = 32'b11111111111111110001001000011100;
assign LUT_2[31425] = 32'b11111111111111101110000000110101;
assign LUT_2[31426] = 32'b11111111111111111000000001011000;
assign LUT_2[31427] = 32'b11111111111111110100111001110001;
assign LUT_2[31428] = 32'b11111111111111101101100110000100;
assign LUT_2[31429] = 32'b11111111111111101010011110011101;
assign LUT_2[31430] = 32'b11111111111111110100011111000000;
assign LUT_2[31431] = 32'b11111111111111110001010111011001;
assign LUT_2[31432] = 32'b11111111111111101011111001111001;
assign LUT_2[31433] = 32'b11111111111111101000110010010010;
assign LUT_2[31434] = 32'b11111111111111110010110010110101;
assign LUT_2[31435] = 32'b11111111111111101111101011001110;
assign LUT_2[31436] = 32'b11111111111111101000010111100001;
assign LUT_2[31437] = 32'b11111111111111100101001111111010;
assign LUT_2[31438] = 32'b11111111111111101111010000011101;
assign LUT_2[31439] = 32'b11111111111111101100001000110110;
assign LUT_2[31440] = 32'b11111111111111101011101100100110;
assign LUT_2[31441] = 32'b11111111111111101000100100111111;
assign LUT_2[31442] = 32'b11111111111111110010100101100010;
assign LUT_2[31443] = 32'b11111111111111101111011101111011;
assign LUT_2[31444] = 32'b11111111111111101000001010001110;
assign LUT_2[31445] = 32'b11111111111111100101000010100111;
assign LUT_2[31446] = 32'b11111111111111101111000011001010;
assign LUT_2[31447] = 32'b11111111111111101011111011100011;
assign LUT_2[31448] = 32'b11111111111111100110011110000011;
assign LUT_2[31449] = 32'b11111111111111100011010110011100;
assign LUT_2[31450] = 32'b11111111111111101101010110111111;
assign LUT_2[31451] = 32'b11111111111111101010001111011000;
assign LUT_2[31452] = 32'b11111111111111100010111011101011;
assign LUT_2[31453] = 32'b11111111111111011111110100000100;
assign LUT_2[31454] = 32'b11111111111111101001110100100111;
assign LUT_2[31455] = 32'b11111111111111100110101101000000;
assign LUT_2[31456] = 32'b11111111111111110001100100000101;
assign LUT_2[31457] = 32'b11111111111111101110011100011110;
assign LUT_2[31458] = 32'b11111111111111111000011101000001;
assign LUT_2[31459] = 32'b11111111111111110101010101011010;
assign LUT_2[31460] = 32'b11111111111111101110000001101101;
assign LUT_2[31461] = 32'b11111111111111101010111010000110;
assign LUT_2[31462] = 32'b11111111111111110100111010101001;
assign LUT_2[31463] = 32'b11111111111111110001110011000010;
assign LUT_2[31464] = 32'b11111111111111101100010101100010;
assign LUT_2[31465] = 32'b11111111111111101001001101111011;
assign LUT_2[31466] = 32'b11111111111111110011001110011110;
assign LUT_2[31467] = 32'b11111111111111110000000110110111;
assign LUT_2[31468] = 32'b11111111111111101000110011001010;
assign LUT_2[31469] = 32'b11111111111111100101101011100011;
assign LUT_2[31470] = 32'b11111111111111101111101100000110;
assign LUT_2[31471] = 32'b11111111111111101100100100011111;
assign LUT_2[31472] = 32'b11111111111111101100001000001111;
assign LUT_2[31473] = 32'b11111111111111101001000000101000;
assign LUT_2[31474] = 32'b11111111111111110011000001001011;
assign LUT_2[31475] = 32'b11111111111111101111111001100100;
assign LUT_2[31476] = 32'b11111111111111101000100101110111;
assign LUT_2[31477] = 32'b11111111111111100101011110010000;
assign LUT_2[31478] = 32'b11111111111111101111011110110011;
assign LUT_2[31479] = 32'b11111111111111101100010111001100;
assign LUT_2[31480] = 32'b11111111111111100110111001101100;
assign LUT_2[31481] = 32'b11111111111111100011110010000101;
assign LUT_2[31482] = 32'b11111111111111101101110010101000;
assign LUT_2[31483] = 32'b11111111111111101010101011000001;
assign LUT_2[31484] = 32'b11111111111111100011010111010100;
assign LUT_2[31485] = 32'b11111111111111100000001111101101;
assign LUT_2[31486] = 32'b11111111111111101010010000010000;
assign LUT_2[31487] = 32'b11111111111111100111001000101001;
assign LUT_2[31488] = 32'b11111111111111111000101010010000;
assign LUT_2[31489] = 32'b11111111111111110101100010101001;
assign LUT_2[31490] = 32'b11111111111111111111100011001100;
assign LUT_2[31491] = 32'b11111111111111111100011011100101;
assign LUT_2[31492] = 32'b11111111111111110101000111111000;
assign LUT_2[31493] = 32'b11111111111111110010000000010001;
assign LUT_2[31494] = 32'b11111111111111111100000000110100;
assign LUT_2[31495] = 32'b11111111111111111000111001001101;
assign LUT_2[31496] = 32'b11111111111111110011011011101101;
assign LUT_2[31497] = 32'b11111111111111110000010100000110;
assign LUT_2[31498] = 32'b11111111111111111010010100101001;
assign LUT_2[31499] = 32'b11111111111111110111001101000010;
assign LUT_2[31500] = 32'b11111111111111101111111001010101;
assign LUT_2[31501] = 32'b11111111111111101100110001101110;
assign LUT_2[31502] = 32'b11111111111111110110110010010001;
assign LUT_2[31503] = 32'b11111111111111110011101010101010;
assign LUT_2[31504] = 32'b11111111111111110011001110011010;
assign LUT_2[31505] = 32'b11111111111111110000000110110011;
assign LUT_2[31506] = 32'b11111111111111111010000111010110;
assign LUT_2[31507] = 32'b11111111111111110110111111101111;
assign LUT_2[31508] = 32'b11111111111111101111101100000010;
assign LUT_2[31509] = 32'b11111111111111101100100100011011;
assign LUT_2[31510] = 32'b11111111111111110110100100111110;
assign LUT_2[31511] = 32'b11111111111111110011011101010111;
assign LUT_2[31512] = 32'b11111111111111101101111111110111;
assign LUT_2[31513] = 32'b11111111111111101010111000010000;
assign LUT_2[31514] = 32'b11111111111111110100111000110011;
assign LUT_2[31515] = 32'b11111111111111110001110001001100;
assign LUT_2[31516] = 32'b11111111111111101010011101011111;
assign LUT_2[31517] = 32'b11111111111111100111010101111000;
assign LUT_2[31518] = 32'b11111111111111110001010110011011;
assign LUT_2[31519] = 32'b11111111111111101110001110110100;
assign LUT_2[31520] = 32'b11111111111111111001000101111001;
assign LUT_2[31521] = 32'b11111111111111110101111110010010;
assign LUT_2[31522] = 32'b11111111111111111111111110110101;
assign LUT_2[31523] = 32'b11111111111111111100110111001110;
assign LUT_2[31524] = 32'b11111111111111110101100011100001;
assign LUT_2[31525] = 32'b11111111111111110010011011111010;
assign LUT_2[31526] = 32'b11111111111111111100011100011101;
assign LUT_2[31527] = 32'b11111111111111111001010100110110;
assign LUT_2[31528] = 32'b11111111111111110011110111010110;
assign LUT_2[31529] = 32'b11111111111111110000101111101111;
assign LUT_2[31530] = 32'b11111111111111111010110000010010;
assign LUT_2[31531] = 32'b11111111111111110111101000101011;
assign LUT_2[31532] = 32'b11111111111111110000010100111110;
assign LUT_2[31533] = 32'b11111111111111101101001101010111;
assign LUT_2[31534] = 32'b11111111111111110111001101111010;
assign LUT_2[31535] = 32'b11111111111111110100000110010011;
assign LUT_2[31536] = 32'b11111111111111110011101010000011;
assign LUT_2[31537] = 32'b11111111111111110000100010011100;
assign LUT_2[31538] = 32'b11111111111111111010100010111111;
assign LUT_2[31539] = 32'b11111111111111110111011011011000;
assign LUT_2[31540] = 32'b11111111111111110000000111101011;
assign LUT_2[31541] = 32'b11111111111111101101000000000100;
assign LUT_2[31542] = 32'b11111111111111110111000000100111;
assign LUT_2[31543] = 32'b11111111111111110011111001000000;
assign LUT_2[31544] = 32'b11111111111111101110011011100000;
assign LUT_2[31545] = 32'b11111111111111101011010011111001;
assign LUT_2[31546] = 32'b11111111111111110101010100011100;
assign LUT_2[31547] = 32'b11111111111111110010001100110101;
assign LUT_2[31548] = 32'b11111111111111101010111001001000;
assign LUT_2[31549] = 32'b11111111111111100111110001100001;
assign LUT_2[31550] = 32'b11111111111111110001110010000100;
assign LUT_2[31551] = 32'b11111111111111101110101010011101;
assign LUT_2[31552] = 32'b11111111111111110000110010110011;
assign LUT_2[31553] = 32'b11111111111111101101101011001100;
assign LUT_2[31554] = 32'b11111111111111110111101011101111;
assign LUT_2[31555] = 32'b11111111111111110100100100001000;
assign LUT_2[31556] = 32'b11111111111111101101010000011011;
assign LUT_2[31557] = 32'b11111111111111101010001000110100;
assign LUT_2[31558] = 32'b11111111111111110100001001010111;
assign LUT_2[31559] = 32'b11111111111111110001000001110000;
assign LUT_2[31560] = 32'b11111111111111101011100100010000;
assign LUT_2[31561] = 32'b11111111111111101000011100101001;
assign LUT_2[31562] = 32'b11111111111111110010011101001100;
assign LUT_2[31563] = 32'b11111111111111101111010101100101;
assign LUT_2[31564] = 32'b11111111111111101000000001111000;
assign LUT_2[31565] = 32'b11111111111111100100111010010001;
assign LUT_2[31566] = 32'b11111111111111101110111010110100;
assign LUT_2[31567] = 32'b11111111111111101011110011001101;
assign LUT_2[31568] = 32'b11111111111111101011010110111101;
assign LUT_2[31569] = 32'b11111111111111101000001111010110;
assign LUT_2[31570] = 32'b11111111111111110010001111111001;
assign LUT_2[31571] = 32'b11111111111111101111001000010010;
assign LUT_2[31572] = 32'b11111111111111100111110100100101;
assign LUT_2[31573] = 32'b11111111111111100100101100111110;
assign LUT_2[31574] = 32'b11111111111111101110101101100001;
assign LUT_2[31575] = 32'b11111111111111101011100101111010;
assign LUT_2[31576] = 32'b11111111111111100110001000011010;
assign LUT_2[31577] = 32'b11111111111111100011000000110011;
assign LUT_2[31578] = 32'b11111111111111101101000001010110;
assign LUT_2[31579] = 32'b11111111111111101001111001101111;
assign LUT_2[31580] = 32'b11111111111111100010100110000010;
assign LUT_2[31581] = 32'b11111111111111011111011110011011;
assign LUT_2[31582] = 32'b11111111111111101001011110111110;
assign LUT_2[31583] = 32'b11111111111111100110010111010111;
assign LUT_2[31584] = 32'b11111111111111110001001110011100;
assign LUT_2[31585] = 32'b11111111111111101110000110110101;
assign LUT_2[31586] = 32'b11111111111111111000000111011000;
assign LUT_2[31587] = 32'b11111111111111110100111111110001;
assign LUT_2[31588] = 32'b11111111111111101101101100000100;
assign LUT_2[31589] = 32'b11111111111111101010100100011101;
assign LUT_2[31590] = 32'b11111111111111110100100101000000;
assign LUT_2[31591] = 32'b11111111111111110001011101011001;
assign LUT_2[31592] = 32'b11111111111111101011111111111001;
assign LUT_2[31593] = 32'b11111111111111101000111000010010;
assign LUT_2[31594] = 32'b11111111111111110010111000110101;
assign LUT_2[31595] = 32'b11111111111111101111110001001110;
assign LUT_2[31596] = 32'b11111111111111101000011101100001;
assign LUT_2[31597] = 32'b11111111111111100101010101111010;
assign LUT_2[31598] = 32'b11111111111111101111010110011101;
assign LUT_2[31599] = 32'b11111111111111101100001110110110;
assign LUT_2[31600] = 32'b11111111111111101011110010100110;
assign LUT_2[31601] = 32'b11111111111111101000101010111111;
assign LUT_2[31602] = 32'b11111111111111110010101011100010;
assign LUT_2[31603] = 32'b11111111111111101111100011111011;
assign LUT_2[31604] = 32'b11111111111111101000010000001110;
assign LUT_2[31605] = 32'b11111111111111100101001000100111;
assign LUT_2[31606] = 32'b11111111111111101111001001001010;
assign LUT_2[31607] = 32'b11111111111111101100000001100011;
assign LUT_2[31608] = 32'b11111111111111100110100100000011;
assign LUT_2[31609] = 32'b11111111111111100011011100011100;
assign LUT_2[31610] = 32'b11111111111111101101011100111111;
assign LUT_2[31611] = 32'b11111111111111101010010101011000;
assign LUT_2[31612] = 32'b11111111111111100011000001101011;
assign LUT_2[31613] = 32'b11111111111111011111111010000100;
assign LUT_2[31614] = 32'b11111111111111101001111010100111;
assign LUT_2[31615] = 32'b11111111111111100110110011000000;
assign LUT_2[31616] = 32'b11111111111111111100111110011111;
assign LUT_2[31617] = 32'b11111111111111111001110110111000;
assign LUT_2[31618] = 32'b00000000000000000011110111011011;
assign LUT_2[31619] = 32'b00000000000000000000101111110100;
assign LUT_2[31620] = 32'b11111111111111111001011100000111;
assign LUT_2[31621] = 32'b11111111111111110110010100100000;
assign LUT_2[31622] = 32'b00000000000000000000010101000011;
assign LUT_2[31623] = 32'b11111111111111111101001101011100;
assign LUT_2[31624] = 32'b11111111111111110111101111111100;
assign LUT_2[31625] = 32'b11111111111111110100101000010101;
assign LUT_2[31626] = 32'b11111111111111111110101000111000;
assign LUT_2[31627] = 32'b11111111111111111011100001010001;
assign LUT_2[31628] = 32'b11111111111111110100001101100100;
assign LUT_2[31629] = 32'b11111111111111110001000101111101;
assign LUT_2[31630] = 32'b11111111111111111011000110100000;
assign LUT_2[31631] = 32'b11111111111111110111111110111001;
assign LUT_2[31632] = 32'b11111111111111110111100010101001;
assign LUT_2[31633] = 32'b11111111111111110100011011000010;
assign LUT_2[31634] = 32'b11111111111111111110011011100101;
assign LUT_2[31635] = 32'b11111111111111111011010011111110;
assign LUT_2[31636] = 32'b11111111111111110100000000010001;
assign LUT_2[31637] = 32'b11111111111111110000111000101010;
assign LUT_2[31638] = 32'b11111111111111111010111001001101;
assign LUT_2[31639] = 32'b11111111111111110111110001100110;
assign LUT_2[31640] = 32'b11111111111111110010010100000110;
assign LUT_2[31641] = 32'b11111111111111101111001100011111;
assign LUT_2[31642] = 32'b11111111111111111001001101000010;
assign LUT_2[31643] = 32'b11111111111111110110000101011011;
assign LUT_2[31644] = 32'b11111111111111101110110001101110;
assign LUT_2[31645] = 32'b11111111111111101011101010000111;
assign LUT_2[31646] = 32'b11111111111111110101101010101010;
assign LUT_2[31647] = 32'b11111111111111110010100011000011;
assign LUT_2[31648] = 32'b11111111111111111101011010001000;
assign LUT_2[31649] = 32'b11111111111111111010010010100001;
assign LUT_2[31650] = 32'b00000000000000000100010011000100;
assign LUT_2[31651] = 32'b00000000000000000001001011011101;
assign LUT_2[31652] = 32'b11111111111111111001110111110000;
assign LUT_2[31653] = 32'b11111111111111110110110000001001;
assign LUT_2[31654] = 32'b00000000000000000000110000101100;
assign LUT_2[31655] = 32'b11111111111111111101101001000101;
assign LUT_2[31656] = 32'b11111111111111111000001011100101;
assign LUT_2[31657] = 32'b11111111111111110101000011111110;
assign LUT_2[31658] = 32'b11111111111111111111000100100001;
assign LUT_2[31659] = 32'b11111111111111111011111100111010;
assign LUT_2[31660] = 32'b11111111111111110100101001001101;
assign LUT_2[31661] = 32'b11111111111111110001100001100110;
assign LUT_2[31662] = 32'b11111111111111111011100010001001;
assign LUT_2[31663] = 32'b11111111111111111000011010100010;
assign LUT_2[31664] = 32'b11111111111111110111111110010010;
assign LUT_2[31665] = 32'b11111111111111110100110110101011;
assign LUT_2[31666] = 32'b11111111111111111110110111001110;
assign LUT_2[31667] = 32'b11111111111111111011101111100111;
assign LUT_2[31668] = 32'b11111111111111110100011011111010;
assign LUT_2[31669] = 32'b11111111111111110001010100010011;
assign LUT_2[31670] = 32'b11111111111111111011010100110110;
assign LUT_2[31671] = 32'b11111111111111111000001101001111;
assign LUT_2[31672] = 32'b11111111111111110010101111101111;
assign LUT_2[31673] = 32'b11111111111111101111101000001000;
assign LUT_2[31674] = 32'b11111111111111111001101000101011;
assign LUT_2[31675] = 32'b11111111111111110110100001000100;
assign LUT_2[31676] = 32'b11111111111111101111001101010111;
assign LUT_2[31677] = 32'b11111111111111101100000101110000;
assign LUT_2[31678] = 32'b11111111111111110110000110010011;
assign LUT_2[31679] = 32'b11111111111111110010111110101100;
assign LUT_2[31680] = 32'b11111111111111110101000111000010;
assign LUT_2[31681] = 32'b11111111111111110001111111011011;
assign LUT_2[31682] = 32'b11111111111111111011111111111110;
assign LUT_2[31683] = 32'b11111111111111111000111000010111;
assign LUT_2[31684] = 32'b11111111111111110001100100101010;
assign LUT_2[31685] = 32'b11111111111111101110011101000011;
assign LUT_2[31686] = 32'b11111111111111111000011101100110;
assign LUT_2[31687] = 32'b11111111111111110101010101111111;
assign LUT_2[31688] = 32'b11111111111111101111111000011111;
assign LUT_2[31689] = 32'b11111111111111101100110000111000;
assign LUT_2[31690] = 32'b11111111111111110110110001011011;
assign LUT_2[31691] = 32'b11111111111111110011101001110100;
assign LUT_2[31692] = 32'b11111111111111101100010110000111;
assign LUT_2[31693] = 32'b11111111111111101001001110100000;
assign LUT_2[31694] = 32'b11111111111111110011001111000011;
assign LUT_2[31695] = 32'b11111111111111110000000111011100;
assign LUT_2[31696] = 32'b11111111111111101111101011001100;
assign LUT_2[31697] = 32'b11111111111111101100100011100101;
assign LUT_2[31698] = 32'b11111111111111110110100100001000;
assign LUT_2[31699] = 32'b11111111111111110011011100100001;
assign LUT_2[31700] = 32'b11111111111111101100001000110100;
assign LUT_2[31701] = 32'b11111111111111101001000001001101;
assign LUT_2[31702] = 32'b11111111111111110011000001110000;
assign LUT_2[31703] = 32'b11111111111111101111111010001001;
assign LUT_2[31704] = 32'b11111111111111101010011100101001;
assign LUT_2[31705] = 32'b11111111111111100111010101000010;
assign LUT_2[31706] = 32'b11111111111111110001010101100101;
assign LUT_2[31707] = 32'b11111111111111101110001101111110;
assign LUT_2[31708] = 32'b11111111111111100110111010010001;
assign LUT_2[31709] = 32'b11111111111111100011110010101010;
assign LUT_2[31710] = 32'b11111111111111101101110011001101;
assign LUT_2[31711] = 32'b11111111111111101010101011100110;
assign LUT_2[31712] = 32'b11111111111111110101100010101011;
assign LUT_2[31713] = 32'b11111111111111110010011011000100;
assign LUT_2[31714] = 32'b11111111111111111100011011100111;
assign LUT_2[31715] = 32'b11111111111111111001010100000000;
assign LUT_2[31716] = 32'b11111111111111110010000000010011;
assign LUT_2[31717] = 32'b11111111111111101110111000101100;
assign LUT_2[31718] = 32'b11111111111111111000111001001111;
assign LUT_2[31719] = 32'b11111111111111110101110001101000;
assign LUT_2[31720] = 32'b11111111111111110000010100001000;
assign LUT_2[31721] = 32'b11111111111111101101001100100001;
assign LUT_2[31722] = 32'b11111111111111110111001101000100;
assign LUT_2[31723] = 32'b11111111111111110100000101011101;
assign LUT_2[31724] = 32'b11111111111111101100110001110000;
assign LUT_2[31725] = 32'b11111111111111101001101010001001;
assign LUT_2[31726] = 32'b11111111111111110011101010101100;
assign LUT_2[31727] = 32'b11111111111111110000100011000101;
assign LUT_2[31728] = 32'b11111111111111110000000110110101;
assign LUT_2[31729] = 32'b11111111111111101100111111001110;
assign LUT_2[31730] = 32'b11111111111111110110111111110001;
assign LUT_2[31731] = 32'b11111111111111110011111000001010;
assign LUT_2[31732] = 32'b11111111111111101100100100011101;
assign LUT_2[31733] = 32'b11111111111111101001011100110110;
assign LUT_2[31734] = 32'b11111111111111110011011101011001;
assign LUT_2[31735] = 32'b11111111111111110000010101110010;
assign LUT_2[31736] = 32'b11111111111111101010111000010010;
assign LUT_2[31737] = 32'b11111111111111100111110000101011;
assign LUT_2[31738] = 32'b11111111111111110001110001001110;
assign LUT_2[31739] = 32'b11111111111111101110101001100111;
assign LUT_2[31740] = 32'b11111111111111100111010101111010;
assign LUT_2[31741] = 32'b11111111111111100100001110010011;
assign LUT_2[31742] = 32'b11111111111111101110001110110110;
assign LUT_2[31743] = 32'b11111111111111101011000111001111;
assign LUT_2[31744] = 32'b11111111111111110110100101111101;
assign LUT_2[31745] = 32'b11111111111111110011011110010110;
assign LUT_2[31746] = 32'b11111111111111111101011110111001;
assign LUT_2[31747] = 32'b11111111111111111010010111010010;
assign LUT_2[31748] = 32'b11111111111111110011000011100101;
assign LUT_2[31749] = 32'b11111111111111101111111011111110;
assign LUT_2[31750] = 32'b11111111111111111001111100100001;
assign LUT_2[31751] = 32'b11111111111111110110110100111010;
assign LUT_2[31752] = 32'b11111111111111110001010111011010;
assign LUT_2[31753] = 32'b11111111111111101110001111110011;
assign LUT_2[31754] = 32'b11111111111111111000010000010110;
assign LUT_2[31755] = 32'b11111111111111110101001000101111;
assign LUT_2[31756] = 32'b11111111111111101101110101000010;
assign LUT_2[31757] = 32'b11111111111111101010101101011011;
assign LUT_2[31758] = 32'b11111111111111110100101101111110;
assign LUT_2[31759] = 32'b11111111111111110001100110010111;
assign LUT_2[31760] = 32'b11111111111111110001001010000111;
assign LUT_2[31761] = 32'b11111111111111101110000010100000;
assign LUT_2[31762] = 32'b11111111111111111000000011000011;
assign LUT_2[31763] = 32'b11111111111111110100111011011100;
assign LUT_2[31764] = 32'b11111111111111101101100111101111;
assign LUT_2[31765] = 32'b11111111111111101010100000001000;
assign LUT_2[31766] = 32'b11111111111111110100100000101011;
assign LUT_2[31767] = 32'b11111111111111110001011001000100;
assign LUT_2[31768] = 32'b11111111111111101011111011100100;
assign LUT_2[31769] = 32'b11111111111111101000110011111101;
assign LUT_2[31770] = 32'b11111111111111110010110100100000;
assign LUT_2[31771] = 32'b11111111111111101111101100111001;
assign LUT_2[31772] = 32'b11111111111111101000011001001100;
assign LUT_2[31773] = 32'b11111111111111100101010001100101;
assign LUT_2[31774] = 32'b11111111111111101111010010001000;
assign LUT_2[31775] = 32'b11111111111111101100001010100001;
assign LUT_2[31776] = 32'b11111111111111110111000001100110;
assign LUT_2[31777] = 32'b11111111111111110011111001111111;
assign LUT_2[31778] = 32'b11111111111111111101111010100010;
assign LUT_2[31779] = 32'b11111111111111111010110010111011;
assign LUT_2[31780] = 32'b11111111111111110011011111001110;
assign LUT_2[31781] = 32'b11111111111111110000010111100111;
assign LUT_2[31782] = 32'b11111111111111111010011000001010;
assign LUT_2[31783] = 32'b11111111111111110111010000100011;
assign LUT_2[31784] = 32'b11111111111111110001110011000011;
assign LUT_2[31785] = 32'b11111111111111101110101011011100;
assign LUT_2[31786] = 32'b11111111111111111000101011111111;
assign LUT_2[31787] = 32'b11111111111111110101100100011000;
assign LUT_2[31788] = 32'b11111111111111101110010000101011;
assign LUT_2[31789] = 32'b11111111111111101011001001000100;
assign LUT_2[31790] = 32'b11111111111111110101001001100111;
assign LUT_2[31791] = 32'b11111111111111110010000010000000;
assign LUT_2[31792] = 32'b11111111111111110001100101110000;
assign LUT_2[31793] = 32'b11111111111111101110011110001001;
assign LUT_2[31794] = 32'b11111111111111111000011110101100;
assign LUT_2[31795] = 32'b11111111111111110101010111000101;
assign LUT_2[31796] = 32'b11111111111111101110000011011000;
assign LUT_2[31797] = 32'b11111111111111101010111011110001;
assign LUT_2[31798] = 32'b11111111111111110100111100010100;
assign LUT_2[31799] = 32'b11111111111111110001110100101101;
assign LUT_2[31800] = 32'b11111111111111101100010111001101;
assign LUT_2[31801] = 32'b11111111111111101001001111100110;
assign LUT_2[31802] = 32'b11111111111111110011010000001001;
assign LUT_2[31803] = 32'b11111111111111110000001000100010;
assign LUT_2[31804] = 32'b11111111111111101000110100110101;
assign LUT_2[31805] = 32'b11111111111111100101101101001110;
assign LUT_2[31806] = 32'b11111111111111101111101101110001;
assign LUT_2[31807] = 32'b11111111111111101100100110001010;
assign LUT_2[31808] = 32'b11111111111111101110101110100000;
assign LUT_2[31809] = 32'b11111111111111101011100110111001;
assign LUT_2[31810] = 32'b11111111111111110101100111011100;
assign LUT_2[31811] = 32'b11111111111111110010011111110101;
assign LUT_2[31812] = 32'b11111111111111101011001100001000;
assign LUT_2[31813] = 32'b11111111111111101000000100100001;
assign LUT_2[31814] = 32'b11111111111111110010000101000100;
assign LUT_2[31815] = 32'b11111111111111101110111101011101;
assign LUT_2[31816] = 32'b11111111111111101001011111111101;
assign LUT_2[31817] = 32'b11111111111111100110011000010110;
assign LUT_2[31818] = 32'b11111111111111110000011000111001;
assign LUT_2[31819] = 32'b11111111111111101101010001010010;
assign LUT_2[31820] = 32'b11111111111111100101111101100101;
assign LUT_2[31821] = 32'b11111111111111100010110101111110;
assign LUT_2[31822] = 32'b11111111111111101100110110100001;
assign LUT_2[31823] = 32'b11111111111111101001101110111010;
assign LUT_2[31824] = 32'b11111111111111101001010010101010;
assign LUT_2[31825] = 32'b11111111111111100110001011000011;
assign LUT_2[31826] = 32'b11111111111111110000001011100110;
assign LUT_2[31827] = 32'b11111111111111101101000011111111;
assign LUT_2[31828] = 32'b11111111111111100101110000010010;
assign LUT_2[31829] = 32'b11111111111111100010101000101011;
assign LUT_2[31830] = 32'b11111111111111101100101001001110;
assign LUT_2[31831] = 32'b11111111111111101001100001100111;
assign LUT_2[31832] = 32'b11111111111111100100000100000111;
assign LUT_2[31833] = 32'b11111111111111100000111100100000;
assign LUT_2[31834] = 32'b11111111111111101010111101000011;
assign LUT_2[31835] = 32'b11111111111111100111110101011100;
assign LUT_2[31836] = 32'b11111111111111100000100001101111;
assign LUT_2[31837] = 32'b11111111111111011101011010001000;
assign LUT_2[31838] = 32'b11111111111111100111011010101011;
assign LUT_2[31839] = 32'b11111111111111100100010011000100;
assign LUT_2[31840] = 32'b11111111111111101111001010001001;
assign LUT_2[31841] = 32'b11111111111111101100000010100010;
assign LUT_2[31842] = 32'b11111111111111110110000011000101;
assign LUT_2[31843] = 32'b11111111111111110010111011011110;
assign LUT_2[31844] = 32'b11111111111111101011100111110001;
assign LUT_2[31845] = 32'b11111111111111101000100000001010;
assign LUT_2[31846] = 32'b11111111111111110010100000101101;
assign LUT_2[31847] = 32'b11111111111111101111011001000110;
assign LUT_2[31848] = 32'b11111111111111101001111011100110;
assign LUT_2[31849] = 32'b11111111111111100110110011111111;
assign LUT_2[31850] = 32'b11111111111111110000110100100010;
assign LUT_2[31851] = 32'b11111111111111101101101100111011;
assign LUT_2[31852] = 32'b11111111111111100110011001001110;
assign LUT_2[31853] = 32'b11111111111111100011010001100111;
assign LUT_2[31854] = 32'b11111111111111101101010010001010;
assign LUT_2[31855] = 32'b11111111111111101010001010100011;
assign LUT_2[31856] = 32'b11111111111111101001101110010011;
assign LUT_2[31857] = 32'b11111111111111100110100110101100;
assign LUT_2[31858] = 32'b11111111111111110000100111001111;
assign LUT_2[31859] = 32'b11111111111111101101011111101000;
assign LUT_2[31860] = 32'b11111111111111100110001011111011;
assign LUT_2[31861] = 32'b11111111111111100011000100010100;
assign LUT_2[31862] = 32'b11111111111111101101000100110111;
assign LUT_2[31863] = 32'b11111111111111101001111101010000;
assign LUT_2[31864] = 32'b11111111111111100100011111110000;
assign LUT_2[31865] = 32'b11111111111111100001011000001001;
assign LUT_2[31866] = 32'b11111111111111101011011000101100;
assign LUT_2[31867] = 32'b11111111111111101000010001000101;
assign LUT_2[31868] = 32'b11111111111111100000111101011000;
assign LUT_2[31869] = 32'b11111111111111011101110101110001;
assign LUT_2[31870] = 32'b11111111111111100111110110010100;
assign LUT_2[31871] = 32'b11111111111111100100101110101101;
assign LUT_2[31872] = 32'b11111111111111111010111010001100;
assign LUT_2[31873] = 32'b11111111111111110111110010100101;
assign LUT_2[31874] = 32'b00000000000000000001110011001000;
assign LUT_2[31875] = 32'b11111111111111111110101011100001;
assign LUT_2[31876] = 32'b11111111111111110111010111110100;
assign LUT_2[31877] = 32'b11111111111111110100010000001101;
assign LUT_2[31878] = 32'b11111111111111111110010000110000;
assign LUT_2[31879] = 32'b11111111111111111011001001001001;
assign LUT_2[31880] = 32'b11111111111111110101101011101001;
assign LUT_2[31881] = 32'b11111111111111110010100100000010;
assign LUT_2[31882] = 32'b11111111111111111100100100100101;
assign LUT_2[31883] = 32'b11111111111111111001011100111110;
assign LUT_2[31884] = 32'b11111111111111110010001001010001;
assign LUT_2[31885] = 32'b11111111111111101111000001101010;
assign LUT_2[31886] = 32'b11111111111111111001000010001101;
assign LUT_2[31887] = 32'b11111111111111110101111010100110;
assign LUT_2[31888] = 32'b11111111111111110101011110010110;
assign LUT_2[31889] = 32'b11111111111111110010010110101111;
assign LUT_2[31890] = 32'b11111111111111111100010111010010;
assign LUT_2[31891] = 32'b11111111111111111001001111101011;
assign LUT_2[31892] = 32'b11111111111111110001111011111110;
assign LUT_2[31893] = 32'b11111111111111101110110100010111;
assign LUT_2[31894] = 32'b11111111111111111000110100111010;
assign LUT_2[31895] = 32'b11111111111111110101101101010011;
assign LUT_2[31896] = 32'b11111111111111110000001111110011;
assign LUT_2[31897] = 32'b11111111111111101101001000001100;
assign LUT_2[31898] = 32'b11111111111111110111001000101111;
assign LUT_2[31899] = 32'b11111111111111110100000001001000;
assign LUT_2[31900] = 32'b11111111111111101100101101011011;
assign LUT_2[31901] = 32'b11111111111111101001100101110100;
assign LUT_2[31902] = 32'b11111111111111110011100110010111;
assign LUT_2[31903] = 32'b11111111111111110000011110110000;
assign LUT_2[31904] = 32'b11111111111111111011010101110101;
assign LUT_2[31905] = 32'b11111111111111111000001110001110;
assign LUT_2[31906] = 32'b00000000000000000010001110110001;
assign LUT_2[31907] = 32'b11111111111111111111000111001010;
assign LUT_2[31908] = 32'b11111111111111110111110011011101;
assign LUT_2[31909] = 32'b11111111111111110100101011110110;
assign LUT_2[31910] = 32'b11111111111111111110101100011001;
assign LUT_2[31911] = 32'b11111111111111111011100100110010;
assign LUT_2[31912] = 32'b11111111111111110110000111010010;
assign LUT_2[31913] = 32'b11111111111111110010111111101011;
assign LUT_2[31914] = 32'b11111111111111111101000000001110;
assign LUT_2[31915] = 32'b11111111111111111001111000100111;
assign LUT_2[31916] = 32'b11111111111111110010100100111010;
assign LUT_2[31917] = 32'b11111111111111101111011101010011;
assign LUT_2[31918] = 32'b11111111111111111001011101110110;
assign LUT_2[31919] = 32'b11111111111111110110010110001111;
assign LUT_2[31920] = 32'b11111111111111110101111001111111;
assign LUT_2[31921] = 32'b11111111111111110010110010011000;
assign LUT_2[31922] = 32'b11111111111111111100110010111011;
assign LUT_2[31923] = 32'b11111111111111111001101011010100;
assign LUT_2[31924] = 32'b11111111111111110010010111100111;
assign LUT_2[31925] = 32'b11111111111111101111010000000000;
assign LUT_2[31926] = 32'b11111111111111111001010000100011;
assign LUT_2[31927] = 32'b11111111111111110110001000111100;
assign LUT_2[31928] = 32'b11111111111111110000101011011100;
assign LUT_2[31929] = 32'b11111111111111101101100011110101;
assign LUT_2[31930] = 32'b11111111111111110111100100011000;
assign LUT_2[31931] = 32'b11111111111111110100011100110001;
assign LUT_2[31932] = 32'b11111111111111101101001001000100;
assign LUT_2[31933] = 32'b11111111111111101010000001011101;
assign LUT_2[31934] = 32'b11111111111111110100000010000000;
assign LUT_2[31935] = 32'b11111111111111110000111010011001;
assign LUT_2[31936] = 32'b11111111111111110011000010101111;
assign LUT_2[31937] = 32'b11111111111111101111111011001000;
assign LUT_2[31938] = 32'b11111111111111111001111011101011;
assign LUT_2[31939] = 32'b11111111111111110110110100000100;
assign LUT_2[31940] = 32'b11111111111111101111100000010111;
assign LUT_2[31941] = 32'b11111111111111101100011000110000;
assign LUT_2[31942] = 32'b11111111111111110110011001010011;
assign LUT_2[31943] = 32'b11111111111111110011010001101100;
assign LUT_2[31944] = 32'b11111111111111101101110100001100;
assign LUT_2[31945] = 32'b11111111111111101010101100100101;
assign LUT_2[31946] = 32'b11111111111111110100101101001000;
assign LUT_2[31947] = 32'b11111111111111110001100101100001;
assign LUT_2[31948] = 32'b11111111111111101010010001110100;
assign LUT_2[31949] = 32'b11111111111111100111001010001101;
assign LUT_2[31950] = 32'b11111111111111110001001010110000;
assign LUT_2[31951] = 32'b11111111111111101110000011001001;
assign LUT_2[31952] = 32'b11111111111111101101100110111001;
assign LUT_2[31953] = 32'b11111111111111101010011111010010;
assign LUT_2[31954] = 32'b11111111111111110100011111110101;
assign LUT_2[31955] = 32'b11111111111111110001011000001110;
assign LUT_2[31956] = 32'b11111111111111101010000100100001;
assign LUT_2[31957] = 32'b11111111111111100110111100111010;
assign LUT_2[31958] = 32'b11111111111111110000111101011101;
assign LUT_2[31959] = 32'b11111111111111101101110101110110;
assign LUT_2[31960] = 32'b11111111111111101000011000010110;
assign LUT_2[31961] = 32'b11111111111111100101010000101111;
assign LUT_2[31962] = 32'b11111111111111101111010001010010;
assign LUT_2[31963] = 32'b11111111111111101100001001101011;
assign LUT_2[31964] = 32'b11111111111111100100110101111110;
assign LUT_2[31965] = 32'b11111111111111100001101110010111;
assign LUT_2[31966] = 32'b11111111111111101011101110111010;
assign LUT_2[31967] = 32'b11111111111111101000100111010011;
assign LUT_2[31968] = 32'b11111111111111110011011110011000;
assign LUT_2[31969] = 32'b11111111111111110000010110110001;
assign LUT_2[31970] = 32'b11111111111111111010010111010100;
assign LUT_2[31971] = 32'b11111111111111110111001111101101;
assign LUT_2[31972] = 32'b11111111111111101111111100000000;
assign LUT_2[31973] = 32'b11111111111111101100110100011001;
assign LUT_2[31974] = 32'b11111111111111110110110100111100;
assign LUT_2[31975] = 32'b11111111111111110011101101010101;
assign LUT_2[31976] = 32'b11111111111111101110001111110101;
assign LUT_2[31977] = 32'b11111111111111101011001000001110;
assign LUT_2[31978] = 32'b11111111111111110101001000110001;
assign LUT_2[31979] = 32'b11111111111111110010000001001010;
assign LUT_2[31980] = 32'b11111111111111101010101101011101;
assign LUT_2[31981] = 32'b11111111111111100111100101110110;
assign LUT_2[31982] = 32'b11111111111111110001100110011001;
assign LUT_2[31983] = 32'b11111111111111101110011110110010;
assign LUT_2[31984] = 32'b11111111111111101110000010100010;
assign LUT_2[31985] = 32'b11111111111111101010111010111011;
assign LUT_2[31986] = 32'b11111111111111110100111011011110;
assign LUT_2[31987] = 32'b11111111111111110001110011110111;
assign LUT_2[31988] = 32'b11111111111111101010100000001010;
assign LUT_2[31989] = 32'b11111111111111100111011000100011;
assign LUT_2[31990] = 32'b11111111111111110001011001000110;
assign LUT_2[31991] = 32'b11111111111111101110010001011111;
assign LUT_2[31992] = 32'b11111111111111101000110011111111;
assign LUT_2[31993] = 32'b11111111111111100101101100011000;
assign LUT_2[31994] = 32'b11111111111111101111101100111011;
assign LUT_2[31995] = 32'b11111111111111101100100101010100;
assign LUT_2[31996] = 32'b11111111111111100101010001100111;
assign LUT_2[31997] = 32'b11111111111111100010001010000000;
assign LUT_2[31998] = 32'b11111111111111101100001010100011;
assign LUT_2[31999] = 32'b11111111111111101001000010111100;
assign LUT_2[32000] = 32'b11111111111111111010100100100011;
assign LUT_2[32001] = 32'b11111111111111110111011100111100;
assign LUT_2[32002] = 32'b00000000000000000001011101011111;
assign LUT_2[32003] = 32'b11111111111111111110010101111000;
assign LUT_2[32004] = 32'b11111111111111110111000010001011;
assign LUT_2[32005] = 32'b11111111111111110011111010100100;
assign LUT_2[32006] = 32'b11111111111111111101111011000111;
assign LUT_2[32007] = 32'b11111111111111111010110011100000;
assign LUT_2[32008] = 32'b11111111111111110101010110000000;
assign LUT_2[32009] = 32'b11111111111111110010001110011001;
assign LUT_2[32010] = 32'b11111111111111111100001110111100;
assign LUT_2[32011] = 32'b11111111111111111001000111010101;
assign LUT_2[32012] = 32'b11111111111111110001110011101000;
assign LUT_2[32013] = 32'b11111111111111101110101100000001;
assign LUT_2[32014] = 32'b11111111111111111000101100100100;
assign LUT_2[32015] = 32'b11111111111111110101100100111101;
assign LUT_2[32016] = 32'b11111111111111110101001000101101;
assign LUT_2[32017] = 32'b11111111111111110010000001000110;
assign LUT_2[32018] = 32'b11111111111111111100000001101001;
assign LUT_2[32019] = 32'b11111111111111111000111010000010;
assign LUT_2[32020] = 32'b11111111111111110001100110010101;
assign LUT_2[32021] = 32'b11111111111111101110011110101110;
assign LUT_2[32022] = 32'b11111111111111111000011111010001;
assign LUT_2[32023] = 32'b11111111111111110101010111101010;
assign LUT_2[32024] = 32'b11111111111111101111111010001010;
assign LUT_2[32025] = 32'b11111111111111101100110010100011;
assign LUT_2[32026] = 32'b11111111111111110110110011000110;
assign LUT_2[32027] = 32'b11111111111111110011101011011111;
assign LUT_2[32028] = 32'b11111111111111101100010111110010;
assign LUT_2[32029] = 32'b11111111111111101001010000001011;
assign LUT_2[32030] = 32'b11111111111111110011010000101110;
assign LUT_2[32031] = 32'b11111111111111110000001001000111;
assign LUT_2[32032] = 32'b11111111111111111011000000001100;
assign LUT_2[32033] = 32'b11111111111111110111111000100101;
assign LUT_2[32034] = 32'b00000000000000000001111001001000;
assign LUT_2[32035] = 32'b11111111111111111110110001100001;
assign LUT_2[32036] = 32'b11111111111111110111011101110100;
assign LUT_2[32037] = 32'b11111111111111110100010110001101;
assign LUT_2[32038] = 32'b11111111111111111110010110110000;
assign LUT_2[32039] = 32'b11111111111111111011001111001001;
assign LUT_2[32040] = 32'b11111111111111110101110001101001;
assign LUT_2[32041] = 32'b11111111111111110010101010000010;
assign LUT_2[32042] = 32'b11111111111111111100101010100101;
assign LUT_2[32043] = 32'b11111111111111111001100010111110;
assign LUT_2[32044] = 32'b11111111111111110010001111010001;
assign LUT_2[32045] = 32'b11111111111111101111000111101010;
assign LUT_2[32046] = 32'b11111111111111111001001000001101;
assign LUT_2[32047] = 32'b11111111111111110110000000100110;
assign LUT_2[32048] = 32'b11111111111111110101100100010110;
assign LUT_2[32049] = 32'b11111111111111110010011100101111;
assign LUT_2[32050] = 32'b11111111111111111100011101010010;
assign LUT_2[32051] = 32'b11111111111111111001010101101011;
assign LUT_2[32052] = 32'b11111111111111110010000001111110;
assign LUT_2[32053] = 32'b11111111111111101110111010010111;
assign LUT_2[32054] = 32'b11111111111111111000111010111010;
assign LUT_2[32055] = 32'b11111111111111110101110011010011;
assign LUT_2[32056] = 32'b11111111111111110000010101110011;
assign LUT_2[32057] = 32'b11111111111111101101001110001100;
assign LUT_2[32058] = 32'b11111111111111110111001110101111;
assign LUT_2[32059] = 32'b11111111111111110100000111001000;
assign LUT_2[32060] = 32'b11111111111111101100110011011011;
assign LUT_2[32061] = 32'b11111111111111101001101011110100;
assign LUT_2[32062] = 32'b11111111111111110011101100010111;
assign LUT_2[32063] = 32'b11111111111111110000100100110000;
assign LUT_2[32064] = 32'b11111111111111110010101101000110;
assign LUT_2[32065] = 32'b11111111111111101111100101011111;
assign LUT_2[32066] = 32'b11111111111111111001100110000010;
assign LUT_2[32067] = 32'b11111111111111110110011110011011;
assign LUT_2[32068] = 32'b11111111111111101111001010101110;
assign LUT_2[32069] = 32'b11111111111111101100000011000111;
assign LUT_2[32070] = 32'b11111111111111110110000011101010;
assign LUT_2[32071] = 32'b11111111111111110010111100000011;
assign LUT_2[32072] = 32'b11111111111111101101011110100011;
assign LUT_2[32073] = 32'b11111111111111101010010110111100;
assign LUT_2[32074] = 32'b11111111111111110100010111011111;
assign LUT_2[32075] = 32'b11111111111111110001001111111000;
assign LUT_2[32076] = 32'b11111111111111101001111100001011;
assign LUT_2[32077] = 32'b11111111111111100110110100100100;
assign LUT_2[32078] = 32'b11111111111111110000110101000111;
assign LUT_2[32079] = 32'b11111111111111101101101101100000;
assign LUT_2[32080] = 32'b11111111111111101101010001010000;
assign LUT_2[32081] = 32'b11111111111111101010001001101001;
assign LUT_2[32082] = 32'b11111111111111110100001010001100;
assign LUT_2[32083] = 32'b11111111111111110001000010100101;
assign LUT_2[32084] = 32'b11111111111111101001101110111000;
assign LUT_2[32085] = 32'b11111111111111100110100111010001;
assign LUT_2[32086] = 32'b11111111111111110000100111110100;
assign LUT_2[32087] = 32'b11111111111111101101100000001101;
assign LUT_2[32088] = 32'b11111111111111101000000010101101;
assign LUT_2[32089] = 32'b11111111111111100100111011000110;
assign LUT_2[32090] = 32'b11111111111111101110111011101001;
assign LUT_2[32091] = 32'b11111111111111101011110100000010;
assign LUT_2[32092] = 32'b11111111111111100100100000010101;
assign LUT_2[32093] = 32'b11111111111111100001011000101110;
assign LUT_2[32094] = 32'b11111111111111101011011001010001;
assign LUT_2[32095] = 32'b11111111111111101000010001101010;
assign LUT_2[32096] = 32'b11111111111111110011001000101111;
assign LUT_2[32097] = 32'b11111111111111110000000001001000;
assign LUT_2[32098] = 32'b11111111111111111010000001101011;
assign LUT_2[32099] = 32'b11111111111111110110111010000100;
assign LUT_2[32100] = 32'b11111111111111101111100110010111;
assign LUT_2[32101] = 32'b11111111111111101100011110110000;
assign LUT_2[32102] = 32'b11111111111111110110011111010011;
assign LUT_2[32103] = 32'b11111111111111110011010111101100;
assign LUT_2[32104] = 32'b11111111111111101101111010001100;
assign LUT_2[32105] = 32'b11111111111111101010110010100101;
assign LUT_2[32106] = 32'b11111111111111110100110011001000;
assign LUT_2[32107] = 32'b11111111111111110001101011100001;
assign LUT_2[32108] = 32'b11111111111111101010010111110100;
assign LUT_2[32109] = 32'b11111111111111100111010000001101;
assign LUT_2[32110] = 32'b11111111111111110001010000110000;
assign LUT_2[32111] = 32'b11111111111111101110001001001001;
assign LUT_2[32112] = 32'b11111111111111101101101100111001;
assign LUT_2[32113] = 32'b11111111111111101010100101010010;
assign LUT_2[32114] = 32'b11111111111111110100100101110101;
assign LUT_2[32115] = 32'b11111111111111110001011110001110;
assign LUT_2[32116] = 32'b11111111111111101010001010100001;
assign LUT_2[32117] = 32'b11111111111111100111000010111010;
assign LUT_2[32118] = 32'b11111111111111110001000011011101;
assign LUT_2[32119] = 32'b11111111111111101101111011110110;
assign LUT_2[32120] = 32'b11111111111111101000011110010110;
assign LUT_2[32121] = 32'b11111111111111100101010110101111;
assign LUT_2[32122] = 32'b11111111111111101111010111010010;
assign LUT_2[32123] = 32'b11111111111111101100001111101011;
assign LUT_2[32124] = 32'b11111111111111100100111011111110;
assign LUT_2[32125] = 32'b11111111111111100001110100010111;
assign LUT_2[32126] = 32'b11111111111111101011110100111010;
assign LUT_2[32127] = 32'b11111111111111101000101101010011;
assign LUT_2[32128] = 32'b11111111111111111110111000110010;
assign LUT_2[32129] = 32'b11111111111111111011110001001011;
assign LUT_2[32130] = 32'b00000000000000000101110001101110;
assign LUT_2[32131] = 32'b00000000000000000010101010000111;
assign LUT_2[32132] = 32'b11111111111111111011010110011010;
assign LUT_2[32133] = 32'b11111111111111111000001110110011;
assign LUT_2[32134] = 32'b00000000000000000010001111010110;
assign LUT_2[32135] = 32'b11111111111111111111000111101111;
assign LUT_2[32136] = 32'b11111111111111111001101010001111;
assign LUT_2[32137] = 32'b11111111111111110110100010101000;
assign LUT_2[32138] = 32'b00000000000000000000100011001011;
assign LUT_2[32139] = 32'b11111111111111111101011011100100;
assign LUT_2[32140] = 32'b11111111111111110110000111110111;
assign LUT_2[32141] = 32'b11111111111111110011000000010000;
assign LUT_2[32142] = 32'b11111111111111111101000000110011;
assign LUT_2[32143] = 32'b11111111111111111001111001001100;
assign LUT_2[32144] = 32'b11111111111111111001011100111100;
assign LUT_2[32145] = 32'b11111111111111110110010101010101;
assign LUT_2[32146] = 32'b00000000000000000000010101111000;
assign LUT_2[32147] = 32'b11111111111111111101001110010001;
assign LUT_2[32148] = 32'b11111111111111110101111010100100;
assign LUT_2[32149] = 32'b11111111111111110010110010111101;
assign LUT_2[32150] = 32'b11111111111111111100110011100000;
assign LUT_2[32151] = 32'b11111111111111111001101011111001;
assign LUT_2[32152] = 32'b11111111111111110100001110011001;
assign LUT_2[32153] = 32'b11111111111111110001000110110010;
assign LUT_2[32154] = 32'b11111111111111111011000111010101;
assign LUT_2[32155] = 32'b11111111111111110111111111101110;
assign LUT_2[32156] = 32'b11111111111111110000101100000001;
assign LUT_2[32157] = 32'b11111111111111101101100100011010;
assign LUT_2[32158] = 32'b11111111111111110111100100111101;
assign LUT_2[32159] = 32'b11111111111111110100011101010110;
assign LUT_2[32160] = 32'b11111111111111111111010100011011;
assign LUT_2[32161] = 32'b11111111111111111100001100110100;
assign LUT_2[32162] = 32'b00000000000000000110001101010111;
assign LUT_2[32163] = 32'b00000000000000000011000101110000;
assign LUT_2[32164] = 32'b11111111111111111011110010000011;
assign LUT_2[32165] = 32'b11111111111111111000101010011100;
assign LUT_2[32166] = 32'b00000000000000000010101010111111;
assign LUT_2[32167] = 32'b11111111111111111111100011011000;
assign LUT_2[32168] = 32'b11111111111111111010000101111000;
assign LUT_2[32169] = 32'b11111111111111110110111110010001;
assign LUT_2[32170] = 32'b00000000000000000000111110110100;
assign LUT_2[32171] = 32'b11111111111111111101110111001101;
assign LUT_2[32172] = 32'b11111111111111110110100011100000;
assign LUT_2[32173] = 32'b11111111111111110011011011111001;
assign LUT_2[32174] = 32'b11111111111111111101011100011100;
assign LUT_2[32175] = 32'b11111111111111111010010100110101;
assign LUT_2[32176] = 32'b11111111111111111001111000100101;
assign LUT_2[32177] = 32'b11111111111111110110110000111110;
assign LUT_2[32178] = 32'b00000000000000000000110001100001;
assign LUT_2[32179] = 32'b11111111111111111101101001111010;
assign LUT_2[32180] = 32'b11111111111111110110010110001101;
assign LUT_2[32181] = 32'b11111111111111110011001110100110;
assign LUT_2[32182] = 32'b11111111111111111101001111001001;
assign LUT_2[32183] = 32'b11111111111111111010000111100010;
assign LUT_2[32184] = 32'b11111111111111110100101010000010;
assign LUT_2[32185] = 32'b11111111111111110001100010011011;
assign LUT_2[32186] = 32'b11111111111111111011100010111110;
assign LUT_2[32187] = 32'b11111111111111111000011011010111;
assign LUT_2[32188] = 32'b11111111111111110001000111101010;
assign LUT_2[32189] = 32'b11111111111111101110000000000011;
assign LUT_2[32190] = 32'b11111111111111111000000000100110;
assign LUT_2[32191] = 32'b11111111111111110100111000111111;
assign LUT_2[32192] = 32'b11111111111111110111000001010101;
assign LUT_2[32193] = 32'b11111111111111110011111001101110;
assign LUT_2[32194] = 32'b11111111111111111101111010010001;
assign LUT_2[32195] = 32'b11111111111111111010110010101010;
assign LUT_2[32196] = 32'b11111111111111110011011110111101;
assign LUT_2[32197] = 32'b11111111111111110000010111010110;
assign LUT_2[32198] = 32'b11111111111111111010010111111001;
assign LUT_2[32199] = 32'b11111111111111110111010000010010;
assign LUT_2[32200] = 32'b11111111111111110001110010110010;
assign LUT_2[32201] = 32'b11111111111111101110101011001011;
assign LUT_2[32202] = 32'b11111111111111111000101011101110;
assign LUT_2[32203] = 32'b11111111111111110101100100000111;
assign LUT_2[32204] = 32'b11111111111111101110010000011010;
assign LUT_2[32205] = 32'b11111111111111101011001000110011;
assign LUT_2[32206] = 32'b11111111111111110101001001010110;
assign LUT_2[32207] = 32'b11111111111111110010000001101111;
assign LUT_2[32208] = 32'b11111111111111110001100101011111;
assign LUT_2[32209] = 32'b11111111111111101110011101111000;
assign LUT_2[32210] = 32'b11111111111111111000011110011011;
assign LUT_2[32211] = 32'b11111111111111110101010110110100;
assign LUT_2[32212] = 32'b11111111111111101110000011000111;
assign LUT_2[32213] = 32'b11111111111111101010111011100000;
assign LUT_2[32214] = 32'b11111111111111110100111100000011;
assign LUT_2[32215] = 32'b11111111111111110001110100011100;
assign LUT_2[32216] = 32'b11111111111111101100010110111100;
assign LUT_2[32217] = 32'b11111111111111101001001111010101;
assign LUT_2[32218] = 32'b11111111111111110011001111111000;
assign LUT_2[32219] = 32'b11111111111111110000001000010001;
assign LUT_2[32220] = 32'b11111111111111101000110100100100;
assign LUT_2[32221] = 32'b11111111111111100101101100111101;
assign LUT_2[32222] = 32'b11111111111111101111101101100000;
assign LUT_2[32223] = 32'b11111111111111101100100101111001;
assign LUT_2[32224] = 32'b11111111111111110111011100111110;
assign LUT_2[32225] = 32'b11111111111111110100010101010111;
assign LUT_2[32226] = 32'b11111111111111111110010101111010;
assign LUT_2[32227] = 32'b11111111111111111011001110010011;
assign LUT_2[32228] = 32'b11111111111111110011111010100110;
assign LUT_2[32229] = 32'b11111111111111110000110010111111;
assign LUT_2[32230] = 32'b11111111111111111010110011100010;
assign LUT_2[32231] = 32'b11111111111111110111101011111011;
assign LUT_2[32232] = 32'b11111111111111110010001110011011;
assign LUT_2[32233] = 32'b11111111111111101111000110110100;
assign LUT_2[32234] = 32'b11111111111111111001000111010111;
assign LUT_2[32235] = 32'b11111111111111110101111111110000;
assign LUT_2[32236] = 32'b11111111111111101110101100000011;
assign LUT_2[32237] = 32'b11111111111111101011100100011100;
assign LUT_2[32238] = 32'b11111111111111110101100100111111;
assign LUT_2[32239] = 32'b11111111111111110010011101011000;
assign LUT_2[32240] = 32'b11111111111111110010000001001000;
assign LUT_2[32241] = 32'b11111111111111101110111001100001;
assign LUT_2[32242] = 32'b11111111111111111000111010000100;
assign LUT_2[32243] = 32'b11111111111111110101110010011101;
assign LUT_2[32244] = 32'b11111111111111101110011110110000;
assign LUT_2[32245] = 32'b11111111111111101011010111001001;
assign LUT_2[32246] = 32'b11111111111111110101010111101100;
assign LUT_2[32247] = 32'b11111111111111110010010000000101;
assign LUT_2[32248] = 32'b11111111111111101100110010100101;
assign LUT_2[32249] = 32'b11111111111111101001101010111110;
assign LUT_2[32250] = 32'b11111111111111110011101011100001;
assign LUT_2[32251] = 32'b11111111111111110000100011111010;
assign LUT_2[32252] = 32'b11111111111111101001010000001101;
assign LUT_2[32253] = 32'b11111111111111100110001000100110;
assign LUT_2[32254] = 32'b11111111111111110000001001001001;
assign LUT_2[32255] = 32'b11111111111111101101000001100010;
assign LUT_2[32256] = 32'b11111111111111111011010111101111;
assign LUT_2[32257] = 32'b11111111111111111000010000001000;
assign LUT_2[32258] = 32'b00000000000000000010010000101011;
assign LUT_2[32259] = 32'b11111111111111111111001001000100;
assign LUT_2[32260] = 32'b11111111111111110111110101010111;
assign LUT_2[32261] = 32'b11111111111111110100101101110000;
assign LUT_2[32262] = 32'b11111111111111111110101110010011;
assign LUT_2[32263] = 32'b11111111111111111011100110101100;
assign LUT_2[32264] = 32'b11111111111111110110001001001100;
assign LUT_2[32265] = 32'b11111111111111110011000001100101;
assign LUT_2[32266] = 32'b11111111111111111101000010001000;
assign LUT_2[32267] = 32'b11111111111111111001111010100001;
assign LUT_2[32268] = 32'b11111111111111110010100110110100;
assign LUT_2[32269] = 32'b11111111111111101111011111001101;
assign LUT_2[32270] = 32'b11111111111111111001011111110000;
assign LUT_2[32271] = 32'b11111111111111110110011000001001;
assign LUT_2[32272] = 32'b11111111111111110101111011111001;
assign LUT_2[32273] = 32'b11111111111111110010110100010010;
assign LUT_2[32274] = 32'b11111111111111111100110100110101;
assign LUT_2[32275] = 32'b11111111111111111001101101001110;
assign LUT_2[32276] = 32'b11111111111111110010011001100001;
assign LUT_2[32277] = 32'b11111111111111101111010001111010;
assign LUT_2[32278] = 32'b11111111111111111001010010011101;
assign LUT_2[32279] = 32'b11111111111111110110001010110110;
assign LUT_2[32280] = 32'b11111111111111110000101101010110;
assign LUT_2[32281] = 32'b11111111111111101101100101101111;
assign LUT_2[32282] = 32'b11111111111111110111100110010010;
assign LUT_2[32283] = 32'b11111111111111110100011110101011;
assign LUT_2[32284] = 32'b11111111111111101101001010111110;
assign LUT_2[32285] = 32'b11111111111111101010000011010111;
assign LUT_2[32286] = 32'b11111111111111110100000011111010;
assign LUT_2[32287] = 32'b11111111111111110000111100010011;
assign LUT_2[32288] = 32'b11111111111111111011110011011000;
assign LUT_2[32289] = 32'b11111111111111111000101011110001;
assign LUT_2[32290] = 32'b00000000000000000010101100010100;
assign LUT_2[32291] = 32'b11111111111111111111100100101101;
assign LUT_2[32292] = 32'b11111111111111111000010001000000;
assign LUT_2[32293] = 32'b11111111111111110101001001011001;
assign LUT_2[32294] = 32'b11111111111111111111001001111100;
assign LUT_2[32295] = 32'b11111111111111111100000010010101;
assign LUT_2[32296] = 32'b11111111111111110110100100110101;
assign LUT_2[32297] = 32'b11111111111111110011011101001110;
assign LUT_2[32298] = 32'b11111111111111111101011101110001;
assign LUT_2[32299] = 32'b11111111111111111010010110001010;
assign LUT_2[32300] = 32'b11111111111111110011000010011101;
assign LUT_2[32301] = 32'b11111111111111101111111010110110;
assign LUT_2[32302] = 32'b11111111111111111001111011011001;
assign LUT_2[32303] = 32'b11111111111111110110110011110010;
assign LUT_2[32304] = 32'b11111111111111110110010111100010;
assign LUT_2[32305] = 32'b11111111111111110011001111111011;
assign LUT_2[32306] = 32'b11111111111111111101010000011110;
assign LUT_2[32307] = 32'b11111111111111111010001000110111;
assign LUT_2[32308] = 32'b11111111111111110010110101001010;
assign LUT_2[32309] = 32'b11111111111111101111101101100011;
assign LUT_2[32310] = 32'b11111111111111111001101110000110;
assign LUT_2[32311] = 32'b11111111111111110110100110011111;
assign LUT_2[32312] = 32'b11111111111111110001001000111111;
assign LUT_2[32313] = 32'b11111111111111101110000001011000;
assign LUT_2[32314] = 32'b11111111111111111000000001111011;
assign LUT_2[32315] = 32'b11111111111111110100111010010100;
assign LUT_2[32316] = 32'b11111111111111101101100110100111;
assign LUT_2[32317] = 32'b11111111111111101010011111000000;
assign LUT_2[32318] = 32'b11111111111111110100011111100011;
assign LUT_2[32319] = 32'b11111111111111110001010111111100;
assign LUT_2[32320] = 32'b11111111111111110011100000010010;
assign LUT_2[32321] = 32'b11111111111111110000011000101011;
assign LUT_2[32322] = 32'b11111111111111111010011001001110;
assign LUT_2[32323] = 32'b11111111111111110111010001100111;
assign LUT_2[32324] = 32'b11111111111111101111111101111010;
assign LUT_2[32325] = 32'b11111111111111101100110110010011;
assign LUT_2[32326] = 32'b11111111111111110110110110110110;
assign LUT_2[32327] = 32'b11111111111111110011101111001111;
assign LUT_2[32328] = 32'b11111111111111101110010001101111;
assign LUT_2[32329] = 32'b11111111111111101011001010001000;
assign LUT_2[32330] = 32'b11111111111111110101001010101011;
assign LUT_2[32331] = 32'b11111111111111110010000011000100;
assign LUT_2[32332] = 32'b11111111111111101010101111010111;
assign LUT_2[32333] = 32'b11111111111111100111100111110000;
assign LUT_2[32334] = 32'b11111111111111110001101000010011;
assign LUT_2[32335] = 32'b11111111111111101110100000101100;
assign LUT_2[32336] = 32'b11111111111111101110000100011100;
assign LUT_2[32337] = 32'b11111111111111101010111100110101;
assign LUT_2[32338] = 32'b11111111111111110100111101011000;
assign LUT_2[32339] = 32'b11111111111111110001110101110001;
assign LUT_2[32340] = 32'b11111111111111101010100010000100;
assign LUT_2[32341] = 32'b11111111111111100111011010011101;
assign LUT_2[32342] = 32'b11111111111111110001011011000000;
assign LUT_2[32343] = 32'b11111111111111101110010011011001;
assign LUT_2[32344] = 32'b11111111111111101000110101111001;
assign LUT_2[32345] = 32'b11111111111111100101101110010010;
assign LUT_2[32346] = 32'b11111111111111101111101110110101;
assign LUT_2[32347] = 32'b11111111111111101100100111001110;
assign LUT_2[32348] = 32'b11111111111111100101010011100001;
assign LUT_2[32349] = 32'b11111111111111100010001011111010;
assign LUT_2[32350] = 32'b11111111111111101100001100011101;
assign LUT_2[32351] = 32'b11111111111111101001000100110110;
assign LUT_2[32352] = 32'b11111111111111110011111011111011;
assign LUT_2[32353] = 32'b11111111111111110000110100010100;
assign LUT_2[32354] = 32'b11111111111111111010110100110111;
assign LUT_2[32355] = 32'b11111111111111110111101101010000;
assign LUT_2[32356] = 32'b11111111111111110000011001100011;
assign LUT_2[32357] = 32'b11111111111111101101010001111100;
assign LUT_2[32358] = 32'b11111111111111110111010010011111;
assign LUT_2[32359] = 32'b11111111111111110100001010111000;
assign LUT_2[32360] = 32'b11111111111111101110101101011000;
assign LUT_2[32361] = 32'b11111111111111101011100101110001;
assign LUT_2[32362] = 32'b11111111111111110101100110010100;
assign LUT_2[32363] = 32'b11111111111111110010011110101101;
assign LUT_2[32364] = 32'b11111111111111101011001011000000;
assign LUT_2[32365] = 32'b11111111111111101000000011011001;
assign LUT_2[32366] = 32'b11111111111111110010000011111100;
assign LUT_2[32367] = 32'b11111111111111101110111100010101;
assign LUT_2[32368] = 32'b11111111111111101110100000000101;
assign LUT_2[32369] = 32'b11111111111111101011011000011110;
assign LUT_2[32370] = 32'b11111111111111110101011001000001;
assign LUT_2[32371] = 32'b11111111111111110010010001011010;
assign LUT_2[32372] = 32'b11111111111111101010111101101101;
assign LUT_2[32373] = 32'b11111111111111100111110110000110;
assign LUT_2[32374] = 32'b11111111111111110001110110101001;
assign LUT_2[32375] = 32'b11111111111111101110101111000010;
assign LUT_2[32376] = 32'b11111111111111101001010001100010;
assign LUT_2[32377] = 32'b11111111111111100110001001111011;
assign LUT_2[32378] = 32'b11111111111111110000001010011110;
assign LUT_2[32379] = 32'b11111111111111101101000010110111;
assign LUT_2[32380] = 32'b11111111111111100101101111001010;
assign LUT_2[32381] = 32'b11111111111111100010100111100011;
assign LUT_2[32382] = 32'b11111111111111101100101000000110;
assign LUT_2[32383] = 32'b11111111111111101001100000011111;
assign LUT_2[32384] = 32'b11111111111111111111101011111110;
assign LUT_2[32385] = 32'b11111111111111111100100100010111;
assign LUT_2[32386] = 32'b00000000000000000110100100111010;
assign LUT_2[32387] = 32'b00000000000000000011011101010011;
assign LUT_2[32388] = 32'b11111111111111111100001001100110;
assign LUT_2[32389] = 32'b11111111111111111001000001111111;
assign LUT_2[32390] = 32'b00000000000000000011000010100010;
assign LUT_2[32391] = 32'b11111111111111111111111010111011;
assign LUT_2[32392] = 32'b11111111111111111010011101011011;
assign LUT_2[32393] = 32'b11111111111111110111010101110100;
assign LUT_2[32394] = 32'b00000000000000000001010110010111;
assign LUT_2[32395] = 32'b11111111111111111110001110110000;
assign LUT_2[32396] = 32'b11111111111111110110111011000011;
assign LUT_2[32397] = 32'b11111111111111110011110011011100;
assign LUT_2[32398] = 32'b11111111111111111101110011111111;
assign LUT_2[32399] = 32'b11111111111111111010101100011000;
assign LUT_2[32400] = 32'b11111111111111111010010000001000;
assign LUT_2[32401] = 32'b11111111111111110111001000100001;
assign LUT_2[32402] = 32'b00000000000000000001001001000100;
assign LUT_2[32403] = 32'b11111111111111111110000001011101;
assign LUT_2[32404] = 32'b11111111111111110110101101110000;
assign LUT_2[32405] = 32'b11111111111111110011100110001001;
assign LUT_2[32406] = 32'b11111111111111111101100110101100;
assign LUT_2[32407] = 32'b11111111111111111010011111000101;
assign LUT_2[32408] = 32'b11111111111111110101000001100101;
assign LUT_2[32409] = 32'b11111111111111110001111001111110;
assign LUT_2[32410] = 32'b11111111111111111011111010100001;
assign LUT_2[32411] = 32'b11111111111111111000110010111010;
assign LUT_2[32412] = 32'b11111111111111110001011111001101;
assign LUT_2[32413] = 32'b11111111111111101110010111100110;
assign LUT_2[32414] = 32'b11111111111111111000011000001001;
assign LUT_2[32415] = 32'b11111111111111110101010000100010;
assign LUT_2[32416] = 32'b00000000000000000000000111100111;
assign LUT_2[32417] = 32'b11111111111111111101000000000000;
assign LUT_2[32418] = 32'b00000000000000000111000000100011;
assign LUT_2[32419] = 32'b00000000000000000011111000111100;
assign LUT_2[32420] = 32'b11111111111111111100100101001111;
assign LUT_2[32421] = 32'b11111111111111111001011101101000;
assign LUT_2[32422] = 32'b00000000000000000011011110001011;
assign LUT_2[32423] = 32'b00000000000000000000010110100100;
assign LUT_2[32424] = 32'b11111111111111111010111001000100;
assign LUT_2[32425] = 32'b11111111111111110111110001011101;
assign LUT_2[32426] = 32'b00000000000000000001110010000000;
assign LUT_2[32427] = 32'b11111111111111111110101010011001;
assign LUT_2[32428] = 32'b11111111111111110111010110101100;
assign LUT_2[32429] = 32'b11111111111111110100001111000101;
assign LUT_2[32430] = 32'b11111111111111111110001111101000;
assign LUT_2[32431] = 32'b11111111111111111011001000000001;
assign LUT_2[32432] = 32'b11111111111111111010101011110001;
assign LUT_2[32433] = 32'b11111111111111110111100100001010;
assign LUT_2[32434] = 32'b00000000000000000001100100101101;
assign LUT_2[32435] = 32'b11111111111111111110011101000110;
assign LUT_2[32436] = 32'b11111111111111110111001001011001;
assign LUT_2[32437] = 32'b11111111111111110100000001110010;
assign LUT_2[32438] = 32'b11111111111111111110000010010101;
assign LUT_2[32439] = 32'b11111111111111111010111010101110;
assign LUT_2[32440] = 32'b11111111111111110101011101001110;
assign LUT_2[32441] = 32'b11111111111111110010010101100111;
assign LUT_2[32442] = 32'b11111111111111111100010110001010;
assign LUT_2[32443] = 32'b11111111111111111001001110100011;
assign LUT_2[32444] = 32'b11111111111111110001111010110110;
assign LUT_2[32445] = 32'b11111111111111101110110011001111;
assign LUT_2[32446] = 32'b11111111111111111000110011110010;
assign LUT_2[32447] = 32'b11111111111111110101101100001011;
assign LUT_2[32448] = 32'b11111111111111110111110100100001;
assign LUT_2[32449] = 32'b11111111111111110100101100111010;
assign LUT_2[32450] = 32'b11111111111111111110101101011101;
assign LUT_2[32451] = 32'b11111111111111111011100101110110;
assign LUT_2[32452] = 32'b11111111111111110100010010001001;
assign LUT_2[32453] = 32'b11111111111111110001001010100010;
assign LUT_2[32454] = 32'b11111111111111111011001011000101;
assign LUT_2[32455] = 32'b11111111111111111000000011011110;
assign LUT_2[32456] = 32'b11111111111111110010100101111110;
assign LUT_2[32457] = 32'b11111111111111101111011110010111;
assign LUT_2[32458] = 32'b11111111111111111001011110111010;
assign LUT_2[32459] = 32'b11111111111111110110010111010011;
assign LUT_2[32460] = 32'b11111111111111101111000011100110;
assign LUT_2[32461] = 32'b11111111111111101011111011111111;
assign LUT_2[32462] = 32'b11111111111111110101111100100010;
assign LUT_2[32463] = 32'b11111111111111110010110100111011;
assign LUT_2[32464] = 32'b11111111111111110010011000101011;
assign LUT_2[32465] = 32'b11111111111111101111010001000100;
assign LUT_2[32466] = 32'b11111111111111111001010001100111;
assign LUT_2[32467] = 32'b11111111111111110110001010000000;
assign LUT_2[32468] = 32'b11111111111111101110110110010011;
assign LUT_2[32469] = 32'b11111111111111101011101110101100;
assign LUT_2[32470] = 32'b11111111111111110101101111001111;
assign LUT_2[32471] = 32'b11111111111111110010100111101000;
assign LUT_2[32472] = 32'b11111111111111101101001010001000;
assign LUT_2[32473] = 32'b11111111111111101010000010100001;
assign LUT_2[32474] = 32'b11111111111111110100000011000100;
assign LUT_2[32475] = 32'b11111111111111110000111011011101;
assign LUT_2[32476] = 32'b11111111111111101001100111110000;
assign LUT_2[32477] = 32'b11111111111111100110100000001001;
assign LUT_2[32478] = 32'b11111111111111110000100000101100;
assign LUT_2[32479] = 32'b11111111111111101101011001000101;
assign LUT_2[32480] = 32'b11111111111111111000010000001010;
assign LUT_2[32481] = 32'b11111111111111110101001000100011;
assign LUT_2[32482] = 32'b11111111111111111111001001000110;
assign LUT_2[32483] = 32'b11111111111111111100000001011111;
assign LUT_2[32484] = 32'b11111111111111110100101101110010;
assign LUT_2[32485] = 32'b11111111111111110001100110001011;
assign LUT_2[32486] = 32'b11111111111111111011100110101110;
assign LUT_2[32487] = 32'b11111111111111111000011111000111;
assign LUT_2[32488] = 32'b11111111111111110011000001100111;
assign LUT_2[32489] = 32'b11111111111111101111111010000000;
assign LUT_2[32490] = 32'b11111111111111111001111010100011;
assign LUT_2[32491] = 32'b11111111111111110110110010111100;
assign LUT_2[32492] = 32'b11111111111111101111011111001111;
assign LUT_2[32493] = 32'b11111111111111101100010111101000;
assign LUT_2[32494] = 32'b11111111111111110110011000001011;
assign LUT_2[32495] = 32'b11111111111111110011010000100100;
assign LUT_2[32496] = 32'b11111111111111110010110100010100;
assign LUT_2[32497] = 32'b11111111111111101111101100101101;
assign LUT_2[32498] = 32'b11111111111111111001101101010000;
assign LUT_2[32499] = 32'b11111111111111110110100101101001;
assign LUT_2[32500] = 32'b11111111111111101111010001111100;
assign LUT_2[32501] = 32'b11111111111111101100001010010101;
assign LUT_2[32502] = 32'b11111111111111110110001010111000;
assign LUT_2[32503] = 32'b11111111111111110011000011010001;
assign LUT_2[32504] = 32'b11111111111111101101100101110001;
assign LUT_2[32505] = 32'b11111111111111101010011110001010;
assign LUT_2[32506] = 32'b11111111111111110100011110101101;
assign LUT_2[32507] = 32'b11111111111111110001010111000110;
assign LUT_2[32508] = 32'b11111111111111101010000011011001;
assign LUT_2[32509] = 32'b11111111111111100110111011110010;
assign LUT_2[32510] = 32'b11111111111111110000111100010101;
assign LUT_2[32511] = 32'b11111111111111101101110100101110;
assign LUT_2[32512] = 32'b11111111111111111111010110010101;
assign LUT_2[32513] = 32'b11111111111111111100001110101110;
assign LUT_2[32514] = 32'b00000000000000000110001111010001;
assign LUT_2[32515] = 32'b00000000000000000011000111101010;
assign LUT_2[32516] = 32'b11111111111111111011110011111101;
assign LUT_2[32517] = 32'b11111111111111111000101100010110;
assign LUT_2[32518] = 32'b00000000000000000010101100111001;
assign LUT_2[32519] = 32'b11111111111111111111100101010010;
assign LUT_2[32520] = 32'b11111111111111111010000111110010;
assign LUT_2[32521] = 32'b11111111111111110111000000001011;
assign LUT_2[32522] = 32'b00000000000000000001000000101110;
assign LUT_2[32523] = 32'b11111111111111111101111001000111;
assign LUT_2[32524] = 32'b11111111111111110110100101011010;
assign LUT_2[32525] = 32'b11111111111111110011011101110011;
assign LUT_2[32526] = 32'b11111111111111111101011110010110;
assign LUT_2[32527] = 32'b11111111111111111010010110101111;
assign LUT_2[32528] = 32'b11111111111111111001111010011111;
assign LUT_2[32529] = 32'b11111111111111110110110010111000;
assign LUT_2[32530] = 32'b00000000000000000000110011011011;
assign LUT_2[32531] = 32'b11111111111111111101101011110100;
assign LUT_2[32532] = 32'b11111111111111110110011000000111;
assign LUT_2[32533] = 32'b11111111111111110011010000100000;
assign LUT_2[32534] = 32'b11111111111111111101010001000011;
assign LUT_2[32535] = 32'b11111111111111111010001001011100;
assign LUT_2[32536] = 32'b11111111111111110100101011111100;
assign LUT_2[32537] = 32'b11111111111111110001100100010101;
assign LUT_2[32538] = 32'b11111111111111111011100100111000;
assign LUT_2[32539] = 32'b11111111111111111000011101010001;
assign LUT_2[32540] = 32'b11111111111111110001001001100100;
assign LUT_2[32541] = 32'b11111111111111101110000001111101;
assign LUT_2[32542] = 32'b11111111111111111000000010100000;
assign LUT_2[32543] = 32'b11111111111111110100111010111001;
assign LUT_2[32544] = 32'b11111111111111111111110001111110;
assign LUT_2[32545] = 32'b11111111111111111100101010010111;
assign LUT_2[32546] = 32'b00000000000000000110101010111010;
assign LUT_2[32547] = 32'b00000000000000000011100011010011;
assign LUT_2[32548] = 32'b11111111111111111100001111100110;
assign LUT_2[32549] = 32'b11111111111111111001000111111111;
assign LUT_2[32550] = 32'b00000000000000000011001000100010;
assign LUT_2[32551] = 32'b00000000000000000000000000111011;
assign LUT_2[32552] = 32'b11111111111111111010100011011011;
assign LUT_2[32553] = 32'b11111111111111110111011011110100;
assign LUT_2[32554] = 32'b00000000000000000001011100010111;
assign LUT_2[32555] = 32'b11111111111111111110010100110000;
assign LUT_2[32556] = 32'b11111111111111110111000001000011;
assign LUT_2[32557] = 32'b11111111111111110011111001011100;
assign LUT_2[32558] = 32'b11111111111111111101111001111111;
assign LUT_2[32559] = 32'b11111111111111111010110010011000;
assign LUT_2[32560] = 32'b11111111111111111010010110001000;
assign LUT_2[32561] = 32'b11111111111111110111001110100001;
assign LUT_2[32562] = 32'b00000000000000000001001111000100;
assign LUT_2[32563] = 32'b11111111111111111110000111011101;
assign LUT_2[32564] = 32'b11111111111111110110110011110000;
assign LUT_2[32565] = 32'b11111111111111110011101100001001;
assign LUT_2[32566] = 32'b11111111111111111101101100101100;
assign LUT_2[32567] = 32'b11111111111111111010100101000101;
assign LUT_2[32568] = 32'b11111111111111110101000111100101;
assign LUT_2[32569] = 32'b11111111111111110001111111111110;
assign LUT_2[32570] = 32'b11111111111111111100000000100001;
assign LUT_2[32571] = 32'b11111111111111111000111000111010;
assign LUT_2[32572] = 32'b11111111111111110001100101001101;
assign LUT_2[32573] = 32'b11111111111111101110011101100110;
assign LUT_2[32574] = 32'b11111111111111111000011110001001;
assign LUT_2[32575] = 32'b11111111111111110101010110100010;
assign LUT_2[32576] = 32'b11111111111111110111011110111000;
assign LUT_2[32577] = 32'b11111111111111110100010111010001;
assign LUT_2[32578] = 32'b11111111111111111110010111110100;
assign LUT_2[32579] = 32'b11111111111111111011010000001101;
assign LUT_2[32580] = 32'b11111111111111110011111100100000;
assign LUT_2[32581] = 32'b11111111111111110000110100111001;
assign LUT_2[32582] = 32'b11111111111111111010110101011100;
assign LUT_2[32583] = 32'b11111111111111110111101101110101;
assign LUT_2[32584] = 32'b11111111111111110010010000010101;
assign LUT_2[32585] = 32'b11111111111111101111001000101110;
assign LUT_2[32586] = 32'b11111111111111111001001001010001;
assign LUT_2[32587] = 32'b11111111111111110110000001101010;
assign LUT_2[32588] = 32'b11111111111111101110101101111101;
assign LUT_2[32589] = 32'b11111111111111101011100110010110;
assign LUT_2[32590] = 32'b11111111111111110101100110111001;
assign LUT_2[32591] = 32'b11111111111111110010011111010010;
assign LUT_2[32592] = 32'b11111111111111110010000011000010;
assign LUT_2[32593] = 32'b11111111111111101110111011011011;
assign LUT_2[32594] = 32'b11111111111111111000111011111110;
assign LUT_2[32595] = 32'b11111111111111110101110100010111;
assign LUT_2[32596] = 32'b11111111111111101110100000101010;
assign LUT_2[32597] = 32'b11111111111111101011011001000011;
assign LUT_2[32598] = 32'b11111111111111110101011001100110;
assign LUT_2[32599] = 32'b11111111111111110010010001111111;
assign LUT_2[32600] = 32'b11111111111111101100110100011111;
assign LUT_2[32601] = 32'b11111111111111101001101100111000;
assign LUT_2[32602] = 32'b11111111111111110011101101011011;
assign LUT_2[32603] = 32'b11111111111111110000100101110100;
assign LUT_2[32604] = 32'b11111111111111101001010010000111;
assign LUT_2[32605] = 32'b11111111111111100110001010100000;
assign LUT_2[32606] = 32'b11111111111111110000001011000011;
assign LUT_2[32607] = 32'b11111111111111101101000011011100;
assign LUT_2[32608] = 32'b11111111111111110111111010100001;
assign LUT_2[32609] = 32'b11111111111111110100110010111010;
assign LUT_2[32610] = 32'b11111111111111111110110011011101;
assign LUT_2[32611] = 32'b11111111111111111011101011110110;
assign LUT_2[32612] = 32'b11111111111111110100011000001001;
assign LUT_2[32613] = 32'b11111111111111110001010000100010;
assign LUT_2[32614] = 32'b11111111111111111011010001000101;
assign LUT_2[32615] = 32'b11111111111111111000001001011110;
assign LUT_2[32616] = 32'b11111111111111110010101011111110;
assign LUT_2[32617] = 32'b11111111111111101111100100010111;
assign LUT_2[32618] = 32'b11111111111111111001100100111010;
assign LUT_2[32619] = 32'b11111111111111110110011101010011;
assign LUT_2[32620] = 32'b11111111111111101111001001100110;
assign LUT_2[32621] = 32'b11111111111111101100000001111111;
assign LUT_2[32622] = 32'b11111111111111110110000010100010;
assign LUT_2[32623] = 32'b11111111111111110010111010111011;
assign LUT_2[32624] = 32'b11111111111111110010011110101011;
assign LUT_2[32625] = 32'b11111111111111101111010111000100;
assign LUT_2[32626] = 32'b11111111111111111001010111100111;
assign LUT_2[32627] = 32'b11111111111111110110010000000000;
assign LUT_2[32628] = 32'b11111111111111101110111100010011;
assign LUT_2[32629] = 32'b11111111111111101011110100101100;
assign LUT_2[32630] = 32'b11111111111111110101110101001111;
assign LUT_2[32631] = 32'b11111111111111110010101101101000;
assign LUT_2[32632] = 32'b11111111111111101101010000001000;
assign LUT_2[32633] = 32'b11111111111111101010001000100001;
assign LUT_2[32634] = 32'b11111111111111110100001001000100;
assign LUT_2[32635] = 32'b11111111111111110001000001011101;
assign LUT_2[32636] = 32'b11111111111111101001101101110000;
assign LUT_2[32637] = 32'b11111111111111100110100110001001;
assign LUT_2[32638] = 32'b11111111111111110000100110101100;
assign LUT_2[32639] = 32'b11111111111111101101011111000101;
assign LUT_2[32640] = 32'b00000000000000000011101010100100;
assign LUT_2[32641] = 32'b00000000000000000000100010111101;
assign LUT_2[32642] = 32'b00000000000000001010100011100000;
assign LUT_2[32643] = 32'b00000000000000000111011011111001;
assign LUT_2[32644] = 32'b00000000000000000000001000001100;
assign LUT_2[32645] = 32'b11111111111111111101000000100101;
assign LUT_2[32646] = 32'b00000000000000000111000001001000;
assign LUT_2[32647] = 32'b00000000000000000011111001100001;
assign LUT_2[32648] = 32'b11111111111111111110011100000001;
assign LUT_2[32649] = 32'b11111111111111111011010100011010;
assign LUT_2[32650] = 32'b00000000000000000101010100111101;
assign LUT_2[32651] = 32'b00000000000000000010001101010110;
assign LUT_2[32652] = 32'b11111111111111111010111001101001;
assign LUT_2[32653] = 32'b11111111111111110111110010000010;
assign LUT_2[32654] = 32'b00000000000000000001110010100101;
assign LUT_2[32655] = 32'b11111111111111111110101010111110;
assign LUT_2[32656] = 32'b11111111111111111110001110101110;
assign LUT_2[32657] = 32'b11111111111111111011000111000111;
assign LUT_2[32658] = 32'b00000000000000000101000111101010;
assign LUT_2[32659] = 32'b00000000000000000010000000000011;
assign LUT_2[32660] = 32'b11111111111111111010101100010110;
assign LUT_2[32661] = 32'b11111111111111110111100100101111;
assign LUT_2[32662] = 32'b00000000000000000001100101010010;
assign LUT_2[32663] = 32'b11111111111111111110011101101011;
assign LUT_2[32664] = 32'b11111111111111111001000000001011;
assign LUT_2[32665] = 32'b11111111111111110101111000100100;
assign LUT_2[32666] = 32'b11111111111111111111111001000111;
assign LUT_2[32667] = 32'b11111111111111111100110001100000;
assign LUT_2[32668] = 32'b11111111111111110101011101110011;
assign LUT_2[32669] = 32'b11111111111111110010010110001100;
assign LUT_2[32670] = 32'b11111111111111111100010110101111;
assign LUT_2[32671] = 32'b11111111111111111001001111001000;
assign LUT_2[32672] = 32'b00000000000000000100000110001101;
assign LUT_2[32673] = 32'b00000000000000000000111110100110;
assign LUT_2[32674] = 32'b00000000000000001010111111001001;
assign LUT_2[32675] = 32'b00000000000000000111110111100010;
assign LUT_2[32676] = 32'b00000000000000000000100011110101;
assign LUT_2[32677] = 32'b11111111111111111101011100001110;
assign LUT_2[32678] = 32'b00000000000000000111011100110001;
assign LUT_2[32679] = 32'b00000000000000000100010101001010;
assign LUT_2[32680] = 32'b11111111111111111110110111101010;
assign LUT_2[32681] = 32'b11111111111111111011110000000011;
assign LUT_2[32682] = 32'b00000000000000000101110000100110;
assign LUT_2[32683] = 32'b00000000000000000010101000111111;
assign LUT_2[32684] = 32'b11111111111111111011010101010010;
assign LUT_2[32685] = 32'b11111111111111111000001101101011;
assign LUT_2[32686] = 32'b00000000000000000010001110001110;
assign LUT_2[32687] = 32'b11111111111111111111000110100111;
assign LUT_2[32688] = 32'b11111111111111111110101010010111;
assign LUT_2[32689] = 32'b11111111111111111011100010110000;
assign LUT_2[32690] = 32'b00000000000000000101100011010011;
assign LUT_2[32691] = 32'b00000000000000000010011011101100;
assign LUT_2[32692] = 32'b11111111111111111011000111111111;
assign LUT_2[32693] = 32'b11111111111111111000000000011000;
assign LUT_2[32694] = 32'b00000000000000000010000000111011;
assign LUT_2[32695] = 32'b11111111111111111110111001010100;
assign LUT_2[32696] = 32'b11111111111111111001011011110100;
assign LUT_2[32697] = 32'b11111111111111110110010100001101;
assign LUT_2[32698] = 32'b00000000000000000000010100110000;
assign LUT_2[32699] = 32'b11111111111111111101001101001001;
assign LUT_2[32700] = 32'b11111111111111110101111001011100;
assign LUT_2[32701] = 32'b11111111111111110010110001110101;
assign LUT_2[32702] = 32'b11111111111111111100110010011000;
assign LUT_2[32703] = 32'b11111111111111111001101010110001;
assign LUT_2[32704] = 32'b11111111111111111011110011000111;
assign LUT_2[32705] = 32'b11111111111111111000101011100000;
assign LUT_2[32706] = 32'b00000000000000000010101100000011;
assign LUT_2[32707] = 32'b11111111111111111111100100011100;
assign LUT_2[32708] = 32'b11111111111111111000010000101111;
assign LUT_2[32709] = 32'b11111111111111110101001001001000;
assign LUT_2[32710] = 32'b11111111111111111111001001101011;
assign LUT_2[32711] = 32'b11111111111111111100000010000100;
assign LUT_2[32712] = 32'b11111111111111110110100100100100;
assign LUT_2[32713] = 32'b11111111111111110011011100111101;
assign LUT_2[32714] = 32'b11111111111111111101011101100000;
assign LUT_2[32715] = 32'b11111111111111111010010101111001;
assign LUT_2[32716] = 32'b11111111111111110011000010001100;
assign LUT_2[32717] = 32'b11111111111111101111111010100101;
assign LUT_2[32718] = 32'b11111111111111111001111011001000;
assign LUT_2[32719] = 32'b11111111111111110110110011100001;
assign LUT_2[32720] = 32'b11111111111111110110010111010001;
assign LUT_2[32721] = 32'b11111111111111110011001111101010;
assign LUT_2[32722] = 32'b11111111111111111101010000001101;
assign LUT_2[32723] = 32'b11111111111111111010001000100110;
assign LUT_2[32724] = 32'b11111111111111110010110100111001;
assign LUT_2[32725] = 32'b11111111111111101111101101010010;
assign LUT_2[32726] = 32'b11111111111111111001101101110101;
assign LUT_2[32727] = 32'b11111111111111110110100110001110;
assign LUT_2[32728] = 32'b11111111111111110001001000101110;
assign LUT_2[32729] = 32'b11111111111111101110000001000111;
assign LUT_2[32730] = 32'b11111111111111111000000001101010;
assign LUT_2[32731] = 32'b11111111111111110100111010000011;
assign LUT_2[32732] = 32'b11111111111111101101100110010110;
assign LUT_2[32733] = 32'b11111111111111101010011110101111;
assign LUT_2[32734] = 32'b11111111111111110100011111010010;
assign LUT_2[32735] = 32'b11111111111111110001010111101011;
assign LUT_2[32736] = 32'b11111111111111111100001110110000;
assign LUT_2[32737] = 32'b11111111111111111001000111001001;
assign LUT_2[32738] = 32'b00000000000000000011000111101100;
assign LUT_2[32739] = 32'b00000000000000000000000000000101;
assign LUT_2[32740] = 32'b11111111111111111000101100011000;
assign LUT_2[32741] = 32'b11111111111111110101100100110001;
assign LUT_2[32742] = 32'b11111111111111111111100101010100;
assign LUT_2[32743] = 32'b11111111111111111100011101101101;
assign LUT_2[32744] = 32'b11111111111111110111000000001101;
assign LUT_2[32745] = 32'b11111111111111110011111000100110;
assign LUT_2[32746] = 32'b11111111111111111101111001001001;
assign LUT_2[32747] = 32'b11111111111111111010110001100010;
assign LUT_2[32748] = 32'b11111111111111110011011101110101;
assign LUT_2[32749] = 32'b11111111111111110000010110001110;
assign LUT_2[32750] = 32'b11111111111111111010010110110001;
assign LUT_2[32751] = 32'b11111111111111110111001111001010;
assign LUT_2[32752] = 32'b11111111111111110110110010111010;
assign LUT_2[32753] = 32'b11111111111111110011101011010011;
assign LUT_2[32754] = 32'b11111111111111111101101011110110;
assign LUT_2[32755] = 32'b11111111111111111010100100001111;
assign LUT_2[32756] = 32'b11111111111111110011010000100010;
assign LUT_2[32757] = 32'b11111111111111110000001000111011;
assign LUT_2[32758] = 32'b11111111111111111010001001011110;
assign LUT_2[32759] = 32'b11111111111111110111000001110111;
assign LUT_2[32760] = 32'b11111111111111110001100100010111;
assign LUT_2[32761] = 32'b11111111111111101110011100110000;
assign LUT_2[32762] = 32'b11111111111111111000011101010011;
assign LUT_2[32763] = 32'b11111111111111110101010101101100;
assign LUT_2[32764] = 32'b11111111111111101110000001111111;
assign LUT_2[32765] = 32'b11111111111111101010111010011000;
assign LUT_2[32766] = 32'b11111111111111110100111010111011;
assign LUT_2[32767] = 32'b11111111111111110001110011010100;
assign LUT_2[32768] = 32'b11111111111111111000011001111111;
assign LUT_2[32769] = 32'b11111111111111110101010010011000;
assign LUT_2[32770] = 32'b11111111111111111111010010111011;
assign LUT_2[32771] = 32'b11111111111111111100001011010100;
assign LUT_2[32772] = 32'b11111111111111110100110111100111;
assign LUT_2[32773] = 32'b11111111111111110001110000000000;
assign LUT_2[32774] = 32'b11111111111111111011110000100011;
assign LUT_2[32775] = 32'b11111111111111111000101000111100;
assign LUT_2[32776] = 32'b11111111111111110011001011011100;
assign LUT_2[32777] = 32'b11111111111111110000000011110101;
assign LUT_2[32778] = 32'b11111111111111111010000100011000;
assign LUT_2[32779] = 32'b11111111111111110110111100110001;
assign LUT_2[32780] = 32'b11111111111111101111101001000100;
assign LUT_2[32781] = 32'b11111111111111101100100001011101;
assign LUT_2[32782] = 32'b11111111111111110110100010000000;
assign LUT_2[32783] = 32'b11111111111111110011011010011001;
assign LUT_2[32784] = 32'b11111111111111110010111110001001;
assign LUT_2[32785] = 32'b11111111111111101111110110100010;
assign LUT_2[32786] = 32'b11111111111111111001110111000101;
assign LUT_2[32787] = 32'b11111111111111110110101111011110;
assign LUT_2[32788] = 32'b11111111111111101111011011110001;
assign LUT_2[32789] = 32'b11111111111111101100010100001010;
assign LUT_2[32790] = 32'b11111111111111110110010100101101;
assign LUT_2[32791] = 32'b11111111111111110011001101000110;
assign LUT_2[32792] = 32'b11111111111111101101101111100110;
assign LUT_2[32793] = 32'b11111111111111101010100111111111;
assign LUT_2[32794] = 32'b11111111111111110100101000100010;
assign LUT_2[32795] = 32'b11111111111111110001100000111011;
assign LUT_2[32796] = 32'b11111111111111101010001101001110;
assign LUT_2[32797] = 32'b11111111111111100111000101100111;
assign LUT_2[32798] = 32'b11111111111111110001000110001010;
assign LUT_2[32799] = 32'b11111111111111101101111110100011;
assign LUT_2[32800] = 32'b11111111111111111000110101101000;
assign LUT_2[32801] = 32'b11111111111111110101101110000001;
assign LUT_2[32802] = 32'b11111111111111111111101110100100;
assign LUT_2[32803] = 32'b11111111111111111100100110111101;
assign LUT_2[32804] = 32'b11111111111111110101010011010000;
assign LUT_2[32805] = 32'b11111111111111110010001011101001;
assign LUT_2[32806] = 32'b11111111111111111100001100001100;
assign LUT_2[32807] = 32'b11111111111111111001000100100101;
assign LUT_2[32808] = 32'b11111111111111110011100111000101;
assign LUT_2[32809] = 32'b11111111111111110000011111011110;
assign LUT_2[32810] = 32'b11111111111111111010100000000001;
assign LUT_2[32811] = 32'b11111111111111110111011000011010;
assign LUT_2[32812] = 32'b11111111111111110000000100101101;
assign LUT_2[32813] = 32'b11111111111111101100111101000110;
assign LUT_2[32814] = 32'b11111111111111110110111101101001;
assign LUT_2[32815] = 32'b11111111111111110011110110000010;
assign LUT_2[32816] = 32'b11111111111111110011011001110010;
assign LUT_2[32817] = 32'b11111111111111110000010010001011;
assign LUT_2[32818] = 32'b11111111111111111010010010101110;
assign LUT_2[32819] = 32'b11111111111111110111001011000111;
assign LUT_2[32820] = 32'b11111111111111101111110111011010;
assign LUT_2[32821] = 32'b11111111111111101100101111110011;
assign LUT_2[32822] = 32'b11111111111111110110110000010110;
assign LUT_2[32823] = 32'b11111111111111110011101000101111;
assign LUT_2[32824] = 32'b11111111111111101110001011001111;
assign LUT_2[32825] = 32'b11111111111111101011000011101000;
assign LUT_2[32826] = 32'b11111111111111110101000100001011;
assign LUT_2[32827] = 32'b11111111111111110001111100100100;
assign LUT_2[32828] = 32'b11111111111111101010101000110111;
assign LUT_2[32829] = 32'b11111111111111100111100001010000;
assign LUT_2[32830] = 32'b11111111111111110001100001110011;
assign LUT_2[32831] = 32'b11111111111111101110011010001100;
assign LUT_2[32832] = 32'b11111111111111110000100010100010;
assign LUT_2[32833] = 32'b11111111111111101101011010111011;
assign LUT_2[32834] = 32'b11111111111111110111011011011110;
assign LUT_2[32835] = 32'b11111111111111110100010011110111;
assign LUT_2[32836] = 32'b11111111111111101101000000001010;
assign LUT_2[32837] = 32'b11111111111111101001111000100011;
assign LUT_2[32838] = 32'b11111111111111110011111001000110;
assign LUT_2[32839] = 32'b11111111111111110000110001011111;
assign LUT_2[32840] = 32'b11111111111111101011010011111111;
assign LUT_2[32841] = 32'b11111111111111101000001100011000;
assign LUT_2[32842] = 32'b11111111111111110010001100111011;
assign LUT_2[32843] = 32'b11111111111111101111000101010100;
assign LUT_2[32844] = 32'b11111111111111100111110001100111;
assign LUT_2[32845] = 32'b11111111111111100100101010000000;
assign LUT_2[32846] = 32'b11111111111111101110101010100011;
assign LUT_2[32847] = 32'b11111111111111101011100010111100;
assign LUT_2[32848] = 32'b11111111111111101011000110101100;
assign LUT_2[32849] = 32'b11111111111111100111111111000101;
assign LUT_2[32850] = 32'b11111111111111110001111111101000;
assign LUT_2[32851] = 32'b11111111111111101110111000000001;
assign LUT_2[32852] = 32'b11111111111111100111100100010100;
assign LUT_2[32853] = 32'b11111111111111100100011100101101;
assign LUT_2[32854] = 32'b11111111111111101110011101010000;
assign LUT_2[32855] = 32'b11111111111111101011010101101001;
assign LUT_2[32856] = 32'b11111111111111100101111000001001;
assign LUT_2[32857] = 32'b11111111111111100010110000100010;
assign LUT_2[32858] = 32'b11111111111111101100110001000101;
assign LUT_2[32859] = 32'b11111111111111101001101001011110;
assign LUT_2[32860] = 32'b11111111111111100010010101110001;
assign LUT_2[32861] = 32'b11111111111111011111001110001010;
assign LUT_2[32862] = 32'b11111111111111101001001110101101;
assign LUT_2[32863] = 32'b11111111111111100110000111000110;
assign LUT_2[32864] = 32'b11111111111111110000111110001011;
assign LUT_2[32865] = 32'b11111111111111101101110110100100;
assign LUT_2[32866] = 32'b11111111111111110111110111000111;
assign LUT_2[32867] = 32'b11111111111111110100101111100000;
assign LUT_2[32868] = 32'b11111111111111101101011011110011;
assign LUT_2[32869] = 32'b11111111111111101010010100001100;
assign LUT_2[32870] = 32'b11111111111111110100010100101111;
assign LUT_2[32871] = 32'b11111111111111110001001101001000;
assign LUT_2[32872] = 32'b11111111111111101011101111101000;
assign LUT_2[32873] = 32'b11111111111111101000101000000001;
assign LUT_2[32874] = 32'b11111111111111110010101000100100;
assign LUT_2[32875] = 32'b11111111111111101111100000111101;
assign LUT_2[32876] = 32'b11111111111111101000001101010000;
assign LUT_2[32877] = 32'b11111111111111100101000101101001;
assign LUT_2[32878] = 32'b11111111111111101111000110001100;
assign LUT_2[32879] = 32'b11111111111111101011111110100101;
assign LUT_2[32880] = 32'b11111111111111101011100010010101;
assign LUT_2[32881] = 32'b11111111111111101000011010101110;
assign LUT_2[32882] = 32'b11111111111111110010011011010001;
assign LUT_2[32883] = 32'b11111111111111101111010011101010;
assign LUT_2[32884] = 32'b11111111111111100111111111111101;
assign LUT_2[32885] = 32'b11111111111111100100111000010110;
assign LUT_2[32886] = 32'b11111111111111101110111000111001;
assign LUT_2[32887] = 32'b11111111111111101011110001010010;
assign LUT_2[32888] = 32'b11111111111111100110010011110010;
assign LUT_2[32889] = 32'b11111111111111100011001100001011;
assign LUT_2[32890] = 32'b11111111111111101101001100101110;
assign LUT_2[32891] = 32'b11111111111111101010000101000111;
assign LUT_2[32892] = 32'b11111111111111100010110001011010;
assign LUT_2[32893] = 32'b11111111111111011111101001110011;
assign LUT_2[32894] = 32'b11111111111111101001101010010110;
assign LUT_2[32895] = 32'b11111111111111100110100010101111;
assign LUT_2[32896] = 32'b11111111111111111100101110001110;
assign LUT_2[32897] = 32'b11111111111111111001100110100111;
assign LUT_2[32898] = 32'b00000000000000000011100111001010;
assign LUT_2[32899] = 32'b00000000000000000000011111100011;
assign LUT_2[32900] = 32'b11111111111111111001001011110110;
assign LUT_2[32901] = 32'b11111111111111110110000100001111;
assign LUT_2[32902] = 32'b00000000000000000000000100110010;
assign LUT_2[32903] = 32'b11111111111111111100111101001011;
assign LUT_2[32904] = 32'b11111111111111110111011111101011;
assign LUT_2[32905] = 32'b11111111111111110100011000000100;
assign LUT_2[32906] = 32'b11111111111111111110011000100111;
assign LUT_2[32907] = 32'b11111111111111111011010001000000;
assign LUT_2[32908] = 32'b11111111111111110011111101010011;
assign LUT_2[32909] = 32'b11111111111111110000110101101100;
assign LUT_2[32910] = 32'b11111111111111111010110110001111;
assign LUT_2[32911] = 32'b11111111111111110111101110101000;
assign LUT_2[32912] = 32'b11111111111111110111010010011000;
assign LUT_2[32913] = 32'b11111111111111110100001010110001;
assign LUT_2[32914] = 32'b11111111111111111110001011010100;
assign LUT_2[32915] = 32'b11111111111111111011000011101101;
assign LUT_2[32916] = 32'b11111111111111110011110000000000;
assign LUT_2[32917] = 32'b11111111111111110000101000011001;
assign LUT_2[32918] = 32'b11111111111111111010101000111100;
assign LUT_2[32919] = 32'b11111111111111110111100001010101;
assign LUT_2[32920] = 32'b11111111111111110010000011110101;
assign LUT_2[32921] = 32'b11111111111111101110111100001110;
assign LUT_2[32922] = 32'b11111111111111111000111100110001;
assign LUT_2[32923] = 32'b11111111111111110101110101001010;
assign LUT_2[32924] = 32'b11111111111111101110100001011101;
assign LUT_2[32925] = 32'b11111111111111101011011001110110;
assign LUT_2[32926] = 32'b11111111111111110101011010011001;
assign LUT_2[32927] = 32'b11111111111111110010010010110010;
assign LUT_2[32928] = 32'b11111111111111111101001001110111;
assign LUT_2[32929] = 32'b11111111111111111010000010010000;
assign LUT_2[32930] = 32'b00000000000000000100000010110011;
assign LUT_2[32931] = 32'b00000000000000000000111011001100;
assign LUT_2[32932] = 32'b11111111111111111001100111011111;
assign LUT_2[32933] = 32'b11111111111111110110011111111000;
assign LUT_2[32934] = 32'b00000000000000000000100000011011;
assign LUT_2[32935] = 32'b11111111111111111101011000110100;
assign LUT_2[32936] = 32'b11111111111111110111111011010100;
assign LUT_2[32937] = 32'b11111111111111110100110011101101;
assign LUT_2[32938] = 32'b11111111111111111110110100010000;
assign LUT_2[32939] = 32'b11111111111111111011101100101001;
assign LUT_2[32940] = 32'b11111111111111110100011000111100;
assign LUT_2[32941] = 32'b11111111111111110001010001010101;
assign LUT_2[32942] = 32'b11111111111111111011010001111000;
assign LUT_2[32943] = 32'b11111111111111111000001010010001;
assign LUT_2[32944] = 32'b11111111111111110111101110000001;
assign LUT_2[32945] = 32'b11111111111111110100100110011010;
assign LUT_2[32946] = 32'b11111111111111111110100110111101;
assign LUT_2[32947] = 32'b11111111111111111011011111010110;
assign LUT_2[32948] = 32'b11111111111111110100001011101001;
assign LUT_2[32949] = 32'b11111111111111110001000100000010;
assign LUT_2[32950] = 32'b11111111111111111011000100100101;
assign LUT_2[32951] = 32'b11111111111111110111111100111110;
assign LUT_2[32952] = 32'b11111111111111110010011111011110;
assign LUT_2[32953] = 32'b11111111111111101111010111110111;
assign LUT_2[32954] = 32'b11111111111111111001011000011010;
assign LUT_2[32955] = 32'b11111111111111110110010000110011;
assign LUT_2[32956] = 32'b11111111111111101110111101000110;
assign LUT_2[32957] = 32'b11111111111111101011110101011111;
assign LUT_2[32958] = 32'b11111111111111110101110110000010;
assign LUT_2[32959] = 32'b11111111111111110010101110011011;
assign LUT_2[32960] = 32'b11111111111111110100110110110001;
assign LUT_2[32961] = 32'b11111111111111110001101111001010;
assign LUT_2[32962] = 32'b11111111111111111011101111101101;
assign LUT_2[32963] = 32'b11111111111111111000101000000110;
assign LUT_2[32964] = 32'b11111111111111110001010100011001;
assign LUT_2[32965] = 32'b11111111111111101110001100110010;
assign LUT_2[32966] = 32'b11111111111111111000001101010101;
assign LUT_2[32967] = 32'b11111111111111110101000101101110;
assign LUT_2[32968] = 32'b11111111111111101111101000001110;
assign LUT_2[32969] = 32'b11111111111111101100100000100111;
assign LUT_2[32970] = 32'b11111111111111110110100001001010;
assign LUT_2[32971] = 32'b11111111111111110011011001100011;
assign LUT_2[32972] = 32'b11111111111111101100000101110110;
assign LUT_2[32973] = 32'b11111111111111101000111110001111;
assign LUT_2[32974] = 32'b11111111111111110010111110110010;
assign LUT_2[32975] = 32'b11111111111111101111110111001011;
assign LUT_2[32976] = 32'b11111111111111101111011010111011;
assign LUT_2[32977] = 32'b11111111111111101100010011010100;
assign LUT_2[32978] = 32'b11111111111111110110010011110111;
assign LUT_2[32979] = 32'b11111111111111110011001100010000;
assign LUT_2[32980] = 32'b11111111111111101011111000100011;
assign LUT_2[32981] = 32'b11111111111111101000110000111100;
assign LUT_2[32982] = 32'b11111111111111110010110001011111;
assign LUT_2[32983] = 32'b11111111111111101111101001111000;
assign LUT_2[32984] = 32'b11111111111111101010001100011000;
assign LUT_2[32985] = 32'b11111111111111100111000100110001;
assign LUT_2[32986] = 32'b11111111111111110001000101010100;
assign LUT_2[32987] = 32'b11111111111111101101111101101101;
assign LUT_2[32988] = 32'b11111111111111100110101010000000;
assign LUT_2[32989] = 32'b11111111111111100011100010011001;
assign LUT_2[32990] = 32'b11111111111111101101100010111100;
assign LUT_2[32991] = 32'b11111111111111101010011011010101;
assign LUT_2[32992] = 32'b11111111111111110101010010011010;
assign LUT_2[32993] = 32'b11111111111111110010001010110011;
assign LUT_2[32994] = 32'b11111111111111111100001011010110;
assign LUT_2[32995] = 32'b11111111111111111001000011101111;
assign LUT_2[32996] = 32'b11111111111111110001110000000010;
assign LUT_2[32997] = 32'b11111111111111101110101000011011;
assign LUT_2[32998] = 32'b11111111111111111000101000111110;
assign LUT_2[32999] = 32'b11111111111111110101100001010111;
assign LUT_2[33000] = 32'b11111111111111110000000011110111;
assign LUT_2[33001] = 32'b11111111111111101100111100010000;
assign LUT_2[33002] = 32'b11111111111111110110111100110011;
assign LUT_2[33003] = 32'b11111111111111110011110101001100;
assign LUT_2[33004] = 32'b11111111111111101100100001011111;
assign LUT_2[33005] = 32'b11111111111111101001011001111000;
assign LUT_2[33006] = 32'b11111111111111110011011010011011;
assign LUT_2[33007] = 32'b11111111111111110000010010110100;
assign LUT_2[33008] = 32'b11111111111111101111110110100100;
assign LUT_2[33009] = 32'b11111111111111101100101110111101;
assign LUT_2[33010] = 32'b11111111111111110110101111100000;
assign LUT_2[33011] = 32'b11111111111111110011100111111001;
assign LUT_2[33012] = 32'b11111111111111101100010100001100;
assign LUT_2[33013] = 32'b11111111111111101001001100100101;
assign LUT_2[33014] = 32'b11111111111111110011001101001000;
assign LUT_2[33015] = 32'b11111111111111110000000101100001;
assign LUT_2[33016] = 32'b11111111111111101010101000000001;
assign LUT_2[33017] = 32'b11111111111111100111100000011010;
assign LUT_2[33018] = 32'b11111111111111110001100000111101;
assign LUT_2[33019] = 32'b11111111111111101110011001010110;
assign LUT_2[33020] = 32'b11111111111111100111000101101001;
assign LUT_2[33021] = 32'b11111111111111100011111110000010;
assign LUT_2[33022] = 32'b11111111111111101101111110100101;
assign LUT_2[33023] = 32'b11111111111111101010110110111110;
assign LUT_2[33024] = 32'b11111111111111111100011000100101;
assign LUT_2[33025] = 32'b11111111111111111001010000111110;
assign LUT_2[33026] = 32'b00000000000000000011010001100001;
assign LUT_2[33027] = 32'b00000000000000000000001001111010;
assign LUT_2[33028] = 32'b11111111111111111000110110001101;
assign LUT_2[33029] = 32'b11111111111111110101101110100110;
assign LUT_2[33030] = 32'b11111111111111111111101111001001;
assign LUT_2[33031] = 32'b11111111111111111100100111100010;
assign LUT_2[33032] = 32'b11111111111111110111001010000010;
assign LUT_2[33033] = 32'b11111111111111110100000010011011;
assign LUT_2[33034] = 32'b11111111111111111110000010111110;
assign LUT_2[33035] = 32'b11111111111111111010111011010111;
assign LUT_2[33036] = 32'b11111111111111110011100111101010;
assign LUT_2[33037] = 32'b11111111111111110000100000000011;
assign LUT_2[33038] = 32'b11111111111111111010100000100110;
assign LUT_2[33039] = 32'b11111111111111110111011000111111;
assign LUT_2[33040] = 32'b11111111111111110110111100101111;
assign LUT_2[33041] = 32'b11111111111111110011110101001000;
assign LUT_2[33042] = 32'b11111111111111111101110101101011;
assign LUT_2[33043] = 32'b11111111111111111010101110000100;
assign LUT_2[33044] = 32'b11111111111111110011011010010111;
assign LUT_2[33045] = 32'b11111111111111110000010010110000;
assign LUT_2[33046] = 32'b11111111111111111010010011010011;
assign LUT_2[33047] = 32'b11111111111111110111001011101100;
assign LUT_2[33048] = 32'b11111111111111110001101110001100;
assign LUT_2[33049] = 32'b11111111111111101110100110100101;
assign LUT_2[33050] = 32'b11111111111111111000100111001000;
assign LUT_2[33051] = 32'b11111111111111110101011111100001;
assign LUT_2[33052] = 32'b11111111111111101110001011110100;
assign LUT_2[33053] = 32'b11111111111111101011000100001101;
assign LUT_2[33054] = 32'b11111111111111110101000100110000;
assign LUT_2[33055] = 32'b11111111111111110001111101001001;
assign LUT_2[33056] = 32'b11111111111111111100110100001110;
assign LUT_2[33057] = 32'b11111111111111111001101100100111;
assign LUT_2[33058] = 32'b00000000000000000011101101001010;
assign LUT_2[33059] = 32'b00000000000000000000100101100011;
assign LUT_2[33060] = 32'b11111111111111111001010001110110;
assign LUT_2[33061] = 32'b11111111111111110110001010001111;
assign LUT_2[33062] = 32'b00000000000000000000001010110010;
assign LUT_2[33063] = 32'b11111111111111111101000011001011;
assign LUT_2[33064] = 32'b11111111111111110111100101101011;
assign LUT_2[33065] = 32'b11111111111111110100011110000100;
assign LUT_2[33066] = 32'b11111111111111111110011110100111;
assign LUT_2[33067] = 32'b11111111111111111011010111000000;
assign LUT_2[33068] = 32'b11111111111111110100000011010011;
assign LUT_2[33069] = 32'b11111111111111110000111011101100;
assign LUT_2[33070] = 32'b11111111111111111010111100001111;
assign LUT_2[33071] = 32'b11111111111111110111110100101000;
assign LUT_2[33072] = 32'b11111111111111110111011000011000;
assign LUT_2[33073] = 32'b11111111111111110100010000110001;
assign LUT_2[33074] = 32'b11111111111111111110010001010100;
assign LUT_2[33075] = 32'b11111111111111111011001001101101;
assign LUT_2[33076] = 32'b11111111111111110011110110000000;
assign LUT_2[33077] = 32'b11111111111111110000101110011001;
assign LUT_2[33078] = 32'b11111111111111111010101110111100;
assign LUT_2[33079] = 32'b11111111111111110111100111010101;
assign LUT_2[33080] = 32'b11111111111111110010001001110101;
assign LUT_2[33081] = 32'b11111111111111101111000010001110;
assign LUT_2[33082] = 32'b11111111111111111001000010110001;
assign LUT_2[33083] = 32'b11111111111111110101111011001010;
assign LUT_2[33084] = 32'b11111111111111101110100111011101;
assign LUT_2[33085] = 32'b11111111111111101011011111110110;
assign LUT_2[33086] = 32'b11111111111111110101100000011001;
assign LUT_2[33087] = 32'b11111111111111110010011000110010;
assign LUT_2[33088] = 32'b11111111111111110100100001001000;
assign LUT_2[33089] = 32'b11111111111111110001011001100001;
assign LUT_2[33090] = 32'b11111111111111111011011010000100;
assign LUT_2[33091] = 32'b11111111111111111000010010011101;
assign LUT_2[33092] = 32'b11111111111111110000111110110000;
assign LUT_2[33093] = 32'b11111111111111101101110111001001;
assign LUT_2[33094] = 32'b11111111111111110111110111101100;
assign LUT_2[33095] = 32'b11111111111111110100110000000101;
assign LUT_2[33096] = 32'b11111111111111101111010010100101;
assign LUT_2[33097] = 32'b11111111111111101100001010111110;
assign LUT_2[33098] = 32'b11111111111111110110001011100001;
assign LUT_2[33099] = 32'b11111111111111110011000011111010;
assign LUT_2[33100] = 32'b11111111111111101011110000001101;
assign LUT_2[33101] = 32'b11111111111111101000101000100110;
assign LUT_2[33102] = 32'b11111111111111110010101001001001;
assign LUT_2[33103] = 32'b11111111111111101111100001100010;
assign LUT_2[33104] = 32'b11111111111111101111000101010010;
assign LUT_2[33105] = 32'b11111111111111101011111101101011;
assign LUT_2[33106] = 32'b11111111111111110101111110001110;
assign LUT_2[33107] = 32'b11111111111111110010110110100111;
assign LUT_2[33108] = 32'b11111111111111101011100010111010;
assign LUT_2[33109] = 32'b11111111111111101000011011010011;
assign LUT_2[33110] = 32'b11111111111111110010011011110110;
assign LUT_2[33111] = 32'b11111111111111101111010100001111;
assign LUT_2[33112] = 32'b11111111111111101001110110101111;
assign LUT_2[33113] = 32'b11111111111111100110101111001000;
assign LUT_2[33114] = 32'b11111111111111110000101111101011;
assign LUT_2[33115] = 32'b11111111111111101101101000000100;
assign LUT_2[33116] = 32'b11111111111111100110010100010111;
assign LUT_2[33117] = 32'b11111111111111100011001100110000;
assign LUT_2[33118] = 32'b11111111111111101101001101010011;
assign LUT_2[33119] = 32'b11111111111111101010000101101100;
assign LUT_2[33120] = 32'b11111111111111110100111100110001;
assign LUT_2[33121] = 32'b11111111111111110001110101001010;
assign LUT_2[33122] = 32'b11111111111111111011110101101101;
assign LUT_2[33123] = 32'b11111111111111111000101110000110;
assign LUT_2[33124] = 32'b11111111111111110001011010011001;
assign LUT_2[33125] = 32'b11111111111111101110010010110010;
assign LUT_2[33126] = 32'b11111111111111111000010011010101;
assign LUT_2[33127] = 32'b11111111111111110101001011101110;
assign LUT_2[33128] = 32'b11111111111111101111101110001110;
assign LUT_2[33129] = 32'b11111111111111101100100110100111;
assign LUT_2[33130] = 32'b11111111111111110110100111001010;
assign LUT_2[33131] = 32'b11111111111111110011011111100011;
assign LUT_2[33132] = 32'b11111111111111101100001011110110;
assign LUT_2[33133] = 32'b11111111111111101001000100001111;
assign LUT_2[33134] = 32'b11111111111111110011000100110010;
assign LUT_2[33135] = 32'b11111111111111101111111101001011;
assign LUT_2[33136] = 32'b11111111111111101111100000111011;
assign LUT_2[33137] = 32'b11111111111111101100011001010100;
assign LUT_2[33138] = 32'b11111111111111110110011001110111;
assign LUT_2[33139] = 32'b11111111111111110011010010010000;
assign LUT_2[33140] = 32'b11111111111111101011111110100011;
assign LUT_2[33141] = 32'b11111111111111101000110110111100;
assign LUT_2[33142] = 32'b11111111111111110010110111011111;
assign LUT_2[33143] = 32'b11111111111111101111101111111000;
assign LUT_2[33144] = 32'b11111111111111101010010010011000;
assign LUT_2[33145] = 32'b11111111111111100111001010110001;
assign LUT_2[33146] = 32'b11111111111111110001001011010100;
assign LUT_2[33147] = 32'b11111111111111101110000011101101;
assign LUT_2[33148] = 32'b11111111111111100110110000000000;
assign LUT_2[33149] = 32'b11111111111111100011101000011001;
assign LUT_2[33150] = 32'b11111111111111101101101000111100;
assign LUT_2[33151] = 32'b11111111111111101010100001010101;
assign LUT_2[33152] = 32'b00000000000000000000101100110100;
assign LUT_2[33153] = 32'b11111111111111111101100101001101;
assign LUT_2[33154] = 32'b00000000000000000111100101110000;
assign LUT_2[33155] = 32'b00000000000000000100011110001001;
assign LUT_2[33156] = 32'b11111111111111111101001010011100;
assign LUT_2[33157] = 32'b11111111111111111010000010110101;
assign LUT_2[33158] = 32'b00000000000000000100000011011000;
assign LUT_2[33159] = 32'b00000000000000000000111011110001;
assign LUT_2[33160] = 32'b11111111111111111011011110010001;
assign LUT_2[33161] = 32'b11111111111111111000010110101010;
assign LUT_2[33162] = 32'b00000000000000000010010111001101;
assign LUT_2[33163] = 32'b11111111111111111111001111100110;
assign LUT_2[33164] = 32'b11111111111111110111111011111001;
assign LUT_2[33165] = 32'b11111111111111110100110100010010;
assign LUT_2[33166] = 32'b11111111111111111110110100110101;
assign LUT_2[33167] = 32'b11111111111111111011101101001110;
assign LUT_2[33168] = 32'b11111111111111111011010000111110;
assign LUT_2[33169] = 32'b11111111111111111000001001010111;
assign LUT_2[33170] = 32'b00000000000000000010001001111010;
assign LUT_2[33171] = 32'b11111111111111111111000010010011;
assign LUT_2[33172] = 32'b11111111111111110111101110100110;
assign LUT_2[33173] = 32'b11111111111111110100100110111111;
assign LUT_2[33174] = 32'b11111111111111111110100111100010;
assign LUT_2[33175] = 32'b11111111111111111011011111111011;
assign LUT_2[33176] = 32'b11111111111111110110000010011011;
assign LUT_2[33177] = 32'b11111111111111110010111010110100;
assign LUT_2[33178] = 32'b11111111111111111100111011010111;
assign LUT_2[33179] = 32'b11111111111111111001110011110000;
assign LUT_2[33180] = 32'b11111111111111110010100000000011;
assign LUT_2[33181] = 32'b11111111111111101111011000011100;
assign LUT_2[33182] = 32'b11111111111111111001011000111111;
assign LUT_2[33183] = 32'b11111111111111110110010001011000;
assign LUT_2[33184] = 32'b00000000000000000001001000011101;
assign LUT_2[33185] = 32'b11111111111111111110000000110110;
assign LUT_2[33186] = 32'b00000000000000001000000001011001;
assign LUT_2[33187] = 32'b00000000000000000100111001110010;
assign LUT_2[33188] = 32'b11111111111111111101100110000101;
assign LUT_2[33189] = 32'b11111111111111111010011110011110;
assign LUT_2[33190] = 32'b00000000000000000100011111000001;
assign LUT_2[33191] = 32'b00000000000000000001010111011010;
assign LUT_2[33192] = 32'b11111111111111111011111001111010;
assign LUT_2[33193] = 32'b11111111111111111000110010010011;
assign LUT_2[33194] = 32'b00000000000000000010110010110110;
assign LUT_2[33195] = 32'b11111111111111111111101011001111;
assign LUT_2[33196] = 32'b11111111111111111000010111100010;
assign LUT_2[33197] = 32'b11111111111111110101001111111011;
assign LUT_2[33198] = 32'b11111111111111111111010000011110;
assign LUT_2[33199] = 32'b11111111111111111100001000110111;
assign LUT_2[33200] = 32'b11111111111111111011101100100111;
assign LUT_2[33201] = 32'b11111111111111111000100101000000;
assign LUT_2[33202] = 32'b00000000000000000010100101100011;
assign LUT_2[33203] = 32'b11111111111111111111011101111100;
assign LUT_2[33204] = 32'b11111111111111111000001010001111;
assign LUT_2[33205] = 32'b11111111111111110101000010101000;
assign LUT_2[33206] = 32'b11111111111111111111000011001011;
assign LUT_2[33207] = 32'b11111111111111111011111011100100;
assign LUT_2[33208] = 32'b11111111111111110110011110000100;
assign LUT_2[33209] = 32'b11111111111111110011010110011101;
assign LUT_2[33210] = 32'b11111111111111111101010111000000;
assign LUT_2[33211] = 32'b11111111111111111010001111011001;
assign LUT_2[33212] = 32'b11111111111111110010111011101100;
assign LUT_2[33213] = 32'b11111111111111101111110100000101;
assign LUT_2[33214] = 32'b11111111111111111001110100101000;
assign LUT_2[33215] = 32'b11111111111111110110101101000001;
assign LUT_2[33216] = 32'b11111111111111111000110101010111;
assign LUT_2[33217] = 32'b11111111111111110101101101110000;
assign LUT_2[33218] = 32'b11111111111111111111101110010011;
assign LUT_2[33219] = 32'b11111111111111111100100110101100;
assign LUT_2[33220] = 32'b11111111111111110101010010111111;
assign LUT_2[33221] = 32'b11111111111111110010001011011000;
assign LUT_2[33222] = 32'b11111111111111111100001011111011;
assign LUT_2[33223] = 32'b11111111111111111001000100010100;
assign LUT_2[33224] = 32'b11111111111111110011100110110100;
assign LUT_2[33225] = 32'b11111111111111110000011111001101;
assign LUT_2[33226] = 32'b11111111111111111010011111110000;
assign LUT_2[33227] = 32'b11111111111111110111011000001001;
assign LUT_2[33228] = 32'b11111111111111110000000100011100;
assign LUT_2[33229] = 32'b11111111111111101100111100110101;
assign LUT_2[33230] = 32'b11111111111111110110111101011000;
assign LUT_2[33231] = 32'b11111111111111110011110101110001;
assign LUT_2[33232] = 32'b11111111111111110011011001100001;
assign LUT_2[33233] = 32'b11111111111111110000010001111010;
assign LUT_2[33234] = 32'b11111111111111111010010010011101;
assign LUT_2[33235] = 32'b11111111111111110111001010110110;
assign LUT_2[33236] = 32'b11111111111111101111110111001001;
assign LUT_2[33237] = 32'b11111111111111101100101111100010;
assign LUT_2[33238] = 32'b11111111111111110110110000000101;
assign LUT_2[33239] = 32'b11111111111111110011101000011110;
assign LUT_2[33240] = 32'b11111111111111101110001010111110;
assign LUT_2[33241] = 32'b11111111111111101011000011010111;
assign LUT_2[33242] = 32'b11111111111111110101000011111010;
assign LUT_2[33243] = 32'b11111111111111110001111100010011;
assign LUT_2[33244] = 32'b11111111111111101010101000100110;
assign LUT_2[33245] = 32'b11111111111111100111100000111111;
assign LUT_2[33246] = 32'b11111111111111110001100001100010;
assign LUT_2[33247] = 32'b11111111111111101110011001111011;
assign LUT_2[33248] = 32'b11111111111111111001010001000000;
assign LUT_2[33249] = 32'b11111111111111110110001001011001;
assign LUT_2[33250] = 32'b00000000000000000000001001111100;
assign LUT_2[33251] = 32'b11111111111111111101000010010101;
assign LUT_2[33252] = 32'b11111111111111110101101110101000;
assign LUT_2[33253] = 32'b11111111111111110010100111000001;
assign LUT_2[33254] = 32'b11111111111111111100100111100100;
assign LUT_2[33255] = 32'b11111111111111111001011111111101;
assign LUT_2[33256] = 32'b11111111111111110100000010011101;
assign LUT_2[33257] = 32'b11111111111111110000111010110110;
assign LUT_2[33258] = 32'b11111111111111111010111011011001;
assign LUT_2[33259] = 32'b11111111111111110111110011110010;
assign LUT_2[33260] = 32'b11111111111111110000100000000101;
assign LUT_2[33261] = 32'b11111111111111101101011000011110;
assign LUT_2[33262] = 32'b11111111111111110111011001000001;
assign LUT_2[33263] = 32'b11111111111111110100010001011010;
assign LUT_2[33264] = 32'b11111111111111110011110101001010;
assign LUT_2[33265] = 32'b11111111111111110000101101100011;
assign LUT_2[33266] = 32'b11111111111111111010101110000110;
assign LUT_2[33267] = 32'b11111111111111110111100110011111;
assign LUT_2[33268] = 32'b11111111111111110000010010110010;
assign LUT_2[33269] = 32'b11111111111111101101001011001011;
assign LUT_2[33270] = 32'b11111111111111110111001011101110;
assign LUT_2[33271] = 32'b11111111111111110100000100000111;
assign LUT_2[33272] = 32'b11111111111111101110100110100111;
assign LUT_2[33273] = 32'b11111111111111101011011111000000;
assign LUT_2[33274] = 32'b11111111111111110101011111100011;
assign LUT_2[33275] = 32'b11111111111111110010010111111100;
assign LUT_2[33276] = 32'b11111111111111101011000100001111;
assign LUT_2[33277] = 32'b11111111111111100111111100101000;
assign LUT_2[33278] = 32'b11111111111111110001111101001011;
assign LUT_2[33279] = 32'b11111111111111101110110101100100;
assign LUT_2[33280] = 32'b11111111111111111101001011110001;
assign LUT_2[33281] = 32'b11111111111111111010000100001010;
assign LUT_2[33282] = 32'b00000000000000000100000100101101;
assign LUT_2[33283] = 32'b00000000000000000000111101000110;
assign LUT_2[33284] = 32'b11111111111111111001101001011001;
assign LUT_2[33285] = 32'b11111111111111110110100001110010;
assign LUT_2[33286] = 32'b00000000000000000000100010010101;
assign LUT_2[33287] = 32'b11111111111111111101011010101110;
assign LUT_2[33288] = 32'b11111111111111110111111101001110;
assign LUT_2[33289] = 32'b11111111111111110100110101100111;
assign LUT_2[33290] = 32'b11111111111111111110110110001010;
assign LUT_2[33291] = 32'b11111111111111111011101110100011;
assign LUT_2[33292] = 32'b11111111111111110100011010110110;
assign LUT_2[33293] = 32'b11111111111111110001010011001111;
assign LUT_2[33294] = 32'b11111111111111111011010011110010;
assign LUT_2[33295] = 32'b11111111111111111000001100001011;
assign LUT_2[33296] = 32'b11111111111111110111101111111011;
assign LUT_2[33297] = 32'b11111111111111110100101000010100;
assign LUT_2[33298] = 32'b11111111111111111110101000110111;
assign LUT_2[33299] = 32'b11111111111111111011100001010000;
assign LUT_2[33300] = 32'b11111111111111110100001101100011;
assign LUT_2[33301] = 32'b11111111111111110001000101111100;
assign LUT_2[33302] = 32'b11111111111111111011000110011111;
assign LUT_2[33303] = 32'b11111111111111110111111110111000;
assign LUT_2[33304] = 32'b11111111111111110010100001011000;
assign LUT_2[33305] = 32'b11111111111111101111011001110001;
assign LUT_2[33306] = 32'b11111111111111111001011010010100;
assign LUT_2[33307] = 32'b11111111111111110110010010101101;
assign LUT_2[33308] = 32'b11111111111111101110111111000000;
assign LUT_2[33309] = 32'b11111111111111101011110111011001;
assign LUT_2[33310] = 32'b11111111111111110101110111111100;
assign LUT_2[33311] = 32'b11111111111111110010110000010101;
assign LUT_2[33312] = 32'b11111111111111111101100111011010;
assign LUT_2[33313] = 32'b11111111111111111010011111110011;
assign LUT_2[33314] = 32'b00000000000000000100100000010110;
assign LUT_2[33315] = 32'b00000000000000000001011000101111;
assign LUT_2[33316] = 32'b11111111111111111010000101000010;
assign LUT_2[33317] = 32'b11111111111111110110111101011011;
assign LUT_2[33318] = 32'b00000000000000000000111101111110;
assign LUT_2[33319] = 32'b11111111111111111101110110010111;
assign LUT_2[33320] = 32'b11111111111111111000011000110111;
assign LUT_2[33321] = 32'b11111111111111110101010001010000;
assign LUT_2[33322] = 32'b11111111111111111111010001110011;
assign LUT_2[33323] = 32'b11111111111111111100001010001100;
assign LUT_2[33324] = 32'b11111111111111110100110110011111;
assign LUT_2[33325] = 32'b11111111111111110001101110111000;
assign LUT_2[33326] = 32'b11111111111111111011101111011011;
assign LUT_2[33327] = 32'b11111111111111111000100111110100;
assign LUT_2[33328] = 32'b11111111111111111000001011100100;
assign LUT_2[33329] = 32'b11111111111111110101000011111101;
assign LUT_2[33330] = 32'b11111111111111111111000100100000;
assign LUT_2[33331] = 32'b11111111111111111011111100111001;
assign LUT_2[33332] = 32'b11111111111111110100101001001100;
assign LUT_2[33333] = 32'b11111111111111110001100001100101;
assign LUT_2[33334] = 32'b11111111111111111011100010001000;
assign LUT_2[33335] = 32'b11111111111111111000011010100001;
assign LUT_2[33336] = 32'b11111111111111110010111101000001;
assign LUT_2[33337] = 32'b11111111111111101111110101011010;
assign LUT_2[33338] = 32'b11111111111111111001110101111101;
assign LUT_2[33339] = 32'b11111111111111110110101110010110;
assign LUT_2[33340] = 32'b11111111111111101111011010101001;
assign LUT_2[33341] = 32'b11111111111111101100010011000010;
assign LUT_2[33342] = 32'b11111111111111110110010011100101;
assign LUT_2[33343] = 32'b11111111111111110011001011111110;
assign LUT_2[33344] = 32'b11111111111111110101010100010100;
assign LUT_2[33345] = 32'b11111111111111110010001100101101;
assign LUT_2[33346] = 32'b11111111111111111100001101010000;
assign LUT_2[33347] = 32'b11111111111111111001000101101001;
assign LUT_2[33348] = 32'b11111111111111110001110001111100;
assign LUT_2[33349] = 32'b11111111111111101110101010010101;
assign LUT_2[33350] = 32'b11111111111111111000101010111000;
assign LUT_2[33351] = 32'b11111111111111110101100011010001;
assign LUT_2[33352] = 32'b11111111111111110000000101110001;
assign LUT_2[33353] = 32'b11111111111111101100111110001010;
assign LUT_2[33354] = 32'b11111111111111110110111110101101;
assign LUT_2[33355] = 32'b11111111111111110011110111000110;
assign LUT_2[33356] = 32'b11111111111111101100100011011001;
assign LUT_2[33357] = 32'b11111111111111101001011011110010;
assign LUT_2[33358] = 32'b11111111111111110011011100010101;
assign LUT_2[33359] = 32'b11111111111111110000010100101110;
assign LUT_2[33360] = 32'b11111111111111101111111000011110;
assign LUT_2[33361] = 32'b11111111111111101100110000110111;
assign LUT_2[33362] = 32'b11111111111111110110110001011010;
assign LUT_2[33363] = 32'b11111111111111110011101001110011;
assign LUT_2[33364] = 32'b11111111111111101100010110000110;
assign LUT_2[33365] = 32'b11111111111111101001001110011111;
assign LUT_2[33366] = 32'b11111111111111110011001111000010;
assign LUT_2[33367] = 32'b11111111111111110000000111011011;
assign LUT_2[33368] = 32'b11111111111111101010101001111011;
assign LUT_2[33369] = 32'b11111111111111100111100010010100;
assign LUT_2[33370] = 32'b11111111111111110001100010110111;
assign LUT_2[33371] = 32'b11111111111111101110011011010000;
assign LUT_2[33372] = 32'b11111111111111100111000111100011;
assign LUT_2[33373] = 32'b11111111111111100011111111111100;
assign LUT_2[33374] = 32'b11111111111111101110000000011111;
assign LUT_2[33375] = 32'b11111111111111101010111000111000;
assign LUT_2[33376] = 32'b11111111111111110101101111111101;
assign LUT_2[33377] = 32'b11111111111111110010101000010110;
assign LUT_2[33378] = 32'b11111111111111111100101000111001;
assign LUT_2[33379] = 32'b11111111111111111001100001010010;
assign LUT_2[33380] = 32'b11111111111111110010001101100101;
assign LUT_2[33381] = 32'b11111111111111101111000101111110;
assign LUT_2[33382] = 32'b11111111111111111001000110100001;
assign LUT_2[33383] = 32'b11111111111111110101111110111010;
assign LUT_2[33384] = 32'b11111111111111110000100001011010;
assign LUT_2[33385] = 32'b11111111111111101101011001110011;
assign LUT_2[33386] = 32'b11111111111111110111011010010110;
assign LUT_2[33387] = 32'b11111111111111110100010010101111;
assign LUT_2[33388] = 32'b11111111111111101100111111000010;
assign LUT_2[33389] = 32'b11111111111111101001110111011011;
assign LUT_2[33390] = 32'b11111111111111110011110111111110;
assign LUT_2[33391] = 32'b11111111111111110000110000010111;
assign LUT_2[33392] = 32'b11111111111111110000010100000111;
assign LUT_2[33393] = 32'b11111111111111101101001100100000;
assign LUT_2[33394] = 32'b11111111111111110111001101000011;
assign LUT_2[33395] = 32'b11111111111111110100000101011100;
assign LUT_2[33396] = 32'b11111111111111101100110001101111;
assign LUT_2[33397] = 32'b11111111111111101001101010001000;
assign LUT_2[33398] = 32'b11111111111111110011101010101011;
assign LUT_2[33399] = 32'b11111111111111110000100011000100;
assign LUT_2[33400] = 32'b11111111111111101011000101100100;
assign LUT_2[33401] = 32'b11111111111111100111111101111101;
assign LUT_2[33402] = 32'b11111111111111110001111110100000;
assign LUT_2[33403] = 32'b11111111111111101110110110111001;
assign LUT_2[33404] = 32'b11111111111111100111100011001100;
assign LUT_2[33405] = 32'b11111111111111100100011011100101;
assign LUT_2[33406] = 32'b11111111111111101110011100001000;
assign LUT_2[33407] = 32'b11111111111111101011010100100001;
assign LUT_2[33408] = 32'b00000000000000000001100000000000;
assign LUT_2[33409] = 32'b11111111111111111110011000011001;
assign LUT_2[33410] = 32'b00000000000000001000011000111100;
assign LUT_2[33411] = 32'b00000000000000000101010001010101;
assign LUT_2[33412] = 32'b11111111111111111101111101101000;
assign LUT_2[33413] = 32'b11111111111111111010110110000001;
assign LUT_2[33414] = 32'b00000000000000000100110110100100;
assign LUT_2[33415] = 32'b00000000000000000001101110111101;
assign LUT_2[33416] = 32'b11111111111111111100010001011101;
assign LUT_2[33417] = 32'b11111111111111111001001001110110;
assign LUT_2[33418] = 32'b00000000000000000011001010011001;
assign LUT_2[33419] = 32'b00000000000000000000000010110010;
assign LUT_2[33420] = 32'b11111111111111111000101111000101;
assign LUT_2[33421] = 32'b11111111111111110101100111011110;
assign LUT_2[33422] = 32'b11111111111111111111101000000001;
assign LUT_2[33423] = 32'b11111111111111111100100000011010;
assign LUT_2[33424] = 32'b11111111111111111100000100001010;
assign LUT_2[33425] = 32'b11111111111111111000111100100011;
assign LUT_2[33426] = 32'b00000000000000000010111101000110;
assign LUT_2[33427] = 32'b11111111111111111111110101011111;
assign LUT_2[33428] = 32'b11111111111111111000100001110010;
assign LUT_2[33429] = 32'b11111111111111110101011010001011;
assign LUT_2[33430] = 32'b11111111111111111111011010101110;
assign LUT_2[33431] = 32'b11111111111111111100010011000111;
assign LUT_2[33432] = 32'b11111111111111110110110101100111;
assign LUT_2[33433] = 32'b11111111111111110011101110000000;
assign LUT_2[33434] = 32'b11111111111111111101101110100011;
assign LUT_2[33435] = 32'b11111111111111111010100110111100;
assign LUT_2[33436] = 32'b11111111111111110011010011001111;
assign LUT_2[33437] = 32'b11111111111111110000001011101000;
assign LUT_2[33438] = 32'b11111111111111111010001100001011;
assign LUT_2[33439] = 32'b11111111111111110111000100100100;
assign LUT_2[33440] = 32'b00000000000000000001111011101001;
assign LUT_2[33441] = 32'b11111111111111111110110100000010;
assign LUT_2[33442] = 32'b00000000000000001000110100100101;
assign LUT_2[33443] = 32'b00000000000000000101101100111110;
assign LUT_2[33444] = 32'b11111111111111111110011001010001;
assign LUT_2[33445] = 32'b11111111111111111011010001101010;
assign LUT_2[33446] = 32'b00000000000000000101010010001101;
assign LUT_2[33447] = 32'b00000000000000000010001010100110;
assign LUT_2[33448] = 32'b11111111111111111100101101000110;
assign LUT_2[33449] = 32'b11111111111111111001100101011111;
assign LUT_2[33450] = 32'b00000000000000000011100110000010;
assign LUT_2[33451] = 32'b00000000000000000000011110011011;
assign LUT_2[33452] = 32'b11111111111111111001001010101110;
assign LUT_2[33453] = 32'b11111111111111110110000011000111;
assign LUT_2[33454] = 32'b00000000000000000000000011101010;
assign LUT_2[33455] = 32'b11111111111111111100111100000011;
assign LUT_2[33456] = 32'b11111111111111111100011111110011;
assign LUT_2[33457] = 32'b11111111111111111001011000001100;
assign LUT_2[33458] = 32'b00000000000000000011011000101111;
assign LUT_2[33459] = 32'b00000000000000000000010001001000;
assign LUT_2[33460] = 32'b11111111111111111000111101011011;
assign LUT_2[33461] = 32'b11111111111111110101110101110100;
assign LUT_2[33462] = 32'b11111111111111111111110110010111;
assign LUT_2[33463] = 32'b11111111111111111100101110110000;
assign LUT_2[33464] = 32'b11111111111111110111010001010000;
assign LUT_2[33465] = 32'b11111111111111110100001001101001;
assign LUT_2[33466] = 32'b11111111111111111110001010001100;
assign LUT_2[33467] = 32'b11111111111111111011000010100101;
assign LUT_2[33468] = 32'b11111111111111110011101110111000;
assign LUT_2[33469] = 32'b11111111111111110000100111010001;
assign LUT_2[33470] = 32'b11111111111111111010100111110100;
assign LUT_2[33471] = 32'b11111111111111110111100000001101;
assign LUT_2[33472] = 32'b11111111111111111001101000100011;
assign LUT_2[33473] = 32'b11111111111111110110100000111100;
assign LUT_2[33474] = 32'b00000000000000000000100001011111;
assign LUT_2[33475] = 32'b11111111111111111101011001111000;
assign LUT_2[33476] = 32'b11111111111111110110000110001011;
assign LUT_2[33477] = 32'b11111111111111110010111110100100;
assign LUT_2[33478] = 32'b11111111111111111100111111000111;
assign LUT_2[33479] = 32'b11111111111111111001110111100000;
assign LUT_2[33480] = 32'b11111111111111110100011010000000;
assign LUT_2[33481] = 32'b11111111111111110001010010011001;
assign LUT_2[33482] = 32'b11111111111111111011010010111100;
assign LUT_2[33483] = 32'b11111111111111111000001011010101;
assign LUT_2[33484] = 32'b11111111111111110000110111101000;
assign LUT_2[33485] = 32'b11111111111111101101110000000001;
assign LUT_2[33486] = 32'b11111111111111110111110000100100;
assign LUT_2[33487] = 32'b11111111111111110100101000111101;
assign LUT_2[33488] = 32'b11111111111111110100001100101101;
assign LUT_2[33489] = 32'b11111111111111110001000101000110;
assign LUT_2[33490] = 32'b11111111111111111011000101101001;
assign LUT_2[33491] = 32'b11111111111111110111111110000010;
assign LUT_2[33492] = 32'b11111111111111110000101010010101;
assign LUT_2[33493] = 32'b11111111111111101101100010101110;
assign LUT_2[33494] = 32'b11111111111111110111100011010001;
assign LUT_2[33495] = 32'b11111111111111110100011011101010;
assign LUT_2[33496] = 32'b11111111111111101110111110001010;
assign LUT_2[33497] = 32'b11111111111111101011110110100011;
assign LUT_2[33498] = 32'b11111111111111110101110111000110;
assign LUT_2[33499] = 32'b11111111111111110010101111011111;
assign LUT_2[33500] = 32'b11111111111111101011011011110010;
assign LUT_2[33501] = 32'b11111111111111101000010100001011;
assign LUT_2[33502] = 32'b11111111111111110010010100101110;
assign LUT_2[33503] = 32'b11111111111111101111001101000111;
assign LUT_2[33504] = 32'b11111111111111111010000100001100;
assign LUT_2[33505] = 32'b11111111111111110110111100100101;
assign LUT_2[33506] = 32'b00000000000000000000111101001000;
assign LUT_2[33507] = 32'b11111111111111111101110101100001;
assign LUT_2[33508] = 32'b11111111111111110110100001110100;
assign LUT_2[33509] = 32'b11111111111111110011011010001101;
assign LUT_2[33510] = 32'b11111111111111111101011010110000;
assign LUT_2[33511] = 32'b11111111111111111010010011001001;
assign LUT_2[33512] = 32'b11111111111111110100110101101001;
assign LUT_2[33513] = 32'b11111111111111110001101110000010;
assign LUT_2[33514] = 32'b11111111111111111011101110100101;
assign LUT_2[33515] = 32'b11111111111111111000100110111110;
assign LUT_2[33516] = 32'b11111111111111110001010011010001;
assign LUT_2[33517] = 32'b11111111111111101110001011101010;
assign LUT_2[33518] = 32'b11111111111111111000001100001101;
assign LUT_2[33519] = 32'b11111111111111110101000100100110;
assign LUT_2[33520] = 32'b11111111111111110100101000010110;
assign LUT_2[33521] = 32'b11111111111111110001100000101111;
assign LUT_2[33522] = 32'b11111111111111111011100001010010;
assign LUT_2[33523] = 32'b11111111111111111000011001101011;
assign LUT_2[33524] = 32'b11111111111111110001000101111110;
assign LUT_2[33525] = 32'b11111111111111101101111110010111;
assign LUT_2[33526] = 32'b11111111111111110111111110111010;
assign LUT_2[33527] = 32'b11111111111111110100110111010011;
assign LUT_2[33528] = 32'b11111111111111101111011001110011;
assign LUT_2[33529] = 32'b11111111111111101100010010001100;
assign LUT_2[33530] = 32'b11111111111111110110010010101111;
assign LUT_2[33531] = 32'b11111111111111110011001011001000;
assign LUT_2[33532] = 32'b11111111111111101011110111011011;
assign LUT_2[33533] = 32'b11111111111111101000101111110100;
assign LUT_2[33534] = 32'b11111111111111110010110000010111;
assign LUT_2[33535] = 32'b11111111111111101111101000110000;
assign LUT_2[33536] = 32'b00000000000000000001001010010111;
assign LUT_2[33537] = 32'b11111111111111111110000010110000;
assign LUT_2[33538] = 32'b00000000000000001000000011010011;
assign LUT_2[33539] = 32'b00000000000000000100111011101100;
assign LUT_2[33540] = 32'b11111111111111111101100111111111;
assign LUT_2[33541] = 32'b11111111111111111010100000011000;
assign LUT_2[33542] = 32'b00000000000000000100100000111011;
assign LUT_2[33543] = 32'b00000000000000000001011001010100;
assign LUT_2[33544] = 32'b11111111111111111011111011110100;
assign LUT_2[33545] = 32'b11111111111111111000110100001101;
assign LUT_2[33546] = 32'b00000000000000000010110100110000;
assign LUT_2[33547] = 32'b11111111111111111111101101001001;
assign LUT_2[33548] = 32'b11111111111111111000011001011100;
assign LUT_2[33549] = 32'b11111111111111110101010001110101;
assign LUT_2[33550] = 32'b11111111111111111111010010011000;
assign LUT_2[33551] = 32'b11111111111111111100001010110001;
assign LUT_2[33552] = 32'b11111111111111111011101110100001;
assign LUT_2[33553] = 32'b11111111111111111000100110111010;
assign LUT_2[33554] = 32'b00000000000000000010100111011101;
assign LUT_2[33555] = 32'b11111111111111111111011111110110;
assign LUT_2[33556] = 32'b11111111111111111000001100001001;
assign LUT_2[33557] = 32'b11111111111111110101000100100010;
assign LUT_2[33558] = 32'b11111111111111111111000101000101;
assign LUT_2[33559] = 32'b11111111111111111011111101011110;
assign LUT_2[33560] = 32'b11111111111111110110011111111110;
assign LUT_2[33561] = 32'b11111111111111110011011000010111;
assign LUT_2[33562] = 32'b11111111111111111101011000111010;
assign LUT_2[33563] = 32'b11111111111111111010010001010011;
assign LUT_2[33564] = 32'b11111111111111110010111101100110;
assign LUT_2[33565] = 32'b11111111111111101111110101111111;
assign LUT_2[33566] = 32'b11111111111111111001110110100010;
assign LUT_2[33567] = 32'b11111111111111110110101110111011;
assign LUT_2[33568] = 32'b00000000000000000001100110000000;
assign LUT_2[33569] = 32'b11111111111111111110011110011001;
assign LUT_2[33570] = 32'b00000000000000001000011110111100;
assign LUT_2[33571] = 32'b00000000000000000101010111010101;
assign LUT_2[33572] = 32'b11111111111111111110000011101000;
assign LUT_2[33573] = 32'b11111111111111111010111100000001;
assign LUT_2[33574] = 32'b00000000000000000100111100100100;
assign LUT_2[33575] = 32'b00000000000000000001110100111101;
assign LUT_2[33576] = 32'b11111111111111111100010111011101;
assign LUT_2[33577] = 32'b11111111111111111001001111110110;
assign LUT_2[33578] = 32'b00000000000000000011010000011001;
assign LUT_2[33579] = 32'b00000000000000000000001000110010;
assign LUT_2[33580] = 32'b11111111111111111000110101000101;
assign LUT_2[33581] = 32'b11111111111111110101101101011110;
assign LUT_2[33582] = 32'b11111111111111111111101110000001;
assign LUT_2[33583] = 32'b11111111111111111100100110011010;
assign LUT_2[33584] = 32'b11111111111111111100001010001010;
assign LUT_2[33585] = 32'b11111111111111111001000010100011;
assign LUT_2[33586] = 32'b00000000000000000011000011000110;
assign LUT_2[33587] = 32'b11111111111111111111111011011111;
assign LUT_2[33588] = 32'b11111111111111111000100111110010;
assign LUT_2[33589] = 32'b11111111111111110101100000001011;
assign LUT_2[33590] = 32'b11111111111111111111100000101110;
assign LUT_2[33591] = 32'b11111111111111111100011001000111;
assign LUT_2[33592] = 32'b11111111111111110110111011100111;
assign LUT_2[33593] = 32'b11111111111111110011110100000000;
assign LUT_2[33594] = 32'b11111111111111111101110100100011;
assign LUT_2[33595] = 32'b11111111111111111010101100111100;
assign LUT_2[33596] = 32'b11111111111111110011011001001111;
assign LUT_2[33597] = 32'b11111111111111110000010001101000;
assign LUT_2[33598] = 32'b11111111111111111010010010001011;
assign LUT_2[33599] = 32'b11111111111111110111001010100100;
assign LUT_2[33600] = 32'b11111111111111111001010010111010;
assign LUT_2[33601] = 32'b11111111111111110110001011010011;
assign LUT_2[33602] = 32'b00000000000000000000001011110110;
assign LUT_2[33603] = 32'b11111111111111111101000100001111;
assign LUT_2[33604] = 32'b11111111111111110101110000100010;
assign LUT_2[33605] = 32'b11111111111111110010101000111011;
assign LUT_2[33606] = 32'b11111111111111111100101001011110;
assign LUT_2[33607] = 32'b11111111111111111001100001110111;
assign LUT_2[33608] = 32'b11111111111111110100000100010111;
assign LUT_2[33609] = 32'b11111111111111110000111100110000;
assign LUT_2[33610] = 32'b11111111111111111010111101010011;
assign LUT_2[33611] = 32'b11111111111111110111110101101100;
assign LUT_2[33612] = 32'b11111111111111110000100001111111;
assign LUT_2[33613] = 32'b11111111111111101101011010011000;
assign LUT_2[33614] = 32'b11111111111111110111011010111011;
assign LUT_2[33615] = 32'b11111111111111110100010011010100;
assign LUT_2[33616] = 32'b11111111111111110011110111000100;
assign LUT_2[33617] = 32'b11111111111111110000101111011101;
assign LUT_2[33618] = 32'b11111111111111111010110000000000;
assign LUT_2[33619] = 32'b11111111111111110111101000011001;
assign LUT_2[33620] = 32'b11111111111111110000010100101100;
assign LUT_2[33621] = 32'b11111111111111101101001101000101;
assign LUT_2[33622] = 32'b11111111111111110111001101101000;
assign LUT_2[33623] = 32'b11111111111111110100000110000001;
assign LUT_2[33624] = 32'b11111111111111101110101000100001;
assign LUT_2[33625] = 32'b11111111111111101011100000111010;
assign LUT_2[33626] = 32'b11111111111111110101100001011101;
assign LUT_2[33627] = 32'b11111111111111110010011001110110;
assign LUT_2[33628] = 32'b11111111111111101011000110001001;
assign LUT_2[33629] = 32'b11111111111111100111111110100010;
assign LUT_2[33630] = 32'b11111111111111110001111111000101;
assign LUT_2[33631] = 32'b11111111111111101110110111011110;
assign LUT_2[33632] = 32'b11111111111111111001101110100011;
assign LUT_2[33633] = 32'b11111111111111110110100110111100;
assign LUT_2[33634] = 32'b00000000000000000000100111011111;
assign LUT_2[33635] = 32'b11111111111111111101011111111000;
assign LUT_2[33636] = 32'b11111111111111110110001100001011;
assign LUT_2[33637] = 32'b11111111111111110011000100100100;
assign LUT_2[33638] = 32'b11111111111111111101000101000111;
assign LUT_2[33639] = 32'b11111111111111111001111101100000;
assign LUT_2[33640] = 32'b11111111111111110100100000000000;
assign LUT_2[33641] = 32'b11111111111111110001011000011001;
assign LUT_2[33642] = 32'b11111111111111111011011000111100;
assign LUT_2[33643] = 32'b11111111111111111000010001010101;
assign LUT_2[33644] = 32'b11111111111111110000111101101000;
assign LUT_2[33645] = 32'b11111111111111101101110110000001;
assign LUT_2[33646] = 32'b11111111111111110111110110100100;
assign LUT_2[33647] = 32'b11111111111111110100101110111101;
assign LUT_2[33648] = 32'b11111111111111110100010010101101;
assign LUT_2[33649] = 32'b11111111111111110001001011000110;
assign LUT_2[33650] = 32'b11111111111111111011001011101001;
assign LUT_2[33651] = 32'b11111111111111111000000100000010;
assign LUT_2[33652] = 32'b11111111111111110000110000010101;
assign LUT_2[33653] = 32'b11111111111111101101101000101110;
assign LUT_2[33654] = 32'b11111111111111110111101001010001;
assign LUT_2[33655] = 32'b11111111111111110100100001101010;
assign LUT_2[33656] = 32'b11111111111111101111000100001010;
assign LUT_2[33657] = 32'b11111111111111101011111100100011;
assign LUT_2[33658] = 32'b11111111111111110101111101000110;
assign LUT_2[33659] = 32'b11111111111111110010110101011111;
assign LUT_2[33660] = 32'b11111111111111101011100001110010;
assign LUT_2[33661] = 32'b11111111111111101000011010001011;
assign LUT_2[33662] = 32'b11111111111111110010011010101110;
assign LUT_2[33663] = 32'b11111111111111101111010011000111;
assign LUT_2[33664] = 32'b00000000000000000101011110100110;
assign LUT_2[33665] = 32'b00000000000000000010010110111111;
assign LUT_2[33666] = 32'b00000000000000001100010111100010;
assign LUT_2[33667] = 32'b00000000000000001001001111111011;
assign LUT_2[33668] = 32'b00000000000000000001111100001110;
assign LUT_2[33669] = 32'b11111111111111111110110100100111;
assign LUT_2[33670] = 32'b00000000000000001000110101001010;
assign LUT_2[33671] = 32'b00000000000000000101101101100011;
assign LUT_2[33672] = 32'b00000000000000000000010000000011;
assign LUT_2[33673] = 32'b11111111111111111101001000011100;
assign LUT_2[33674] = 32'b00000000000000000111001000111111;
assign LUT_2[33675] = 32'b00000000000000000100000001011000;
assign LUT_2[33676] = 32'b11111111111111111100101101101011;
assign LUT_2[33677] = 32'b11111111111111111001100110000100;
assign LUT_2[33678] = 32'b00000000000000000011100110100111;
assign LUT_2[33679] = 32'b00000000000000000000011111000000;
assign LUT_2[33680] = 32'b00000000000000000000000010110000;
assign LUT_2[33681] = 32'b11111111111111111100111011001001;
assign LUT_2[33682] = 32'b00000000000000000110111011101100;
assign LUT_2[33683] = 32'b00000000000000000011110100000101;
assign LUT_2[33684] = 32'b11111111111111111100100000011000;
assign LUT_2[33685] = 32'b11111111111111111001011000110001;
assign LUT_2[33686] = 32'b00000000000000000011011001010100;
assign LUT_2[33687] = 32'b00000000000000000000010001101101;
assign LUT_2[33688] = 32'b11111111111111111010110100001101;
assign LUT_2[33689] = 32'b11111111111111110111101100100110;
assign LUT_2[33690] = 32'b00000000000000000001101101001001;
assign LUT_2[33691] = 32'b11111111111111111110100101100010;
assign LUT_2[33692] = 32'b11111111111111110111010001110101;
assign LUT_2[33693] = 32'b11111111111111110100001010001110;
assign LUT_2[33694] = 32'b11111111111111111110001010110001;
assign LUT_2[33695] = 32'b11111111111111111011000011001010;
assign LUT_2[33696] = 32'b00000000000000000101111010001111;
assign LUT_2[33697] = 32'b00000000000000000010110010101000;
assign LUT_2[33698] = 32'b00000000000000001100110011001011;
assign LUT_2[33699] = 32'b00000000000000001001101011100100;
assign LUT_2[33700] = 32'b00000000000000000010010111110111;
assign LUT_2[33701] = 32'b11111111111111111111010000010000;
assign LUT_2[33702] = 32'b00000000000000001001010000110011;
assign LUT_2[33703] = 32'b00000000000000000110001001001100;
assign LUT_2[33704] = 32'b00000000000000000000101011101100;
assign LUT_2[33705] = 32'b11111111111111111101100100000101;
assign LUT_2[33706] = 32'b00000000000000000111100100101000;
assign LUT_2[33707] = 32'b00000000000000000100011101000001;
assign LUT_2[33708] = 32'b11111111111111111101001001010100;
assign LUT_2[33709] = 32'b11111111111111111010000001101101;
assign LUT_2[33710] = 32'b00000000000000000100000010010000;
assign LUT_2[33711] = 32'b00000000000000000000111010101001;
assign LUT_2[33712] = 32'b00000000000000000000011110011001;
assign LUT_2[33713] = 32'b11111111111111111101010110110010;
assign LUT_2[33714] = 32'b00000000000000000111010111010101;
assign LUT_2[33715] = 32'b00000000000000000100001111101110;
assign LUT_2[33716] = 32'b11111111111111111100111100000001;
assign LUT_2[33717] = 32'b11111111111111111001110100011010;
assign LUT_2[33718] = 32'b00000000000000000011110100111101;
assign LUT_2[33719] = 32'b00000000000000000000101101010110;
assign LUT_2[33720] = 32'b11111111111111111011001111110110;
assign LUT_2[33721] = 32'b11111111111111111000001000001111;
assign LUT_2[33722] = 32'b00000000000000000010001000110010;
assign LUT_2[33723] = 32'b11111111111111111111000001001011;
assign LUT_2[33724] = 32'b11111111111111110111101101011110;
assign LUT_2[33725] = 32'b11111111111111110100100101110111;
assign LUT_2[33726] = 32'b11111111111111111110100110011010;
assign LUT_2[33727] = 32'b11111111111111111011011110110011;
assign LUT_2[33728] = 32'b11111111111111111101100111001001;
assign LUT_2[33729] = 32'b11111111111111111010011111100010;
assign LUT_2[33730] = 32'b00000000000000000100100000000101;
assign LUT_2[33731] = 32'b00000000000000000001011000011110;
assign LUT_2[33732] = 32'b11111111111111111010000100110001;
assign LUT_2[33733] = 32'b11111111111111110110111101001010;
assign LUT_2[33734] = 32'b00000000000000000000111101101101;
assign LUT_2[33735] = 32'b11111111111111111101110110000110;
assign LUT_2[33736] = 32'b11111111111111111000011000100110;
assign LUT_2[33737] = 32'b11111111111111110101010000111111;
assign LUT_2[33738] = 32'b11111111111111111111010001100010;
assign LUT_2[33739] = 32'b11111111111111111100001001111011;
assign LUT_2[33740] = 32'b11111111111111110100110110001110;
assign LUT_2[33741] = 32'b11111111111111110001101110100111;
assign LUT_2[33742] = 32'b11111111111111111011101111001010;
assign LUT_2[33743] = 32'b11111111111111111000100111100011;
assign LUT_2[33744] = 32'b11111111111111111000001011010011;
assign LUT_2[33745] = 32'b11111111111111110101000011101100;
assign LUT_2[33746] = 32'b11111111111111111111000100001111;
assign LUT_2[33747] = 32'b11111111111111111011111100101000;
assign LUT_2[33748] = 32'b11111111111111110100101000111011;
assign LUT_2[33749] = 32'b11111111111111110001100001010100;
assign LUT_2[33750] = 32'b11111111111111111011100001110111;
assign LUT_2[33751] = 32'b11111111111111111000011010010000;
assign LUT_2[33752] = 32'b11111111111111110010111100110000;
assign LUT_2[33753] = 32'b11111111111111101111110101001001;
assign LUT_2[33754] = 32'b11111111111111111001110101101100;
assign LUT_2[33755] = 32'b11111111111111110110101110000101;
assign LUT_2[33756] = 32'b11111111111111101111011010011000;
assign LUT_2[33757] = 32'b11111111111111101100010010110001;
assign LUT_2[33758] = 32'b11111111111111110110010011010100;
assign LUT_2[33759] = 32'b11111111111111110011001011101101;
assign LUT_2[33760] = 32'b11111111111111111110000010110010;
assign LUT_2[33761] = 32'b11111111111111111010111011001011;
assign LUT_2[33762] = 32'b00000000000000000100111011101110;
assign LUT_2[33763] = 32'b00000000000000000001110100000111;
assign LUT_2[33764] = 32'b11111111111111111010100000011010;
assign LUT_2[33765] = 32'b11111111111111110111011000110011;
assign LUT_2[33766] = 32'b00000000000000000001011001010110;
assign LUT_2[33767] = 32'b11111111111111111110010001101111;
assign LUT_2[33768] = 32'b11111111111111111000110100001111;
assign LUT_2[33769] = 32'b11111111111111110101101100101000;
assign LUT_2[33770] = 32'b11111111111111111111101101001011;
assign LUT_2[33771] = 32'b11111111111111111100100101100100;
assign LUT_2[33772] = 32'b11111111111111110101010001110111;
assign LUT_2[33773] = 32'b11111111111111110010001010010000;
assign LUT_2[33774] = 32'b11111111111111111100001010110011;
assign LUT_2[33775] = 32'b11111111111111111001000011001100;
assign LUT_2[33776] = 32'b11111111111111111000100110111100;
assign LUT_2[33777] = 32'b11111111111111110101011111010101;
assign LUT_2[33778] = 32'b11111111111111111111011111111000;
assign LUT_2[33779] = 32'b11111111111111111100011000010001;
assign LUT_2[33780] = 32'b11111111111111110101000100100100;
assign LUT_2[33781] = 32'b11111111111111110001111100111101;
assign LUT_2[33782] = 32'b11111111111111111011111101100000;
assign LUT_2[33783] = 32'b11111111111111111000110101111001;
assign LUT_2[33784] = 32'b11111111111111110011011000011001;
assign LUT_2[33785] = 32'b11111111111111110000010000110010;
assign LUT_2[33786] = 32'b11111111111111111010010001010101;
assign LUT_2[33787] = 32'b11111111111111110111001001101110;
assign LUT_2[33788] = 32'b11111111111111101111110110000001;
assign LUT_2[33789] = 32'b11111111111111101100101110011010;
assign LUT_2[33790] = 32'b11111111111111110110101110111101;
assign LUT_2[33791] = 32'b11111111111111110011100111010110;
assign LUT_2[33792] = 32'b11111111111111111111000110000100;
assign LUT_2[33793] = 32'b11111111111111111011111110011101;
assign LUT_2[33794] = 32'b00000000000000000101111111000000;
assign LUT_2[33795] = 32'b00000000000000000010110111011001;
assign LUT_2[33796] = 32'b11111111111111111011100011101100;
assign LUT_2[33797] = 32'b11111111111111111000011100000101;
assign LUT_2[33798] = 32'b00000000000000000010011100101000;
assign LUT_2[33799] = 32'b11111111111111111111010101000001;
assign LUT_2[33800] = 32'b11111111111111111001110111100001;
assign LUT_2[33801] = 32'b11111111111111110110101111111010;
assign LUT_2[33802] = 32'b00000000000000000000110000011101;
assign LUT_2[33803] = 32'b11111111111111111101101000110110;
assign LUT_2[33804] = 32'b11111111111111110110010101001001;
assign LUT_2[33805] = 32'b11111111111111110011001101100010;
assign LUT_2[33806] = 32'b11111111111111111101001110000101;
assign LUT_2[33807] = 32'b11111111111111111010000110011110;
assign LUT_2[33808] = 32'b11111111111111111001101010001110;
assign LUT_2[33809] = 32'b11111111111111110110100010100111;
assign LUT_2[33810] = 32'b00000000000000000000100011001010;
assign LUT_2[33811] = 32'b11111111111111111101011011100011;
assign LUT_2[33812] = 32'b11111111111111110110000111110110;
assign LUT_2[33813] = 32'b11111111111111110011000000001111;
assign LUT_2[33814] = 32'b11111111111111111101000000110010;
assign LUT_2[33815] = 32'b11111111111111111001111001001011;
assign LUT_2[33816] = 32'b11111111111111110100011011101011;
assign LUT_2[33817] = 32'b11111111111111110001010100000100;
assign LUT_2[33818] = 32'b11111111111111111011010100100111;
assign LUT_2[33819] = 32'b11111111111111111000001101000000;
assign LUT_2[33820] = 32'b11111111111111110000111001010011;
assign LUT_2[33821] = 32'b11111111111111101101110001101100;
assign LUT_2[33822] = 32'b11111111111111110111110010001111;
assign LUT_2[33823] = 32'b11111111111111110100101010101000;
assign LUT_2[33824] = 32'b11111111111111111111100001101101;
assign LUT_2[33825] = 32'b11111111111111111100011010000110;
assign LUT_2[33826] = 32'b00000000000000000110011010101001;
assign LUT_2[33827] = 32'b00000000000000000011010011000010;
assign LUT_2[33828] = 32'b11111111111111111011111111010101;
assign LUT_2[33829] = 32'b11111111111111111000110111101110;
assign LUT_2[33830] = 32'b00000000000000000010111000010001;
assign LUT_2[33831] = 32'b11111111111111111111110000101010;
assign LUT_2[33832] = 32'b11111111111111111010010011001010;
assign LUT_2[33833] = 32'b11111111111111110111001011100011;
assign LUT_2[33834] = 32'b00000000000000000001001100000110;
assign LUT_2[33835] = 32'b11111111111111111110000100011111;
assign LUT_2[33836] = 32'b11111111111111110110110000110010;
assign LUT_2[33837] = 32'b11111111111111110011101001001011;
assign LUT_2[33838] = 32'b11111111111111111101101001101110;
assign LUT_2[33839] = 32'b11111111111111111010100010000111;
assign LUT_2[33840] = 32'b11111111111111111010000101110111;
assign LUT_2[33841] = 32'b11111111111111110110111110010000;
assign LUT_2[33842] = 32'b00000000000000000000111110110011;
assign LUT_2[33843] = 32'b11111111111111111101110111001100;
assign LUT_2[33844] = 32'b11111111111111110110100011011111;
assign LUT_2[33845] = 32'b11111111111111110011011011111000;
assign LUT_2[33846] = 32'b11111111111111111101011100011011;
assign LUT_2[33847] = 32'b11111111111111111010010100110100;
assign LUT_2[33848] = 32'b11111111111111110100110111010100;
assign LUT_2[33849] = 32'b11111111111111110001101111101101;
assign LUT_2[33850] = 32'b11111111111111111011110000010000;
assign LUT_2[33851] = 32'b11111111111111111000101000101001;
assign LUT_2[33852] = 32'b11111111111111110001010100111100;
assign LUT_2[33853] = 32'b11111111111111101110001101010101;
assign LUT_2[33854] = 32'b11111111111111111000001101111000;
assign LUT_2[33855] = 32'b11111111111111110101000110010001;
assign LUT_2[33856] = 32'b11111111111111110111001110100111;
assign LUT_2[33857] = 32'b11111111111111110100000111000000;
assign LUT_2[33858] = 32'b11111111111111111110000111100011;
assign LUT_2[33859] = 32'b11111111111111111010111111111100;
assign LUT_2[33860] = 32'b11111111111111110011101100001111;
assign LUT_2[33861] = 32'b11111111111111110000100100101000;
assign LUT_2[33862] = 32'b11111111111111111010100101001011;
assign LUT_2[33863] = 32'b11111111111111110111011101100100;
assign LUT_2[33864] = 32'b11111111111111110010000000000100;
assign LUT_2[33865] = 32'b11111111111111101110111000011101;
assign LUT_2[33866] = 32'b11111111111111111000111001000000;
assign LUT_2[33867] = 32'b11111111111111110101110001011001;
assign LUT_2[33868] = 32'b11111111111111101110011101101100;
assign LUT_2[33869] = 32'b11111111111111101011010110000101;
assign LUT_2[33870] = 32'b11111111111111110101010110101000;
assign LUT_2[33871] = 32'b11111111111111110010001111000001;
assign LUT_2[33872] = 32'b11111111111111110001110010110001;
assign LUT_2[33873] = 32'b11111111111111101110101011001010;
assign LUT_2[33874] = 32'b11111111111111111000101011101101;
assign LUT_2[33875] = 32'b11111111111111110101100100000110;
assign LUT_2[33876] = 32'b11111111111111101110010000011001;
assign LUT_2[33877] = 32'b11111111111111101011001000110010;
assign LUT_2[33878] = 32'b11111111111111110101001001010101;
assign LUT_2[33879] = 32'b11111111111111110010000001101110;
assign LUT_2[33880] = 32'b11111111111111101100100100001110;
assign LUT_2[33881] = 32'b11111111111111101001011100100111;
assign LUT_2[33882] = 32'b11111111111111110011011101001010;
assign LUT_2[33883] = 32'b11111111111111110000010101100011;
assign LUT_2[33884] = 32'b11111111111111101001000001110110;
assign LUT_2[33885] = 32'b11111111111111100101111010001111;
assign LUT_2[33886] = 32'b11111111111111101111111010110010;
assign LUT_2[33887] = 32'b11111111111111101100110011001011;
assign LUT_2[33888] = 32'b11111111111111110111101010010000;
assign LUT_2[33889] = 32'b11111111111111110100100010101001;
assign LUT_2[33890] = 32'b11111111111111111110100011001100;
assign LUT_2[33891] = 32'b11111111111111111011011011100101;
assign LUT_2[33892] = 32'b11111111111111110100000111111000;
assign LUT_2[33893] = 32'b11111111111111110001000000010001;
assign LUT_2[33894] = 32'b11111111111111111011000000110100;
assign LUT_2[33895] = 32'b11111111111111110111111001001101;
assign LUT_2[33896] = 32'b11111111111111110010011011101101;
assign LUT_2[33897] = 32'b11111111111111101111010100000110;
assign LUT_2[33898] = 32'b11111111111111111001010100101001;
assign LUT_2[33899] = 32'b11111111111111110110001101000010;
assign LUT_2[33900] = 32'b11111111111111101110111001010101;
assign LUT_2[33901] = 32'b11111111111111101011110001101110;
assign LUT_2[33902] = 32'b11111111111111110101110010010001;
assign LUT_2[33903] = 32'b11111111111111110010101010101010;
assign LUT_2[33904] = 32'b11111111111111110010001110011010;
assign LUT_2[33905] = 32'b11111111111111101111000110110011;
assign LUT_2[33906] = 32'b11111111111111111001000111010110;
assign LUT_2[33907] = 32'b11111111111111110101111111101111;
assign LUT_2[33908] = 32'b11111111111111101110101100000010;
assign LUT_2[33909] = 32'b11111111111111101011100100011011;
assign LUT_2[33910] = 32'b11111111111111110101100100111110;
assign LUT_2[33911] = 32'b11111111111111110010011101010111;
assign LUT_2[33912] = 32'b11111111111111101100111111110111;
assign LUT_2[33913] = 32'b11111111111111101001111000010000;
assign LUT_2[33914] = 32'b11111111111111110011111000110011;
assign LUT_2[33915] = 32'b11111111111111110000110001001100;
assign LUT_2[33916] = 32'b11111111111111101001011101011111;
assign LUT_2[33917] = 32'b11111111111111100110010101111000;
assign LUT_2[33918] = 32'b11111111111111110000010110011011;
assign LUT_2[33919] = 32'b11111111111111101101001110110100;
assign LUT_2[33920] = 32'b00000000000000000011011010010011;
assign LUT_2[33921] = 32'b00000000000000000000010010101100;
assign LUT_2[33922] = 32'b00000000000000001010010011001111;
assign LUT_2[33923] = 32'b00000000000000000111001011101000;
assign LUT_2[33924] = 32'b11111111111111111111110111111011;
assign LUT_2[33925] = 32'b11111111111111111100110000010100;
assign LUT_2[33926] = 32'b00000000000000000110110000110111;
assign LUT_2[33927] = 32'b00000000000000000011101001010000;
assign LUT_2[33928] = 32'b11111111111111111110001011110000;
assign LUT_2[33929] = 32'b11111111111111111011000100001001;
assign LUT_2[33930] = 32'b00000000000000000101000100101100;
assign LUT_2[33931] = 32'b00000000000000000001111101000101;
assign LUT_2[33932] = 32'b11111111111111111010101001011000;
assign LUT_2[33933] = 32'b11111111111111110111100001110001;
assign LUT_2[33934] = 32'b00000000000000000001100010010100;
assign LUT_2[33935] = 32'b11111111111111111110011010101101;
assign LUT_2[33936] = 32'b11111111111111111101111110011101;
assign LUT_2[33937] = 32'b11111111111111111010110110110110;
assign LUT_2[33938] = 32'b00000000000000000100110111011001;
assign LUT_2[33939] = 32'b00000000000000000001101111110010;
assign LUT_2[33940] = 32'b11111111111111111010011100000101;
assign LUT_2[33941] = 32'b11111111111111110111010100011110;
assign LUT_2[33942] = 32'b00000000000000000001010101000001;
assign LUT_2[33943] = 32'b11111111111111111110001101011010;
assign LUT_2[33944] = 32'b11111111111111111000101111111010;
assign LUT_2[33945] = 32'b11111111111111110101101000010011;
assign LUT_2[33946] = 32'b11111111111111111111101000110110;
assign LUT_2[33947] = 32'b11111111111111111100100001001111;
assign LUT_2[33948] = 32'b11111111111111110101001101100010;
assign LUT_2[33949] = 32'b11111111111111110010000101111011;
assign LUT_2[33950] = 32'b11111111111111111100000110011110;
assign LUT_2[33951] = 32'b11111111111111111000111110110111;
assign LUT_2[33952] = 32'b00000000000000000011110101111100;
assign LUT_2[33953] = 32'b00000000000000000000101110010101;
assign LUT_2[33954] = 32'b00000000000000001010101110111000;
assign LUT_2[33955] = 32'b00000000000000000111100111010001;
assign LUT_2[33956] = 32'b00000000000000000000010011100100;
assign LUT_2[33957] = 32'b11111111111111111101001011111101;
assign LUT_2[33958] = 32'b00000000000000000111001100100000;
assign LUT_2[33959] = 32'b00000000000000000100000100111001;
assign LUT_2[33960] = 32'b11111111111111111110100111011001;
assign LUT_2[33961] = 32'b11111111111111111011011111110010;
assign LUT_2[33962] = 32'b00000000000000000101100000010101;
assign LUT_2[33963] = 32'b00000000000000000010011000101110;
assign LUT_2[33964] = 32'b11111111111111111011000101000001;
assign LUT_2[33965] = 32'b11111111111111110111111101011010;
assign LUT_2[33966] = 32'b00000000000000000001111101111101;
assign LUT_2[33967] = 32'b11111111111111111110110110010110;
assign LUT_2[33968] = 32'b11111111111111111110011010000110;
assign LUT_2[33969] = 32'b11111111111111111011010010011111;
assign LUT_2[33970] = 32'b00000000000000000101010011000010;
assign LUT_2[33971] = 32'b00000000000000000010001011011011;
assign LUT_2[33972] = 32'b11111111111111111010110111101110;
assign LUT_2[33973] = 32'b11111111111111110111110000000111;
assign LUT_2[33974] = 32'b00000000000000000001110000101010;
assign LUT_2[33975] = 32'b11111111111111111110101001000011;
assign LUT_2[33976] = 32'b11111111111111111001001011100011;
assign LUT_2[33977] = 32'b11111111111111110110000011111100;
assign LUT_2[33978] = 32'b00000000000000000000000100011111;
assign LUT_2[33979] = 32'b11111111111111111100111100111000;
assign LUT_2[33980] = 32'b11111111111111110101101001001011;
assign LUT_2[33981] = 32'b11111111111111110010100001100100;
assign LUT_2[33982] = 32'b11111111111111111100100010000111;
assign LUT_2[33983] = 32'b11111111111111111001011010100000;
assign LUT_2[33984] = 32'b11111111111111111011100010110110;
assign LUT_2[33985] = 32'b11111111111111111000011011001111;
assign LUT_2[33986] = 32'b00000000000000000010011011110010;
assign LUT_2[33987] = 32'b11111111111111111111010100001011;
assign LUT_2[33988] = 32'b11111111111111111000000000011110;
assign LUT_2[33989] = 32'b11111111111111110100111000110111;
assign LUT_2[33990] = 32'b11111111111111111110111001011010;
assign LUT_2[33991] = 32'b11111111111111111011110001110011;
assign LUT_2[33992] = 32'b11111111111111110110010100010011;
assign LUT_2[33993] = 32'b11111111111111110011001100101100;
assign LUT_2[33994] = 32'b11111111111111111101001101001111;
assign LUT_2[33995] = 32'b11111111111111111010000101101000;
assign LUT_2[33996] = 32'b11111111111111110010110001111011;
assign LUT_2[33997] = 32'b11111111111111101111101010010100;
assign LUT_2[33998] = 32'b11111111111111111001101010110111;
assign LUT_2[33999] = 32'b11111111111111110110100011010000;
assign LUT_2[34000] = 32'b11111111111111110110000111000000;
assign LUT_2[34001] = 32'b11111111111111110010111111011001;
assign LUT_2[34002] = 32'b11111111111111111100111111111100;
assign LUT_2[34003] = 32'b11111111111111111001111000010101;
assign LUT_2[34004] = 32'b11111111111111110010100100101000;
assign LUT_2[34005] = 32'b11111111111111101111011101000001;
assign LUT_2[34006] = 32'b11111111111111111001011101100100;
assign LUT_2[34007] = 32'b11111111111111110110010101111101;
assign LUT_2[34008] = 32'b11111111111111110000111000011101;
assign LUT_2[34009] = 32'b11111111111111101101110000110110;
assign LUT_2[34010] = 32'b11111111111111110111110001011001;
assign LUT_2[34011] = 32'b11111111111111110100101001110010;
assign LUT_2[34012] = 32'b11111111111111101101010110000101;
assign LUT_2[34013] = 32'b11111111111111101010001110011110;
assign LUT_2[34014] = 32'b11111111111111110100001111000001;
assign LUT_2[34015] = 32'b11111111111111110001000111011010;
assign LUT_2[34016] = 32'b11111111111111111011111110011111;
assign LUT_2[34017] = 32'b11111111111111111000110110111000;
assign LUT_2[34018] = 32'b00000000000000000010110111011011;
assign LUT_2[34019] = 32'b11111111111111111111101111110100;
assign LUT_2[34020] = 32'b11111111111111111000011100000111;
assign LUT_2[34021] = 32'b11111111111111110101010100100000;
assign LUT_2[34022] = 32'b11111111111111111111010101000011;
assign LUT_2[34023] = 32'b11111111111111111100001101011100;
assign LUT_2[34024] = 32'b11111111111111110110101111111100;
assign LUT_2[34025] = 32'b11111111111111110011101000010101;
assign LUT_2[34026] = 32'b11111111111111111101101000111000;
assign LUT_2[34027] = 32'b11111111111111111010100001010001;
assign LUT_2[34028] = 32'b11111111111111110011001101100100;
assign LUT_2[34029] = 32'b11111111111111110000000101111101;
assign LUT_2[34030] = 32'b11111111111111111010000110100000;
assign LUT_2[34031] = 32'b11111111111111110110111110111001;
assign LUT_2[34032] = 32'b11111111111111110110100010101001;
assign LUT_2[34033] = 32'b11111111111111110011011011000010;
assign LUT_2[34034] = 32'b11111111111111111101011011100101;
assign LUT_2[34035] = 32'b11111111111111111010010011111110;
assign LUT_2[34036] = 32'b11111111111111110011000000010001;
assign LUT_2[34037] = 32'b11111111111111101111111000101010;
assign LUT_2[34038] = 32'b11111111111111111001111001001101;
assign LUT_2[34039] = 32'b11111111111111110110110001100110;
assign LUT_2[34040] = 32'b11111111111111110001010100000110;
assign LUT_2[34041] = 32'b11111111111111101110001100011111;
assign LUT_2[34042] = 32'b11111111111111111000001101000010;
assign LUT_2[34043] = 32'b11111111111111110101000101011011;
assign LUT_2[34044] = 32'b11111111111111101101110001101110;
assign LUT_2[34045] = 32'b11111111111111101010101010000111;
assign LUT_2[34046] = 32'b11111111111111110100101010101010;
assign LUT_2[34047] = 32'b11111111111111110001100011000011;
assign LUT_2[34048] = 32'b00000000000000000011000100101010;
assign LUT_2[34049] = 32'b11111111111111111111111101000011;
assign LUT_2[34050] = 32'b00000000000000001001111101100110;
assign LUT_2[34051] = 32'b00000000000000000110110101111111;
assign LUT_2[34052] = 32'b11111111111111111111100010010010;
assign LUT_2[34053] = 32'b11111111111111111100011010101011;
assign LUT_2[34054] = 32'b00000000000000000110011011001110;
assign LUT_2[34055] = 32'b00000000000000000011010011100111;
assign LUT_2[34056] = 32'b11111111111111111101110110000111;
assign LUT_2[34057] = 32'b11111111111111111010101110100000;
assign LUT_2[34058] = 32'b00000000000000000100101111000011;
assign LUT_2[34059] = 32'b00000000000000000001100111011100;
assign LUT_2[34060] = 32'b11111111111111111010010011101111;
assign LUT_2[34061] = 32'b11111111111111110111001100001000;
assign LUT_2[34062] = 32'b00000000000000000001001100101011;
assign LUT_2[34063] = 32'b11111111111111111110000101000100;
assign LUT_2[34064] = 32'b11111111111111111101101000110100;
assign LUT_2[34065] = 32'b11111111111111111010100001001101;
assign LUT_2[34066] = 32'b00000000000000000100100001110000;
assign LUT_2[34067] = 32'b00000000000000000001011010001001;
assign LUT_2[34068] = 32'b11111111111111111010000110011100;
assign LUT_2[34069] = 32'b11111111111111110110111110110101;
assign LUT_2[34070] = 32'b00000000000000000000111111011000;
assign LUT_2[34071] = 32'b11111111111111111101110111110001;
assign LUT_2[34072] = 32'b11111111111111111000011010010001;
assign LUT_2[34073] = 32'b11111111111111110101010010101010;
assign LUT_2[34074] = 32'b11111111111111111111010011001101;
assign LUT_2[34075] = 32'b11111111111111111100001011100110;
assign LUT_2[34076] = 32'b11111111111111110100110111111001;
assign LUT_2[34077] = 32'b11111111111111110001110000010010;
assign LUT_2[34078] = 32'b11111111111111111011110000110101;
assign LUT_2[34079] = 32'b11111111111111111000101001001110;
assign LUT_2[34080] = 32'b00000000000000000011100000010011;
assign LUT_2[34081] = 32'b00000000000000000000011000101100;
assign LUT_2[34082] = 32'b00000000000000001010011001001111;
assign LUT_2[34083] = 32'b00000000000000000111010001101000;
assign LUT_2[34084] = 32'b11111111111111111111111101111011;
assign LUT_2[34085] = 32'b11111111111111111100110110010100;
assign LUT_2[34086] = 32'b00000000000000000110110110110111;
assign LUT_2[34087] = 32'b00000000000000000011101111010000;
assign LUT_2[34088] = 32'b11111111111111111110010001110000;
assign LUT_2[34089] = 32'b11111111111111111011001010001001;
assign LUT_2[34090] = 32'b00000000000000000101001010101100;
assign LUT_2[34091] = 32'b00000000000000000010000011000101;
assign LUT_2[34092] = 32'b11111111111111111010101111011000;
assign LUT_2[34093] = 32'b11111111111111110111100111110001;
assign LUT_2[34094] = 32'b00000000000000000001101000010100;
assign LUT_2[34095] = 32'b11111111111111111110100000101101;
assign LUT_2[34096] = 32'b11111111111111111110000100011101;
assign LUT_2[34097] = 32'b11111111111111111010111100110110;
assign LUT_2[34098] = 32'b00000000000000000100111101011001;
assign LUT_2[34099] = 32'b00000000000000000001110101110010;
assign LUT_2[34100] = 32'b11111111111111111010100010000101;
assign LUT_2[34101] = 32'b11111111111111110111011010011110;
assign LUT_2[34102] = 32'b00000000000000000001011011000001;
assign LUT_2[34103] = 32'b11111111111111111110010011011010;
assign LUT_2[34104] = 32'b11111111111111111000110101111010;
assign LUT_2[34105] = 32'b11111111111111110101101110010011;
assign LUT_2[34106] = 32'b11111111111111111111101110110110;
assign LUT_2[34107] = 32'b11111111111111111100100111001111;
assign LUT_2[34108] = 32'b11111111111111110101010011100010;
assign LUT_2[34109] = 32'b11111111111111110010001011111011;
assign LUT_2[34110] = 32'b11111111111111111100001100011110;
assign LUT_2[34111] = 32'b11111111111111111001000100110111;
assign LUT_2[34112] = 32'b11111111111111111011001101001101;
assign LUT_2[34113] = 32'b11111111111111111000000101100110;
assign LUT_2[34114] = 32'b00000000000000000010000110001001;
assign LUT_2[34115] = 32'b11111111111111111110111110100010;
assign LUT_2[34116] = 32'b11111111111111110111101010110101;
assign LUT_2[34117] = 32'b11111111111111110100100011001110;
assign LUT_2[34118] = 32'b11111111111111111110100011110001;
assign LUT_2[34119] = 32'b11111111111111111011011100001010;
assign LUT_2[34120] = 32'b11111111111111110101111110101010;
assign LUT_2[34121] = 32'b11111111111111110010110111000011;
assign LUT_2[34122] = 32'b11111111111111111100110111100110;
assign LUT_2[34123] = 32'b11111111111111111001101111111111;
assign LUT_2[34124] = 32'b11111111111111110010011100010010;
assign LUT_2[34125] = 32'b11111111111111101111010100101011;
assign LUT_2[34126] = 32'b11111111111111111001010101001110;
assign LUT_2[34127] = 32'b11111111111111110110001101100111;
assign LUT_2[34128] = 32'b11111111111111110101110001010111;
assign LUT_2[34129] = 32'b11111111111111110010101001110000;
assign LUT_2[34130] = 32'b11111111111111111100101010010011;
assign LUT_2[34131] = 32'b11111111111111111001100010101100;
assign LUT_2[34132] = 32'b11111111111111110010001110111111;
assign LUT_2[34133] = 32'b11111111111111101111000111011000;
assign LUT_2[34134] = 32'b11111111111111111001000111111011;
assign LUT_2[34135] = 32'b11111111111111110110000000010100;
assign LUT_2[34136] = 32'b11111111111111110000100010110100;
assign LUT_2[34137] = 32'b11111111111111101101011011001101;
assign LUT_2[34138] = 32'b11111111111111110111011011110000;
assign LUT_2[34139] = 32'b11111111111111110100010100001001;
assign LUT_2[34140] = 32'b11111111111111101101000000011100;
assign LUT_2[34141] = 32'b11111111111111101001111000110101;
assign LUT_2[34142] = 32'b11111111111111110011111001011000;
assign LUT_2[34143] = 32'b11111111111111110000110001110001;
assign LUT_2[34144] = 32'b11111111111111111011101000110110;
assign LUT_2[34145] = 32'b11111111111111111000100001001111;
assign LUT_2[34146] = 32'b00000000000000000010100001110010;
assign LUT_2[34147] = 32'b11111111111111111111011010001011;
assign LUT_2[34148] = 32'b11111111111111111000000110011110;
assign LUT_2[34149] = 32'b11111111111111110100111110110111;
assign LUT_2[34150] = 32'b11111111111111111110111111011010;
assign LUT_2[34151] = 32'b11111111111111111011110111110011;
assign LUT_2[34152] = 32'b11111111111111110110011010010011;
assign LUT_2[34153] = 32'b11111111111111110011010010101100;
assign LUT_2[34154] = 32'b11111111111111111101010011001111;
assign LUT_2[34155] = 32'b11111111111111111010001011101000;
assign LUT_2[34156] = 32'b11111111111111110010110111111011;
assign LUT_2[34157] = 32'b11111111111111101111110000010100;
assign LUT_2[34158] = 32'b11111111111111111001110000110111;
assign LUT_2[34159] = 32'b11111111111111110110101001010000;
assign LUT_2[34160] = 32'b11111111111111110110001101000000;
assign LUT_2[34161] = 32'b11111111111111110011000101011001;
assign LUT_2[34162] = 32'b11111111111111111101000101111100;
assign LUT_2[34163] = 32'b11111111111111111001111110010101;
assign LUT_2[34164] = 32'b11111111111111110010101010101000;
assign LUT_2[34165] = 32'b11111111111111101111100011000001;
assign LUT_2[34166] = 32'b11111111111111111001100011100100;
assign LUT_2[34167] = 32'b11111111111111110110011011111101;
assign LUT_2[34168] = 32'b11111111111111110000111110011101;
assign LUT_2[34169] = 32'b11111111111111101101110110110110;
assign LUT_2[34170] = 32'b11111111111111110111110111011001;
assign LUT_2[34171] = 32'b11111111111111110100101111110010;
assign LUT_2[34172] = 32'b11111111111111101101011100000101;
assign LUT_2[34173] = 32'b11111111111111101010010100011110;
assign LUT_2[34174] = 32'b11111111111111110100010101000001;
assign LUT_2[34175] = 32'b11111111111111110001001101011010;
assign LUT_2[34176] = 32'b00000000000000000111011000111001;
assign LUT_2[34177] = 32'b00000000000000000100010001010010;
assign LUT_2[34178] = 32'b00000000000000001110010001110101;
assign LUT_2[34179] = 32'b00000000000000001011001010001110;
assign LUT_2[34180] = 32'b00000000000000000011110110100001;
assign LUT_2[34181] = 32'b00000000000000000000101110111010;
assign LUT_2[34182] = 32'b00000000000000001010101111011101;
assign LUT_2[34183] = 32'b00000000000000000111100111110110;
assign LUT_2[34184] = 32'b00000000000000000010001010010110;
assign LUT_2[34185] = 32'b11111111111111111111000010101111;
assign LUT_2[34186] = 32'b00000000000000001001000011010010;
assign LUT_2[34187] = 32'b00000000000000000101111011101011;
assign LUT_2[34188] = 32'b11111111111111111110100111111110;
assign LUT_2[34189] = 32'b11111111111111111011100000010111;
assign LUT_2[34190] = 32'b00000000000000000101100000111010;
assign LUT_2[34191] = 32'b00000000000000000010011001010011;
assign LUT_2[34192] = 32'b00000000000000000001111101000011;
assign LUT_2[34193] = 32'b11111111111111111110110101011100;
assign LUT_2[34194] = 32'b00000000000000001000110101111111;
assign LUT_2[34195] = 32'b00000000000000000101101110011000;
assign LUT_2[34196] = 32'b11111111111111111110011010101011;
assign LUT_2[34197] = 32'b11111111111111111011010011000100;
assign LUT_2[34198] = 32'b00000000000000000101010011100111;
assign LUT_2[34199] = 32'b00000000000000000010001100000000;
assign LUT_2[34200] = 32'b11111111111111111100101110100000;
assign LUT_2[34201] = 32'b11111111111111111001100110111001;
assign LUT_2[34202] = 32'b00000000000000000011100111011100;
assign LUT_2[34203] = 32'b00000000000000000000011111110101;
assign LUT_2[34204] = 32'b11111111111111111001001100001000;
assign LUT_2[34205] = 32'b11111111111111110110000100100001;
assign LUT_2[34206] = 32'b00000000000000000000000101000100;
assign LUT_2[34207] = 32'b11111111111111111100111101011101;
assign LUT_2[34208] = 32'b00000000000000000111110100100010;
assign LUT_2[34209] = 32'b00000000000000000100101100111011;
assign LUT_2[34210] = 32'b00000000000000001110101101011110;
assign LUT_2[34211] = 32'b00000000000000001011100101110111;
assign LUT_2[34212] = 32'b00000000000000000100010010001010;
assign LUT_2[34213] = 32'b00000000000000000001001010100011;
assign LUT_2[34214] = 32'b00000000000000001011001011000110;
assign LUT_2[34215] = 32'b00000000000000001000000011011111;
assign LUT_2[34216] = 32'b00000000000000000010100101111111;
assign LUT_2[34217] = 32'b11111111111111111111011110011000;
assign LUT_2[34218] = 32'b00000000000000001001011110111011;
assign LUT_2[34219] = 32'b00000000000000000110010111010100;
assign LUT_2[34220] = 32'b11111111111111111111000011100111;
assign LUT_2[34221] = 32'b11111111111111111011111100000000;
assign LUT_2[34222] = 32'b00000000000000000101111100100011;
assign LUT_2[34223] = 32'b00000000000000000010110100111100;
assign LUT_2[34224] = 32'b00000000000000000010011000101100;
assign LUT_2[34225] = 32'b11111111111111111111010001000101;
assign LUT_2[34226] = 32'b00000000000000001001010001101000;
assign LUT_2[34227] = 32'b00000000000000000110001010000001;
assign LUT_2[34228] = 32'b11111111111111111110110110010100;
assign LUT_2[34229] = 32'b11111111111111111011101110101101;
assign LUT_2[34230] = 32'b00000000000000000101101111010000;
assign LUT_2[34231] = 32'b00000000000000000010100111101001;
assign LUT_2[34232] = 32'b11111111111111111101001010001001;
assign LUT_2[34233] = 32'b11111111111111111010000010100010;
assign LUT_2[34234] = 32'b00000000000000000100000011000101;
assign LUT_2[34235] = 32'b00000000000000000000111011011110;
assign LUT_2[34236] = 32'b11111111111111111001100111110001;
assign LUT_2[34237] = 32'b11111111111111110110100000001010;
assign LUT_2[34238] = 32'b00000000000000000000100000101101;
assign LUT_2[34239] = 32'b11111111111111111101011001000110;
assign LUT_2[34240] = 32'b11111111111111111111100001011100;
assign LUT_2[34241] = 32'b11111111111111111100011001110101;
assign LUT_2[34242] = 32'b00000000000000000110011010011000;
assign LUT_2[34243] = 32'b00000000000000000011010010110001;
assign LUT_2[34244] = 32'b11111111111111111011111111000100;
assign LUT_2[34245] = 32'b11111111111111111000110111011101;
assign LUT_2[34246] = 32'b00000000000000000010111000000000;
assign LUT_2[34247] = 32'b11111111111111111111110000011001;
assign LUT_2[34248] = 32'b11111111111111111010010010111001;
assign LUT_2[34249] = 32'b11111111111111110111001011010010;
assign LUT_2[34250] = 32'b00000000000000000001001011110101;
assign LUT_2[34251] = 32'b11111111111111111110000100001110;
assign LUT_2[34252] = 32'b11111111111111110110110000100001;
assign LUT_2[34253] = 32'b11111111111111110011101000111010;
assign LUT_2[34254] = 32'b11111111111111111101101001011101;
assign LUT_2[34255] = 32'b11111111111111111010100001110110;
assign LUT_2[34256] = 32'b11111111111111111010000101100110;
assign LUT_2[34257] = 32'b11111111111111110110111101111111;
assign LUT_2[34258] = 32'b00000000000000000000111110100010;
assign LUT_2[34259] = 32'b11111111111111111101110110111011;
assign LUT_2[34260] = 32'b11111111111111110110100011001110;
assign LUT_2[34261] = 32'b11111111111111110011011011100111;
assign LUT_2[34262] = 32'b11111111111111111101011100001010;
assign LUT_2[34263] = 32'b11111111111111111010010100100011;
assign LUT_2[34264] = 32'b11111111111111110100110111000011;
assign LUT_2[34265] = 32'b11111111111111110001101111011100;
assign LUT_2[34266] = 32'b11111111111111111011101111111111;
assign LUT_2[34267] = 32'b11111111111111111000101000011000;
assign LUT_2[34268] = 32'b11111111111111110001010100101011;
assign LUT_2[34269] = 32'b11111111111111101110001101000100;
assign LUT_2[34270] = 32'b11111111111111111000001101100111;
assign LUT_2[34271] = 32'b11111111111111110101000110000000;
assign LUT_2[34272] = 32'b11111111111111111111111101000101;
assign LUT_2[34273] = 32'b11111111111111111100110101011110;
assign LUT_2[34274] = 32'b00000000000000000110110110000001;
assign LUT_2[34275] = 32'b00000000000000000011101110011010;
assign LUT_2[34276] = 32'b11111111111111111100011010101101;
assign LUT_2[34277] = 32'b11111111111111111001010011000110;
assign LUT_2[34278] = 32'b00000000000000000011010011101001;
assign LUT_2[34279] = 32'b00000000000000000000001100000010;
assign LUT_2[34280] = 32'b11111111111111111010101110100010;
assign LUT_2[34281] = 32'b11111111111111110111100110111011;
assign LUT_2[34282] = 32'b00000000000000000001100111011110;
assign LUT_2[34283] = 32'b11111111111111111110011111110111;
assign LUT_2[34284] = 32'b11111111111111110111001100001010;
assign LUT_2[34285] = 32'b11111111111111110100000100100011;
assign LUT_2[34286] = 32'b11111111111111111110000101000110;
assign LUT_2[34287] = 32'b11111111111111111010111101011111;
assign LUT_2[34288] = 32'b11111111111111111010100001001111;
assign LUT_2[34289] = 32'b11111111111111110111011001101000;
assign LUT_2[34290] = 32'b00000000000000000001011010001011;
assign LUT_2[34291] = 32'b11111111111111111110010010100100;
assign LUT_2[34292] = 32'b11111111111111110110111110110111;
assign LUT_2[34293] = 32'b11111111111111110011110111010000;
assign LUT_2[34294] = 32'b11111111111111111101110111110011;
assign LUT_2[34295] = 32'b11111111111111111010110000001100;
assign LUT_2[34296] = 32'b11111111111111110101010010101100;
assign LUT_2[34297] = 32'b11111111111111110010001011000101;
assign LUT_2[34298] = 32'b11111111111111111100001011101000;
assign LUT_2[34299] = 32'b11111111111111111001000100000001;
assign LUT_2[34300] = 32'b11111111111111110001110000010100;
assign LUT_2[34301] = 32'b11111111111111101110101000101101;
assign LUT_2[34302] = 32'b11111111111111111000101001010000;
assign LUT_2[34303] = 32'b11111111111111110101100001101001;
assign LUT_2[34304] = 32'b00000000000000000011110111110110;
assign LUT_2[34305] = 32'b00000000000000000000110000001111;
assign LUT_2[34306] = 32'b00000000000000001010110000110010;
assign LUT_2[34307] = 32'b00000000000000000111101001001011;
assign LUT_2[34308] = 32'b00000000000000000000010101011110;
assign LUT_2[34309] = 32'b11111111111111111101001101110111;
assign LUT_2[34310] = 32'b00000000000000000111001110011010;
assign LUT_2[34311] = 32'b00000000000000000100000110110011;
assign LUT_2[34312] = 32'b11111111111111111110101001010011;
assign LUT_2[34313] = 32'b11111111111111111011100001101100;
assign LUT_2[34314] = 32'b00000000000000000101100010001111;
assign LUT_2[34315] = 32'b00000000000000000010011010101000;
assign LUT_2[34316] = 32'b11111111111111111011000110111011;
assign LUT_2[34317] = 32'b11111111111111110111111111010100;
assign LUT_2[34318] = 32'b00000000000000000001111111110111;
assign LUT_2[34319] = 32'b11111111111111111110111000010000;
assign LUT_2[34320] = 32'b11111111111111111110011100000000;
assign LUT_2[34321] = 32'b11111111111111111011010100011001;
assign LUT_2[34322] = 32'b00000000000000000101010100111100;
assign LUT_2[34323] = 32'b00000000000000000010001101010101;
assign LUT_2[34324] = 32'b11111111111111111010111001101000;
assign LUT_2[34325] = 32'b11111111111111110111110010000001;
assign LUT_2[34326] = 32'b00000000000000000001110010100100;
assign LUT_2[34327] = 32'b11111111111111111110101010111101;
assign LUT_2[34328] = 32'b11111111111111111001001101011101;
assign LUT_2[34329] = 32'b11111111111111110110000101110110;
assign LUT_2[34330] = 32'b00000000000000000000000110011001;
assign LUT_2[34331] = 32'b11111111111111111100111110110010;
assign LUT_2[34332] = 32'b11111111111111110101101011000101;
assign LUT_2[34333] = 32'b11111111111111110010100011011110;
assign LUT_2[34334] = 32'b11111111111111111100100100000001;
assign LUT_2[34335] = 32'b11111111111111111001011100011010;
assign LUT_2[34336] = 32'b00000000000000000100010011011111;
assign LUT_2[34337] = 32'b00000000000000000001001011111000;
assign LUT_2[34338] = 32'b00000000000000001011001100011011;
assign LUT_2[34339] = 32'b00000000000000001000000100110100;
assign LUT_2[34340] = 32'b00000000000000000000110001000111;
assign LUT_2[34341] = 32'b11111111111111111101101001100000;
assign LUT_2[34342] = 32'b00000000000000000111101010000011;
assign LUT_2[34343] = 32'b00000000000000000100100010011100;
assign LUT_2[34344] = 32'b11111111111111111111000100111100;
assign LUT_2[34345] = 32'b11111111111111111011111101010101;
assign LUT_2[34346] = 32'b00000000000000000101111101111000;
assign LUT_2[34347] = 32'b00000000000000000010110110010001;
assign LUT_2[34348] = 32'b11111111111111111011100010100100;
assign LUT_2[34349] = 32'b11111111111111111000011010111101;
assign LUT_2[34350] = 32'b00000000000000000010011011100000;
assign LUT_2[34351] = 32'b11111111111111111111010011111001;
assign LUT_2[34352] = 32'b11111111111111111110110111101001;
assign LUT_2[34353] = 32'b11111111111111111011110000000010;
assign LUT_2[34354] = 32'b00000000000000000101110000100101;
assign LUT_2[34355] = 32'b00000000000000000010101000111110;
assign LUT_2[34356] = 32'b11111111111111111011010101010001;
assign LUT_2[34357] = 32'b11111111111111111000001101101010;
assign LUT_2[34358] = 32'b00000000000000000010001110001101;
assign LUT_2[34359] = 32'b11111111111111111111000110100110;
assign LUT_2[34360] = 32'b11111111111111111001101001000110;
assign LUT_2[34361] = 32'b11111111111111110110100001011111;
assign LUT_2[34362] = 32'b00000000000000000000100010000010;
assign LUT_2[34363] = 32'b11111111111111111101011010011011;
assign LUT_2[34364] = 32'b11111111111111110110000110101110;
assign LUT_2[34365] = 32'b11111111111111110010111111000111;
assign LUT_2[34366] = 32'b11111111111111111100111111101010;
assign LUT_2[34367] = 32'b11111111111111111001111000000011;
assign LUT_2[34368] = 32'b11111111111111111100000000011001;
assign LUT_2[34369] = 32'b11111111111111111000111000110010;
assign LUT_2[34370] = 32'b00000000000000000010111001010101;
assign LUT_2[34371] = 32'b11111111111111111111110001101110;
assign LUT_2[34372] = 32'b11111111111111111000011110000001;
assign LUT_2[34373] = 32'b11111111111111110101010110011010;
assign LUT_2[34374] = 32'b11111111111111111111010110111101;
assign LUT_2[34375] = 32'b11111111111111111100001111010110;
assign LUT_2[34376] = 32'b11111111111111110110110001110110;
assign LUT_2[34377] = 32'b11111111111111110011101010001111;
assign LUT_2[34378] = 32'b11111111111111111101101010110010;
assign LUT_2[34379] = 32'b11111111111111111010100011001011;
assign LUT_2[34380] = 32'b11111111111111110011001111011110;
assign LUT_2[34381] = 32'b11111111111111110000000111110111;
assign LUT_2[34382] = 32'b11111111111111111010001000011010;
assign LUT_2[34383] = 32'b11111111111111110111000000110011;
assign LUT_2[34384] = 32'b11111111111111110110100100100011;
assign LUT_2[34385] = 32'b11111111111111110011011100111100;
assign LUT_2[34386] = 32'b11111111111111111101011101011111;
assign LUT_2[34387] = 32'b11111111111111111010010101111000;
assign LUT_2[34388] = 32'b11111111111111110011000010001011;
assign LUT_2[34389] = 32'b11111111111111101111111010100100;
assign LUT_2[34390] = 32'b11111111111111111001111011000111;
assign LUT_2[34391] = 32'b11111111111111110110110011100000;
assign LUT_2[34392] = 32'b11111111111111110001010110000000;
assign LUT_2[34393] = 32'b11111111111111101110001110011001;
assign LUT_2[34394] = 32'b11111111111111111000001110111100;
assign LUT_2[34395] = 32'b11111111111111110101000111010101;
assign LUT_2[34396] = 32'b11111111111111101101110011101000;
assign LUT_2[34397] = 32'b11111111111111101010101100000001;
assign LUT_2[34398] = 32'b11111111111111110100101100100100;
assign LUT_2[34399] = 32'b11111111111111110001100100111101;
assign LUT_2[34400] = 32'b11111111111111111100011100000010;
assign LUT_2[34401] = 32'b11111111111111111001010100011011;
assign LUT_2[34402] = 32'b00000000000000000011010100111110;
assign LUT_2[34403] = 32'b00000000000000000000001101010111;
assign LUT_2[34404] = 32'b11111111111111111000111001101010;
assign LUT_2[34405] = 32'b11111111111111110101110010000011;
assign LUT_2[34406] = 32'b11111111111111111111110010100110;
assign LUT_2[34407] = 32'b11111111111111111100101010111111;
assign LUT_2[34408] = 32'b11111111111111110111001101011111;
assign LUT_2[34409] = 32'b11111111111111110100000101111000;
assign LUT_2[34410] = 32'b11111111111111111110000110011011;
assign LUT_2[34411] = 32'b11111111111111111010111110110100;
assign LUT_2[34412] = 32'b11111111111111110011101011000111;
assign LUT_2[34413] = 32'b11111111111111110000100011100000;
assign LUT_2[34414] = 32'b11111111111111111010100100000011;
assign LUT_2[34415] = 32'b11111111111111110111011100011100;
assign LUT_2[34416] = 32'b11111111111111110111000000001100;
assign LUT_2[34417] = 32'b11111111111111110011111000100101;
assign LUT_2[34418] = 32'b11111111111111111101111001001000;
assign LUT_2[34419] = 32'b11111111111111111010110001100001;
assign LUT_2[34420] = 32'b11111111111111110011011101110100;
assign LUT_2[34421] = 32'b11111111111111110000010110001101;
assign LUT_2[34422] = 32'b11111111111111111010010110110000;
assign LUT_2[34423] = 32'b11111111111111110111001111001001;
assign LUT_2[34424] = 32'b11111111111111110001110001101001;
assign LUT_2[34425] = 32'b11111111111111101110101010000010;
assign LUT_2[34426] = 32'b11111111111111111000101010100101;
assign LUT_2[34427] = 32'b11111111111111110101100010111110;
assign LUT_2[34428] = 32'b11111111111111101110001111010001;
assign LUT_2[34429] = 32'b11111111111111101011000111101010;
assign LUT_2[34430] = 32'b11111111111111110101001000001101;
assign LUT_2[34431] = 32'b11111111111111110010000000100110;
assign LUT_2[34432] = 32'b00000000000000001000001100000101;
assign LUT_2[34433] = 32'b00000000000000000101000100011110;
assign LUT_2[34434] = 32'b00000000000000001111000101000001;
assign LUT_2[34435] = 32'b00000000000000001011111101011010;
assign LUT_2[34436] = 32'b00000000000000000100101001101101;
assign LUT_2[34437] = 32'b00000000000000000001100010000110;
assign LUT_2[34438] = 32'b00000000000000001011100010101001;
assign LUT_2[34439] = 32'b00000000000000001000011011000010;
assign LUT_2[34440] = 32'b00000000000000000010111101100010;
assign LUT_2[34441] = 32'b11111111111111111111110101111011;
assign LUT_2[34442] = 32'b00000000000000001001110110011110;
assign LUT_2[34443] = 32'b00000000000000000110101110110111;
assign LUT_2[34444] = 32'b11111111111111111111011011001010;
assign LUT_2[34445] = 32'b11111111111111111100010011100011;
assign LUT_2[34446] = 32'b00000000000000000110010100000110;
assign LUT_2[34447] = 32'b00000000000000000011001100011111;
assign LUT_2[34448] = 32'b00000000000000000010110000001111;
assign LUT_2[34449] = 32'b11111111111111111111101000101000;
assign LUT_2[34450] = 32'b00000000000000001001101001001011;
assign LUT_2[34451] = 32'b00000000000000000110100001100100;
assign LUT_2[34452] = 32'b11111111111111111111001101110111;
assign LUT_2[34453] = 32'b11111111111111111100000110010000;
assign LUT_2[34454] = 32'b00000000000000000110000110110011;
assign LUT_2[34455] = 32'b00000000000000000010111111001100;
assign LUT_2[34456] = 32'b11111111111111111101100001101100;
assign LUT_2[34457] = 32'b11111111111111111010011010000101;
assign LUT_2[34458] = 32'b00000000000000000100011010101000;
assign LUT_2[34459] = 32'b00000000000000000001010011000001;
assign LUT_2[34460] = 32'b11111111111111111001111111010100;
assign LUT_2[34461] = 32'b11111111111111110110110111101101;
assign LUT_2[34462] = 32'b00000000000000000000111000010000;
assign LUT_2[34463] = 32'b11111111111111111101110000101001;
assign LUT_2[34464] = 32'b00000000000000001000100111101110;
assign LUT_2[34465] = 32'b00000000000000000101100000000111;
assign LUT_2[34466] = 32'b00000000000000001111100000101010;
assign LUT_2[34467] = 32'b00000000000000001100011001000011;
assign LUT_2[34468] = 32'b00000000000000000101000101010110;
assign LUT_2[34469] = 32'b00000000000000000001111101101111;
assign LUT_2[34470] = 32'b00000000000000001011111110010010;
assign LUT_2[34471] = 32'b00000000000000001000110110101011;
assign LUT_2[34472] = 32'b00000000000000000011011001001011;
assign LUT_2[34473] = 32'b00000000000000000000010001100100;
assign LUT_2[34474] = 32'b00000000000000001010010010000111;
assign LUT_2[34475] = 32'b00000000000000000111001010100000;
assign LUT_2[34476] = 32'b11111111111111111111110110110011;
assign LUT_2[34477] = 32'b11111111111111111100101111001100;
assign LUT_2[34478] = 32'b00000000000000000110101111101111;
assign LUT_2[34479] = 32'b00000000000000000011101000001000;
assign LUT_2[34480] = 32'b00000000000000000011001011111000;
assign LUT_2[34481] = 32'b00000000000000000000000100010001;
assign LUT_2[34482] = 32'b00000000000000001010000100110100;
assign LUT_2[34483] = 32'b00000000000000000110111101001101;
assign LUT_2[34484] = 32'b11111111111111111111101001100000;
assign LUT_2[34485] = 32'b11111111111111111100100001111001;
assign LUT_2[34486] = 32'b00000000000000000110100010011100;
assign LUT_2[34487] = 32'b00000000000000000011011010110101;
assign LUT_2[34488] = 32'b11111111111111111101111101010101;
assign LUT_2[34489] = 32'b11111111111111111010110101101110;
assign LUT_2[34490] = 32'b00000000000000000100110110010001;
assign LUT_2[34491] = 32'b00000000000000000001101110101010;
assign LUT_2[34492] = 32'b11111111111111111010011010111101;
assign LUT_2[34493] = 32'b11111111111111110111010011010110;
assign LUT_2[34494] = 32'b00000000000000000001010011111001;
assign LUT_2[34495] = 32'b11111111111111111110001100010010;
assign LUT_2[34496] = 32'b00000000000000000000010100101000;
assign LUT_2[34497] = 32'b11111111111111111101001101000001;
assign LUT_2[34498] = 32'b00000000000000000111001101100100;
assign LUT_2[34499] = 32'b00000000000000000100000101111101;
assign LUT_2[34500] = 32'b11111111111111111100110010010000;
assign LUT_2[34501] = 32'b11111111111111111001101010101001;
assign LUT_2[34502] = 32'b00000000000000000011101011001100;
assign LUT_2[34503] = 32'b00000000000000000000100011100101;
assign LUT_2[34504] = 32'b11111111111111111011000110000101;
assign LUT_2[34505] = 32'b11111111111111110111111110011110;
assign LUT_2[34506] = 32'b00000000000000000001111111000001;
assign LUT_2[34507] = 32'b11111111111111111110110111011010;
assign LUT_2[34508] = 32'b11111111111111110111100011101101;
assign LUT_2[34509] = 32'b11111111111111110100011100000110;
assign LUT_2[34510] = 32'b11111111111111111110011100101001;
assign LUT_2[34511] = 32'b11111111111111111011010101000010;
assign LUT_2[34512] = 32'b11111111111111111010111000110010;
assign LUT_2[34513] = 32'b11111111111111110111110001001011;
assign LUT_2[34514] = 32'b00000000000000000001110001101110;
assign LUT_2[34515] = 32'b11111111111111111110101010000111;
assign LUT_2[34516] = 32'b11111111111111110111010110011010;
assign LUT_2[34517] = 32'b11111111111111110100001110110011;
assign LUT_2[34518] = 32'b11111111111111111110001111010110;
assign LUT_2[34519] = 32'b11111111111111111011000111101111;
assign LUT_2[34520] = 32'b11111111111111110101101010001111;
assign LUT_2[34521] = 32'b11111111111111110010100010101000;
assign LUT_2[34522] = 32'b11111111111111111100100011001011;
assign LUT_2[34523] = 32'b11111111111111111001011011100100;
assign LUT_2[34524] = 32'b11111111111111110010000111110111;
assign LUT_2[34525] = 32'b11111111111111101111000000010000;
assign LUT_2[34526] = 32'b11111111111111111001000000110011;
assign LUT_2[34527] = 32'b11111111111111110101111001001100;
assign LUT_2[34528] = 32'b00000000000000000000110000010001;
assign LUT_2[34529] = 32'b11111111111111111101101000101010;
assign LUT_2[34530] = 32'b00000000000000000111101001001101;
assign LUT_2[34531] = 32'b00000000000000000100100001100110;
assign LUT_2[34532] = 32'b11111111111111111101001101111001;
assign LUT_2[34533] = 32'b11111111111111111010000110010010;
assign LUT_2[34534] = 32'b00000000000000000100000110110101;
assign LUT_2[34535] = 32'b00000000000000000000111111001110;
assign LUT_2[34536] = 32'b11111111111111111011100001101110;
assign LUT_2[34537] = 32'b11111111111111111000011010000111;
assign LUT_2[34538] = 32'b00000000000000000010011010101010;
assign LUT_2[34539] = 32'b11111111111111111111010011000011;
assign LUT_2[34540] = 32'b11111111111111110111111111010110;
assign LUT_2[34541] = 32'b11111111111111110100110111101111;
assign LUT_2[34542] = 32'b11111111111111111110111000010010;
assign LUT_2[34543] = 32'b11111111111111111011110000101011;
assign LUT_2[34544] = 32'b11111111111111111011010100011011;
assign LUT_2[34545] = 32'b11111111111111111000001100110100;
assign LUT_2[34546] = 32'b00000000000000000010001101010111;
assign LUT_2[34547] = 32'b11111111111111111111000101110000;
assign LUT_2[34548] = 32'b11111111111111110111110010000011;
assign LUT_2[34549] = 32'b11111111111111110100101010011100;
assign LUT_2[34550] = 32'b11111111111111111110101010111111;
assign LUT_2[34551] = 32'b11111111111111111011100011011000;
assign LUT_2[34552] = 32'b11111111111111110110000101111000;
assign LUT_2[34553] = 32'b11111111111111110010111110010001;
assign LUT_2[34554] = 32'b11111111111111111100111110110100;
assign LUT_2[34555] = 32'b11111111111111111001110111001101;
assign LUT_2[34556] = 32'b11111111111111110010100011100000;
assign LUT_2[34557] = 32'b11111111111111101111011011111001;
assign LUT_2[34558] = 32'b11111111111111111001011100011100;
assign LUT_2[34559] = 32'b11111111111111110110010100110101;
assign LUT_2[34560] = 32'b00000000000000000111110110011100;
assign LUT_2[34561] = 32'b00000000000000000100101110110101;
assign LUT_2[34562] = 32'b00000000000000001110101111011000;
assign LUT_2[34563] = 32'b00000000000000001011100111110001;
assign LUT_2[34564] = 32'b00000000000000000100010100000100;
assign LUT_2[34565] = 32'b00000000000000000001001100011101;
assign LUT_2[34566] = 32'b00000000000000001011001101000000;
assign LUT_2[34567] = 32'b00000000000000001000000101011001;
assign LUT_2[34568] = 32'b00000000000000000010100111111001;
assign LUT_2[34569] = 32'b11111111111111111111100000010010;
assign LUT_2[34570] = 32'b00000000000000001001100000110101;
assign LUT_2[34571] = 32'b00000000000000000110011001001110;
assign LUT_2[34572] = 32'b11111111111111111111000101100001;
assign LUT_2[34573] = 32'b11111111111111111011111101111010;
assign LUT_2[34574] = 32'b00000000000000000101111110011101;
assign LUT_2[34575] = 32'b00000000000000000010110110110110;
assign LUT_2[34576] = 32'b00000000000000000010011010100110;
assign LUT_2[34577] = 32'b11111111111111111111010010111111;
assign LUT_2[34578] = 32'b00000000000000001001010011100010;
assign LUT_2[34579] = 32'b00000000000000000110001011111011;
assign LUT_2[34580] = 32'b11111111111111111110111000001110;
assign LUT_2[34581] = 32'b11111111111111111011110000100111;
assign LUT_2[34582] = 32'b00000000000000000101110001001010;
assign LUT_2[34583] = 32'b00000000000000000010101001100011;
assign LUT_2[34584] = 32'b11111111111111111101001100000011;
assign LUT_2[34585] = 32'b11111111111111111010000100011100;
assign LUT_2[34586] = 32'b00000000000000000100000100111111;
assign LUT_2[34587] = 32'b00000000000000000000111101011000;
assign LUT_2[34588] = 32'b11111111111111111001101001101011;
assign LUT_2[34589] = 32'b11111111111111110110100010000100;
assign LUT_2[34590] = 32'b00000000000000000000100010100111;
assign LUT_2[34591] = 32'b11111111111111111101011011000000;
assign LUT_2[34592] = 32'b00000000000000001000010010000101;
assign LUT_2[34593] = 32'b00000000000000000101001010011110;
assign LUT_2[34594] = 32'b00000000000000001111001011000001;
assign LUT_2[34595] = 32'b00000000000000001100000011011010;
assign LUT_2[34596] = 32'b00000000000000000100101111101101;
assign LUT_2[34597] = 32'b00000000000000000001101000000110;
assign LUT_2[34598] = 32'b00000000000000001011101000101001;
assign LUT_2[34599] = 32'b00000000000000001000100001000010;
assign LUT_2[34600] = 32'b00000000000000000011000011100010;
assign LUT_2[34601] = 32'b11111111111111111111111011111011;
assign LUT_2[34602] = 32'b00000000000000001001111100011110;
assign LUT_2[34603] = 32'b00000000000000000110110100110111;
assign LUT_2[34604] = 32'b11111111111111111111100001001010;
assign LUT_2[34605] = 32'b11111111111111111100011001100011;
assign LUT_2[34606] = 32'b00000000000000000110011010000110;
assign LUT_2[34607] = 32'b00000000000000000011010010011111;
assign LUT_2[34608] = 32'b00000000000000000010110110001111;
assign LUT_2[34609] = 32'b11111111111111111111101110101000;
assign LUT_2[34610] = 32'b00000000000000001001101111001011;
assign LUT_2[34611] = 32'b00000000000000000110100111100100;
assign LUT_2[34612] = 32'b11111111111111111111010011110111;
assign LUT_2[34613] = 32'b11111111111111111100001100010000;
assign LUT_2[34614] = 32'b00000000000000000110001100110011;
assign LUT_2[34615] = 32'b00000000000000000011000101001100;
assign LUT_2[34616] = 32'b11111111111111111101100111101100;
assign LUT_2[34617] = 32'b11111111111111111010100000000101;
assign LUT_2[34618] = 32'b00000000000000000100100000101000;
assign LUT_2[34619] = 32'b00000000000000000001011001000001;
assign LUT_2[34620] = 32'b11111111111111111010000101010100;
assign LUT_2[34621] = 32'b11111111111111110110111101101101;
assign LUT_2[34622] = 32'b00000000000000000000111110010000;
assign LUT_2[34623] = 32'b11111111111111111101110110101001;
assign LUT_2[34624] = 32'b11111111111111111111111110111111;
assign LUT_2[34625] = 32'b11111111111111111100110111011000;
assign LUT_2[34626] = 32'b00000000000000000110110111111011;
assign LUT_2[34627] = 32'b00000000000000000011110000010100;
assign LUT_2[34628] = 32'b11111111111111111100011100100111;
assign LUT_2[34629] = 32'b11111111111111111001010101000000;
assign LUT_2[34630] = 32'b00000000000000000011010101100011;
assign LUT_2[34631] = 32'b00000000000000000000001101111100;
assign LUT_2[34632] = 32'b11111111111111111010110000011100;
assign LUT_2[34633] = 32'b11111111111111110111101000110101;
assign LUT_2[34634] = 32'b00000000000000000001101001011000;
assign LUT_2[34635] = 32'b11111111111111111110100001110001;
assign LUT_2[34636] = 32'b11111111111111110111001110000100;
assign LUT_2[34637] = 32'b11111111111111110100000110011101;
assign LUT_2[34638] = 32'b11111111111111111110000111000000;
assign LUT_2[34639] = 32'b11111111111111111010111111011001;
assign LUT_2[34640] = 32'b11111111111111111010100011001001;
assign LUT_2[34641] = 32'b11111111111111110111011011100010;
assign LUT_2[34642] = 32'b00000000000000000001011100000101;
assign LUT_2[34643] = 32'b11111111111111111110010100011110;
assign LUT_2[34644] = 32'b11111111111111110111000000110001;
assign LUT_2[34645] = 32'b11111111111111110011111001001010;
assign LUT_2[34646] = 32'b11111111111111111101111001101101;
assign LUT_2[34647] = 32'b11111111111111111010110010000110;
assign LUT_2[34648] = 32'b11111111111111110101010100100110;
assign LUT_2[34649] = 32'b11111111111111110010001100111111;
assign LUT_2[34650] = 32'b11111111111111111100001101100010;
assign LUT_2[34651] = 32'b11111111111111111001000101111011;
assign LUT_2[34652] = 32'b11111111111111110001110010001110;
assign LUT_2[34653] = 32'b11111111111111101110101010100111;
assign LUT_2[34654] = 32'b11111111111111111000101011001010;
assign LUT_2[34655] = 32'b11111111111111110101100011100011;
assign LUT_2[34656] = 32'b00000000000000000000011010101000;
assign LUT_2[34657] = 32'b11111111111111111101010011000001;
assign LUT_2[34658] = 32'b00000000000000000111010011100100;
assign LUT_2[34659] = 32'b00000000000000000100001011111101;
assign LUT_2[34660] = 32'b11111111111111111100111000010000;
assign LUT_2[34661] = 32'b11111111111111111001110000101001;
assign LUT_2[34662] = 32'b00000000000000000011110001001100;
assign LUT_2[34663] = 32'b00000000000000000000101001100101;
assign LUT_2[34664] = 32'b11111111111111111011001100000101;
assign LUT_2[34665] = 32'b11111111111111111000000100011110;
assign LUT_2[34666] = 32'b00000000000000000010000101000001;
assign LUT_2[34667] = 32'b11111111111111111110111101011010;
assign LUT_2[34668] = 32'b11111111111111110111101001101101;
assign LUT_2[34669] = 32'b11111111111111110100100010000110;
assign LUT_2[34670] = 32'b11111111111111111110100010101001;
assign LUT_2[34671] = 32'b11111111111111111011011011000010;
assign LUT_2[34672] = 32'b11111111111111111010111110110010;
assign LUT_2[34673] = 32'b11111111111111110111110111001011;
assign LUT_2[34674] = 32'b00000000000000000001110111101110;
assign LUT_2[34675] = 32'b11111111111111111110110000000111;
assign LUT_2[34676] = 32'b11111111111111110111011100011010;
assign LUT_2[34677] = 32'b11111111111111110100010100110011;
assign LUT_2[34678] = 32'b11111111111111111110010101010110;
assign LUT_2[34679] = 32'b11111111111111111011001101101111;
assign LUT_2[34680] = 32'b11111111111111110101110000001111;
assign LUT_2[34681] = 32'b11111111111111110010101000101000;
assign LUT_2[34682] = 32'b11111111111111111100101001001011;
assign LUT_2[34683] = 32'b11111111111111111001100001100100;
assign LUT_2[34684] = 32'b11111111111111110010001101110111;
assign LUT_2[34685] = 32'b11111111111111101111000110010000;
assign LUT_2[34686] = 32'b11111111111111111001000110110011;
assign LUT_2[34687] = 32'b11111111111111110101111111001100;
assign LUT_2[34688] = 32'b00000000000000001100001010101011;
assign LUT_2[34689] = 32'b00000000000000001001000011000100;
assign LUT_2[34690] = 32'b00000000000000010011000011100111;
assign LUT_2[34691] = 32'b00000000000000001111111100000000;
assign LUT_2[34692] = 32'b00000000000000001000101000010011;
assign LUT_2[34693] = 32'b00000000000000000101100000101100;
assign LUT_2[34694] = 32'b00000000000000001111100001001111;
assign LUT_2[34695] = 32'b00000000000000001100011001101000;
assign LUT_2[34696] = 32'b00000000000000000110111100001000;
assign LUT_2[34697] = 32'b00000000000000000011110100100001;
assign LUT_2[34698] = 32'b00000000000000001101110101000100;
assign LUT_2[34699] = 32'b00000000000000001010101101011101;
assign LUT_2[34700] = 32'b00000000000000000011011001110000;
assign LUT_2[34701] = 32'b00000000000000000000010010001001;
assign LUT_2[34702] = 32'b00000000000000001010010010101100;
assign LUT_2[34703] = 32'b00000000000000000111001011000101;
assign LUT_2[34704] = 32'b00000000000000000110101110110101;
assign LUT_2[34705] = 32'b00000000000000000011100111001110;
assign LUT_2[34706] = 32'b00000000000000001101100111110001;
assign LUT_2[34707] = 32'b00000000000000001010100000001010;
assign LUT_2[34708] = 32'b00000000000000000011001100011101;
assign LUT_2[34709] = 32'b00000000000000000000000100110110;
assign LUT_2[34710] = 32'b00000000000000001010000101011001;
assign LUT_2[34711] = 32'b00000000000000000110111101110010;
assign LUT_2[34712] = 32'b00000000000000000001100000010010;
assign LUT_2[34713] = 32'b11111111111111111110011000101011;
assign LUT_2[34714] = 32'b00000000000000001000011001001110;
assign LUT_2[34715] = 32'b00000000000000000101010001100111;
assign LUT_2[34716] = 32'b11111111111111111101111101111010;
assign LUT_2[34717] = 32'b11111111111111111010110110010011;
assign LUT_2[34718] = 32'b00000000000000000100110110110110;
assign LUT_2[34719] = 32'b00000000000000000001101111001111;
assign LUT_2[34720] = 32'b00000000000000001100100110010100;
assign LUT_2[34721] = 32'b00000000000000001001011110101101;
assign LUT_2[34722] = 32'b00000000000000010011011111010000;
assign LUT_2[34723] = 32'b00000000000000010000010111101001;
assign LUT_2[34724] = 32'b00000000000000001001000011111100;
assign LUT_2[34725] = 32'b00000000000000000101111100010101;
assign LUT_2[34726] = 32'b00000000000000001111111100111000;
assign LUT_2[34727] = 32'b00000000000000001100110101010001;
assign LUT_2[34728] = 32'b00000000000000000111010111110001;
assign LUT_2[34729] = 32'b00000000000000000100010000001010;
assign LUT_2[34730] = 32'b00000000000000001110010000101101;
assign LUT_2[34731] = 32'b00000000000000001011001001000110;
assign LUT_2[34732] = 32'b00000000000000000011110101011001;
assign LUT_2[34733] = 32'b00000000000000000000101101110010;
assign LUT_2[34734] = 32'b00000000000000001010101110010101;
assign LUT_2[34735] = 32'b00000000000000000111100110101110;
assign LUT_2[34736] = 32'b00000000000000000111001010011110;
assign LUT_2[34737] = 32'b00000000000000000100000010110111;
assign LUT_2[34738] = 32'b00000000000000001110000011011010;
assign LUT_2[34739] = 32'b00000000000000001010111011110011;
assign LUT_2[34740] = 32'b00000000000000000011101000000110;
assign LUT_2[34741] = 32'b00000000000000000000100000011111;
assign LUT_2[34742] = 32'b00000000000000001010100001000010;
assign LUT_2[34743] = 32'b00000000000000000111011001011011;
assign LUT_2[34744] = 32'b00000000000000000001111011111011;
assign LUT_2[34745] = 32'b11111111111111111110110100010100;
assign LUT_2[34746] = 32'b00000000000000001000110100110111;
assign LUT_2[34747] = 32'b00000000000000000101101101010000;
assign LUT_2[34748] = 32'b11111111111111111110011001100011;
assign LUT_2[34749] = 32'b11111111111111111011010001111100;
assign LUT_2[34750] = 32'b00000000000000000101010010011111;
assign LUT_2[34751] = 32'b00000000000000000010001010111000;
assign LUT_2[34752] = 32'b00000000000000000100010011001110;
assign LUT_2[34753] = 32'b00000000000000000001001011100111;
assign LUT_2[34754] = 32'b00000000000000001011001100001010;
assign LUT_2[34755] = 32'b00000000000000001000000100100011;
assign LUT_2[34756] = 32'b00000000000000000000110000110110;
assign LUT_2[34757] = 32'b11111111111111111101101001001111;
assign LUT_2[34758] = 32'b00000000000000000111101001110010;
assign LUT_2[34759] = 32'b00000000000000000100100010001011;
assign LUT_2[34760] = 32'b11111111111111111111000100101011;
assign LUT_2[34761] = 32'b11111111111111111011111101000100;
assign LUT_2[34762] = 32'b00000000000000000101111101100111;
assign LUT_2[34763] = 32'b00000000000000000010110110000000;
assign LUT_2[34764] = 32'b11111111111111111011100010010011;
assign LUT_2[34765] = 32'b11111111111111111000011010101100;
assign LUT_2[34766] = 32'b00000000000000000010011011001111;
assign LUT_2[34767] = 32'b11111111111111111111010011101000;
assign LUT_2[34768] = 32'b11111111111111111110110111011000;
assign LUT_2[34769] = 32'b11111111111111111011101111110001;
assign LUT_2[34770] = 32'b00000000000000000101110000010100;
assign LUT_2[34771] = 32'b00000000000000000010101000101101;
assign LUT_2[34772] = 32'b11111111111111111011010101000000;
assign LUT_2[34773] = 32'b11111111111111111000001101011001;
assign LUT_2[34774] = 32'b00000000000000000010001101111100;
assign LUT_2[34775] = 32'b11111111111111111111000110010101;
assign LUT_2[34776] = 32'b11111111111111111001101000110101;
assign LUT_2[34777] = 32'b11111111111111110110100001001110;
assign LUT_2[34778] = 32'b00000000000000000000100001110001;
assign LUT_2[34779] = 32'b11111111111111111101011010001010;
assign LUT_2[34780] = 32'b11111111111111110110000110011101;
assign LUT_2[34781] = 32'b11111111111111110010111110110110;
assign LUT_2[34782] = 32'b11111111111111111100111111011001;
assign LUT_2[34783] = 32'b11111111111111111001110111110010;
assign LUT_2[34784] = 32'b00000000000000000100101110110111;
assign LUT_2[34785] = 32'b00000000000000000001100111010000;
assign LUT_2[34786] = 32'b00000000000000001011100111110011;
assign LUT_2[34787] = 32'b00000000000000001000100000001100;
assign LUT_2[34788] = 32'b00000000000000000001001100011111;
assign LUT_2[34789] = 32'b11111111111111111110000100111000;
assign LUT_2[34790] = 32'b00000000000000001000000101011011;
assign LUT_2[34791] = 32'b00000000000000000100111101110100;
assign LUT_2[34792] = 32'b11111111111111111111100000010100;
assign LUT_2[34793] = 32'b11111111111111111100011000101101;
assign LUT_2[34794] = 32'b00000000000000000110011001010000;
assign LUT_2[34795] = 32'b00000000000000000011010001101001;
assign LUT_2[34796] = 32'b11111111111111111011111101111100;
assign LUT_2[34797] = 32'b11111111111111111000110110010101;
assign LUT_2[34798] = 32'b00000000000000000010110110111000;
assign LUT_2[34799] = 32'b11111111111111111111101111010001;
assign LUT_2[34800] = 32'b11111111111111111111010011000001;
assign LUT_2[34801] = 32'b11111111111111111100001011011010;
assign LUT_2[34802] = 32'b00000000000000000110001011111101;
assign LUT_2[34803] = 32'b00000000000000000011000100010110;
assign LUT_2[34804] = 32'b11111111111111111011110000101001;
assign LUT_2[34805] = 32'b11111111111111111000101001000010;
assign LUT_2[34806] = 32'b00000000000000000010101001100101;
assign LUT_2[34807] = 32'b11111111111111111111100001111110;
assign LUT_2[34808] = 32'b11111111111111111010000100011110;
assign LUT_2[34809] = 32'b11111111111111110110111100110111;
assign LUT_2[34810] = 32'b00000000000000000000111101011010;
assign LUT_2[34811] = 32'b11111111111111111101110101110011;
assign LUT_2[34812] = 32'b11111111111111110110100010000110;
assign LUT_2[34813] = 32'b11111111111111110011011010011111;
assign LUT_2[34814] = 32'b11111111111111111101011011000010;
assign LUT_2[34815] = 32'b11111111111111111010010011011011;
assign LUT_2[34816] = 32'b11111111111111110100001111111011;
assign LUT_2[34817] = 32'b11111111111111110001001000010100;
assign LUT_2[34818] = 32'b11111111111111111011001000110111;
assign LUT_2[34819] = 32'b11111111111111111000000001010000;
assign LUT_2[34820] = 32'b11111111111111110000101101100011;
assign LUT_2[34821] = 32'b11111111111111101101100101111100;
assign LUT_2[34822] = 32'b11111111111111110111100110011111;
assign LUT_2[34823] = 32'b11111111111111110100011110111000;
assign LUT_2[34824] = 32'b11111111111111101111000001011000;
assign LUT_2[34825] = 32'b11111111111111101011111001110001;
assign LUT_2[34826] = 32'b11111111111111110101111010010100;
assign LUT_2[34827] = 32'b11111111111111110010110010101101;
assign LUT_2[34828] = 32'b11111111111111101011011111000000;
assign LUT_2[34829] = 32'b11111111111111101000010111011001;
assign LUT_2[34830] = 32'b11111111111111110010010111111100;
assign LUT_2[34831] = 32'b11111111111111101111010000010101;
assign LUT_2[34832] = 32'b11111111111111101110110100000101;
assign LUT_2[34833] = 32'b11111111111111101011101100011110;
assign LUT_2[34834] = 32'b11111111111111110101101101000001;
assign LUT_2[34835] = 32'b11111111111111110010100101011010;
assign LUT_2[34836] = 32'b11111111111111101011010001101101;
assign LUT_2[34837] = 32'b11111111111111101000001010000110;
assign LUT_2[34838] = 32'b11111111111111110010001010101001;
assign LUT_2[34839] = 32'b11111111111111101111000011000010;
assign LUT_2[34840] = 32'b11111111111111101001100101100010;
assign LUT_2[34841] = 32'b11111111111111100110011101111011;
assign LUT_2[34842] = 32'b11111111111111110000011110011110;
assign LUT_2[34843] = 32'b11111111111111101101010110110111;
assign LUT_2[34844] = 32'b11111111111111100110000011001010;
assign LUT_2[34845] = 32'b11111111111111100010111011100011;
assign LUT_2[34846] = 32'b11111111111111101100111100000110;
assign LUT_2[34847] = 32'b11111111111111101001110100011111;
assign LUT_2[34848] = 32'b11111111111111110100101011100100;
assign LUT_2[34849] = 32'b11111111111111110001100011111101;
assign LUT_2[34850] = 32'b11111111111111111011100100100000;
assign LUT_2[34851] = 32'b11111111111111111000011100111001;
assign LUT_2[34852] = 32'b11111111111111110001001001001100;
assign LUT_2[34853] = 32'b11111111111111101110000001100101;
assign LUT_2[34854] = 32'b11111111111111111000000010001000;
assign LUT_2[34855] = 32'b11111111111111110100111010100001;
assign LUT_2[34856] = 32'b11111111111111101111011101000001;
assign LUT_2[34857] = 32'b11111111111111101100010101011010;
assign LUT_2[34858] = 32'b11111111111111110110010101111101;
assign LUT_2[34859] = 32'b11111111111111110011001110010110;
assign LUT_2[34860] = 32'b11111111111111101011111010101001;
assign LUT_2[34861] = 32'b11111111111111101000110011000010;
assign LUT_2[34862] = 32'b11111111111111110010110011100101;
assign LUT_2[34863] = 32'b11111111111111101111101011111110;
assign LUT_2[34864] = 32'b11111111111111101111001111101110;
assign LUT_2[34865] = 32'b11111111111111101100001000000111;
assign LUT_2[34866] = 32'b11111111111111110110001000101010;
assign LUT_2[34867] = 32'b11111111111111110011000001000011;
assign LUT_2[34868] = 32'b11111111111111101011101101010110;
assign LUT_2[34869] = 32'b11111111111111101000100101101111;
assign LUT_2[34870] = 32'b11111111111111110010100110010010;
assign LUT_2[34871] = 32'b11111111111111101111011110101011;
assign LUT_2[34872] = 32'b11111111111111101010000001001011;
assign LUT_2[34873] = 32'b11111111111111100110111001100100;
assign LUT_2[34874] = 32'b11111111111111110000111010000111;
assign LUT_2[34875] = 32'b11111111111111101101110010100000;
assign LUT_2[34876] = 32'b11111111111111100110011110110011;
assign LUT_2[34877] = 32'b11111111111111100011010111001100;
assign LUT_2[34878] = 32'b11111111111111101101010111101111;
assign LUT_2[34879] = 32'b11111111111111101010010000001000;
assign LUT_2[34880] = 32'b11111111111111101100011000011110;
assign LUT_2[34881] = 32'b11111111111111101001010000110111;
assign LUT_2[34882] = 32'b11111111111111110011010001011010;
assign LUT_2[34883] = 32'b11111111111111110000001001110011;
assign LUT_2[34884] = 32'b11111111111111101000110110000110;
assign LUT_2[34885] = 32'b11111111111111100101101110011111;
assign LUT_2[34886] = 32'b11111111111111101111101111000010;
assign LUT_2[34887] = 32'b11111111111111101100100111011011;
assign LUT_2[34888] = 32'b11111111111111100111001001111011;
assign LUT_2[34889] = 32'b11111111111111100100000010010100;
assign LUT_2[34890] = 32'b11111111111111101110000010110111;
assign LUT_2[34891] = 32'b11111111111111101010111011010000;
assign LUT_2[34892] = 32'b11111111111111100011100111100011;
assign LUT_2[34893] = 32'b11111111111111100000011111111100;
assign LUT_2[34894] = 32'b11111111111111101010100000011111;
assign LUT_2[34895] = 32'b11111111111111100111011000111000;
assign LUT_2[34896] = 32'b11111111111111100110111100101000;
assign LUT_2[34897] = 32'b11111111111111100011110101000001;
assign LUT_2[34898] = 32'b11111111111111101101110101100100;
assign LUT_2[34899] = 32'b11111111111111101010101101111101;
assign LUT_2[34900] = 32'b11111111111111100011011010010000;
assign LUT_2[34901] = 32'b11111111111111100000010010101001;
assign LUT_2[34902] = 32'b11111111111111101010010011001100;
assign LUT_2[34903] = 32'b11111111111111100111001011100101;
assign LUT_2[34904] = 32'b11111111111111100001101110000101;
assign LUT_2[34905] = 32'b11111111111111011110100110011110;
assign LUT_2[34906] = 32'b11111111111111101000100111000001;
assign LUT_2[34907] = 32'b11111111111111100101011111011010;
assign LUT_2[34908] = 32'b11111111111111011110001011101101;
assign LUT_2[34909] = 32'b11111111111111011011000100000110;
assign LUT_2[34910] = 32'b11111111111111100101000100101001;
assign LUT_2[34911] = 32'b11111111111111100001111101000010;
assign LUT_2[34912] = 32'b11111111111111101100110100000111;
assign LUT_2[34913] = 32'b11111111111111101001101100100000;
assign LUT_2[34914] = 32'b11111111111111110011101101000011;
assign LUT_2[34915] = 32'b11111111111111110000100101011100;
assign LUT_2[34916] = 32'b11111111111111101001010001101111;
assign LUT_2[34917] = 32'b11111111111111100110001010001000;
assign LUT_2[34918] = 32'b11111111111111110000001010101011;
assign LUT_2[34919] = 32'b11111111111111101101000011000100;
assign LUT_2[34920] = 32'b11111111111111100111100101100100;
assign LUT_2[34921] = 32'b11111111111111100100011101111101;
assign LUT_2[34922] = 32'b11111111111111101110011110100000;
assign LUT_2[34923] = 32'b11111111111111101011010110111001;
assign LUT_2[34924] = 32'b11111111111111100100000011001100;
assign LUT_2[34925] = 32'b11111111111111100000111011100101;
assign LUT_2[34926] = 32'b11111111111111101010111100001000;
assign LUT_2[34927] = 32'b11111111111111100111110100100001;
assign LUT_2[34928] = 32'b11111111111111100111011000010001;
assign LUT_2[34929] = 32'b11111111111111100100010000101010;
assign LUT_2[34930] = 32'b11111111111111101110010001001101;
assign LUT_2[34931] = 32'b11111111111111101011001001100110;
assign LUT_2[34932] = 32'b11111111111111100011110101111001;
assign LUT_2[34933] = 32'b11111111111111100000101110010010;
assign LUT_2[34934] = 32'b11111111111111101010101110110101;
assign LUT_2[34935] = 32'b11111111111111100111100111001110;
assign LUT_2[34936] = 32'b11111111111111100010001001101110;
assign LUT_2[34937] = 32'b11111111111111011111000010000111;
assign LUT_2[34938] = 32'b11111111111111101001000010101010;
assign LUT_2[34939] = 32'b11111111111111100101111011000011;
assign LUT_2[34940] = 32'b11111111111111011110100111010110;
assign LUT_2[34941] = 32'b11111111111111011011011111101111;
assign LUT_2[34942] = 32'b11111111111111100101100000010010;
assign LUT_2[34943] = 32'b11111111111111100010011000101011;
assign LUT_2[34944] = 32'b11111111111111111000100100001010;
assign LUT_2[34945] = 32'b11111111111111110101011100100011;
assign LUT_2[34946] = 32'b11111111111111111111011101000110;
assign LUT_2[34947] = 32'b11111111111111111100010101011111;
assign LUT_2[34948] = 32'b11111111111111110101000001110010;
assign LUT_2[34949] = 32'b11111111111111110001111010001011;
assign LUT_2[34950] = 32'b11111111111111111011111010101110;
assign LUT_2[34951] = 32'b11111111111111111000110011000111;
assign LUT_2[34952] = 32'b11111111111111110011010101100111;
assign LUT_2[34953] = 32'b11111111111111110000001110000000;
assign LUT_2[34954] = 32'b11111111111111111010001110100011;
assign LUT_2[34955] = 32'b11111111111111110111000110111100;
assign LUT_2[34956] = 32'b11111111111111101111110011001111;
assign LUT_2[34957] = 32'b11111111111111101100101011101000;
assign LUT_2[34958] = 32'b11111111111111110110101100001011;
assign LUT_2[34959] = 32'b11111111111111110011100100100100;
assign LUT_2[34960] = 32'b11111111111111110011001000010100;
assign LUT_2[34961] = 32'b11111111111111110000000000101101;
assign LUT_2[34962] = 32'b11111111111111111010000001010000;
assign LUT_2[34963] = 32'b11111111111111110110111001101001;
assign LUT_2[34964] = 32'b11111111111111101111100101111100;
assign LUT_2[34965] = 32'b11111111111111101100011110010101;
assign LUT_2[34966] = 32'b11111111111111110110011110111000;
assign LUT_2[34967] = 32'b11111111111111110011010111010001;
assign LUT_2[34968] = 32'b11111111111111101101111001110001;
assign LUT_2[34969] = 32'b11111111111111101010110010001010;
assign LUT_2[34970] = 32'b11111111111111110100110010101101;
assign LUT_2[34971] = 32'b11111111111111110001101011000110;
assign LUT_2[34972] = 32'b11111111111111101010010111011001;
assign LUT_2[34973] = 32'b11111111111111100111001111110010;
assign LUT_2[34974] = 32'b11111111111111110001010000010101;
assign LUT_2[34975] = 32'b11111111111111101110001000101110;
assign LUT_2[34976] = 32'b11111111111111111000111111110011;
assign LUT_2[34977] = 32'b11111111111111110101111000001100;
assign LUT_2[34978] = 32'b11111111111111111111111000101111;
assign LUT_2[34979] = 32'b11111111111111111100110001001000;
assign LUT_2[34980] = 32'b11111111111111110101011101011011;
assign LUT_2[34981] = 32'b11111111111111110010010101110100;
assign LUT_2[34982] = 32'b11111111111111111100010110010111;
assign LUT_2[34983] = 32'b11111111111111111001001110110000;
assign LUT_2[34984] = 32'b11111111111111110011110001010000;
assign LUT_2[34985] = 32'b11111111111111110000101001101001;
assign LUT_2[34986] = 32'b11111111111111111010101010001100;
assign LUT_2[34987] = 32'b11111111111111110111100010100101;
assign LUT_2[34988] = 32'b11111111111111110000001110111000;
assign LUT_2[34989] = 32'b11111111111111101101000111010001;
assign LUT_2[34990] = 32'b11111111111111110111000111110100;
assign LUT_2[34991] = 32'b11111111111111110100000000001101;
assign LUT_2[34992] = 32'b11111111111111110011100011111101;
assign LUT_2[34993] = 32'b11111111111111110000011100010110;
assign LUT_2[34994] = 32'b11111111111111111010011100111001;
assign LUT_2[34995] = 32'b11111111111111110111010101010010;
assign LUT_2[34996] = 32'b11111111111111110000000001100101;
assign LUT_2[34997] = 32'b11111111111111101100111001111110;
assign LUT_2[34998] = 32'b11111111111111110110111010100001;
assign LUT_2[34999] = 32'b11111111111111110011110010111010;
assign LUT_2[35000] = 32'b11111111111111101110010101011010;
assign LUT_2[35001] = 32'b11111111111111101011001101110011;
assign LUT_2[35002] = 32'b11111111111111110101001110010110;
assign LUT_2[35003] = 32'b11111111111111110010000110101111;
assign LUT_2[35004] = 32'b11111111111111101010110011000010;
assign LUT_2[35005] = 32'b11111111111111100111101011011011;
assign LUT_2[35006] = 32'b11111111111111110001101011111110;
assign LUT_2[35007] = 32'b11111111111111101110100100010111;
assign LUT_2[35008] = 32'b11111111111111110000101100101101;
assign LUT_2[35009] = 32'b11111111111111101101100101000110;
assign LUT_2[35010] = 32'b11111111111111110111100101101001;
assign LUT_2[35011] = 32'b11111111111111110100011110000010;
assign LUT_2[35012] = 32'b11111111111111101101001010010101;
assign LUT_2[35013] = 32'b11111111111111101010000010101110;
assign LUT_2[35014] = 32'b11111111111111110100000011010001;
assign LUT_2[35015] = 32'b11111111111111110000111011101010;
assign LUT_2[35016] = 32'b11111111111111101011011110001010;
assign LUT_2[35017] = 32'b11111111111111101000010110100011;
assign LUT_2[35018] = 32'b11111111111111110010010111000110;
assign LUT_2[35019] = 32'b11111111111111101111001111011111;
assign LUT_2[35020] = 32'b11111111111111100111111011110010;
assign LUT_2[35021] = 32'b11111111111111100100110100001011;
assign LUT_2[35022] = 32'b11111111111111101110110100101110;
assign LUT_2[35023] = 32'b11111111111111101011101101000111;
assign LUT_2[35024] = 32'b11111111111111101011010000110111;
assign LUT_2[35025] = 32'b11111111111111101000001001010000;
assign LUT_2[35026] = 32'b11111111111111110010001001110011;
assign LUT_2[35027] = 32'b11111111111111101111000010001100;
assign LUT_2[35028] = 32'b11111111111111100111101110011111;
assign LUT_2[35029] = 32'b11111111111111100100100110111000;
assign LUT_2[35030] = 32'b11111111111111101110100111011011;
assign LUT_2[35031] = 32'b11111111111111101011011111110100;
assign LUT_2[35032] = 32'b11111111111111100110000010010100;
assign LUT_2[35033] = 32'b11111111111111100010111010101101;
assign LUT_2[35034] = 32'b11111111111111101100111011010000;
assign LUT_2[35035] = 32'b11111111111111101001110011101001;
assign LUT_2[35036] = 32'b11111111111111100010011111111100;
assign LUT_2[35037] = 32'b11111111111111011111011000010101;
assign LUT_2[35038] = 32'b11111111111111101001011000111000;
assign LUT_2[35039] = 32'b11111111111111100110010001010001;
assign LUT_2[35040] = 32'b11111111111111110001001000010110;
assign LUT_2[35041] = 32'b11111111111111101110000000101111;
assign LUT_2[35042] = 32'b11111111111111111000000001010010;
assign LUT_2[35043] = 32'b11111111111111110100111001101011;
assign LUT_2[35044] = 32'b11111111111111101101100101111110;
assign LUT_2[35045] = 32'b11111111111111101010011110010111;
assign LUT_2[35046] = 32'b11111111111111110100011110111010;
assign LUT_2[35047] = 32'b11111111111111110001010111010011;
assign LUT_2[35048] = 32'b11111111111111101011111001110011;
assign LUT_2[35049] = 32'b11111111111111101000110010001100;
assign LUT_2[35050] = 32'b11111111111111110010110010101111;
assign LUT_2[35051] = 32'b11111111111111101111101011001000;
assign LUT_2[35052] = 32'b11111111111111101000010111011011;
assign LUT_2[35053] = 32'b11111111111111100101001111110100;
assign LUT_2[35054] = 32'b11111111111111101111010000010111;
assign LUT_2[35055] = 32'b11111111111111101100001000110000;
assign LUT_2[35056] = 32'b11111111111111101011101100100000;
assign LUT_2[35057] = 32'b11111111111111101000100100111001;
assign LUT_2[35058] = 32'b11111111111111110010100101011100;
assign LUT_2[35059] = 32'b11111111111111101111011101110101;
assign LUT_2[35060] = 32'b11111111111111101000001010001000;
assign LUT_2[35061] = 32'b11111111111111100101000010100001;
assign LUT_2[35062] = 32'b11111111111111101111000011000100;
assign LUT_2[35063] = 32'b11111111111111101011111011011101;
assign LUT_2[35064] = 32'b11111111111111100110011101111101;
assign LUT_2[35065] = 32'b11111111111111100011010110010110;
assign LUT_2[35066] = 32'b11111111111111101101010110111001;
assign LUT_2[35067] = 32'b11111111111111101010001111010010;
assign LUT_2[35068] = 32'b11111111111111100010111011100101;
assign LUT_2[35069] = 32'b11111111111111011111110011111110;
assign LUT_2[35070] = 32'b11111111111111101001110100100001;
assign LUT_2[35071] = 32'b11111111111111100110101100111010;
assign LUT_2[35072] = 32'b11111111111111111000001110100001;
assign LUT_2[35073] = 32'b11111111111111110101000110111010;
assign LUT_2[35074] = 32'b11111111111111111111000111011101;
assign LUT_2[35075] = 32'b11111111111111111011111111110110;
assign LUT_2[35076] = 32'b11111111111111110100101100001001;
assign LUT_2[35077] = 32'b11111111111111110001100100100010;
assign LUT_2[35078] = 32'b11111111111111111011100101000101;
assign LUT_2[35079] = 32'b11111111111111111000011101011110;
assign LUT_2[35080] = 32'b11111111111111110010111111111110;
assign LUT_2[35081] = 32'b11111111111111101111111000010111;
assign LUT_2[35082] = 32'b11111111111111111001111000111010;
assign LUT_2[35083] = 32'b11111111111111110110110001010011;
assign LUT_2[35084] = 32'b11111111111111101111011101100110;
assign LUT_2[35085] = 32'b11111111111111101100010101111111;
assign LUT_2[35086] = 32'b11111111111111110110010110100010;
assign LUT_2[35087] = 32'b11111111111111110011001110111011;
assign LUT_2[35088] = 32'b11111111111111110010110010101011;
assign LUT_2[35089] = 32'b11111111111111101111101011000100;
assign LUT_2[35090] = 32'b11111111111111111001101011100111;
assign LUT_2[35091] = 32'b11111111111111110110100100000000;
assign LUT_2[35092] = 32'b11111111111111101111010000010011;
assign LUT_2[35093] = 32'b11111111111111101100001000101100;
assign LUT_2[35094] = 32'b11111111111111110110001001001111;
assign LUT_2[35095] = 32'b11111111111111110011000001101000;
assign LUT_2[35096] = 32'b11111111111111101101100100001000;
assign LUT_2[35097] = 32'b11111111111111101010011100100001;
assign LUT_2[35098] = 32'b11111111111111110100011101000100;
assign LUT_2[35099] = 32'b11111111111111110001010101011101;
assign LUT_2[35100] = 32'b11111111111111101010000001110000;
assign LUT_2[35101] = 32'b11111111111111100110111010001001;
assign LUT_2[35102] = 32'b11111111111111110000111010101100;
assign LUT_2[35103] = 32'b11111111111111101101110011000101;
assign LUT_2[35104] = 32'b11111111111111111000101010001010;
assign LUT_2[35105] = 32'b11111111111111110101100010100011;
assign LUT_2[35106] = 32'b11111111111111111111100011000110;
assign LUT_2[35107] = 32'b11111111111111111100011011011111;
assign LUT_2[35108] = 32'b11111111111111110101000111110010;
assign LUT_2[35109] = 32'b11111111111111110010000000001011;
assign LUT_2[35110] = 32'b11111111111111111100000000101110;
assign LUT_2[35111] = 32'b11111111111111111000111001000111;
assign LUT_2[35112] = 32'b11111111111111110011011011100111;
assign LUT_2[35113] = 32'b11111111111111110000010100000000;
assign LUT_2[35114] = 32'b11111111111111111010010100100011;
assign LUT_2[35115] = 32'b11111111111111110111001100111100;
assign LUT_2[35116] = 32'b11111111111111101111111001001111;
assign LUT_2[35117] = 32'b11111111111111101100110001101000;
assign LUT_2[35118] = 32'b11111111111111110110110010001011;
assign LUT_2[35119] = 32'b11111111111111110011101010100100;
assign LUT_2[35120] = 32'b11111111111111110011001110010100;
assign LUT_2[35121] = 32'b11111111111111110000000110101101;
assign LUT_2[35122] = 32'b11111111111111111010000111010000;
assign LUT_2[35123] = 32'b11111111111111110110111111101001;
assign LUT_2[35124] = 32'b11111111111111101111101011111100;
assign LUT_2[35125] = 32'b11111111111111101100100100010101;
assign LUT_2[35126] = 32'b11111111111111110110100100111000;
assign LUT_2[35127] = 32'b11111111111111110011011101010001;
assign LUT_2[35128] = 32'b11111111111111101101111111110001;
assign LUT_2[35129] = 32'b11111111111111101010111000001010;
assign LUT_2[35130] = 32'b11111111111111110100111000101101;
assign LUT_2[35131] = 32'b11111111111111110001110001000110;
assign LUT_2[35132] = 32'b11111111111111101010011101011001;
assign LUT_2[35133] = 32'b11111111111111100111010101110010;
assign LUT_2[35134] = 32'b11111111111111110001010110010101;
assign LUT_2[35135] = 32'b11111111111111101110001110101110;
assign LUT_2[35136] = 32'b11111111111111110000010111000100;
assign LUT_2[35137] = 32'b11111111111111101101001111011101;
assign LUT_2[35138] = 32'b11111111111111110111010000000000;
assign LUT_2[35139] = 32'b11111111111111110100001000011001;
assign LUT_2[35140] = 32'b11111111111111101100110100101100;
assign LUT_2[35141] = 32'b11111111111111101001101101000101;
assign LUT_2[35142] = 32'b11111111111111110011101101101000;
assign LUT_2[35143] = 32'b11111111111111110000100110000001;
assign LUT_2[35144] = 32'b11111111111111101011001000100001;
assign LUT_2[35145] = 32'b11111111111111101000000000111010;
assign LUT_2[35146] = 32'b11111111111111110010000001011101;
assign LUT_2[35147] = 32'b11111111111111101110111001110110;
assign LUT_2[35148] = 32'b11111111111111100111100110001001;
assign LUT_2[35149] = 32'b11111111111111100100011110100010;
assign LUT_2[35150] = 32'b11111111111111101110011111000101;
assign LUT_2[35151] = 32'b11111111111111101011010111011110;
assign LUT_2[35152] = 32'b11111111111111101010111011001110;
assign LUT_2[35153] = 32'b11111111111111100111110011100111;
assign LUT_2[35154] = 32'b11111111111111110001110100001010;
assign LUT_2[35155] = 32'b11111111111111101110101100100011;
assign LUT_2[35156] = 32'b11111111111111100111011000110110;
assign LUT_2[35157] = 32'b11111111111111100100010001001111;
assign LUT_2[35158] = 32'b11111111111111101110010001110010;
assign LUT_2[35159] = 32'b11111111111111101011001010001011;
assign LUT_2[35160] = 32'b11111111111111100101101100101011;
assign LUT_2[35161] = 32'b11111111111111100010100101000100;
assign LUT_2[35162] = 32'b11111111111111101100100101100111;
assign LUT_2[35163] = 32'b11111111111111101001011110000000;
assign LUT_2[35164] = 32'b11111111111111100010001010010011;
assign LUT_2[35165] = 32'b11111111111111011111000010101100;
assign LUT_2[35166] = 32'b11111111111111101001000011001111;
assign LUT_2[35167] = 32'b11111111111111100101111011101000;
assign LUT_2[35168] = 32'b11111111111111110000110010101101;
assign LUT_2[35169] = 32'b11111111111111101101101011000110;
assign LUT_2[35170] = 32'b11111111111111110111101011101001;
assign LUT_2[35171] = 32'b11111111111111110100100100000010;
assign LUT_2[35172] = 32'b11111111111111101101010000010101;
assign LUT_2[35173] = 32'b11111111111111101010001000101110;
assign LUT_2[35174] = 32'b11111111111111110100001001010001;
assign LUT_2[35175] = 32'b11111111111111110001000001101010;
assign LUT_2[35176] = 32'b11111111111111101011100100001010;
assign LUT_2[35177] = 32'b11111111111111101000011100100011;
assign LUT_2[35178] = 32'b11111111111111110010011101000110;
assign LUT_2[35179] = 32'b11111111111111101111010101011111;
assign LUT_2[35180] = 32'b11111111111111101000000001110010;
assign LUT_2[35181] = 32'b11111111111111100100111010001011;
assign LUT_2[35182] = 32'b11111111111111101110111010101110;
assign LUT_2[35183] = 32'b11111111111111101011110011000111;
assign LUT_2[35184] = 32'b11111111111111101011010110110111;
assign LUT_2[35185] = 32'b11111111111111101000001111010000;
assign LUT_2[35186] = 32'b11111111111111110010001111110011;
assign LUT_2[35187] = 32'b11111111111111101111001000001100;
assign LUT_2[35188] = 32'b11111111111111100111110100011111;
assign LUT_2[35189] = 32'b11111111111111100100101100111000;
assign LUT_2[35190] = 32'b11111111111111101110101101011011;
assign LUT_2[35191] = 32'b11111111111111101011100101110100;
assign LUT_2[35192] = 32'b11111111111111100110001000010100;
assign LUT_2[35193] = 32'b11111111111111100011000000101101;
assign LUT_2[35194] = 32'b11111111111111101101000001010000;
assign LUT_2[35195] = 32'b11111111111111101001111001101001;
assign LUT_2[35196] = 32'b11111111111111100010100101111100;
assign LUT_2[35197] = 32'b11111111111111011111011110010101;
assign LUT_2[35198] = 32'b11111111111111101001011110111000;
assign LUT_2[35199] = 32'b11111111111111100110010111010001;
assign LUT_2[35200] = 32'b11111111111111111100100010110000;
assign LUT_2[35201] = 32'b11111111111111111001011011001001;
assign LUT_2[35202] = 32'b00000000000000000011011011101100;
assign LUT_2[35203] = 32'b00000000000000000000010100000101;
assign LUT_2[35204] = 32'b11111111111111111001000000011000;
assign LUT_2[35205] = 32'b11111111111111110101111000110001;
assign LUT_2[35206] = 32'b11111111111111111111111001010100;
assign LUT_2[35207] = 32'b11111111111111111100110001101101;
assign LUT_2[35208] = 32'b11111111111111110111010100001101;
assign LUT_2[35209] = 32'b11111111111111110100001100100110;
assign LUT_2[35210] = 32'b11111111111111111110001101001001;
assign LUT_2[35211] = 32'b11111111111111111011000101100010;
assign LUT_2[35212] = 32'b11111111111111110011110001110101;
assign LUT_2[35213] = 32'b11111111111111110000101010001110;
assign LUT_2[35214] = 32'b11111111111111111010101010110001;
assign LUT_2[35215] = 32'b11111111111111110111100011001010;
assign LUT_2[35216] = 32'b11111111111111110111000110111010;
assign LUT_2[35217] = 32'b11111111111111110011111111010011;
assign LUT_2[35218] = 32'b11111111111111111101111111110110;
assign LUT_2[35219] = 32'b11111111111111111010111000001111;
assign LUT_2[35220] = 32'b11111111111111110011100100100010;
assign LUT_2[35221] = 32'b11111111111111110000011100111011;
assign LUT_2[35222] = 32'b11111111111111111010011101011110;
assign LUT_2[35223] = 32'b11111111111111110111010101110111;
assign LUT_2[35224] = 32'b11111111111111110001111000010111;
assign LUT_2[35225] = 32'b11111111111111101110110000110000;
assign LUT_2[35226] = 32'b11111111111111111000110001010011;
assign LUT_2[35227] = 32'b11111111111111110101101001101100;
assign LUT_2[35228] = 32'b11111111111111101110010101111111;
assign LUT_2[35229] = 32'b11111111111111101011001110011000;
assign LUT_2[35230] = 32'b11111111111111110101001110111011;
assign LUT_2[35231] = 32'b11111111111111110010000111010100;
assign LUT_2[35232] = 32'b11111111111111111100111110011001;
assign LUT_2[35233] = 32'b11111111111111111001110110110010;
assign LUT_2[35234] = 32'b00000000000000000011110111010101;
assign LUT_2[35235] = 32'b00000000000000000000101111101110;
assign LUT_2[35236] = 32'b11111111111111111001011100000001;
assign LUT_2[35237] = 32'b11111111111111110110010100011010;
assign LUT_2[35238] = 32'b00000000000000000000010100111101;
assign LUT_2[35239] = 32'b11111111111111111101001101010110;
assign LUT_2[35240] = 32'b11111111111111110111101111110110;
assign LUT_2[35241] = 32'b11111111111111110100101000001111;
assign LUT_2[35242] = 32'b11111111111111111110101000110010;
assign LUT_2[35243] = 32'b11111111111111111011100001001011;
assign LUT_2[35244] = 32'b11111111111111110100001101011110;
assign LUT_2[35245] = 32'b11111111111111110001000101110111;
assign LUT_2[35246] = 32'b11111111111111111011000110011010;
assign LUT_2[35247] = 32'b11111111111111110111111110110011;
assign LUT_2[35248] = 32'b11111111111111110111100010100011;
assign LUT_2[35249] = 32'b11111111111111110100011010111100;
assign LUT_2[35250] = 32'b11111111111111111110011011011111;
assign LUT_2[35251] = 32'b11111111111111111011010011111000;
assign LUT_2[35252] = 32'b11111111111111110100000000001011;
assign LUT_2[35253] = 32'b11111111111111110000111000100100;
assign LUT_2[35254] = 32'b11111111111111111010111001000111;
assign LUT_2[35255] = 32'b11111111111111110111110001100000;
assign LUT_2[35256] = 32'b11111111111111110010010100000000;
assign LUT_2[35257] = 32'b11111111111111101111001100011001;
assign LUT_2[35258] = 32'b11111111111111111001001100111100;
assign LUT_2[35259] = 32'b11111111111111110110000101010101;
assign LUT_2[35260] = 32'b11111111111111101110110001101000;
assign LUT_2[35261] = 32'b11111111111111101011101010000001;
assign LUT_2[35262] = 32'b11111111111111110101101010100100;
assign LUT_2[35263] = 32'b11111111111111110010100010111101;
assign LUT_2[35264] = 32'b11111111111111110100101011010011;
assign LUT_2[35265] = 32'b11111111111111110001100011101100;
assign LUT_2[35266] = 32'b11111111111111111011100100001111;
assign LUT_2[35267] = 32'b11111111111111111000011100101000;
assign LUT_2[35268] = 32'b11111111111111110001001000111011;
assign LUT_2[35269] = 32'b11111111111111101110000001010100;
assign LUT_2[35270] = 32'b11111111111111111000000001110111;
assign LUT_2[35271] = 32'b11111111111111110100111010010000;
assign LUT_2[35272] = 32'b11111111111111101111011100110000;
assign LUT_2[35273] = 32'b11111111111111101100010101001001;
assign LUT_2[35274] = 32'b11111111111111110110010101101100;
assign LUT_2[35275] = 32'b11111111111111110011001110000101;
assign LUT_2[35276] = 32'b11111111111111101011111010011000;
assign LUT_2[35277] = 32'b11111111111111101000110010110001;
assign LUT_2[35278] = 32'b11111111111111110010110011010100;
assign LUT_2[35279] = 32'b11111111111111101111101011101101;
assign LUT_2[35280] = 32'b11111111111111101111001111011101;
assign LUT_2[35281] = 32'b11111111111111101100000111110110;
assign LUT_2[35282] = 32'b11111111111111110110001000011001;
assign LUT_2[35283] = 32'b11111111111111110011000000110010;
assign LUT_2[35284] = 32'b11111111111111101011101101000101;
assign LUT_2[35285] = 32'b11111111111111101000100101011110;
assign LUT_2[35286] = 32'b11111111111111110010100110000001;
assign LUT_2[35287] = 32'b11111111111111101111011110011010;
assign LUT_2[35288] = 32'b11111111111111101010000000111010;
assign LUT_2[35289] = 32'b11111111111111100110111001010011;
assign LUT_2[35290] = 32'b11111111111111110000111001110110;
assign LUT_2[35291] = 32'b11111111111111101101110010001111;
assign LUT_2[35292] = 32'b11111111111111100110011110100010;
assign LUT_2[35293] = 32'b11111111111111100011010110111011;
assign LUT_2[35294] = 32'b11111111111111101101010111011110;
assign LUT_2[35295] = 32'b11111111111111101010001111110111;
assign LUT_2[35296] = 32'b11111111111111110101000110111100;
assign LUT_2[35297] = 32'b11111111111111110001111111010101;
assign LUT_2[35298] = 32'b11111111111111111011111111111000;
assign LUT_2[35299] = 32'b11111111111111111000111000010001;
assign LUT_2[35300] = 32'b11111111111111110001100100100100;
assign LUT_2[35301] = 32'b11111111111111101110011100111101;
assign LUT_2[35302] = 32'b11111111111111111000011101100000;
assign LUT_2[35303] = 32'b11111111111111110101010101111001;
assign LUT_2[35304] = 32'b11111111111111101111111000011001;
assign LUT_2[35305] = 32'b11111111111111101100110000110010;
assign LUT_2[35306] = 32'b11111111111111110110110001010101;
assign LUT_2[35307] = 32'b11111111111111110011101001101110;
assign LUT_2[35308] = 32'b11111111111111101100010110000001;
assign LUT_2[35309] = 32'b11111111111111101001001110011010;
assign LUT_2[35310] = 32'b11111111111111110011001110111101;
assign LUT_2[35311] = 32'b11111111111111110000000111010110;
assign LUT_2[35312] = 32'b11111111111111101111101011000110;
assign LUT_2[35313] = 32'b11111111111111101100100011011111;
assign LUT_2[35314] = 32'b11111111111111110110100100000010;
assign LUT_2[35315] = 32'b11111111111111110011011100011011;
assign LUT_2[35316] = 32'b11111111111111101100001000101110;
assign LUT_2[35317] = 32'b11111111111111101001000001000111;
assign LUT_2[35318] = 32'b11111111111111110011000001101010;
assign LUT_2[35319] = 32'b11111111111111101111111010000011;
assign LUT_2[35320] = 32'b11111111111111101010011100100011;
assign LUT_2[35321] = 32'b11111111111111100111010100111100;
assign LUT_2[35322] = 32'b11111111111111110001010101011111;
assign LUT_2[35323] = 32'b11111111111111101110001101111000;
assign LUT_2[35324] = 32'b11111111111111100110111010001011;
assign LUT_2[35325] = 32'b11111111111111100011110010100100;
assign LUT_2[35326] = 32'b11111111111111101101110011000111;
assign LUT_2[35327] = 32'b11111111111111101010101011100000;
assign LUT_2[35328] = 32'b11111111111111111001000001101101;
assign LUT_2[35329] = 32'b11111111111111110101111010000110;
assign LUT_2[35330] = 32'b11111111111111111111111010101001;
assign LUT_2[35331] = 32'b11111111111111111100110011000010;
assign LUT_2[35332] = 32'b11111111111111110101011111010101;
assign LUT_2[35333] = 32'b11111111111111110010010111101110;
assign LUT_2[35334] = 32'b11111111111111111100011000010001;
assign LUT_2[35335] = 32'b11111111111111111001010000101010;
assign LUT_2[35336] = 32'b11111111111111110011110011001010;
assign LUT_2[35337] = 32'b11111111111111110000101011100011;
assign LUT_2[35338] = 32'b11111111111111111010101100000110;
assign LUT_2[35339] = 32'b11111111111111110111100100011111;
assign LUT_2[35340] = 32'b11111111111111110000010000110010;
assign LUT_2[35341] = 32'b11111111111111101101001001001011;
assign LUT_2[35342] = 32'b11111111111111110111001001101110;
assign LUT_2[35343] = 32'b11111111111111110100000010000111;
assign LUT_2[35344] = 32'b11111111111111110011100101110111;
assign LUT_2[35345] = 32'b11111111111111110000011110010000;
assign LUT_2[35346] = 32'b11111111111111111010011110110011;
assign LUT_2[35347] = 32'b11111111111111110111010111001100;
assign LUT_2[35348] = 32'b11111111111111110000000011011111;
assign LUT_2[35349] = 32'b11111111111111101100111011111000;
assign LUT_2[35350] = 32'b11111111111111110110111100011011;
assign LUT_2[35351] = 32'b11111111111111110011110100110100;
assign LUT_2[35352] = 32'b11111111111111101110010111010100;
assign LUT_2[35353] = 32'b11111111111111101011001111101101;
assign LUT_2[35354] = 32'b11111111111111110101010000010000;
assign LUT_2[35355] = 32'b11111111111111110010001000101001;
assign LUT_2[35356] = 32'b11111111111111101010110100111100;
assign LUT_2[35357] = 32'b11111111111111100111101101010101;
assign LUT_2[35358] = 32'b11111111111111110001101101111000;
assign LUT_2[35359] = 32'b11111111111111101110100110010001;
assign LUT_2[35360] = 32'b11111111111111111001011101010110;
assign LUT_2[35361] = 32'b11111111111111110110010101101111;
assign LUT_2[35362] = 32'b00000000000000000000010110010010;
assign LUT_2[35363] = 32'b11111111111111111101001110101011;
assign LUT_2[35364] = 32'b11111111111111110101111010111110;
assign LUT_2[35365] = 32'b11111111111111110010110011010111;
assign LUT_2[35366] = 32'b11111111111111111100110011111010;
assign LUT_2[35367] = 32'b11111111111111111001101100010011;
assign LUT_2[35368] = 32'b11111111111111110100001110110011;
assign LUT_2[35369] = 32'b11111111111111110001000111001100;
assign LUT_2[35370] = 32'b11111111111111111011000111101111;
assign LUT_2[35371] = 32'b11111111111111111000000000001000;
assign LUT_2[35372] = 32'b11111111111111110000101100011011;
assign LUT_2[35373] = 32'b11111111111111101101100100110100;
assign LUT_2[35374] = 32'b11111111111111110111100101010111;
assign LUT_2[35375] = 32'b11111111111111110100011101110000;
assign LUT_2[35376] = 32'b11111111111111110100000001100000;
assign LUT_2[35377] = 32'b11111111111111110000111001111001;
assign LUT_2[35378] = 32'b11111111111111111010111010011100;
assign LUT_2[35379] = 32'b11111111111111110111110010110101;
assign LUT_2[35380] = 32'b11111111111111110000011111001000;
assign LUT_2[35381] = 32'b11111111111111101101010111100001;
assign LUT_2[35382] = 32'b11111111111111110111011000000100;
assign LUT_2[35383] = 32'b11111111111111110100010000011101;
assign LUT_2[35384] = 32'b11111111111111101110110010111101;
assign LUT_2[35385] = 32'b11111111111111101011101011010110;
assign LUT_2[35386] = 32'b11111111111111110101101011111001;
assign LUT_2[35387] = 32'b11111111111111110010100100010010;
assign LUT_2[35388] = 32'b11111111111111101011010000100101;
assign LUT_2[35389] = 32'b11111111111111101000001000111110;
assign LUT_2[35390] = 32'b11111111111111110010001001100001;
assign LUT_2[35391] = 32'b11111111111111101111000001111010;
assign LUT_2[35392] = 32'b11111111111111110001001010010000;
assign LUT_2[35393] = 32'b11111111111111101110000010101001;
assign LUT_2[35394] = 32'b11111111111111111000000011001100;
assign LUT_2[35395] = 32'b11111111111111110100111011100101;
assign LUT_2[35396] = 32'b11111111111111101101100111111000;
assign LUT_2[35397] = 32'b11111111111111101010100000010001;
assign LUT_2[35398] = 32'b11111111111111110100100000110100;
assign LUT_2[35399] = 32'b11111111111111110001011001001101;
assign LUT_2[35400] = 32'b11111111111111101011111011101101;
assign LUT_2[35401] = 32'b11111111111111101000110100000110;
assign LUT_2[35402] = 32'b11111111111111110010110100101001;
assign LUT_2[35403] = 32'b11111111111111101111101101000010;
assign LUT_2[35404] = 32'b11111111111111101000011001010101;
assign LUT_2[35405] = 32'b11111111111111100101010001101110;
assign LUT_2[35406] = 32'b11111111111111101111010010010001;
assign LUT_2[35407] = 32'b11111111111111101100001010101010;
assign LUT_2[35408] = 32'b11111111111111101011101110011010;
assign LUT_2[35409] = 32'b11111111111111101000100110110011;
assign LUT_2[35410] = 32'b11111111111111110010100111010110;
assign LUT_2[35411] = 32'b11111111111111101111011111101111;
assign LUT_2[35412] = 32'b11111111111111101000001100000010;
assign LUT_2[35413] = 32'b11111111111111100101000100011011;
assign LUT_2[35414] = 32'b11111111111111101111000100111110;
assign LUT_2[35415] = 32'b11111111111111101011111101010111;
assign LUT_2[35416] = 32'b11111111111111100110011111110111;
assign LUT_2[35417] = 32'b11111111111111100011011000010000;
assign LUT_2[35418] = 32'b11111111111111101101011000110011;
assign LUT_2[35419] = 32'b11111111111111101010010001001100;
assign LUT_2[35420] = 32'b11111111111111100010111101011111;
assign LUT_2[35421] = 32'b11111111111111011111110101111000;
assign LUT_2[35422] = 32'b11111111111111101001110110011011;
assign LUT_2[35423] = 32'b11111111111111100110101110110100;
assign LUT_2[35424] = 32'b11111111111111110001100101111001;
assign LUT_2[35425] = 32'b11111111111111101110011110010010;
assign LUT_2[35426] = 32'b11111111111111111000011110110101;
assign LUT_2[35427] = 32'b11111111111111110101010111001110;
assign LUT_2[35428] = 32'b11111111111111101110000011100001;
assign LUT_2[35429] = 32'b11111111111111101010111011111010;
assign LUT_2[35430] = 32'b11111111111111110100111100011101;
assign LUT_2[35431] = 32'b11111111111111110001110100110110;
assign LUT_2[35432] = 32'b11111111111111101100010111010110;
assign LUT_2[35433] = 32'b11111111111111101001001111101111;
assign LUT_2[35434] = 32'b11111111111111110011010000010010;
assign LUT_2[35435] = 32'b11111111111111110000001000101011;
assign LUT_2[35436] = 32'b11111111111111101000110100111110;
assign LUT_2[35437] = 32'b11111111111111100101101101010111;
assign LUT_2[35438] = 32'b11111111111111101111101101111010;
assign LUT_2[35439] = 32'b11111111111111101100100110010011;
assign LUT_2[35440] = 32'b11111111111111101100001010000011;
assign LUT_2[35441] = 32'b11111111111111101001000010011100;
assign LUT_2[35442] = 32'b11111111111111110011000010111111;
assign LUT_2[35443] = 32'b11111111111111101111111011011000;
assign LUT_2[35444] = 32'b11111111111111101000100111101011;
assign LUT_2[35445] = 32'b11111111111111100101100000000100;
assign LUT_2[35446] = 32'b11111111111111101111100000100111;
assign LUT_2[35447] = 32'b11111111111111101100011001000000;
assign LUT_2[35448] = 32'b11111111111111100110111011100000;
assign LUT_2[35449] = 32'b11111111111111100011110011111001;
assign LUT_2[35450] = 32'b11111111111111101101110100011100;
assign LUT_2[35451] = 32'b11111111111111101010101100110101;
assign LUT_2[35452] = 32'b11111111111111100011011001001000;
assign LUT_2[35453] = 32'b11111111111111100000010001100001;
assign LUT_2[35454] = 32'b11111111111111101010010010000100;
assign LUT_2[35455] = 32'b11111111111111100111001010011101;
assign LUT_2[35456] = 32'b11111111111111111101010101111100;
assign LUT_2[35457] = 32'b11111111111111111010001110010101;
assign LUT_2[35458] = 32'b00000000000000000100001110111000;
assign LUT_2[35459] = 32'b00000000000000000001000111010001;
assign LUT_2[35460] = 32'b11111111111111111001110011100100;
assign LUT_2[35461] = 32'b11111111111111110110101011111101;
assign LUT_2[35462] = 32'b00000000000000000000101100100000;
assign LUT_2[35463] = 32'b11111111111111111101100100111001;
assign LUT_2[35464] = 32'b11111111111111111000000111011001;
assign LUT_2[35465] = 32'b11111111111111110100111111110010;
assign LUT_2[35466] = 32'b11111111111111111111000000010101;
assign LUT_2[35467] = 32'b11111111111111111011111000101110;
assign LUT_2[35468] = 32'b11111111111111110100100101000001;
assign LUT_2[35469] = 32'b11111111111111110001011101011010;
assign LUT_2[35470] = 32'b11111111111111111011011101111101;
assign LUT_2[35471] = 32'b11111111111111111000010110010110;
assign LUT_2[35472] = 32'b11111111111111110111111010000110;
assign LUT_2[35473] = 32'b11111111111111110100110010011111;
assign LUT_2[35474] = 32'b11111111111111111110110011000010;
assign LUT_2[35475] = 32'b11111111111111111011101011011011;
assign LUT_2[35476] = 32'b11111111111111110100010111101110;
assign LUT_2[35477] = 32'b11111111111111110001010000000111;
assign LUT_2[35478] = 32'b11111111111111111011010000101010;
assign LUT_2[35479] = 32'b11111111111111111000001001000011;
assign LUT_2[35480] = 32'b11111111111111110010101011100011;
assign LUT_2[35481] = 32'b11111111111111101111100011111100;
assign LUT_2[35482] = 32'b11111111111111111001100100011111;
assign LUT_2[35483] = 32'b11111111111111110110011100111000;
assign LUT_2[35484] = 32'b11111111111111101111001001001011;
assign LUT_2[35485] = 32'b11111111111111101100000001100100;
assign LUT_2[35486] = 32'b11111111111111110110000010000111;
assign LUT_2[35487] = 32'b11111111111111110010111010100000;
assign LUT_2[35488] = 32'b11111111111111111101110001100101;
assign LUT_2[35489] = 32'b11111111111111111010101001111110;
assign LUT_2[35490] = 32'b00000000000000000100101010100001;
assign LUT_2[35491] = 32'b00000000000000000001100010111010;
assign LUT_2[35492] = 32'b11111111111111111010001111001101;
assign LUT_2[35493] = 32'b11111111111111110111000111100110;
assign LUT_2[35494] = 32'b00000000000000000001001000001001;
assign LUT_2[35495] = 32'b11111111111111111110000000100010;
assign LUT_2[35496] = 32'b11111111111111111000100011000010;
assign LUT_2[35497] = 32'b11111111111111110101011011011011;
assign LUT_2[35498] = 32'b11111111111111111111011011111110;
assign LUT_2[35499] = 32'b11111111111111111100010100010111;
assign LUT_2[35500] = 32'b11111111111111110101000000101010;
assign LUT_2[35501] = 32'b11111111111111110001111001000011;
assign LUT_2[35502] = 32'b11111111111111111011111001100110;
assign LUT_2[35503] = 32'b11111111111111111000110001111111;
assign LUT_2[35504] = 32'b11111111111111111000010101101111;
assign LUT_2[35505] = 32'b11111111111111110101001110001000;
assign LUT_2[35506] = 32'b11111111111111111111001110101011;
assign LUT_2[35507] = 32'b11111111111111111100000111000100;
assign LUT_2[35508] = 32'b11111111111111110100110011010111;
assign LUT_2[35509] = 32'b11111111111111110001101011110000;
assign LUT_2[35510] = 32'b11111111111111111011101100010011;
assign LUT_2[35511] = 32'b11111111111111111000100100101100;
assign LUT_2[35512] = 32'b11111111111111110011000111001100;
assign LUT_2[35513] = 32'b11111111111111101111111111100101;
assign LUT_2[35514] = 32'b11111111111111111010000000001000;
assign LUT_2[35515] = 32'b11111111111111110110111000100001;
assign LUT_2[35516] = 32'b11111111111111101111100100110100;
assign LUT_2[35517] = 32'b11111111111111101100011101001101;
assign LUT_2[35518] = 32'b11111111111111110110011101110000;
assign LUT_2[35519] = 32'b11111111111111110011010110001001;
assign LUT_2[35520] = 32'b11111111111111110101011110011111;
assign LUT_2[35521] = 32'b11111111111111110010010110111000;
assign LUT_2[35522] = 32'b11111111111111111100010111011011;
assign LUT_2[35523] = 32'b11111111111111111001001111110100;
assign LUT_2[35524] = 32'b11111111111111110001111100000111;
assign LUT_2[35525] = 32'b11111111111111101110110100100000;
assign LUT_2[35526] = 32'b11111111111111111000110101000011;
assign LUT_2[35527] = 32'b11111111111111110101101101011100;
assign LUT_2[35528] = 32'b11111111111111110000001111111100;
assign LUT_2[35529] = 32'b11111111111111101101001000010101;
assign LUT_2[35530] = 32'b11111111111111110111001000111000;
assign LUT_2[35531] = 32'b11111111111111110100000001010001;
assign LUT_2[35532] = 32'b11111111111111101100101101100100;
assign LUT_2[35533] = 32'b11111111111111101001100101111101;
assign LUT_2[35534] = 32'b11111111111111110011100110100000;
assign LUT_2[35535] = 32'b11111111111111110000011110111001;
assign LUT_2[35536] = 32'b11111111111111110000000010101001;
assign LUT_2[35537] = 32'b11111111111111101100111011000010;
assign LUT_2[35538] = 32'b11111111111111110110111011100101;
assign LUT_2[35539] = 32'b11111111111111110011110011111110;
assign LUT_2[35540] = 32'b11111111111111101100100000010001;
assign LUT_2[35541] = 32'b11111111111111101001011000101010;
assign LUT_2[35542] = 32'b11111111111111110011011001001101;
assign LUT_2[35543] = 32'b11111111111111110000010001100110;
assign LUT_2[35544] = 32'b11111111111111101010110100000110;
assign LUT_2[35545] = 32'b11111111111111100111101100011111;
assign LUT_2[35546] = 32'b11111111111111110001101101000010;
assign LUT_2[35547] = 32'b11111111111111101110100101011011;
assign LUT_2[35548] = 32'b11111111111111100111010001101110;
assign LUT_2[35549] = 32'b11111111111111100100001010000111;
assign LUT_2[35550] = 32'b11111111111111101110001010101010;
assign LUT_2[35551] = 32'b11111111111111101011000011000011;
assign LUT_2[35552] = 32'b11111111111111110101111010001000;
assign LUT_2[35553] = 32'b11111111111111110010110010100001;
assign LUT_2[35554] = 32'b11111111111111111100110011000100;
assign LUT_2[35555] = 32'b11111111111111111001101011011101;
assign LUT_2[35556] = 32'b11111111111111110010010111110000;
assign LUT_2[35557] = 32'b11111111111111101111010000001001;
assign LUT_2[35558] = 32'b11111111111111111001010000101100;
assign LUT_2[35559] = 32'b11111111111111110110001001000101;
assign LUT_2[35560] = 32'b11111111111111110000101011100101;
assign LUT_2[35561] = 32'b11111111111111101101100011111110;
assign LUT_2[35562] = 32'b11111111111111110111100100100001;
assign LUT_2[35563] = 32'b11111111111111110100011100111010;
assign LUT_2[35564] = 32'b11111111111111101101001001001101;
assign LUT_2[35565] = 32'b11111111111111101010000001100110;
assign LUT_2[35566] = 32'b11111111111111110100000010001001;
assign LUT_2[35567] = 32'b11111111111111110000111010100010;
assign LUT_2[35568] = 32'b11111111111111110000011110010010;
assign LUT_2[35569] = 32'b11111111111111101101010110101011;
assign LUT_2[35570] = 32'b11111111111111110111010111001110;
assign LUT_2[35571] = 32'b11111111111111110100001111100111;
assign LUT_2[35572] = 32'b11111111111111101100111011111010;
assign LUT_2[35573] = 32'b11111111111111101001110100010011;
assign LUT_2[35574] = 32'b11111111111111110011110100110110;
assign LUT_2[35575] = 32'b11111111111111110000101101001111;
assign LUT_2[35576] = 32'b11111111111111101011001111101111;
assign LUT_2[35577] = 32'b11111111111111101000001000001000;
assign LUT_2[35578] = 32'b11111111111111110010001000101011;
assign LUT_2[35579] = 32'b11111111111111101111000001000100;
assign LUT_2[35580] = 32'b11111111111111100111101101010111;
assign LUT_2[35581] = 32'b11111111111111100100100101110000;
assign LUT_2[35582] = 32'b11111111111111101110100110010011;
assign LUT_2[35583] = 32'b11111111111111101011011110101100;
assign LUT_2[35584] = 32'b11111111111111111101000000010011;
assign LUT_2[35585] = 32'b11111111111111111001111000101100;
assign LUT_2[35586] = 32'b00000000000000000011111001001111;
assign LUT_2[35587] = 32'b00000000000000000000110001101000;
assign LUT_2[35588] = 32'b11111111111111111001011101111011;
assign LUT_2[35589] = 32'b11111111111111110110010110010100;
assign LUT_2[35590] = 32'b00000000000000000000010110110111;
assign LUT_2[35591] = 32'b11111111111111111101001111010000;
assign LUT_2[35592] = 32'b11111111111111110111110001110000;
assign LUT_2[35593] = 32'b11111111111111110100101010001001;
assign LUT_2[35594] = 32'b11111111111111111110101010101100;
assign LUT_2[35595] = 32'b11111111111111111011100011000101;
assign LUT_2[35596] = 32'b11111111111111110100001111011000;
assign LUT_2[35597] = 32'b11111111111111110001000111110001;
assign LUT_2[35598] = 32'b11111111111111111011001000010100;
assign LUT_2[35599] = 32'b11111111111111111000000000101101;
assign LUT_2[35600] = 32'b11111111111111110111100100011101;
assign LUT_2[35601] = 32'b11111111111111110100011100110110;
assign LUT_2[35602] = 32'b11111111111111111110011101011001;
assign LUT_2[35603] = 32'b11111111111111111011010101110010;
assign LUT_2[35604] = 32'b11111111111111110100000010000101;
assign LUT_2[35605] = 32'b11111111111111110000111010011110;
assign LUT_2[35606] = 32'b11111111111111111010111011000001;
assign LUT_2[35607] = 32'b11111111111111110111110011011010;
assign LUT_2[35608] = 32'b11111111111111110010010101111010;
assign LUT_2[35609] = 32'b11111111111111101111001110010011;
assign LUT_2[35610] = 32'b11111111111111111001001110110110;
assign LUT_2[35611] = 32'b11111111111111110110000111001111;
assign LUT_2[35612] = 32'b11111111111111101110110011100010;
assign LUT_2[35613] = 32'b11111111111111101011101011111011;
assign LUT_2[35614] = 32'b11111111111111110101101100011110;
assign LUT_2[35615] = 32'b11111111111111110010100100110111;
assign LUT_2[35616] = 32'b11111111111111111101011011111100;
assign LUT_2[35617] = 32'b11111111111111111010010100010101;
assign LUT_2[35618] = 32'b00000000000000000100010100111000;
assign LUT_2[35619] = 32'b00000000000000000001001101010001;
assign LUT_2[35620] = 32'b11111111111111111001111001100100;
assign LUT_2[35621] = 32'b11111111111111110110110001111101;
assign LUT_2[35622] = 32'b00000000000000000000110010100000;
assign LUT_2[35623] = 32'b11111111111111111101101010111001;
assign LUT_2[35624] = 32'b11111111111111111000001101011001;
assign LUT_2[35625] = 32'b11111111111111110101000101110010;
assign LUT_2[35626] = 32'b11111111111111111111000110010101;
assign LUT_2[35627] = 32'b11111111111111111011111110101110;
assign LUT_2[35628] = 32'b11111111111111110100101011000001;
assign LUT_2[35629] = 32'b11111111111111110001100011011010;
assign LUT_2[35630] = 32'b11111111111111111011100011111101;
assign LUT_2[35631] = 32'b11111111111111111000011100010110;
assign LUT_2[35632] = 32'b11111111111111111000000000000110;
assign LUT_2[35633] = 32'b11111111111111110100111000011111;
assign LUT_2[35634] = 32'b11111111111111111110111001000010;
assign LUT_2[35635] = 32'b11111111111111111011110001011011;
assign LUT_2[35636] = 32'b11111111111111110100011101101110;
assign LUT_2[35637] = 32'b11111111111111110001010110000111;
assign LUT_2[35638] = 32'b11111111111111111011010110101010;
assign LUT_2[35639] = 32'b11111111111111111000001111000011;
assign LUT_2[35640] = 32'b11111111111111110010110001100011;
assign LUT_2[35641] = 32'b11111111111111101111101001111100;
assign LUT_2[35642] = 32'b11111111111111111001101010011111;
assign LUT_2[35643] = 32'b11111111111111110110100010111000;
assign LUT_2[35644] = 32'b11111111111111101111001111001011;
assign LUT_2[35645] = 32'b11111111111111101100000111100100;
assign LUT_2[35646] = 32'b11111111111111110110001000000111;
assign LUT_2[35647] = 32'b11111111111111110011000000100000;
assign LUT_2[35648] = 32'b11111111111111110101001000110110;
assign LUT_2[35649] = 32'b11111111111111110010000001001111;
assign LUT_2[35650] = 32'b11111111111111111100000001110010;
assign LUT_2[35651] = 32'b11111111111111111000111010001011;
assign LUT_2[35652] = 32'b11111111111111110001100110011110;
assign LUT_2[35653] = 32'b11111111111111101110011110110111;
assign LUT_2[35654] = 32'b11111111111111111000011111011010;
assign LUT_2[35655] = 32'b11111111111111110101010111110011;
assign LUT_2[35656] = 32'b11111111111111101111111010010011;
assign LUT_2[35657] = 32'b11111111111111101100110010101100;
assign LUT_2[35658] = 32'b11111111111111110110110011001111;
assign LUT_2[35659] = 32'b11111111111111110011101011101000;
assign LUT_2[35660] = 32'b11111111111111101100010111111011;
assign LUT_2[35661] = 32'b11111111111111101001010000010100;
assign LUT_2[35662] = 32'b11111111111111110011010000110111;
assign LUT_2[35663] = 32'b11111111111111110000001001010000;
assign LUT_2[35664] = 32'b11111111111111101111101101000000;
assign LUT_2[35665] = 32'b11111111111111101100100101011001;
assign LUT_2[35666] = 32'b11111111111111110110100101111100;
assign LUT_2[35667] = 32'b11111111111111110011011110010101;
assign LUT_2[35668] = 32'b11111111111111101100001010101000;
assign LUT_2[35669] = 32'b11111111111111101001000011000001;
assign LUT_2[35670] = 32'b11111111111111110011000011100100;
assign LUT_2[35671] = 32'b11111111111111101111111011111101;
assign LUT_2[35672] = 32'b11111111111111101010011110011101;
assign LUT_2[35673] = 32'b11111111111111100111010110110110;
assign LUT_2[35674] = 32'b11111111111111110001010111011001;
assign LUT_2[35675] = 32'b11111111111111101110001111110010;
assign LUT_2[35676] = 32'b11111111111111100110111100000101;
assign LUT_2[35677] = 32'b11111111111111100011110100011110;
assign LUT_2[35678] = 32'b11111111111111101101110101000001;
assign LUT_2[35679] = 32'b11111111111111101010101101011010;
assign LUT_2[35680] = 32'b11111111111111110101100100011111;
assign LUT_2[35681] = 32'b11111111111111110010011100111000;
assign LUT_2[35682] = 32'b11111111111111111100011101011011;
assign LUT_2[35683] = 32'b11111111111111111001010101110100;
assign LUT_2[35684] = 32'b11111111111111110010000010000111;
assign LUT_2[35685] = 32'b11111111111111101110111010100000;
assign LUT_2[35686] = 32'b11111111111111111000111011000011;
assign LUT_2[35687] = 32'b11111111111111110101110011011100;
assign LUT_2[35688] = 32'b11111111111111110000010101111100;
assign LUT_2[35689] = 32'b11111111111111101101001110010101;
assign LUT_2[35690] = 32'b11111111111111110111001110111000;
assign LUT_2[35691] = 32'b11111111111111110100000111010001;
assign LUT_2[35692] = 32'b11111111111111101100110011100100;
assign LUT_2[35693] = 32'b11111111111111101001101011111101;
assign LUT_2[35694] = 32'b11111111111111110011101100100000;
assign LUT_2[35695] = 32'b11111111111111110000100100111001;
assign LUT_2[35696] = 32'b11111111111111110000001000101001;
assign LUT_2[35697] = 32'b11111111111111101101000001000010;
assign LUT_2[35698] = 32'b11111111111111110111000001100101;
assign LUT_2[35699] = 32'b11111111111111110011111001111110;
assign LUT_2[35700] = 32'b11111111111111101100100110010001;
assign LUT_2[35701] = 32'b11111111111111101001011110101010;
assign LUT_2[35702] = 32'b11111111111111110011011111001101;
assign LUT_2[35703] = 32'b11111111111111110000010111100110;
assign LUT_2[35704] = 32'b11111111111111101010111010000110;
assign LUT_2[35705] = 32'b11111111111111100111110010011111;
assign LUT_2[35706] = 32'b11111111111111110001110011000010;
assign LUT_2[35707] = 32'b11111111111111101110101011011011;
assign LUT_2[35708] = 32'b11111111111111100111010111101110;
assign LUT_2[35709] = 32'b11111111111111100100010000000111;
assign LUT_2[35710] = 32'b11111111111111101110010000101010;
assign LUT_2[35711] = 32'b11111111111111101011001001000011;
assign LUT_2[35712] = 32'b00000000000000000001010100100010;
assign LUT_2[35713] = 32'b11111111111111111110001100111011;
assign LUT_2[35714] = 32'b00000000000000001000001101011110;
assign LUT_2[35715] = 32'b00000000000000000101000101110111;
assign LUT_2[35716] = 32'b11111111111111111101110010001010;
assign LUT_2[35717] = 32'b11111111111111111010101010100011;
assign LUT_2[35718] = 32'b00000000000000000100101011000110;
assign LUT_2[35719] = 32'b00000000000000000001100011011111;
assign LUT_2[35720] = 32'b11111111111111111100000101111111;
assign LUT_2[35721] = 32'b11111111111111111000111110011000;
assign LUT_2[35722] = 32'b00000000000000000010111110111011;
assign LUT_2[35723] = 32'b11111111111111111111110111010100;
assign LUT_2[35724] = 32'b11111111111111111000100011100111;
assign LUT_2[35725] = 32'b11111111111111110101011100000000;
assign LUT_2[35726] = 32'b11111111111111111111011100100011;
assign LUT_2[35727] = 32'b11111111111111111100010100111100;
assign LUT_2[35728] = 32'b11111111111111111011111000101100;
assign LUT_2[35729] = 32'b11111111111111111000110001000101;
assign LUT_2[35730] = 32'b00000000000000000010110001101000;
assign LUT_2[35731] = 32'b11111111111111111111101010000001;
assign LUT_2[35732] = 32'b11111111111111111000010110010100;
assign LUT_2[35733] = 32'b11111111111111110101001110101101;
assign LUT_2[35734] = 32'b11111111111111111111001111010000;
assign LUT_2[35735] = 32'b11111111111111111100000111101001;
assign LUT_2[35736] = 32'b11111111111111110110101010001001;
assign LUT_2[35737] = 32'b11111111111111110011100010100010;
assign LUT_2[35738] = 32'b11111111111111111101100011000101;
assign LUT_2[35739] = 32'b11111111111111111010011011011110;
assign LUT_2[35740] = 32'b11111111111111110011000111110001;
assign LUT_2[35741] = 32'b11111111111111110000000000001010;
assign LUT_2[35742] = 32'b11111111111111111010000000101101;
assign LUT_2[35743] = 32'b11111111111111110110111001000110;
assign LUT_2[35744] = 32'b00000000000000000001110000001011;
assign LUT_2[35745] = 32'b11111111111111111110101000100100;
assign LUT_2[35746] = 32'b00000000000000001000101001000111;
assign LUT_2[35747] = 32'b00000000000000000101100001100000;
assign LUT_2[35748] = 32'b11111111111111111110001101110011;
assign LUT_2[35749] = 32'b11111111111111111011000110001100;
assign LUT_2[35750] = 32'b00000000000000000101000110101111;
assign LUT_2[35751] = 32'b00000000000000000001111111001000;
assign LUT_2[35752] = 32'b11111111111111111100100001101000;
assign LUT_2[35753] = 32'b11111111111111111001011010000001;
assign LUT_2[35754] = 32'b00000000000000000011011010100100;
assign LUT_2[35755] = 32'b00000000000000000000010010111101;
assign LUT_2[35756] = 32'b11111111111111111000111111010000;
assign LUT_2[35757] = 32'b11111111111111110101110111101001;
assign LUT_2[35758] = 32'b11111111111111111111111000001100;
assign LUT_2[35759] = 32'b11111111111111111100110000100101;
assign LUT_2[35760] = 32'b11111111111111111100010100010101;
assign LUT_2[35761] = 32'b11111111111111111001001100101110;
assign LUT_2[35762] = 32'b00000000000000000011001101010001;
assign LUT_2[35763] = 32'b00000000000000000000000101101010;
assign LUT_2[35764] = 32'b11111111111111111000110001111101;
assign LUT_2[35765] = 32'b11111111111111110101101010010110;
assign LUT_2[35766] = 32'b11111111111111111111101010111001;
assign LUT_2[35767] = 32'b11111111111111111100100011010010;
assign LUT_2[35768] = 32'b11111111111111110111000101110010;
assign LUT_2[35769] = 32'b11111111111111110011111110001011;
assign LUT_2[35770] = 32'b11111111111111111101111110101110;
assign LUT_2[35771] = 32'b11111111111111111010110111000111;
assign LUT_2[35772] = 32'b11111111111111110011100011011010;
assign LUT_2[35773] = 32'b11111111111111110000011011110011;
assign LUT_2[35774] = 32'b11111111111111111010011100010110;
assign LUT_2[35775] = 32'b11111111111111110111010100101111;
assign LUT_2[35776] = 32'b11111111111111111001011101000101;
assign LUT_2[35777] = 32'b11111111111111110110010101011110;
assign LUT_2[35778] = 32'b00000000000000000000010110000001;
assign LUT_2[35779] = 32'b11111111111111111101001110011010;
assign LUT_2[35780] = 32'b11111111111111110101111010101101;
assign LUT_2[35781] = 32'b11111111111111110010110011000110;
assign LUT_2[35782] = 32'b11111111111111111100110011101001;
assign LUT_2[35783] = 32'b11111111111111111001101100000010;
assign LUT_2[35784] = 32'b11111111111111110100001110100010;
assign LUT_2[35785] = 32'b11111111111111110001000110111011;
assign LUT_2[35786] = 32'b11111111111111111011000111011110;
assign LUT_2[35787] = 32'b11111111111111110111111111110111;
assign LUT_2[35788] = 32'b11111111111111110000101100001010;
assign LUT_2[35789] = 32'b11111111111111101101100100100011;
assign LUT_2[35790] = 32'b11111111111111110111100101000110;
assign LUT_2[35791] = 32'b11111111111111110100011101011111;
assign LUT_2[35792] = 32'b11111111111111110100000001001111;
assign LUT_2[35793] = 32'b11111111111111110000111001101000;
assign LUT_2[35794] = 32'b11111111111111111010111010001011;
assign LUT_2[35795] = 32'b11111111111111110111110010100100;
assign LUT_2[35796] = 32'b11111111111111110000011110110111;
assign LUT_2[35797] = 32'b11111111111111101101010111010000;
assign LUT_2[35798] = 32'b11111111111111110111010111110011;
assign LUT_2[35799] = 32'b11111111111111110100010000001100;
assign LUT_2[35800] = 32'b11111111111111101110110010101100;
assign LUT_2[35801] = 32'b11111111111111101011101011000101;
assign LUT_2[35802] = 32'b11111111111111110101101011101000;
assign LUT_2[35803] = 32'b11111111111111110010100100000001;
assign LUT_2[35804] = 32'b11111111111111101011010000010100;
assign LUT_2[35805] = 32'b11111111111111101000001000101101;
assign LUT_2[35806] = 32'b11111111111111110010001001010000;
assign LUT_2[35807] = 32'b11111111111111101111000001101001;
assign LUT_2[35808] = 32'b11111111111111111001111000101110;
assign LUT_2[35809] = 32'b11111111111111110110110001000111;
assign LUT_2[35810] = 32'b00000000000000000000110001101010;
assign LUT_2[35811] = 32'b11111111111111111101101010000011;
assign LUT_2[35812] = 32'b11111111111111110110010110010110;
assign LUT_2[35813] = 32'b11111111111111110011001110101111;
assign LUT_2[35814] = 32'b11111111111111111101001111010010;
assign LUT_2[35815] = 32'b11111111111111111010000111101011;
assign LUT_2[35816] = 32'b11111111111111110100101010001011;
assign LUT_2[35817] = 32'b11111111111111110001100010100100;
assign LUT_2[35818] = 32'b11111111111111111011100011000111;
assign LUT_2[35819] = 32'b11111111111111111000011011100000;
assign LUT_2[35820] = 32'b11111111111111110001000111110011;
assign LUT_2[35821] = 32'b11111111111111101110000000001100;
assign LUT_2[35822] = 32'b11111111111111111000000000101111;
assign LUT_2[35823] = 32'b11111111111111110100111001001000;
assign LUT_2[35824] = 32'b11111111111111110100011100111000;
assign LUT_2[35825] = 32'b11111111111111110001010101010001;
assign LUT_2[35826] = 32'b11111111111111111011010101110100;
assign LUT_2[35827] = 32'b11111111111111111000001110001101;
assign LUT_2[35828] = 32'b11111111111111110000111010100000;
assign LUT_2[35829] = 32'b11111111111111101101110010111001;
assign LUT_2[35830] = 32'b11111111111111110111110011011100;
assign LUT_2[35831] = 32'b11111111111111110100101011110101;
assign LUT_2[35832] = 32'b11111111111111101111001110010101;
assign LUT_2[35833] = 32'b11111111111111101100000110101110;
assign LUT_2[35834] = 32'b11111111111111110110000111010001;
assign LUT_2[35835] = 32'b11111111111111110010111111101010;
assign LUT_2[35836] = 32'b11111111111111101011101011111101;
assign LUT_2[35837] = 32'b11111111111111101000100100010110;
assign LUT_2[35838] = 32'b11111111111111110010100100111001;
assign LUT_2[35839] = 32'b11111111111111101111011101010010;
assign LUT_2[35840] = 32'b11111111111111111010111100000000;
assign LUT_2[35841] = 32'b11111111111111110111110100011001;
assign LUT_2[35842] = 32'b00000000000000000001110100111100;
assign LUT_2[35843] = 32'b11111111111111111110101101010101;
assign LUT_2[35844] = 32'b11111111111111110111011001101000;
assign LUT_2[35845] = 32'b11111111111111110100010010000001;
assign LUT_2[35846] = 32'b11111111111111111110010010100100;
assign LUT_2[35847] = 32'b11111111111111111011001010111101;
assign LUT_2[35848] = 32'b11111111111111110101101101011101;
assign LUT_2[35849] = 32'b11111111111111110010100101110110;
assign LUT_2[35850] = 32'b11111111111111111100100110011001;
assign LUT_2[35851] = 32'b11111111111111111001011110110010;
assign LUT_2[35852] = 32'b11111111111111110010001011000101;
assign LUT_2[35853] = 32'b11111111111111101111000011011110;
assign LUT_2[35854] = 32'b11111111111111111001000100000001;
assign LUT_2[35855] = 32'b11111111111111110101111100011010;
assign LUT_2[35856] = 32'b11111111111111110101100000001010;
assign LUT_2[35857] = 32'b11111111111111110010011000100011;
assign LUT_2[35858] = 32'b11111111111111111100011001000110;
assign LUT_2[35859] = 32'b11111111111111111001010001011111;
assign LUT_2[35860] = 32'b11111111111111110001111101110010;
assign LUT_2[35861] = 32'b11111111111111101110110110001011;
assign LUT_2[35862] = 32'b11111111111111111000110110101110;
assign LUT_2[35863] = 32'b11111111111111110101101111000111;
assign LUT_2[35864] = 32'b11111111111111110000010001100111;
assign LUT_2[35865] = 32'b11111111111111101101001010000000;
assign LUT_2[35866] = 32'b11111111111111110111001010100011;
assign LUT_2[35867] = 32'b11111111111111110100000010111100;
assign LUT_2[35868] = 32'b11111111111111101100101111001111;
assign LUT_2[35869] = 32'b11111111111111101001100111101000;
assign LUT_2[35870] = 32'b11111111111111110011101000001011;
assign LUT_2[35871] = 32'b11111111111111110000100000100100;
assign LUT_2[35872] = 32'b11111111111111111011010111101001;
assign LUT_2[35873] = 32'b11111111111111111000010000000010;
assign LUT_2[35874] = 32'b00000000000000000010010000100101;
assign LUT_2[35875] = 32'b11111111111111111111001000111110;
assign LUT_2[35876] = 32'b11111111111111110111110101010001;
assign LUT_2[35877] = 32'b11111111111111110100101101101010;
assign LUT_2[35878] = 32'b11111111111111111110101110001101;
assign LUT_2[35879] = 32'b11111111111111111011100110100110;
assign LUT_2[35880] = 32'b11111111111111110110001001000110;
assign LUT_2[35881] = 32'b11111111111111110011000001011111;
assign LUT_2[35882] = 32'b11111111111111111101000010000010;
assign LUT_2[35883] = 32'b11111111111111111001111010011011;
assign LUT_2[35884] = 32'b11111111111111110010100110101110;
assign LUT_2[35885] = 32'b11111111111111101111011111000111;
assign LUT_2[35886] = 32'b11111111111111111001011111101010;
assign LUT_2[35887] = 32'b11111111111111110110011000000011;
assign LUT_2[35888] = 32'b11111111111111110101111011110011;
assign LUT_2[35889] = 32'b11111111111111110010110100001100;
assign LUT_2[35890] = 32'b11111111111111111100110100101111;
assign LUT_2[35891] = 32'b11111111111111111001101101001000;
assign LUT_2[35892] = 32'b11111111111111110010011001011011;
assign LUT_2[35893] = 32'b11111111111111101111010001110100;
assign LUT_2[35894] = 32'b11111111111111111001010010010111;
assign LUT_2[35895] = 32'b11111111111111110110001010110000;
assign LUT_2[35896] = 32'b11111111111111110000101101010000;
assign LUT_2[35897] = 32'b11111111111111101101100101101001;
assign LUT_2[35898] = 32'b11111111111111110111100110001100;
assign LUT_2[35899] = 32'b11111111111111110100011110100101;
assign LUT_2[35900] = 32'b11111111111111101101001010111000;
assign LUT_2[35901] = 32'b11111111111111101010000011010001;
assign LUT_2[35902] = 32'b11111111111111110100000011110100;
assign LUT_2[35903] = 32'b11111111111111110000111100001101;
assign LUT_2[35904] = 32'b11111111111111110011000100100011;
assign LUT_2[35905] = 32'b11111111111111101111111100111100;
assign LUT_2[35906] = 32'b11111111111111111001111101011111;
assign LUT_2[35907] = 32'b11111111111111110110110101111000;
assign LUT_2[35908] = 32'b11111111111111101111100010001011;
assign LUT_2[35909] = 32'b11111111111111101100011010100100;
assign LUT_2[35910] = 32'b11111111111111110110011011000111;
assign LUT_2[35911] = 32'b11111111111111110011010011100000;
assign LUT_2[35912] = 32'b11111111111111101101110110000000;
assign LUT_2[35913] = 32'b11111111111111101010101110011001;
assign LUT_2[35914] = 32'b11111111111111110100101110111100;
assign LUT_2[35915] = 32'b11111111111111110001100111010101;
assign LUT_2[35916] = 32'b11111111111111101010010011101000;
assign LUT_2[35917] = 32'b11111111111111100111001100000001;
assign LUT_2[35918] = 32'b11111111111111110001001100100100;
assign LUT_2[35919] = 32'b11111111111111101110000100111101;
assign LUT_2[35920] = 32'b11111111111111101101101000101101;
assign LUT_2[35921] = 32'b11111111111111101010100001000110;
assign LUT_2[35922] = 32'b11111111111111110100100001101001;
assign LUT_2[35923] = 32'b11111111111111110001011010000010;
assign LUT_2[35924] = 32'b11111111111111101010000110010101;
assign LUT_2[35925] = 32'b11111111111111100110111110101110;
assign LUT_2[35926] = 32'b11111111111111110000111111010001;
assign LUT_2[35927] = 32'b11111111111111101101110111101010;
assign LUT_2[35928] = 32'b11111111111111101000011010001010;
assign LUT_2[35929] = 32'b11111111111111100101010010100011;
assign LUT_2[35930] = 32'b11111111111111101111010011000110;
assign LUT_2[35931] = 32'b11111111111111101100001011011111;
assign LUT_2[35932] = 32'b11111111111111100100110111110010;
assign LUT_2[35933] = 32'b11111111111111100001110000001011;
assign LUT_2[35934] = 32'b11111111111111101011110000101110;
assign LUT_2[35935] = 32'b11111111111111101000101001000111;
assign LUT_2[35936] = 32'b11111111111111110011100000001100;
assign LUT_2[35937] = 32'b11111111111111110000011000100101;
assign LUT_2[35938] = 32'b11111111111111111010011001001000;
assign LUT_2[35939] = 32'b11111111111111110111010001100001;
assign LUT_2[35940] = 32'b11111111111111101111111101110100;
assign LUT_2[35941] = 32'b11111111111111101100110110001101;
assign LUT_2[35942] = 32'b11111111111111110110110110110000;
assign LUT_2[35943] = 32'b11111111111111110011101111001001;
assign LUT_2[35944] = 32'b11111111111111101110010001101001;
assign LUT_2[35945] = 32'b11111111111111101011001010000010;
assign LUT_2[35946] = 32'b11111111111111110101001010100101;
assign LUT_2[35947] = 32'b11111111111111110010000010111110;
assign LUT_2[35948] = 32'b11111111111111101010101111010001;
assign LUT_2[35949] = 32'b11111111111111100111100111101010;
assign LUT_2[35950] = 32'b11111111111111110001101000001101;
assign LUT_2[35951] = 32'b11111111111111101110100000100110;
assign LUT_2[35952] = 32'b11111111111111101110000100010110;
assign LUT_2[35953] = 32'b11111111111111101010111100101111;
assign LUT_2[35954] = 32'b11111111111111110100111101010010;
assign LUT_2[35955] = 32'b11111111111111110001110101101011;
assign LUT_2[35956] = 32'b11111111111111101010100001111110;
assign LUT_2[35957] = 32'b11111111111111100111011010010111;
assign LUT_2[35958] = 32'b11111111111111110001011010111010;
assign LUT_2[35959] = 32'b11111111111111101110010011010011;
assign LUT_2[35960] = 32'b11111111111111101000110101110011;
assign LUT_2[35961] = 32'b11111111111111100101101110001100;
assign LUT_2[35962] = 32'b11111111111111101111101110101111;
assign LUT_2[35963] = 32'b11111111111111101100100111001000;
assign LUT_2[35964] = 32'b11111111111111100101010011011011;
assign LUT_2[35965] = 32'b11111111111111100010001011110100;
assign LUT_2[35966] = 32'b11111111111111101100001100010111;
assign LUT_2[35967] = 32'b11111111111111101001000100110000;
assign LUT_2[35968] = 32'b11111111111111111111010000001111;
assign LUT_2[35969] = 32'b11111111111111111100001000101000;
assign LUT_2[35970] = 32'b00000000000000000110001001001011;
assign LUT_2[35971] = 32'b00000000000000000011000001100100;
assign LUT_2[35972] = 32'b11111111111111111011101101110111;
assign LUT_2[35973] = 32'b11111111111111111000100110010000;
assign LUT_2[35974] = 32'b00000000000000000010100110110011;
assign LUT_2[35975] = 32'b11111111111111111111011111001100;
assign LUT_2[35976] = 32'b11111111111111111010000001101100;
assign LUT_2[35977] = 32'b11111111111111110110111010000101;
assign LUT_2[35978] = 32'b00000000000000000000111010101000;
assign LUT_2[35979] = 32'b11111111111111111101110011000001;
assign LUT_2[35980] = 32'b11111111111111110110011111010100;
assign LUT_2[35981] = 32'b11111111111111110011010111101101;
assign LUT_2[35982] = 32'b11111111111111111101011000010000;
assign LUT_2[35983] = 32'b11111111111111111010010000101001;
assign LUT_2[35984] = 32'b11111111111111111001110100011001;
assign LUT_2[35985] = 32'b11111111111111110110101100110010;
assign LUT_2[35986] = 32'b00000000000000000000101101010101;
assign LUT_2[35987] = 32'b11111111111111111101100101101110;
assign LUT_2[35988] = 32'b11111111111111110110010010000001;
assign LUT_2[35989] = 32'b11111111111111110011001010011010;
assign LUT_2[35990] = 32'b11111111111111111101001010111101;
assign LUT_2[35991] = 32'b11111111111111111010000011010110;
assign LUT_2[35992] = 32'b11111111111111110100100101110110;
assign LUT_2[35993] = 32'b11111111111111110001011110001111;
assign LUT_2[35994] = 32'b11111111111111111011011110110010;
assign LUT_2[35995] = 32'b11111111111111111000010111001011;
assign LUT_2[35996] = 32'b11111111111111110001000011011110;
assign LUT_2[35997] = 32'b11111111111111101101111011110111;
assign LUT_2[35998] = 32'b11111111111111110111111100011010;
assign LUT_2[35999] = 32'b11111111111111110100110100110011;
assign LUT_2[36000] = 32'b11111111111111111111101011111000;
assign LUT_2[36001] = 32'b11111111111111111100100100010001;
assign LUT_2[36002] = 32'b00000000000000000110100100110100;
assign LUT_2[36003] = 32'b00000000000000000011011101001101;
assign LUT_2[36004] = 32'b11111111111111111100001001100000;
assign LUT_2[36005] = 32'b11111111111111111001000001111001;
assign LUT_2[36006] = 32'b00000000000000000011000010011100;
assign LUT_2[36007] = 32'b11111111111111111111111010110101;
assign LUT_2[36008] = 32'b11111111111111111010011101010101;
assign LUT_2[36009] = 32'b11111111111111110111010101101110;
assign LUT_2[36010] = 32'b00000000000000000001010110010001;
assign LUT_2[36011] = 32'b11111111111111111110001110101010;
assign LUT_2[36012] = 32'b11111111111111110110111010111101;
assign LUT_2[36013] = 32'b11111111111111110011110011010110;
assign LUT_2[36014] = 32'b11111111111111111101110011111001;
assign LUT_2[36015] = 32'b11111111111111111010101100010010;
assign LUT_2[36016] = 32'b11111111111111111010010000000010;
assign LUT_2[36017] = 32'b11111111111111110111001000011011;
assign LUT_2[36018] = 32'b00000000000000000001001000111110;
assign LUT_2[36019] = 32'b11111111111111111110000001010111;
assign LUT_2[36020] = 32'b11111111111111110110101101101010;
assign LUT_2[36021] = 32'b11111111111111110011100110000011;
assign LUT_2[36022] = 32'b11111111111111111101100110100110;
assign LUT_2[36023] = 32'b11111111111111111010011110111111;
assign LUT_2[36024] = 32'b11111111111111110101000001011111;
assign LUT_2[36025] = 32'b11111111111111110001111001111000;
assign LUT_2[36026] = 32'b11111111111111111011111010011011;
assign LUT_2[36027] = 32'b11111111111111111000110010110100;
assign LUT_2[36028] = 32'b11111111111111110001011111000111;
assign LUT_2[36029] = 32'b11111111111111101110010111100000;
assign LUT_2[36030] = 32'b11111111111111111000011000000011;
assign LUT_2[36031] = 32'b11111111111111110101010000011100;
assign LUT_2[36032] = 32'b11111111111111110111011000110010;
assign LUT_2[36033] = 32'b11111111111111110100010001001011;
assign LUT_2[36034] = 32'b11111111111111111110010001101110;
assign LUT_2[36035] = 32'b11111111111111111011001010000111;
assign LUT_2[36036] = 32'b11111111111111110011110110011010;
assign LUT_2[36037] = 32'b11111111111111110000101110110011;
assign LUT_2[36038] = 32'b11111111111111111010101111010110;
assign LUT_2[36039] = 32'b11111111111111110111100111101111;
assign LUT_2[36040] = 32'b11111111111111110010001010001111;
assign LUT_2[36041] = 32'b11111111111111101111000010101000;
assign LUT_2[36042] = 32'b11111111111111111001000011001011;
assign LUT_2[36043] = 32'b11111111111111110101111011100100;
assign LUT_2[36044] = 32'b11111111111111101110100111110111;
assign LUT_2[36045] = 32'b11111111111111101011100000010000;
assign LUT_2[36046] = 32'b11111111111111110101100000110011;
assign LUT_2[36047] = 32'b11111111111111110010011001001100;
assign LUT_2[36048] = 32'b11111111111111110001111100111100;
assign LUT_2[36049] = 32'b11111111111111101110110101010101;
assign LUT_2[36050] = 32'b11111111111111111000110101111000;
assign LUT_2[36051] = 32'b11111111111111110101101110010001;
assign LUT_2[36052] = 32'b11111111111111101110011010100100;
assign LUT_2[36053] = 32'b11111111111111101011010010111101;
assign LUT_2[36054] = 32'b11111111111111110101010011100000;
assign LUT_2[36055] = 32'b11111111111111110010001011111001;
assign LUT_2[36056] = 32'b11111111111111101100101110011001;
assign LUT_2[36057] = 32'b11111111111111101001100110110010;
assign LUT_2[36058] = 32'b11111111111111110011100111010101;
assign LUT_2[36059] = 32'b11111111111111110000011111101110;
assign LUT_2[36060] = 32'b11111111111111101001001100000001;
assign LUT_2[36061] = 32'b11111111111111100110000100011010;
assign LUT_2[36062] = 32'b11111111111111110000000100111101;
assign LUT_2[36063] = 32'b11111111111111101100111101010110;
assign LUT_2[36064] = 32'b11111111111111110111110100011011;
assign LUT_2[36065] = 32'b11111111111111110100101100110100;
assign LUT_2[36066] = 32'b11111111111111111110101101010111;
assign LUT_2[36067] = 32'b11111111111111111011100101110000;
assign LUT_2[36068] = 32'b11111111111111110100010010000011;
assign LUT_2[36069] = 32'b11111111111111110001001010011100;
assign LUT_2[36070] = 32'b11111111111111111011001010111111;
assign LUT_2[36071] = 32'b11111111111111111000000011011000;
assign LUT_2[36072] = 32'b11111111111111110010100101111000;
assign LUT_2[36073] = 32'b11111111111111101111011110010001;
assign LUT_2[36074] = 32'b11111111111111111001011110110100;
assign LUT_2[36075] = 32'b11111111111111110110010111001101;
assign LUT_2[36076] = 32'b11111111111111101111000011100000;
assign LUT_2[36077] = 32'b11111111111111101011111011111001;
assign LUT_2[36078] = 32'b11111111111111110101111100011100;
assign LUT_2[36079] = 32'b11111111111111110010110100110101;
assign LUT_2[36080] = 32'b11111111111111110010011000100101;
assign LUT_2[36081] = 32'b11111111111111101111010000111110;
assign LUT_2[36082] = 32'b11111111111111111001010001100001;
assign LUT_2[36083] = 32'b11111111111111110110001001111010;
assign LUT_2[36084] = 32'b11111111111111101110110110001101;
assign LUT_2[36085] = 32'b11111111111111101011101110100110;
assign LUT_2[36086] = 32'b11111111111111110101101111001001;
assign LUT_2[36087] = 32'b11111111111111110010100111100010;
assign LUT_2[36088] = 32'b11111111111111101101001010000010;
assign LUT_2[36089] = 32'b11111111111111101010000010011011;
assign LUT_2[36090] = 32'b11111111111111110100000010111110;
assign LUT_2[36091] = 32'b11111111111111110000111011010111;
assign LUT_2[36092] = 32'b11111111111111101001100111101010;
assign LUT_2[36093] = 32'b11111111111111100110100000000011;
assign LUT_2[36094] = 32'b11111111111111110000100000100110;
assign LUT_2[36095] = 32'b11111111111111101101011000111111;
assign LUT_2[36096] = 32'b11111111111111111110111010100110;
assign LUT_2[36097] = 32'b11111111111111111011110010111111;
assign LUT_2[36098] = 32'b00000000000000000101110011100010;
assign LUT_2[36099] = 32'b00000000000000000010101011111011;
assign LUT_2[36100] = 32'b11111111111111111011011000001110;
assign LUT_2[36101] = 32'b11111111111111111000010000100111;
assign LUT_2[36102] = 32'b00000000000000000010010001001010;
assign LUT_2[36103] = 32'b11111111111111111111001001100011;
assign LUT_2[36104] = 32'b11111111111111111001101100000011;
assign LUT_2[36105] = 32'b11111111111111110110100100011100;
assign LUT_2[36106] = 32'b00000000000000000000100100111111;
assign LUT_2[36107] = 32'b11111111111111111101011101011000;
assign LUT_2[36108] = 32'b11111111111111110110001001101011;
assign LUT_2[36109] = 32'b11111111111111110011000010000100;
assign LUT_2[36110] = 32'b11111111111111111101000010100111;
assign LUT_2[36111] = 32'b11111111111111111001111011000000;
assign LUT_2[36112] = 32'b11111111111111111001011110110000;
assign LUT_2[36113] = 32'b11111111111111110110010111001001;
assign LUT_2[36114] = 32'b00000000000000000000010111101100;
assign LUT_2[36115] = 32'b11111111111111111101010000000101;
assign LUT_2[36116] = 32'b11111111111111110101111100011000;
assign LUT_2[36117] = 32'b11111111111111110010110100110001;
assign LUT_2[36118] = 32'b11111111111111111100110101010100;
assign LUT_2[36119] = 32'b11111111111111111001101101101101;
assign LUT_2[36120] = 32'b11111111111111110100010000001101;
assign LUT_2[36121] = 32'b11111111111111110001001000100110;
assign LUT_2[36122] = 32'b11111111111111111011001001001001;
assign LUT_2[36123] = 32'b11111111111111111000000001100010;
assign LUT_2[36124] = 32'b11111111111111110000101101110101;
assign LUT_2[36125] = 32'b11111111111111101101100110001110;
assign LUT_2[36126] = 32'b11111111111111110111100110110001;
assign LUT_2[36127] = 32'b11111111111111110100011111001010;
assign LUT_2[36128] = 32'b11111111111111111111010110001111;
assign LUT_2[36129] = 32'b11111111111111111100001110101000;
assign LUT_2[36130] = 32'b00000000000000000110001111001011;
assign LUT_2[36131] = 32'b00000000000000000011000111100100;
assign LUT_2[36132] = 32'b11111111111111111011110011110111;
assign LUT_2[36133] = 32'b11111111111111111000101100010000;
assign LUT_2[36134] = 32'b00000000000000000010101100110011;
assign LUT_2[36135] = 32'b11111111111111111111100101001100;
assign LUT_2[36136] = 32'b11111111111111111010000111101100;
assign LUT_2[36137] = 32'b11111111111111110111000000000101;
assign LUT_2[36138] = 32'b00000000000000000001000000101000;
assign LUT_2[36139] = 32'b11111111111111111101111001000001;
assign LUT_2[36140] = 32'b11111111111111110110100101010100;
assign LUT_2[36141] = 32'b11111111111111110011011101101101;
assign LUT_2[36142] = 32'b11111111111111111101011110010000;
assign LUT_2[36143] = 32'b11111111111111111010010110101001;
assign LUT_2[36144] = 32'b11111111111111111001111010011001;
assign LUT_2[36145] = 32'b11111111111111110110110010110010;
assign LUT_2[36146] = 32'b00000000000000000000110011010101;
assign LUT_2[36147] = 32'b11111111111111111101101011101110;
assign LUT_2[36148] = 32'b11111111111111110110011000000001;
assign LUT_2[36149] = 32'b11111111111111110011010000011010;
assign LUT_2[36150] = 32'b11111111111111111101010000111101;
assign LUT_2[36151] = 32'b11111111111111111010001001010110;
assign LUT_2[36152] = 32'b11111111111111110100101011110110;
assign LUT_2[36153] = 32'b11111111111111110001100100001111;
assign LUT_2[36154] = 32'b11111111111111111011100100110010;
assign LUT_2[36155] = 32'b11111111111111111000011101001011;
assign LUT_2[36156] = 32'b11111111111111110001001001011110;
assign LUT_2[36157] = 32'b11111111111111101110000001110111;
assign LUT_2[36158] = 32'b11111111111111111000000010011010;
assign LUT_2[36159] = 32'b11111111111111110100111010110011;
assign LUT_2[36160] = 32'b11111111111111110111000011001001;
assign LUT_2[36161] = 32'b11111111111111110011111011100010;
assign LUT_2[36162] = 32'b11111111111111111101111100000101;
assign LUT_2[36163] = 32'b11111111111111111010110100011110;
assign LUT_2[36164] = 32'b11111111111111110011100000110001;
assign LUT_2[36165] = 32'b11111111111111110000011001001010;
assign LUT_2[36166] = 32'b11111111111111111010011001101101;
assign LUT_2[36167] = 32'b11111111111111110111010010000110;
assign LUT_2[36168] = 32'b11111111111111110001110100100110;
assign LUT_2[36169] = 32'b11111111111111101110101100111111;
assign LUT_2[36170] = 32'b11111111111111111000101101100010;
assign LUT_2[36171] = 32'b11111111111111110101100101111011;
assign LUT_2[36172] = 32'b11111111111111101110010010001110;
assign LUT_2[36173] = 32'b11111111111111101011001010100111;
assign LUT_2[36174] = 32'b11111111111111110101001011001010;
assign LUT_2[36175] = 32'b11111111111111110010000011100011;
assign LUT_2[36176] = 32'b11111111111111110001100111010011;
assign LUT_2[36177] = 32'b11111111111111101110011111101100;
assign LUT_2[36178] = 32'b11111111111111111000100000001111;
assign LUT_2[36179] = 32'b11111111111111110101011000101000;
assign LUT_2[36180] = 32'b11111111111111101110000100111011;
assign LUT_2[36181] = 32'b11111111111111101010111101010100;
assign LUT_2[36182] = 32'b11111111111111110100111101110111;
assign LUT_2[36183] = 32'b11111111111111110001110110010000;
assign LUT_2[36184] = 32'b11111111111111101100011000110000;
assign LUT_2[36185] = 32'b11111111111111101001010001001001;
assign LUT_2[36186] = 32'b11111111111111110011010001101100;
assign LUT_2[36187] = 32'b11111111111111110000001010000101;
assign LUT_2[36188] = 32'b11111111111111101000110110011000;
assign LUT_2[36189] = 32'b11111111111111100101101110110001;
assign LUT_2[36190] = 32'b11111111111111101111101111010100;
assign LUT_2[36191] = 32'b11111111111111101100100111101101;
assign LUT_2[36192] = 32'b11111111111111110111011110110010;
assign LUT_2[36193] = 32'b11111111111111110100010111001011;
assign LUT_2[36194] = 32'b11111111111111111110010111101110;
assign LUT_2[36195] = 32'b11111111111111111011010000000111;
assign LUT_2[36196] = 32'b11111111111111110011111100011010;
assign LUT_2[36197] = 32'b11111111111111110000110100110011;
assign LUT_2[36198] = 32'b11111111111111111010110101010110;
assign LUT_2[36199] = 32'b11111111111111110111101101101111;
assign LUT_2[36200] = 32'b11111111111111110010010000001111;
assign LUT_2[36201] = 32'b11111111111111101111001000101000;
assign LUT_2[36202] = 32'b11111111111111111001001001001011;
assign LUT_2[36203] = 32'b11111111111111110110000001100100;
assign LUT_2[36204] = 32'b11111111111111101110101101110111;
assign LUT_2[36205] = 32'b11111111111111101011100110010000;
assign LUT_2[36206] = 32'b11111111111111110101100110110011;
assign LUT_2[36207] = 32'b11111111111111110010011111001100;
assign LUT_2[36208] = 32'b11111111111111110010000010111100;
assign LUT_2[36209] = 32'b11111111111111101110111011010101;
assign LUT_2[36210] = 32'b11111111111111111000111011111000;
assign LUT_2[36211] = 32'b11111111111111110101110100010001;
assign LUT_2[36212] = 32'b11111111111111101110100000100100;
assign LUT_2[36213] = 32'b11111111111111101011011000111101;
assign LUT_2[36214] = 32'b11111111111111110101011001100000;
assign LUT_2[36215] = 32'b11111111111111110010010001111001;
assign LUT_2[36216] = 32'b11111111111111101100110100011001;
assign LUT_2[36217] = 32'b11111111111111101001101100110010;
assign LUT_2[36218] = 32'b11111111111111110011101101010101;
assign LUT_2[36219] = 32'b11111111111111110000100101101110;
assign LUT_2[36220] = 32'b11111111111111101001010010000001;
assign LUT_2[36221] = 32'b11111111111111100110001010011010;
assign LUT_2[36222] = 32'b11111111111111110000001010111101;
assign LUT_2[36223] = 32'b11111111111111101101000011010110;
assign LUT_2[36224] = 32'b00000000000000000011001110110101;
assign LUT_2[36225] = 32'b00000000000000000000000111001110;
assign LUT_2[36226] = 32'b00000000000000001010000111110001;
assign LUT_2[36227] = 32'b00000000000000000111000000001010;
assign LUT_2[36228] = 32'b11111111111111111111101100011101;
assign LUT_2[36229] = 32'b11111111111111111100100100110110;
assign LUT_2[36230] = 32'b00000000000000000110100101011001;
assign LUT_2[36231] = 32'b00000000000000000011011101110010;
assign LUT_2[36232] = 32'b11111111111111111110000000010010;
assign LUT_2[36233] = 32'b11111111111111111010111000101011;
assign LUT_2[36234] = 32'b00000000000000000100111001001110;
assign LUT_2[36235] = 32'b00000000000000000001110001100111;
assign LUT_2[36236] = 32'b11111111111111111010011101111010;
assign LUT_2[36237] = 32'b11111111111111110111010110010011;
assign LUT_2[36238] = 32'b00000000000000000001010110110110;
assign LUT_2[36239] = 32'b11111111111111111110001111001111;
assign LUT_2[36240] = 32'b11111111111111111101110010111111;
assign LUT_2[36241] = 32'b11111111111111111010101011011000;
assign LUT_2[36242] = 32'b00000000000000000100101011111011;
assign LUT_2[36243] = 32'b00000000000000000001100100010100;
assign LUT_2[36244] = 32'b11111111111111111010010000100111;
assign LUT_2[36245] = 32'b11111111111111110111001001000000;
assign LUT_2[36246] = 32'b00000000000000000001001001100011;
assign LUT_2[36247] = 32'b11111111111111111110000001111100;
assign LUT_2[36248] = 32'b11111111111111111000100100011100;
assign LUT_2[36249] = 32'b11111111111111110101011100110101;
assign LUT_2[36250] = 32'b11111111111111111111011101011000;
assign LUT_2[36251] = 32'b11111111111111111100010101110001;
assign LUT_2[36252] = 32'b11111111111111110101000010000100;
assign LUT_2[36253] = 32'b11111111111111110001111010011101;
assign LUT_2[36254] = 32'b11111111111111111011111011000000;
assign LUT_2[36255] = 32'b11111111111111111000110011011001;
assign LUT_2[36256] = 32'b00000000000000000011101010011110;
assign LUT_2[36257] = 32'b00000000000000000000100010110111;
assign LUT_2[36258] = 32'b00000000000000001010100011011010;
assign LUT_2[36259] = 32'b00000000000000000111011011110011;
assign LUT_2[36260] = 32'b00000000000000000000001000000110;
assign LUT_2[36261] = 32'b11111111111111111101000000011111;
assign LUT_2[36262] = 32'b00000000000000000111000001000010;
assign LUT_2[36263] = 32'b00000000000000000011111001011011;
assign LUT_2[36264] = 32'b11111111111111111110011011111011;
assign LUT_2[36265] = 32'b11111111111111111011010100010100;
assign LUT_2[36266] = 32'b00000000000000000101010100110111;
assign LUT_2[36267] = 32'b00000000000000000010001101010000;
assign LUT_2[36268] = 32'b11111111111111111010111001100011;
assign LUT_2[36269] = 32'b11111111111111110111110001111100;
assign LUT_2[36270] = 32'b00000000000000000001110010011111;
assign LUT_2[36271] = 32'b11111111111111111110101010111000;
assign LUT_2[36272] = 32'b11111111111111111110001110101000;
assign LUT_2[36273] = 32'b11111111111111111011000111000001;
assign LUT_2[36274] = 32'b00000000000000000101000111100100;
assign LUT_2[36275] = 32'b00000000000000000001111111111101;
assign LUT_2[36276] = 32'b11111111111111111010101100010000;
assign LUT_2[36277] = 32'b11111111111111110111100100101001;
assign LUT_2[36278] = 32'b00000000000000000001100101001100;
assign LUT_2[36279] = 32'b11111111111111111110011101100101;
assign LUT_2[36280] = 32'b11111111111111111001000000000101;
assign LUT_2[36281] = 32'b11111111111111110101111000011110;
assign LUT_2[36282] = 32'b11111111111111111111111001000001;
assign LUT_2[36283] = 32'b11111111111111111100110001011010;
assign LUT_2[36284] = 32'b11111111111111110101011101101101;
assign LUT_2[36285] = 32'b11111111111111110010010110000110;
assign LUT_2[36286] = 32'b11111111111111111100010110101001;
assign LUT_2[36287] = 32'b11111111111111111001001111000010;
assign LUT_2[36288] = 32'b11111111111111111011010111011000;
assign LUT_2[36289] = 32'b11111111111111111000001111110001;
assign LUT_2[36290] = 32'b00000000000000000010010000010100;
assign LUT_2[36291] = 32'b11111111111111111111001000101101;
assign LUT_2[36292] = 32'b11111111111111110111110101000000;
assign LUT_2[36293] = 32'b11111111111111110100101101011001;
assign LUT_2[36294] = 32'b11111111111111111110101101111100;
assign LUT_2[36295] = 32'b11111111111111111011100110010101;
assign LUT_2[36296] = 32'b11111111111111110110001000110101;
assign LUT_2[36297] = 32'b11111111111111110011000001001110;
assign LUT_2[36298] = 32'b11111111111111111101000001110001;
assign LUT_2[36299] = 32'b11111111111111111001111010001010;
assign LUT_2[36300] = 32'b11111111111111110010100110011101;
assign LUT_2[36301] = 32'b11111111111111101111011110110110;
assign LUT_2[36302] = 32'b11111111111111111001011111011001;
assign LUT_2[36303] = 32'b11111111111111110110010111110010;
assign LUT_2[36304] = 32'b11111111111111110101111011100010;
assign LUT_2[36305] = 32'b11111111111111110010110011111011;
assign LUT_2[36306] = 32'b11111111111111111100110100011110;
assign LUT_2[36307] = 32'b11111111111111111001101100110111;
assign LUT_2[36308] = 32'b11111111111111110010011001001010;
assign LUT_2[36309] = 32'b11111111111111101111010001100011;
assign LUT_2[36310] = 32'b11111111111111111001010010000110;
assign LUT_2[36311] = 32'b11111111111111110110001010011111;
assign LUT_2[36312] = 32'b11111111111111110000101100111111;
assign LUT_2[36313] = 32'b11111111111111101101100101011000;
assign LUT_2[36314] = 32'b11111111111111110111100101111011;
assign LUT_2[36315] = 32'b11111111111111110100011110010100;
assign LUT_2[36316] = 32'b11111111111111101101001010100111;
assign LUT_2[36317] = 32'b11111111111111101010000011000000;
assign LUT_2[36318] = 32'b11111111111111110100000011100011;
assign LUT_2[36319] = 32'b11111111111111110000111011111100;
assign LUT_2[36320] = 32'b11111111111111111011110011000001;
assign LUT_2[36321] = 32'b11111111111111111000101011011010;
assign LUT_2[36322] = 32'b00000000000000000010101011111101;
assign LUT_2[36323] = 32'b11111111111111111111100100010110;
assign LUT_2[36324] = 32'b11111111111111111000010000101001;
assign LUT_2[36325] = 32'b11111111111111110101001001000010;
assign LUT_2[36326] = 32'b11111111111111111111001001100101;
assign LUT_2[36327] = 32'b11111111111111111100000001111110;
assign LUT_2[36328] = 32'b11111111111111110110100100011110;
assign LUT_2[36329] = 32'b11111111111111110011011100110111;
assign LUT_2[36330] = 32'b11111111111111111101011101011010;
assign LUT_2[36331] = 32'b11111111111111111010010101110011;
assign LUT_2[36332] = 32'b11111111111111110011000010000110;
assign LUT_2[36333] = 32'b11111111111111101111111010011111;
assign LUT_2[36334] = 32'b11111111111111111001111011000010;
assign LUT_2[36335] = 32'b11111111111111110110110011011011;
assign LUT_2[36336] = 32'b11111111111111110110010111001011;
assign LUT_2[36337] = 32'b11111111111111110011001111100100;
assign LUT_2[36338] = 32'b11111111111111111101010000000111;
assign LUT_2[36339] = 32'b11111111111111111010001000100000;
assign LUT_2[36340] = 32'b11111111111111110010110100110011;
assign LUT_2[36341] = 32'b11111111111111101111101101001100;
assign LUT_2[36342] = 32'b11111111111111111001101101101111;
assign LUT_2[36343] = 32'b11111111111111110110100110001000;
assign LUT_2[36344] = 32'b11111111111111110001001000101000;
assign LUT_2[36345] = 32'b11111111111111101110000001000001;
assign LUT_2[36346] = 32'b11111111111111111000000001100100;
assign LUT_2[36347] = 32'b11111111111111110100111001111101;
assign LUT_2[36348] = 32'b11111111111111101101100110010000;
assign LUT_2[36349] = 32'b11111111111111101010011110101001;
assign LUT_2[36350] = 32'b11111111111111110100011111001100;
assign LUT_2[36351] = 32'b11111111111111110001010111100101;
assign LUT_2[36352] = 32'b11111111111111111111101101110010;
assign LUT_2[36353] = 32'b11111111111111111100100110001011;
assign LUT_2[36354] = 32'b00000000000000000110100110101110;
assign LUT_2[36355] = 32'b00000000000000000011011111000111;
assign LUT_2[36356] = 32'b11111111111111111100001011011010;
assign LUT_2[36357] = 32'b11111111111111111001000011110011;
assign LUT_2[36358] = 32'b00000000000000000011000100010110;
assign LUT_2[36359] = 32'b11111111111111111111111100101111;
assign LUT_2[36360] = 32'b11111111111111111010011111001111;
assign LUT_2[36361] = 32'b11111111111111110111010111101000;
assign LUT_2[36362] = 32'b00000000000000000001011000001011;
assign LUT_2[36363] = 32'b11111111111111111110010000100100;
assign LUT_2[36364] = 32'b11111111111111110110111100110111;
assign LUT_2[36365] = 32'b11111111111111110011110101010000;
assign LUT_2[36366] = 32'b11111111111111111101110101110011;
assign LUT_2[36367] = 32'b11111111111111111010101110001100;
assign LUT_2[36368] = 32'b11111111111111111010010001111100;
assign LUT_2[36369] = 32'b11111111111111110111001010010101;
assign LUT_2[36370] = 32'b00000000000000000001001010111000;
assign LUT_2[36371] = 32'b11111111111111111110000011010001;
assign LUT_2[36372] = 32'b11111111111111110110101111100100;
assign LUT_2[36373] = 32'b11111111111111110011100111111101;
assign LUT_2[36374] = 32'b11111111111111111101101000100000;
assign LUT_2[36375] = 32'b11111111111111111010100000111001;
assign LUT_2[36376] = 32'b11111111111111110101000011011001;
assign LUT_2[36377] = 32'b11111111111111110001111011110010;
assign LUT_2[36378] = 32'b11111111111111111011111100010101;
assign LUT_2[36379] = 32'b11111111111111111000110100101110;
assign LUT_2[36380] = 32'b11111111111111110001100001000001;
assign LUT_2[36381] = 32'b11111111111111101110011001011010;
assign LUT_2[36382] = 32'b11111111111111111000011001111101;
assign LUT_2[36383] = 32'b11111111111111110101010010010110;
assign LUT_2[36384] = 32'b00000000000000000000001001011011;
assign LUT_2[36385] = 32'b11111111111111111101000001110100;
assign LUT_2[36386] = 32'b00000000000000000111000010010111;
assign LUT_2[36387] = 32'b00000000000000000011111010110000;
assign LUT_2[36388] = 32'b11111111111111111100100111000011;
assign LUT_2[36389] = 32'b11111111111111111001011111011100;
assign LUT_2[36390] = 32'b00000000000000000011011111111111;
assign LUT_2[36391] = 32'b00000000000000000000011000011000;
assign LUT_2[36392] = 32'b11111111111111111010111010111000;
assign LUT_2[36393] = 32'b11111111111111110111110011010001;
assign LUT_2[36394] = 32'b00000000000000000001110011110100;
assign LUT_2[36395] = 32'b11111111111111111110101100001101;
assign LUT_2[36396] = 32'b11111111111111110111011000100000;
assign LUT_2[36397] = 32'b11111111111111110100010000111001;
assign LUT_2[36398] = 32'b11111111111111111110010001011100;
assign LUT_2[36399] = 32'b11111111111111111011001001110101;
assign LUT_2[36400] = 32'b11111111111111111010101101100101;
assign LUT_2[36401] = 32'b11111111111111110111100101111110;
assign LUT_2[36402] = 32'b00000000000000000001100110100001;
assign LUT_2[36403] = 32'b11111111111111111110011110111010;
assign LUT_2[36404] = 32'b11111111111111110111001011001101;
assign LUT_2[36405] = 32'b11111111111111110100000011100110;
assign LUT_2[36406] = 32'b11111111111111111110000100001001;
assign LUT_2[36407] = 32'b11111111111111111010111100100010;
assign LUT_2[36408] = 32'b11111111111111110101011111000010;
assign LUT_2[36409] = 32'b11111111111111110010010111011011;
assign LUT_2[36410] = 32'b11111111111111111100010111111110;
assign LUT_2[36411] = 32'b11111111111111111001010000010111;
assign LUT_2[36412] = 32'b11111111111111110001111100101010;
assign LUT_2[36413] = 32'b11111111111111101110110101000011;
assign LUT_2[36414] = 32'b11111111111111111000110101100110;
assign LUT_2[36415] = 32'b11111111111111110101101101111111;
assign LUT_2[36416] = 32'b11111111111111110111110110010101;
assign LUT_2[36417] = 32'b11111111111111110100101110101110;
assign LUT_2[36418] = 32'b11111111111111111110101111010001;
assign LUT_2[36419] = 32'b11111111111111111011100111101010;
assign LUT_2[36420] = 32'b11111111111111110100010011111101;
assign LUT_2[36421] = 32'b11111111111111110001001100010110;
assign LUT_2[36422] = 32'b11111111111111111011001100111001;
assign LUT_2[36423] = 32'b11111111111111111000000101010010;
assign LUT_2[36424] = 32'b11111111111111110010100111110010;
assign LUT_2[36425] = 32'b11111111111111101111100000001011;
assign LUT_2[36426] = 32'b11111111111111111001100000101110;
assign LUT_2[36427] = 32'b11111111111111110110011001000111;
assign LUT_2[36428] = 32'b11111111111111101111000101011010;
assign LUT_2[36429] = 32'b11111111111111101011111101110011;
assign LUT_2[36430] = 32'b11111111111111110101111110010110;
assign LUT_2[36431] = 32'b11111111111111110010110110101111;
assign LUT_2[36432] = 32'b11111111111111110010011010011111;
assign LUT_2[36433] = 32'b11111111111111101111010010111000;
assign LUT_2[36434] = 32'b11111111111111111001010011011011;
assign LUT_2[36435] = 32'b11111111111111110110001011110100;
assign LUT_2[36436] = 32'b11111111111111101110111000000111;
assign LUT_2[36437] = 32'b11111111111111101011110000100000;
assign LUT_2[36438] = 32'b11111111111111110101110001000011;
assign LUT_2[36439] = 32'b11111111111111110010101001011100;
assign LUT_2[36440] = 32'b11111111111111101101001011111100;
assign LUT_2[36441] = 32'b11111111111111101010000100010101;
assign LUT_2[36442] = 32'b11111111111111110100000100111000;
assign LUT_2[36443] = 32'b11111111111111110000111101010001;
assign LUT_2[36444] = 32'b11111111111111101001101001100100;
assign LUT_2[36445] = 32'b11111111111111100110100001111101;
assign LUT_2[36446] = 32'b11111111111111110000100010100000;
assign LUT_2[36447] = 32'b11111111111111101101011010111001;
assign LUT_2[36448] = 32'b11111111111111111000010001111110;
assign LUT_2[36449] = 32'b11111111111111110101001010010111;
assign LUT_2[36450] = 32'b11111111111111111111001010111010;
assign LUT_2[36451] = 32'b11111111111111111100000011010011;
assign LUT_2[36452] = 32'b11111111111111110100101111100110;
assign LUT_2[36453] = 32'b11111111111111110001100111111111;
assign LUT_2[36454] = 32'b11111111111111111011101000100010;
assign LUT_2[36455] = 32'b11111111111111111000100000111011;
assign LUT_2[36456] = 32'b11111111111111110011000011011011;
assign LUT_2[36457] = 32'b11111111111111101111111011110100;
assign LUT_2[36458] = 32'b11111111111111111001111100010111;
assign LUT_2[36459] = 32'b11111111111111110110110100110000;
assign LUT_2[36460] = 32'b11111111111111101111100001000011;
assign LUT_2[36461] = 32'b11111111111111101100011001011100;
assign LUT_2[36462] = 32'b11111111111111110110011001111111;
assign LUT_2[36463] = 32'b11111111111111110011010010011000;
assign LUT_2[36464] = 32'b11111111111111110010110110001000;
assign LUT_2[36465] = 32'b11111111111111101111101110100001;
assign LUT_2[36466] = 32'b11111111111111111001101111000100;
assign LUT_2[36467] = 32'b11111111111111110110100111011101;
assign LUT_2[36468] = 32'b11111111111111101111010011110000;
assign LUT_2[36469] = 32'b11111111111111101100001100001001;
assign LUT_2[36470] = 32'b11111111111111110110001100101100;
assign LUT_2[36471] = 32'b11111111111111110011000101000101;
assign LUT_2[36472] = 32'b11111111111111101101100111100101;
assign LUT_2[36473] = 32'b11111111111111101010011111111110;
assign LUT_2[36474] = 32'b11111111111111110100100000100001;
assign LUT_2[36475] = 32'b11111111111111110001011000111010;
assign LUT_2[36476] = 32'b11111111111111101010000101001101;
assign LUT_2[36477] = 32'b11111111111111100110111101100110;
assign LUT_2[36478] = 32'b11111111111111110000111110001001;
assign LUT_2[36479] = 32'b11111111111111101101110110100010;
assign LUT_2[36480] = 32'b00000000000000000100000010000001;
assign LUT_2[36481] = 32'b00000000000000000000111010011010;
assign LUT_2[36482] = 32'b00000000000000001010111010111101;
assign LUT_2[36483] = 32'b00000000000000000111110011010110;
assign LUT_2[36484] = 32'b00000000000000000000011111101001;
assign LUT_2[36485] = 32'b11111111111111111101011000000010;
assign LUT_2[36486] = 32'b00000000000000000111011000100101;
assign LUT_2[36487] = 32'b00000000000000000100010000111110;
assign LUT_2[36488] = 32'b11111111111111111110110011011110;
assign LUT_2[36489] = 32'b11111111111111111011101011110111;
assign LUT_2[36490] = 32'b00000000000000000101101100011010;
assign LUT_2[36491] = 32'b00000000000000000010100100110011;
assign LUT_2[36492] = 32'b11111111111111111011010001000110;
assign LUT_2[36493] = 32'b11111111111111111000001001011111;
assign LUT_2[36494] = 32'b00000000000000000010001010000010;
assign LUT_2[36495] = 32'b11111111111111111111000010011011;
assign LUT_2[36496] = 32'b11111111111111111110100110001011;
assign LUT_2[36497] = 32'b11111111111111111011011110100100;
assign LUT_2[36498] = 32'b00000000000000000101011111000111;
assign LUT_2[36499] = 32'b00000000000000000010010111100000;
assign LUT_2[36500] = 32'b11111111111111111011000011110011;
assign LUT_2[36501] = 32'b11111111111111110111111100001100;
assign LUT_2[36502] = 32'b00000000000000000001111100101111;
assign LUT_2[36503] = 32'b11111111111111111110110101001000;
assign LUT_2[36504] = 32'b11111111111111111001010111101000;
assign LUT_2[36505] = 32'b11111111111111110110010000000001;
assign LUT_2[36506] = 32'b00000000000000000000010000100100;
assign LUT_2[36507] = 32'b11111111111111111101001000111101;
assign LUT_2[36508] = 32'b11111111111111110101110101010000;
assign LUT_2[36509] = 32'b11111111111111110010101101101001;
assign LUT_2[36510] = 32'b11111111111111111100101110001100;
assign LUT_2[36511] = 32'b11111111111111111001100110100101;
assign LUT_2[36512] = 32'b00000000000000000100011101101010;
assign LUT_2[36513] = 32'b00000000000000000001010110000011;
assign LUT_2[36514] = 32'b00000000000000001011010110100110;
assign LUT_2[36515] = 32'b00000000000000001000001110111111;
assign LUT_2[36516] = 32'b00000000000000000000111011010010;
assign LUT_2[36517] = 32'b11111111111111111101110011101011;
assign LUT_2[36518] = 32'b00000000000000000111110100001110;
assign LUT_2[36519] = 32'b00000000000000000100101100100111;
assign LUT_2[36520] = 32'b11111111111111111111001111000111;
assign LUT_2[36521] = 32'b11111111111111111100000111100000;
assign LUT_2[36522] = 32'b00000000000000000110001000000011;
assign LUT_2[36523] = 32'b00000000000000000011000000011100;
assign LUT_2[36524] = 32'b11111111111111111011101100101111;
assign LUT_2[36525] = 32'b11111111111111111000100101001000;
assign LUT_2[36526] = 32'b00000000000000000010100101101011;
assign LUT_2[36527] = 32'b11111111111111111111011110000100;
assign LUT_2[36528] = 32'b11111111111111111111000001110100;
assign LUT_2[36529] = 32'b11111111111111111011111010001101;
assign LUT_2[36530] = 32'b00000000000000000101111010110000;
assign LUT_2[36531] = 32'b00000000000000000010110011001001;
assign LUT_2[36532] = 32'b11111111111111111011011111011100;
assign LUT_2[36533] = 32'b11111111111111111000010111110101;
assign LUT_2[36534] = 32'b00000000000000000010011000011000;
assign LUT_2[36535] = 32'b11111111111111111111010000110001;
assign LUT_2[36536] = 32'b11111111111111111001110011010001;
assign LUT_2[36537] = 32'b11111111111111110110101011101010;
assign LUT_2[36538] = 32'b00000000000000000000101100001101;
assign LUT_2[36539] = 32'b11111111111111111101100100100110;
assign LUT_2[36540] = 32'b11111111111111110110010000111001;
assign LUT_2[36541] = 32'b11111111111111110011001001010010;
assign LUT_2[36542] = 32'b11111111111111111101001001110101;
assign LUT_2[36543] = 32'b11111111111111111010000010001110;
assign LUT_2[36544] = 32'b11111111111111111100001010100100;
assign LUT_2[36545] = 32'b11111111111111111001000010111101;
assign LUT_2[36546] = 32'b00000000000000000011000011100000;
assign LUT_2[36547] = 32'b11111111111111111111111011111001;
assign LUT_2[36548] = 32'b11111111111111111000101000001100;
assign LUT_2[36549] = 32'b11111111111111110101100000100101;
assign LUT_2[36550] = 32'b11111111111111111111100001001000;
assign LUT_2[36551] = 32'b11111111111111111100011001100001;
assign LUT_2[36552] = 32'b11111111111111110110111100000001;
assign LUT_2[36553] = 32'b11111111111111110011110100011010;
assign LUT_2[36554] = 32'b11111111111111111101110100111101;
assign LUT_2[36555] = 32'b11111111111111111010101101010110;
assign LUT_2[36556] = 32'b11111111111111110011011001101001;
assign LUT_2[36557] = 32'b11111111111111110000010010000010;
assign LUT_2[36558] = 32'b11111111111111111010010010100101;
assign LUT_2[36559] = 32'b11111111111111110111001010111110;
assign LUT_2[36560] = 32'b11111111111111110110101110101110;
assign LUT_2[36561] = 32'b11111111111111110011100111000111;
assign LUT_2[36562] = 32'b11111111111111111101100111101010;
assign LUT_2[36563] = 32'b11111111111111111010100000000011;
assign LUT_2[36564] = 32'b11111111111111110011001100010110;
assign LUT_2[36565] = 32'b11111111111111110000000100101111;
assign LUT_2[36566] = 32'b11111111111111111010000101010010;
assign LUT_2[36567] = 32'b11111111111111110110111101101011;
assign LUT_2[36568] = 32'b11111111111111110001100000001011;
assign LUT_2[36569] = 32'b11111111111111101110011000100100;
assign LUT_2[36570] = 32'b11111111111111111000011001000111;
assign LUT_2[36571] = 32'b11111111111111110101010001100000;
assign LUT_2[36572] = 32'b11111111111111101101111101110011;
assign LUT_2[36573] = 32'b11111111111111101010110110001100;
assign LUT_2[36574] = 32'b11111111111111110100110110101111;
assign LUT_2[36575] = 32'b11111111111111110001101111001000;
assign LUT_2[36576] = 32'b11111111111111111100100110001101;
assign LUT_2[36577] = 32'b11111111111111111001011110100110;
assign LUT_2[36578] = 32'b00000000000000000011011111001001;
assign LUT_2[36579] = 32'b00000000000000000000010111100010;
assign LUT_2[36580] = 32'b11111111111111111001000011110101;
assign LUT_2[36581] = 32'b11111111111111110101111100001110;
assign LUT_2[36582] = 32'b11111111111111111111111100110001;
assign LUT_2[36583] = 32'b11111111111111111100110101001010;
assign LUT_2[36584] = 32'b11111111111111110111010111101010;
assign LUT_2[36585] = 32'b11111111111111110100010000000011;
assign LUT_2[36586] = 32'b11111111111111111110010000100110;
assign LUT_2[36587] = 32'b11111111111111111011001000111111;
assign LUT_2[36588] = 32'b11111111111111110011110101010010;
assign LUT_2[36589] = 32'b11111111111111110000101101101011;
assign LUT_2[36590] = 32'b11111111111111111010101110001110;
assign LUT_2[36591] = 32'b11111111111111110111100110100111;
assign LUT_2[36592] = 32'b11111111111111110111001010010111;
assign LUT_2[36593] = 32'b11111111111111110100000010110000;
assign LUT_2[36594] = 32'b11111111111111111110000011010011;
assign LUT_2[36595] = 32'b11111111111111111010111011101100;
assign LUT_2[36596] = 32'b11111111111111110011100111111111;
assign LUT_2[36597] = 32'b11111111111111110000100000011000;
assign LUT_2[36598] = 32'b11111111111111111010100000111011;
assign LUT_2[36599] = 32'b11111111111111110111011001010100;
assign LUT_2[36600] = 32'b11111111111111110001111011110100;
assign LUT_2[36601] = 32'b11111111111111101110110100001101;
assign LUT_2[36602] = 32'b11111111111111111000110100110000;
assign LUT_2[36603] = 32'b11111111111111110101101101001001;
assign LUT_2[36604] = 32'b11111111111111101110011001011100;
assign LUT_2[36605] = 32'b11111111111111101011010001110101;
assign LUT_2[36606] = 32'b11111111111111110101010010011000;
assign LUT_2[36607] = 32'b11111111111111110010001010110001;
assign LUT_2[36608] = 32'b00000000000000000011101100011000;
assign LUT_2[36609] = 32'b00000000000000000000100100110001;
assign LUT_2[36610] = 32'b00000000000000001010100101010100;
assign LUT_2[36611] = 32'b00000000000000000111011101101101;
assign LUT_2[36612] = 32'b00000000000000000000001010000000;
assign LUT_2[36613] = 32'b11111111111111111101000010011001;
assign LUT_2[36614] = 32'b00000000000000000111000010111100;
assign LUT_2[36615] = 32'b00000000000000000011111011010101;
assign LUT_2[36616] = 32'b11111111111111111110011101110101;
assign LUT_2[36617] = 32'b11111111111111111011010110001110;
assign LUT_2[36618] = 32'b00000000000000000101010110110001;
assign LUT_2[36619] = 32'b00000000000000000010001111001010;
assign LUT_2[36620] = 32'b11111111111111111010111011011101;
assign LUT_2[36621] = 32'b11111111111111110111110011110110;
assign LUT_2[36622] = 32'b00000000000000000001110100011001;
assign LUT_2[36623] = 32'b11111111111111111110101100110010;
assign LUT_2[36624] = 32'b11111111111111111110010000100010;
assign LUT_2[36625] = 32'b11111111111111111011001000111011;
assign LUT_2[36626] = 32'b00000000000000000101001001011110;
assign LUT_2[36627] = 32'b00000000000000000010000001110111;
assign LUT_2[36628] = 32'b11111111111111111010101110001010;
assign LUT_2[36629] = 32'b11111111111111110111100110100011;
assign LUT_2[36630] = 32'b00000000000000000001100111000110;
assign LUT_2[36631] = 32'b11111111111111111110011111011111;
assign LUT_2[36632] = 32'b11111111111111111001000001111111;
assign LUT_2[36633] = 32'b11111111111111110101111010011000;
assign LUT_2[36634] = 32'b11111111111111111111111010111011;
assign LUT_2[36635] = 32'b11111111111111111100110011010100;
assign LUT_2[36636] = 32'b11111111111111110101011111100111;
assign LUT_2[36637] = 32'b11111111111111110010011000000000;
assign LUT_2[36638] = 32'b11111111111111111100011000100011;
assign LUT_2[36639] = 32'b11111111111111111001010000111100;
assign LUT_2[36640] = 32'b00000000000000000100001000000001;
assign LUT_2[36641] = 32'b00000000000000000001000000011010;
assign LUT_2[36642] = 32'b00000000000000001011000000111101;
assign LUT_2[36643] = 32'b00000000000000000111111001010110;
assign LUT_2[36644] = 32'b00000000000000000000100101101001;
assign LUT_2[36645] = 32'b11111111111111111101011110000010;
assign LUT_2[36646] = 32'b00000000000000000111011110100101;
assign LUT_2[36647] = 32'b00000000000000000100010110111110;
assign LUT_2[36648] = 32'b11111111111111111110111001011110;
assign LUT_2[36649] = 32'b11111111111111111011110001110111;
assign LUT_2[36650] = 32'b00000000000000000101110010011010;
assign LUT_2[36651] = 32'b00000000000000000010101010110011;
assign LUT_2[36652] = 32'b11111111111111111011010111000110;
assign LUT_2[36653] = 32'b11111111111111111000001111011111;
assign LUT_2[36654] = 32'b00000000000000000010010000000010;
assign LUT_2[36655] = 32'b11111111111111111111001000011011;
assign LUT_2[36656] = 32'b11111111111111111110101100001011;
assign LUT_2[36657] = 32'b11111111111111111011100100100100;
assign LUT_2[36658] = 32'b00000000000000000101100101000111;
assign LUT_2[36659] = 32'b00000000000000000010011101100000;
assign LUT_2[36660] = 32'b11111111111111111011001001110011;
assign LUT_2[36661] = 32'b11111111111111111000000010001100;
assign LUT_2[36662] = 32'b00000000000000000010000010101111;
assign LUT_2[36663] = 32'b11111111111111111110111011001000;
assign LUT_2[36664] = 32'b11111111111111111001011101101000;
assign LUT_2[36665] = 32'b11111111111111110110010110000001;
assign LUT_2[36666] = 32'b00000000000000000000010110100100;
assign LUT_2[36667] = 32'b11111111111111111101001110111101;
assign LUT_2[36668] = 32'b11111111111111110101111011010000;
assign LUT_2[36669] = 32'b11111111111111110010110011101001;
assign LUT_2[36670] = 32'b11111111111111111100110100001100;
assign LUT_2[36671] = 32'b11111111111111111001101100100101;
assign LUT_2[36672] = 32'b11111111111111111011110100111011;
assign LUT_2[36673] = 32'b11111111111111111000101101010100;
assign LUT_2[36674] = 32'b00000000000000000010101101110111;
assign LUT_2[36675] = 32'b11111111111111111111100110010000;
assign LUT_2[36676] = 32'b11111111111111111000010010100011;
assign LUT_2[36677] = 32'b11111111111111110101001010111100;
assign LUT_2[36678] = 32'b11111111111111111111001011011111;
assign LUT_2[36679] = 32'b11111111111111111100000011111000;
assign LUT_2[36680] = 32'b11111111111111110110100110011000;
assign LUT_2[36681] = 32'b11111111111111110011011110110001;
assign LUT_2[36682] = 32'b11111111111111111101011111010100;
assign LUT_2[36683] = 32'b11111111111111111010010111101101;
assign LUT_2[36684] = 32'b11111111111111110011000100000000;
assign LUT_2[36685] = 32'b11111111111111101111111100011001;
assign LUT_2[36686] = 32'b11111111111111111001111100111100;
assign LUT_2[36687] = 32'b11111111111111110110110101010101;
assign LUT_2[36688] = 32'b11111111111111110110011001000101;
assign LUT_2[36689] = 32'b11111111111111110011010001011110;
assign LUT_2[36690] = 32'b11111111111111111101010010000001;
assign LUT_2[36691] = 32'b11111111111111111010001010011010;
assign LUT_2[36692] = 32'b11111111111111110010110110101101;
assign LUT_2[36693] = 32'b11111111111111101111101111000110;
assign LUT_2[36694] = 32'b11111111111111111001101111101001;
assign LUT_2[36695] = 32'b11111111111111110110101000000010;
assign LUT_2[36696] = 32'b11111111111111110001001010100010;
assign LUT_2[36697] = 32'b11111111111111101110000010111011;
assign LUT_2[36698] = 32'b11111111111111111000000011011110;
assign LUT_2[36699] = 32'b11111111111111110100111011110111;
assign LUT_2[36700] = 32'b11111111111111101101101000001010;
assign LUT_2[36701] = 32'b11111111111111101010100000100011;
assign LUT_2[36702] = 32'b11111111111111110100100001000110;
assign LUT_2[36703] = 32'b11111111111111110001011001011111;
assign LUT_2[36704] = 32'b11111111111111111100010000100100;
assign LUT_2[36705] = 32'b11111111111111111001001000111101;
assign LUT_2[36706] = 32'b00000000000000000011001001100000;
assign LUT_2[36707] = 32'b00000000000000000000000001111001;
assign LUT_2[36708] = 32'b11111111111111111000101110001100;
assign LUT_2[36709] = 32'b11111111111111110101100110100101;
assign LUT_2[36710] = 32'b11111111111111111111100111001000;
assign LUT_2[36711] = 32'b11111111111111111100011111100001;
assign LUT_2[36712] = 32'b11111111111111110111000010000001;
assign LUT_2[36713] = 32'b11111111111111110011111010011010;
assign LUT_2[36714] = 32'b11111111111111111101111010111101;
assign LUT_2[36715] = 32'b11111111111111111010110011010110;
assign LUT_2[36716] = 32'b11111111111111110011011111101001;
assign LUT_2[36717] = 32'b11111111111111110000011000000010;
assign LUT_2[36718] = 32'b11111111111111111010011000100101;
assign LUT_2[36719] = 32'b11111111111111110111010000111110;
assign LUT_2[36720] = 32'b11111111111111110110110100101110;
assign LUT_2[36721] = 32'b11111111111111110011101101000111;
assign LUT_2[36722] = 32'b11111111111111111101101101101010;
assign LUT_2[36723] = 32'b11111111111111111010100110000011;
assign LUT_2[36724] = 32'b11111111111111110011010010010110;
assign LUT_2[36725] = 32'b11111111111111110000001010101111;
assign LUT_2[36726] = 32'b11111111111111111010001011010010;
assign LUT_2[36727] = 32'b11111111111111110111000011101011;
assign LUT_2[36728] = 32'b11111111111111110001100110001011;
assign LUT_2[36729] = 32'b11111111111111101110011110100100;
assign LUT_2[36730] = 32'b11111111111111111000011111000111;
assign LUT_2[36731] = 32'b11111111111111110101010111100000;
assign LUT_2[36732] = 32'b11111111111111101110000011110011;
assign LUT_2[36733] = 32'b11111111111111101010111100001100;
assign LUT_2[36734] = 32'b11111111111111110100111100101111;
assign LUT_2[36735] = 32'b11111111111111110001110101001000;
assign LUT_2[36736] = 32'b00000000000000001000000000100111;
assign LUT_2[36737] = 32'b00000000000000000100111001000000;
assign LUT_2[36738] = 32'b00000000000000001110111001100011;
assign LUT_2[36739] = 32'b00000000000000001011110001111100;
assign LUT_2[36740] = 32'b00000000000000000100011110001111;
assign LUT_2[36741] = 32'b00000000000000000001010110101000;
assign LUT_2[36742] = 32'b00000000000000001011010111001011;
assign LUT_2[36743] = 32'b00000000000000001000001111100100;
assign LUT_2[36744] = 32'b00000000000000000010110010000100;
assign LUT_2[36745] = 32'b11111111111111111111101010011101;
assign LUT_2[36746] = 32'b00000000000000001001101011000000;
assign LUT_2[36747] = 32'b00000000000000000110100011011001;
assign LUT_2[36748] = 32'b11111111111111111111001111101100;
assign LUT_2[36749] = 32'b11111111111111111100001000000101;
assign LUT_2[36750] = 32'b00000000000000000110001000101000;
assign LUT_2[36751] = 32'b00000000000000000011000001000001;
assign LUT_2[36752] = 32'b00000000000000000010100100110001;
assign LUT_2[36753] = 32'b11111111111111111111011101001010;
assign LUT_2[36754] = 32'b00000000000000001001011101101101;
assign LUT_2[36755] = 32'b00000000000000000110010110000110;
assign LUT_2[36756] = 32'b11111111111111111111000010011001;
assign LUT_2[36757] = 32'b11111111111111111011111010110010;
assign LUT_2[36758] = 32'b00000000000000000101111011010101;
assign LUT_2[36759] = 32'b00000000000000000010110011101110;
assign LUT_2[36760] = 32'b11111111111111111101010110001110;
assign LUT_2[36761] = 32'b11111111111111111010001110100111;
assign LUT_2[36762] = 32'b00000000000000000100001111001010;
assign LUT_2[36763] = 32'b00000000000000000001000111100011;
assign LUT_2[36764] = 32'b11111111111111111001110011110110;
assign LUT_2[36765] = 32'b11111111111111110110101100001111;
assign LUT_2[36766] = 32'b00000000000000000000101100110010;
assign LUT_2[36767] = 32'b11111111111111111101100101001011;
assign LUT_2[36768] = 32'b00000000000000001000011100010000;
assign LUT_2[36769] = 32'b00000000000000000101010100101001;
assign LUT_2[36770] = 32'b00000000000000001111010101001100;
assign LUT_2[36771] = 32'b00000000000000001100001101100101;
assign LUT_2[36772] = 32'b00000000000000000100111001111000;
assign LUT_2[36773] = 32'b00000000000000000001110010010001;
assign LUT_2[36774] = 32'b00000000000000001011110010110100;
assign LUT_2[36775] = 32'b00000000000000001000101011001101;
assign LUT_2[36776] = 32'b00000000000000000011001101101101;
assign LUT_2[36777] = 32'b00000000000000000000000110000110;
assign LUT_2[36778] = 32'b00000000000000001010000110101001;
assign LUT_2[36779] = 32'b00000000000000000110111111000010;
assign LUT_2[36780] = 32'b11111111111111111111101011010101;
assign LUT_2[36781] = 32'b11111111111111111100100011101110;
assign LUT_2[36782] = 32'b00000000000000000110100100010001;
assign LUT_2[36783] = 32'b00000000000000000011011100101010;
assign LUT_2[36784] = 32'b00000000000000000011000000011010;
assign LUT_2[36785] = 32'b11111111111111111111111000110011;
assign LUT_2[36786] = 32'b00000000000000001001111001010110;
assign LUT_2[36787] = 32'b00000000000000000110110001101111;
assign LUT_2[36788] = 32'b11111111111111111111011110000010;
assign LUT_2[36789] = 32'b11111111111111111100010110011011;
assign LUT_2[36790] = 32'b00000000000000000110010110111110;
assign LUT_2[36791] = 32'b00000000000000000011001111010111;
assign LUT_2[36792] = 32'b11111111111111111101110001110111;
assign LUT_2[36793] = 32'b11111111111111111010101010010000;
assign LUT_2[36794] = 32'b00000000000000000100101010110011;
assign LUT_2[36795] = 32'b00000000000000000001100011001100;
assign LUT_2[36796] = 32'b11111111111111111010001111011111;
assign LUT_2[36797] = 32'b11111111111111110111000111111000;
assign LUT_2[36798] = 32'b00000000000000000001001000011011;
assign LUT_2[36799] = 32'b11111111111111111110000000110100;
assign LUT_2[36800] = 32'b00000000000000000000001001001010;
assign LUT_2[36801] = 32'b11111111111111111101000001100011;
assign LUT_2[36802] = 32'b00000000000000000111000010000110;
assign LUT_2[36803] = 32'b00000000000000000011111010011111;
assign LUT_2[36804] = 32'b11111111111111111100100110110010;
assign LUT_2[36805] = 32'b11111111111111111001011111001011;
assign LUT_2[36806] = 32'b00000000000000000011011111101110;
assign LUT_2[36807] = 32'b00000000000000000000011000000111;
assign LUT_2[36808] = 32'b11111111111111111010111010100111;
assign LUT_2[36809] = 32'b11111111111111110111110011000000;
assign LUT_2[36810] = 32'b00000000000000000001110011100011;
assign LUT_2[36811] = 32'b11111111111111111110101011111100;
assign LUT_2[36812] = 32'b11111111111111110111011000001111;
assign LUT_2[36813] = 32'b11111111111111110100010000101000;
assign LUT_2[36814] = 32'b11111111111111111110010001001011;
assign LUT_2[36815] = 32'b11111111111111111011001001100100;
assign LUT_2[36816] = 32'b11111111111111111010101101010100;
assign LUT_2[36817] = 32'b11111111111111110111100101101101;
assign LUT_2[36818] = 32'b00000000000000000001100110010000;
assign LUT_2[36819] = 32'b11111111111111111110011110101001;
assign LUT_2[36820] = 32'b11111111111111110111001010111100;
assign LUT_2[36821] = 32'b11111111111111110100000011010101;
assign LUT_2[36822] = 32'b11111111111111111110000011111000;
assign LUT_2[36823] = 32'b11111111111111111010111100010001;
assign LUT_2[36824] = 32'b11111111111111110101011110110001;
assign LUT_2[36825] = 32'b11111111111111110010010111001010;
assign LUT_2[36826] = 32'b11111111111111111100010111101101;
assign LUT_2[36827] = 32'b11111111111111111001010000000110;
assign LUT_2[36828] = 32'b11111111111111110001111100011001;
assign LUT_2[36829] = 32'b11111111111111101110110100110010;
assign LUT_2[36830] = 32'b11111111111111111000110101010101;
assign LUT_2[36831] = 32'b11111111111111110101101101101110;
assign LUT_2[36832] = 32'b00000000000000000000100100110011;
assign LUT_2[36833] = 32'b11111111111111111101011101001100;
assign LUT_2[36834] = 32'b00000000000000000111011101101111;
assign LUT_2[36835] = 32'b00000000000000000100010110001000;
assign LUT_2[36836] = 32'b11111111111111111101000010011011;
assign LUT_2[36837] = 32'b11111111111111111001111010110100;
assign LUT_2[36838] = 32'b00000000000000000011111011010111;
assign LUT_2[36839] = 32'b00000000000000000000110011110000;
assign LUT_2[36840] = 32'b11111111111111111011010110010000;
assign LUT_2[36841] = 32'b11111111111111111000001110101001;
assign LUT_2[36842] = 32'b00000000000000000010001111001100;
assign LUT_2[36843] = 32'b11111111111111111111000111100101;
assign LUT_2[36844] = 32'b11111111111111110111110011111000;
assign LUT_2[36845] = 32'b11111111111111110100101100010001;
assign LUT_2[36846] = 32'b11111111111111111110101100110100;
assign LUT_2[36847] = 32'b11111111111111111011100101001101;
assign LUT_2[36848] = 32'b11111111111111111011001000111101;
assign LUT_2[36849] = 32'b11111111111111111000000001010110;
assign LUT_2[36850] = 32'b00000000000000000010000001111001;
assign LUT_2[36851] = 32'b11111111111111111110111010010010;
assign LUT_2[36852] = 32'b11111111111111110111100110100101;
assign LUT_2[36853] = 32'b11111111111111110100011110111110;
assign LUT_2[36854] = 32'b11111111111111111110011111100001;
assign LUT_2[36855] = 32'b11111111111111111011010111111010;
assign LUT_2[36856] = 32'b11111111111111110101111010011010;
assign LUT_2[36857] = 32'b11111111111111110010110010110011;
assign LUT_2[36858] = 32'b11111111111111111100110011010110;
assign LUT_2[36859] = 32'b11111111111111111001101011101111;
assign LUT_2[36860] = 32'b11111111111111110010011000000010;
assign LUT_2[36861] = 32'b11111111111111101111010000011011;
assign LUT_2[36862] = 32'b11111111111111111001010000111110;
assign LUT_2[36863] = 32'b11111111111111110110001001010111;
assign LUT_2[36864] = 32'b11111111111111110111011110001010;
assign LUT_2[36865] = 32'b11111111111111110100010110100011;
assign LUT_2[36866] = 32'b11111111111111111110010111000110;
assign LUT_2[36867] = 32'b11111111111111111011001111011111;
assign LUT_2[36868] = 32'b11111111111111110011111011110010;
assign LUT_2[36869] = 32'b11111111111111110000110100001011;
assign LUT_2[36870] = 32'b11111111111111111010110100101110;
assign LUT_2[36871] = 32'b11111111111111110111101101000111;
assign LUT_2[36872] = 32'b11111111111111110010001111100111;
assign LUT_2[36873] = 32'b11111111111111101111001000000000;
assign LUT_2[36874] = 32'b11111111111111111001001000100011;
assign LUT_2[36875] = 32'b11111111111111110110000000111100;
assign LUT_2[36876] = 32'b11111111111111101110101101001111;
assign LUT_2[36877] = 32'b11111111111111101011100101101000;
assign LUT_2[36878] = 32'b11111111111111110101100110001011;
assign LUT_2[36879] = 32'b11111111111111110010011110100100;
assign LUT_2[36880] = 32'b11111111111111110010000010010100;
assign LUT_2[36881] = 32'b11111111111111101110111010101101;
assign LUT_2[36882] = 32'b11111111111111111000111011010000;
assign LUT_2[36883] = 32'b11111111111111110101110011101001;
assign LUT_2[36884] = 32'b11111111111111101110011111111100;
assign LUT_2[36885] = 32'b11111111111111101011011000010101;
assign LUT_2[36886] = 32'b11111111111111110101011000111000;
assign LUT_2[36887] = 32'b11111111111111110010010001010001;
assign LUT_2[36888] = 32'b11111111111111101100110011110001;
assign LUT_2[36889] = 32'b11111111111111101001101100001010;
assign LUT_2[36890] = 32'b11111111111111110011101100101101;
assign LUT_2[36891] = 32'b11111111111111110000100101000110;
assign LUT_2[36892] = 32'b11111111111111101001010001011001;
assign LUT_2[36893] = 32'b11111111111111100110001001110010;
assign LUT_2[36894] = 32'b11111111111111110000001010010101;
assign LUT_2[36895] = 32'b11111111111111101101000010101110;
assign LUT_2[36896] = 32'b11111111111111110111111001110011;
assign LUT_2[36897] = 32'b11111111111111110100110010001100;
assign LUT_2[36898] = 32'b11111111111111111110110010101111;
assign LUT_2[36899] = 32'b11111111111111111011101011001000;
assign LUT_2[36900] = 32'b11111111111111110100010111011011;
assign LUT_2[36901] = 32'b11111111111111110001001111110100;
assign LUT_2[36902] = 32'b11111111111111111011010000010111;
assign LUT_2[36903] = 32'b11111111111111111000001000110000;
assign LUT_2[36904] = 32'b11111111111111110010101011010000;
assign LUT_2[36905] = 32'b11111111111111101111100011101001;
assign LUT_2[36906] = 32'b11111111111111111001100100001100;
assign LUT_2[36907] = 32'b11111111111111110110011100100101;
assign LUT_2[36908] = 32'b11111111111111101111001000111000;
assign LUT_2[36909] = 32'b11111111111111101100000001010001;
assign LUT_2[36910] = 32'b11111111111111110110000001110100;
assign LUT_2[36911] = 32'b11111111111111110010111010001101;
assign LUT_2[36912] = 32'b11111111111111110010011101111101;
assign LUT_2[36913] = 32'b11111111111111101111010110010110;
assign LUT_2[36914] = 32'b11111111111111111001010110111001;
assign LUT_2[36915] = 32'b11111111111111110110001111010010;
assign LUT_2[36916] = 32'b11111111111111101110111011100101;
assign LUT_2[36917] = 32'b11111111111111101011110011111110;
assign LUT_2[36918] = 32'b11111111111111110101110100100001;
assign LUT_2[36919] = 32'b11111111111111110010101100111010;
assign LUT_2[36920] = 32'b11111111111111101101001111011010;
assign LUT_2[36921] = 32'b11111111111111101010000111110011;
assign LUT_2[36922] = 32'b11111111111111110100001000010110;
assign LUT_2[36923] = 32'b11111111111111110001000000101111;
assign LUT_2[36924] = 32'b11111111111111101001101101000010;
assign LUT_2[36925] = 32'b11111111111111100110100101011011;
assign LUT_2[36926] = 32'b11111111111111110000100101111110;
assign LUT_2[36927] = 32'b11111111111111101101011110010111;
assign LUT_2[36928] = 32'b11111111111111101111100110101101;
assign LUT_2[36929] = 32'b11111111111111101100011111000110;
assign LUT_2[36930] = 32'b11111111111111110110011111101001;
assign LUT_2[36931] = 32'b11111111111111110011011000000010;
assign LUT_2[36932] = 32'b11111111111111101100000100010101;
assign LUT_2[36933] = 32'b11111111111111101000111100101110;
assign LUT_2[36934] = 32'b11111111111111110010111101010001;
assign LUT_2[36935] = 32'b11111111111111101111110101101010;
assign LUT_2[36936] = 32'b11111111111111101010011000001010;
assign LUT_2[36937] = 32'b11111111111111100111010000100011;
assign LUT_2[36938] = 32'b11111111111111110001010001000110;
assign LUT_2[36939] = 32'b11111111111111101110001001011111;
assign LUT_2[36940] = 32'b11111111111111100110110101110010;
assign LUT_2[36941] = 32'b11111111111111100011101110001011;
assign LUT_2[36942] = 32'b11111111111111101101101110101110;
assign LUT_2[36943] = 32'b11111111111111101010100111000111;
assign LUT_2[36944] = 32'b11111111111111101010001010110111;
assign LUT_2[36945] = 32'b11111111111111100111000011010000;
assign LUT_2[36946] = 32'b11111111111111110001000011110011;
assign LUT_2[36947] = 32'b11111111111111101101111100001100;
assign LUT_2[36948] = 32'b11111111111111100110101000011111;
assign LUT_2[36949] = 32'b11111111111111100011100000111000;
assign LUT_2[36950] = 32'b11111111111111101101100001011011;
assign LUT_2[36951] = 32'b11111111111111101010011001110100;
assign LUT_2[36952] = 32'b11111111111111100100111100010100;
assign LUT_2[36953] = 32'b11111111111111100001110100101101;
assign LUT_2[36954] = 32'b11111111111111101011110101010000;
assign LUT_2[36955] = 32'b11111111111111101000101101101001;
assign LUT_2[36956] = 32'b11111111111111100001011001111100;
assign LUT_2[36957] = 32'b11111111111111011110010010010101;
assign LUT_2[36958] = 32'b11111111111111101000010010111000;
assign LUT_2[36959] = 32'b11111111111111100101001011010001;
assign LUT_2[36960] = 32'b11111111111111110000000010010110;
assign LUT_2[36961] = 32'b11111111111111101100111010101111;
assign LUT_2[36962] = 32'b11111111111111110110111011010010;
assign LUT_2[36963] = 32'b11111111111111110011110011101011;
assign LUT_2[36964] = 32'b11111111111111101100011111111110;
assign LUT_2[36965] = 32'b11111111111111101001011000010111;
assign LUT_2[36966] = 32'b11111111111111110011011000111010;
assign LUT_2[36967] = 32'b11111111111111110000010001010011;
assign LUT_2[36968] = 32'b11111111111111101010110011110011;
assign LUT_2[36969] = 32'b11111111111111100111101100001100;
assign LUT_2[36970] = 32'b11111111111111110001101100101111;
assign LUT_2[36971] = 32'b11111111111111101110100101001000;
assign LUT_2[36972] = 32'b11111111111111100111010001011011;
assign LUT_2[36973] = 32'b11111111111111100100001001110100;
assign LUT_2[36974] = 32'b11111111111111101110001010010111;
assign LUT_2[36975] = 32'b11111111111111101011000010110000;
assign LUT_2[36976] = 32'b11111111111111101010100110100000;
assign LUT_2[36977] = 32'b11111111111111100111011110111001;
assign LUT_2[36978] = 32'b11111111111111110001011111011100;
assign LUT_2[36979] = 32'b11111111111111101110010111110101;
assign LUT_2[36980] = 32'b11111111111111100111000100001000;
assign LUT_2[36981] = 32'b11111111111111100011111100100001;
assign LUT_2[36982] = 32'b11111111111111101101111101000100;
assign LUT_2[36983] = 32'b11111111111111101010110101011101;
assign LUT_2[36984] = 32'b11111111111111100101010111111101;
assign LUT_2[36985] = 32'b11111111111111100010010000010110;
assign LUT_2[36986] = 32'b11111111111111101100010000111001;
assign LUT_2[36987] = 32'b11111111111111101001001001010010;
assign LUT_2[36988] = 32'b11111111111111100001110101100101;
assign LUT_2[36989] = 32'b11111111111111011110101101111110;
assign LUT_2[36990] = 32'b11111111111111101000101110100001;
assign LUT_2[36991] = 32'b11111111111111100101100110111010;
assign LUT_2[36992] = 32'b11111111111111111011110010011001;
assign LUT_2[36993] = 32'b11111111111111111000101010110010;
assign LUT_2[36994] = 32'b00000000000000000010101011010101;
assign LUT_2[36995] = 32'b11111111111111111111100011101110;
assign LUT_2[36996] = 32'b11111111111111111000010000000001;
assign LUT_2[36997] = 32'b11111111111111110101001000011010;
assign LUT_2[36998] = 32'b11111111111111111111001000111101;
assign LUT_2[36999] = 32'b11111111111111111100000001010110;
assign LUT_2[37000] = 32'b11111111111111110110100011110110;
assign LUT_2[37001] = 32'b11111111111111110011011100001111;
assign LUT_2[37002] = 32'b11111111111111111101011100110010;
assign LUT_2[37003] = 32'b11111111111111111010010101001011;
assign LUT_2[37004] = 32'b11111111111111110011000001011110;
assign LUT_2[37005] = 32'b11111111111111101111111001110111;
assign LUT_2[37006] = 32'b11111111111111111001111010011010;
assign LUT_2[37007] = 32'b11111111111111110110110010110011;
assign LUT_2[37008] = 32'b11111111111111110110010110100011;
assign LUT_2[37009] = 32'b11111111111111110011001110111100;
assign LUT_2[37010] = 32'b11111111111111111101001111011111;
assign LUT_2[37011] = 32'b11111111111111111010000111111000;
assign LUT_2[37012] = 32'b11111111111111110010110100001011;
assign LUT_2[37013] = 32'b11111111111111101111101100100100;
assign LUT_2[37014] = 32'b11111111111111111001101101000111;
assign LUT_2[37015] = 32'b11111111111111110110100101100000;
assign LUT_2[37016] = 32'b11111111111111110001001000000000;
assign LUT_2[37017] = 32'b11111111111111101110000000011001;
assign LUT_2[37018] = 32'b11111111111111111000000000111100;
assign LUT_2[37019] = 32'b11111111111111110100111001010101;
assign LUT_2[37020] = 32'b11111111111111101101100101101000;
assign LUT_2[37021] = 32'b11111111111111101010011110000001;
assign LUT_2[37022] = 32'b11111111111111110100011110100100;
assign LUT_2[37023] = 32'b11111111111111110001010110111101;
assign LUT_2[37024] = 32'b11111111111111111100001110000010;
assign LUT_2[37025] = 32'b11111111111111111001000110011011;
assign LUT_2[37026] = 32'b00000000000000000011000110111110;
assign LUT_2[37027] = 32'b11111111111111111111111111010111;
assign LUT_2[37028] = 32'b11111111111111111000101011101010;
assign LUT_2[37029] = 32'b11111111111111110101100100000011;
assign LUT_2[37030] = 32'b11111111111111111111100100100110;
assign LUT_2[37031] = 32'b11111111111111111100011100111111;
assign LUT_2[37032] = 32'b11111111111111110110111111011111;
assign LUT_2[37033] = 32'b11111111111111110011110111111000;
assign LUT_2[37034] = 32'b11111111111111111101111000011011;
assign LUT_2[37035] = 32'b11111111111111111010110000110100;
assign LUT_2[37036] = 32'b11111111111111110011011101000111;
assign LUT_2[37037] = 32'b11111111111111110000010101100000;
assign LUT_2[37038] = 32'b11111111111111111010010110000011;
assign LUT_2[37039] = 32'b11111111111111110111001110011100;
assign LUT_2[37040] = 32'b11111111111111110110110010001100;
assign LUT_2[37041] = 32'b11111111111111110011101010100101;
assign LUT_2[37042] = 32'b11111111111111111101101011001000;
assign LUT_2[37043] = 32'b11111111111111111010100011100001;
assign LUT_2[37044] = 32'b11111111111111110011001111110100;
assign LUT_2[37045] = 32'b11111111111111110000001000001101;
assign LUT_2[37046] = 32'b11111111111111111010001000110000;
assign LUT_2[37047] = 32'b11111111111111110111000001001001;
assign LUT_2[37048] = 32'b11111111111111110001100011101001;
assign LUT_2[37049] = 32'b11111111111111101110011100000010;
assign LUT_2[37050] = 32'b11111111111111111000011100100101;
assign LUT_2[37051] = 32'b11111111111111110101010100111110;
assign LUT_2[37052] = 32'b11111111111111101110000001010001;
assign LUT_2[37053] = 32'b11111111111111101010111001101010;
assign LUT_2[37054] = 32'b11111111111111110100111010001101;
assign LUT_2[37055] = 32'b11111111111111110001110010100110;
assign LUT_2[37056] = 32'b11111111111111110011111010111100;
assign LUT_2[37057] = 32'b11111111111111110000110011010101;
assign LUT_2[37058] = 32'b11111111111111111010110011111000;
assign LUT_2[37059] = 32'b11111111111111110111101100010001;
assign LUT_2[37060] = 32'b11111111111111110000011000100100;
assign LUT_2[37061] = 32'b11111111111111101101010000111101;
assign LUT_2[37062] = 32'b11111111111111110111010001100000;
assign LUT_2[37063] = 32'b11111111111111110100001001111001;
assign LUT_2[37064] = 32'b11111111111111101110101100011001;
assign LUT_2[37065] = 32'b11111111111111101011100100110010;
assign LUT_2[37066] = 32'b11111111111111110101100101010101;
assign LUT_2[37067] = 32'b11111111111111110010011101101110;
assign LUT_2[37068] = 32'b11111111111111101011001010000001;
assign LUT_2[37069] = 32'b11111111111111101000000010011010;
assign LUT_2[37070] = 32'b11111111111111110010000010111101;
assign LUT_2[37071] = 32'b11111111111111101110111011010110;
assign LUT_2[37072] = 32'b11111111111111101110011111000110;
assign LUT_2[37073] = 32'b11111111111111101011010111011111;
assign LUT_2[37074] = 32'b11111111111111110101011000000010;
assign LUT_2[37075] = 32'b11111111111111110010010000011011;
assign LUT_2[37076] = 32'b11111111111111101010111100101110;
assign LUT_2[37077] = 32'b11111111111111100111110101000111;
assign LUT_2[37078] = 32'b11111111111111110001110101101010;
assign LUT_2[37079] = 32'b11111111111111101110101110000011;
assign LUT_2[37080] = 32'b11111111111111101001010000100011;
assign LUT_2[37081] = 32'b11111111111111100110001000111100;
assign LUT_2[37082] = 32'b11111111111111110000001001011111;
assign LUT_2[37083] = 32'b11111111111111101101000001111000;
assign LUT_2[37084] = 32'b11111111111111100101101110001011;
assign LUT_2[37085] = 32'b11111111111111100010100110100100;
assign LUT_2[37086] = 32'b11111111111111101100100111000111;
assign LUT_2[37087] = 32'b11111111111111101001011111100000;
assign LUT_2[37088] = 32'b11111111111111110100010110100101;
assign LUT_2[37089] = 32'b11111111111111110001001110111110;
assign LUT_2[37090] = 32'b11111111111111111011001111100001;
assign LUT_2[37091] = 32'b11111111111111111000000111111010;
assign LUT_2[37092] = 32'b11111111111111110000110100001101;
assign LUT_2[37093] = 32'b11111111111111101101101100100110;
assign LUT_2[37094] = 32'b11111111111111110111101101001001;
assign LUT_2[37095] = 32'b11111111111111110100100101100010;
assign LUT_2[37096] = 32'b11111111111111101111001000000010;
assign LUT_2[37097] = 32'b11111111111111101100000000011011;
assign LUT_2[37098] = 32'b11111111111111110110000000111110;
assign LUT_2[37099] = 32'b11111111111111110010111001010111;
assign LUT_2[37100] = 32'b11111111111111101011100101101010;
assign LUT_2[37101] = 32'b11111111111111101000011110000011;
assign LUT_2[37102] = 32'b11111111111111110010011110100110;
assign LUT_2[37103] = 32'b11111111111111101111010110111111;
assign LUT_2[37104] = 32'b11111111111111101110111010101111;
assign LUT_2[37105] = 32'b11111111111111101011110011001000;
assign LUT_2[37106] = 32'b11111111111111110101110011101011;
assign LUT_2[37107] = 32'b11111111111111110010101100000100;
assign LUT_2[37108] = 32'b11111111111111101011011000010111;
assign LUT_2[37109] = 32'b11111111111111101000010000110000;
assign LUT_2[37110] = 32'b11111111111111110010010001010011;
assign LUT_2[37111] = 32'b11111111111111101111001001101100;
assign LUT_2[37112] = 32'b11111111111111101001101100001100;
assign LUT_2[37113] = 32'b11111111111111100110100100100101;
assign LUT_2[37114] = 32'b11111111111111110000100101001000;
assign LUT_2[37115] = 32'b11111111111111101101011101100001;
assign LUT_2[37116] = 32'b11111111111111100110001001110100;
assign LUT_2[37117] = 32'b11111111111111100011000010001101;
assign LUT_2[37118] = 32'b11111111111111101101000010110000;
assign LUT_2[37119] = 32'b11111111111111101001111011001001;
assign LUT_2[37120] = 32'b11111111111111111011011100110000;
assign LUT_2[37121] = 32'b11111111111111111000010101001001;
assign LUT_2[37122] = 32'b00000000000000000010010101101100;
assign LUT_2[37123] = 32'b11111111111111111111001110000101;
assign LUT_2[37124] = 32'b11111111111111110111111010011000;
assign LUT_2[37125] = 32'b11111111111111110100110010110001;
assign LUT_2[37126] = 32'b11111111111111111110110011010100;
assign LUT_2[37127] = 32'b11111111111111111011101011101101;
assign LUT_2[37128] = 32'b11111111111111110110001110001101;
assign LUT_2[37129] = 32'b11111111111111110011000110100110;
assign LUT_2[37130] = 32'b11111111111111111101000111001001;
assign LUT_2[37131] = 32'b11111111111111111001111111100010;
assign LUT_2[37132] = 32'b11111111111111110010101011110101;
assign LUT_2[37133] = 32'b11111111111111101111100100001110;
assign LUT_2[37134] = 32'b11111111111111111001100100110001;
assign LUT_2[37135] = 32'b11111111111111110110011101001010;
assign LUT_2[37136] = 32'b11111111111111110110000000111010;
assign LUT_2[37137] = 32'b11111111111111110010111001010011;
assign LUT_2[37138] = 32'b11111111111111111100111001110110;
assign LUT_2[37139] = 32'b11111111111111111001110010001111;
assign LUT_2[37140] = 32'b11111111111111110010011110100010;
assign LUT_2[37141] = 32'b11111111111111101111010110111011;
assign LUT_2[37142] = 32'b11111111111111111001010111011110;
assign LUT_2[37143] = 32'b11111111111111110110001111110111;
assign LUT_2[37144] = 32'b11111111111111110000110010010111;
assign LUT_2[37145] = 32'b11111111111111101101101010110000;
assign LUT_2[37146] = 32'b11111111111111110111101011010011;
assign LUT_2[37147] = 32'b11111111111111110100100011101100;
assign LUT_2[37148] = 32'b11111111111111101101001111111111;
assign LUT_2[37149] = 32'b11111111111111101010001000011000;
assign LUT_2[37150] = 32'b11111111111111110100001000111011;
assign LUT_2[37151] = 32'b11111111111111110001000001010100;
assign LUT_2[37152] = 32'b11111111111111111011111000011001;
assign LUT_2[37153] = 32'b11111111111111111000110000110010;
assign LUT_2[37154] = 32'b00000000000000000010110001010101;
assign LUT_2[37155] = 32'b11111111111111111111101001101110;
assign LUT_2[37156] = 32'b11111111111111111000010110000001;
assign LUT_2[37157] = 32'b11111111111111110101001110011010;
assign LUT_2[37158] = 32'b11111111111111111111001110111101;
assign LUT_2[37159] = 32'b11111111111111111100000111010110;
assign LUT_2[37160] = 32'b11111111111111110110101001110110;
assign LUT_2[37161] = 32'b11111111111111110011100010001111;
assign LUT_2[37162] = 32'b11111111111111111101100010110010;
assign LUT_2[37163] = 32'b11111111111111111010011011001011;
assign LUT_2[37164] = 32'b11111111111111110011000111011110;
assign LUT_2[37165] = 32'b11111111111111101111111111110111;
assign LUT_2[37166] = 32'b11111111111111111010000000011010;
assign LUT_2[37167] = 32'b11111111111111110110111000110011;
assign LUT_2[37168] = 32'b11111111111111110110011100100011;
assign LUT_2[37169] = 32'b11111111111111110011010100111100;
assign LUT_2[37170] = 32'b11111111111111111101010101011111;
assign LUT_2[37171] = 32'b11111111111111111010001101111000;
assign LUT_2[37172] = 32'b11111111111111110010111010001011;
assign LUT_2[37173] = 32'b11111111111111101111110010100100;
assign LUT_2[37174] = 32'b11111111111111111001110011000111;
assign LUT_2[37175] = 32'b11111111111111110110101011100000;
assign LUT_2[37176] = 32'b11111111111111110001001110000000;
assign LUT_2[37177] = 32'b11111111111111101110000110011001;
assign LUT_2[37178] = 32'b11111111111111111000000110111100;
assign LUT_2[37179] = 32'b11111111111111110100111111010101;
assign LUT_2[37180] = 32'b11111111111111101101101011101000;
assign LUT_2[37181] = 32'b11111111111111101010100100000001;
assign LUT_2[37182] = 32'b11111111111111110100100100100100;
assign LUT_2[37183] = 32'b11111111111111110001011100111101;
assign LUT_2[37184] = 32'b11111111111111110011100101010011;
assign LUT_2[37185] = 32'b11111111111111110000011101101100;
assign LUT_2[37186] = 32'b11111111111111111010011110001111;
assign LUT_2[37187] = 32'b11111111111111110111010110101000;
assign LUT_2[37188] = 32'b11111111111111110000000010111011;
assign LUT_2[37189] = 32'b11111111111111101100111011010100;
assign LUT_2[37190] = 32'b11111111111111110110111011110111;
assign LUT_2[37191] = 32'b11111111111111110011110100010000;
assign LUT_2[37192] = 32'b11111111111111101110010110110000;
assign LUT_2[37193] = 32'b11111111111111101011001111001001;
assign LUT_2[37194] = 32'b11111111111111110101001111101100;
assign LUT_2[37195] = 32'b11111111111111110010001000000101;
assign LUT_2[37196] = 32'b11111111111111101010110100011000;
assign LUT_2[37197] = 32'b11111111111111100111101100110001;
assign LUT_2[37198] = 32'b11111111111111110001101101010100;
assign LUT_2[37199] = 32'b11111111111111101110100101101101;
assign LUT_2[37200] = 32'b11111111111111101110001001011101;
assign LUT_2[37201] = 32'b11111111111111101011000001110110;
assign LUT_2[37202] = 32'b11111111111111110101000010011001;
assign LUT_2[37203] = 32'b11111111111111110001111010110010;
assign LUT_2[37204] = 32'b11111111111111101010100111000101;
assign LUT_2[37205] = 32'b11111111111111100111011111011110;
assign LUT_2[37206] = 32'b11111111111111110001100000000001;
assign LUT_2[37207] = 32'b11111111111111101110011000011010;
assign LUT_2[37208] = 32'b11111111111111101000111010111010;
assign LUT_2[37209] = 32'b11111111111111100101110011010011;
assign LUT_2[37210] = 32'b11111111111111101111110011110110;
assign LUT_2[37211] = 32'b11111111111111101100101100001111;
assign LUT_2[37212] = 32'b11111111111111100101011000100010;
assign LUT_2[37213] = 32'b11111111111111100010010000111011;
assign LUT_2[37214] = 32'b11111111111111101100010001011110;
assign LUT_2[37215] = 32'b11111111111111101001001001110111;
assign LUT_2[37216] = 32'b11111111111111110100000000111100;
assign LUT_2[37217] = 32'b11111111111111110000111001010101;
assign LUT_2[37218] = 32'b11111111111111111010111001111000;
assign LUT_2[37219] = 32'b11111111111111110111110010010001;
assign LUT_2[37220] = 32'b11111111111111110000011110100100;
assign LUT_2[37221] = 32'b11111111111111101101010110111101;
assign LUT_2[37222] = 32'b11111111111111110111010111100000;
assign LUT_2[37223] = 32'b11111111111111110100001111111001;
assign LUT_2[37224] = 32'b11111111111111101110110010011001;
assign LUT_2[37225] = 32'b11111111111111101011101010110010;
assign LUT_2[37226] = 32'b11111111111111110101101011010101;
assign LUT_2[37227] = 32'b11111111111111110010100011101110;
assign LUT_2[37228] = 32'b11111111111111101011010000000001;
assign LUT_2[37229] = 32'b11111111111111101000001000011010;
assign LUT_2[37230] = 32'b11111111111111110010001000111101;
assign LUT_2[37231] = 32'b11111111111111101111000001010110;
assign LUT_2[37232] = 32'b11111111111111101110100101000110;
assign LUT_2[37233] = 32'b11111111111111101011011101011111;
assign LUT_2[37234] = 32'b11111111111111110101011110000010;
assign LUT_2[37235] = 32'b11111111111111110010010110011011;
assign LUT_2[37236] = 32'b11111111111111101011000010101110;
assign LUT_2[37237] = 32'b11111111111111100111111011000111;
assign LUT_2[37238] = 32'b11111111111111110001111011101010;
assign LUT_2[37239] = 32'b11111111111111101110110100000011;
assign LUT_2[37240] = 32'b11111111111111101001010110100011;
assign LUT_2[37241] = 32'b11111111111111100110001110111100;
assign LUT_2[37242] = 32'b11111111111111110000001111011111;
assign LUT_2[37243] = 32'b11111111111111101101000111111000;
assign LUT_2[37244] = 32'b11111111111111100101110100001011;
assign LUT_2[37245] = 32'b11111111111111100010101100100100;
assign LUT_2[37246] = 32'b11111111111111101100101101000111;
assign LUT_2[37247] = 32'b11111111111111101001100101100000;
assign LUT_2[37248] = 32'b11111111111111111111110000111111;
assign LUT_2[37249] = 32'b11111111111111111100101001011000;
assign LUT_2[37250] = 32'b00000000000000000110101001111011;
assign LUT_2[37251] = 32'b00000000000000000011100010010100;
assign LUT_2[37252] = 32'b11111111111111111100001110100111;
assign LUT_2[37253] = 32'b11111111111111111001000111000000;
assign LUT_2[37254] = 32'b00000000000000000011000111100011;
assign LUT_2[37255] = 32'b11111111111111111111111111111100;
assign LUT_2[37256] = 32'b11111111111111111010100010011100;
assign LUT_2[37257] = 32'b11111111111111110111011010110101;
assign LUT_2[37258] = 32'b00000000000000000001011011011000;
assign LUT_2[37259] = 32'b11111111111111111110010011110001;
assign LUT_2[37260] = 32'b11111111111111110111000000000100;
assign LUT_2[37261] = 32'b11111111111111110011111000011101;
assign LUT_2[37262] = 32'b11111111111111111101111001000000;
assign LUT_2[37263] = 32'b11111111111111111010110001011001;
assign LUT_2[37264] = 32'b11111111111111111010010101001001;
assign LUT_2[37265] = 32'b11111111111111110111001101100010;
assign LUT_2[37266] = 32'b00000000000000000001001110000101;
assign LUT_2[37267] = 32'b11111111111111111110000110011110;
assign LUT_2[37268] = 32'b11111111111111110110110010110001;
assign LUT_2[37269] = 32'b11111111111111110011101011001010;
assign LUT_2[37270] = 32'b11111111111111111101101011101101;
assign LUT_2[37271] = 32'b11111111111111111010100100000110;
assign LUT_2[37272] = 32'b11111111111111110101000110100110;
assign LUT_2[37273] = 32'b11111111111111110001111110111111;
assign LUT_2[37274] = 32'b11111111111111111011111111100010;
assign LUT_2[37275] = 32'b11111111111111111000110111111011;
assign LUT_2[37276] = 32'b11111111111111110001100100001110;
assign LUT_2[37277] = 32'b11111111111111101110011100100111;
assign LUT_2[37278] = 32'b11111111111111111000011101001010;
assign LUT_2[37279] = 32'b11111111111111110101010101100011;
assign LUT_2[37280] = 32'b00000000000000000000001100101000;
assign LUT_2[37281] = 32'b11111111111111111101000101000001;
assign LUT_2[37282] = 32'b00000000000000000111000101100100;
assign LUT_2[37283] = 32'b00000000000000000011111101111101;
assign LUT_2[37284] = 32'b11111111111111111100101010010000;
assign LUT_2[37285] = 32'b11111111111111111001100010101001;
assign LUT_2[37286] = 32'b00000000000000000011100011001100;
assign LUT_2[37287] = 32'b00000000000000000000011011100101;
assign LUT_2[37288] = 32'b11111111111111111010111110000101;
assign LUT_2[37289] = 32'b11111111111111110111110110011110;
assign LUT_2[37290] = 32'b00000000000000000001110111000001;
assign LUT_2[37291] = 32'b11111111111111111110101111011010;
assign LUT_2[37292] = 32'b11111111111111110111011011101101;
assign LUT_2[37293] = 32'b11111111111111110100010100000110;
assign LUT_2[37294] = 32'b11111111111111111110010100101001;
assign LUT_2[37295] = 32'b11111111111111111011001101000010;
assign LUT_2[37296] = 32'b11111111111111111010110000110010;
assign LUT_2[37297] = 32'b11111111111111110111101001001011;
assign LUT_2[37298] = 32'b00000000000000000001101001101110;
assign LUT_2[37299] = 32'b11111111111111111110100010000111;
assign LUT_2[37300] = 32'b11111111111111110111001110011010;
assign LUT_2[37301] = 32'b11111111111111110100000110110011;
assign LUT_2[37302] = 32'b11111111111111111110000111010110;
assign LUT_2[37303] = 32'b11111111111111111010111111101111;
assign LUT_2[37304] = 32'b11111111111111110101100010001111;
assign LUT_2[37305] = 32'b11111111111111110010011010101000;
assign LUT_2[37306] = 32'b11111111111111111100011011001011;
assign LUT_2[37307] = 32'b11111111111111111001010011100100;
assign LUT_2[37308] = 32'b11111111111111110001111111110111;
assign LUT_2[37309] = 32'b11111111111111101110111000010000;
assign LUT_2[37310] = 32'b11111111111111111000111000110011;
assign LUT_2[37311] = 32'b11111111111111110101110001001100;
assign LUT_2[37312] = 32'b11111111111111110111111001100010;
assign LUT_2[37313] = 32'b11111111111111110100110001111011;
assign LUT_2[37314] = 32'b11111111111111111110110010011110;
assign LUT_2[37315] = 32'b11111111111111111011101010110111;
assign LUT_2[37316] = 32'b11111111111111110100010111001010;
assign LUT_2[37317] = 32'b11111111111111110001001111100011;
assign LUT_2[37318] = 32'b11111111111111111011010000000110;
assign LUT_2[37319] = 32'b11111111111111111000001000011111;
assign LUT_2[37320] = 32'b11111111111111110010101010111111;
assign LUT_2[37321] = 32'b11111111111111101111100011011000;
assign LUT_2[37322] = 32'b11111111111111111001100011111011;
assign LUT_2[37323] = 32'b11111111111111110110011100010100;
assign LUT_2[37324] = 32'b11111111111111101111001000100111;
assign LUT_2[37325] = 32'b11111111111111101100000001000000;
assign LUT_2[37326] = 32'b11111111111111110110000001100011;
assign LUT_2[37327] = 32'b11111111111111110010111001111100;
assign LUT_2[37328] = 32'b11111111111111110010011101101100;
assign LUT_2[37329] = 32'b11111111111111101111010110000101;
assign LUT_2[37330] = 32'b11111111111111111001010110101000;
assign LUT_2[37331] = 32'b11111111111111110110001111000001;
assign LUT_2[37332] = 32'b11111111111111101110111011010100;
assign LUT_2[37333] = 32'b11111111111111101011110011101101;
assign LUT_2[37334] = 32'b11111111111111110101110100010000;
assign LUT_2[37335] = 32'b11111111111111110010101100101001;
assign LUT_2[37336] = 32'b11111111111111101101001111001001;
assign LUT_2[37337] = 32'b11111111111111101010000111100010;
assign LUT_2[37338] = 32'b11111111111111110100001000000101;
assign LUT_2[37339] = 32'b11111111111111110001000000011110;
assign LUT_2[37340] = 32'b11111111111111101001101100110001;
assign LUT_2[37341] = 32'b11111111111111100110100101001010;
assign LUT_2[37342] = 32'b11111111111111110000100101101101;
assign LUT_2[37343] = 32'b11111111111111101101011110000110;
assign LUT_2[37344] = 32'b11111111111111111000010101001011;
assign LUT_2[37345] = 32'b11111111111111110101001101100100;
assign LUT_2[37346] = 32'b11111111111111111111001110000111;
assign LUT_2[37347] = 32'b11111111111111111100000110100000;
assign LUT_2[37348] = 32'b11111111111111110100110010110011;
assign LUT_2[37349] = 32'b11111111111111110001101011001100;
assign LUT_2[37350] = 32'b11111111111111111011101011101111;
assign LUT_2[37351] = 32'b11111111111111111000100100001000;
assign LUT_2[37352] = 32'b11111111111111110011000110101000;
assign LUT_2[37353] = 32'b11111111111111101111111111000001;
assign LUT_2[37354] = 32'b11111111111111111001111111100100;
assign LUT_2[37355] = 32'b11111111111111110110110111111101;
assign LUT_2[37356] = 32'b11111111111111101111100100010000;
assign LUT_2[37357] = 32'b11111111111111101100011100101001;
assign LUT_2[37358] = 32'b11111111111111110110011101001100;
assign LUT_2[37359] = 32'b11111111111111110011010101100101;
assign LUT_2[37360] = 32'b11111111111111110010111001010101;
assign LUT_2[37361] = 32'b11111111111111101111110001101110;
assign LUT_2[37362] = 32'b11111111111111111001110010010001;
assign LUT_2[37363] = 32'b11111111111111110110101010101010;
assign LUT_2[37364] = 32'b11111111111111101111010110111101;
assign LUT_2[37365] = 32'b11111111111111101100001111010110;
assign LUT_2[37366] = 32'b11111111111111110110001111111001;
assign LUT_2[37367] = 32'b11111111111111110011001000010010;
assign LUT_2[37368] = 32'b11111111111111101101101010110010;
assign LUT_2[37369] = 32'b11111111111111101010100011001011;
assign LUT_2[37370] = 32'b11111111111111110100100011101110;
assign LUT_2[37371] = 32'b11111111111111110001011100000111;
assign LUT_2[37372] = 32'b11111111111111101010001000011010;
assign LUT_2[37373] = 32'b11111111111111100111000000110011;
assign LUT_2[37374] = 32'b11111111111111110001000001010110;
assign LUT_2[37375] = 32'b11111111111111101101111001101111;
assign LUT_2[37376] = 32'b11111111111111111100001111111100;
assign LUT_2[37377] = 32'b11111111111111111001001000010101;
assign LUT_2[37378] = 32'b00000000000000000011001000111000;
assign LUT_2[37379] = 32'b00000000000000000000000001010001;
assign LUT_2[37380] = 32'b11111111111111111000101101100100;
assign LUT_2[37381] = 32'b11111111111111110101100101111101;
assign LUT_2[37382] = 32'b11111111111111111111100110100000;
assign LUT_2[37383] = 32'b11111111111111111100011110111001;
assign LUT_2[37384] = 32'b11111111111111110111000001011001;
assign LUT_2[37385] = 32'b11111111111111110011111001110010;
assign LUT_2[37386] = 32'b11111111111111111101111010010101;
assign LUT_2[37387] = 32'b11111111111111111010110010101110;
assign LUT_2[37388] = 32'b11111111111111110011011111000001;
assign LUT_2[37389] = 32'b11111111111111110000010111011010;
assign LUT_2[37390] = 32'b11111111111111111010010111111101;
assign LUT_2[37391] = 32'b11111111111111110111010000010110;
assign LUT_2[37392] = 32'b11111111111111110110110100000110;
assign LUT_2[37393] = 32'b11111111111111110011101100011111;
assign LUT_2[37394] = 32'b11111111111111111101101101000010;
assign LUT_2[37395] = 32'b11111111111111111010100101011011;
assign LUT_2[37396] = 32'b11111111111111110011010001101110;
assign LUT_2[37397] = 32'b11111111111111110000001010000111;
assign LUT_2[37398] = 32'b11111111111111111010001010101010;
assign LUT_2[37399] = 32'b11111111111111110111000011000011;
assign LUT_2[37400] = 32'b11111111111111110001100101100011;
assign LUT_2[37401] = 32'b11111111111111101110011101111100;
assign LUT_2[37402] = 32'b11111111111111111000011110011111;
assign LUT_2[37403] = 32'b11111111111111110101010110111000;
assign LUT_2[37404] = 32'b11111111111111101110000011001011;
assign LUT_2[37405] = 32'b11111111111111101010111011100100;
assign LUT_2[37406] = 32'b11111111111111110100111100000111;
assign LUT_2[37407] = 32'b11111111111111110001110100100000;
assign LUT_2[37408] = 32'b11111111111111111100101011100101;
assign LUT_2[37409] = 32'b11111111111111111001100011111110;
assign LUT_2[37410] = 32'b00000000000000000011100100100001;
assign LUT_2[37411] = 32'b00000000000000000000011100111010;
assign LUT_2[37412] = 32'b11111111111111111001001001001101;
assign LUT_2[37413] = 32'b11111111111111110110000001100110;
assign LUT_2[37414] = 32'b00000000000000000000000010001001;
assign LUT_2[37415] = 32'b11111111111111111100111010100010;
assign LUT_2[37416] = 32'b11111111111111110111011101000010;
assign LUT_2[37417] = 32'b11111111111111110100010101011011;
assign LUT_2[37418] = 32'b11111111111111111110010101111110;
assign LUT_2[37419] = 32'b11111111111111111011001110010111;
assign LUT_2[37420] = 32'b11111111111111110011111010101010;
assign LUT_2[37421] = 32'b11111111111111110000110011000011;
assign LUT_2[37422] = 32'b11111111111111111010110011100110;
assign LUT_2[37423] = 32'b11111111111111110111101011111111;
assign LUT_2[37424] = 32'b11111111111111110111001111101111;
assign LUT_2[37425] = 32'b11111111111111110100001000001000;
assign LUT_2[37426] = 32'b11111111111111111110001000101011;
assign LUT_2[37427] = 32'b11111111111111111011000001000100;
assign LUT_2[37428] = 32'b11111111111111110011101101010111;
assign LUT_2[37429] = 32'b11111111111111110000100101110000;
assign LUT_2[37430] = 32'b11111111111111111010100110010011;
assign LUT_2[37431] = 32'b11111111111111110111011110101100;
assign LUT_2[37432] = 32'b11111111111111110010000001001100;
assign LUT_2[37433] = 32'b11111111111111101110111001100101;
assign LUT_2[37434] = 32'b11111111111111111000111010001000;
assign LUT_2[37435] = 32'b11111111111111110101110010100001;
assign LUT_2[37436] = 32'b11111111111111101110011110110100;
assign LUT_2[37437] = 32'b11111111111111101011010111001101;
assign LUT_2[37438] = 32'b11111111111111110101010111110000;
assign LUT_2[37439] = 32'b11111111111111110010010000001001;
assign LUT_2[37440] = 32'b11111111111111110100011000011111;
assign LUT_2[37441] = 32'b11111111111111110001010000111000;
assign LUT_2[37442] = 32'b11111111111111111011010001011011;
assign LUT_2[37443] = 32'b11111111111111111000001001110100;
assign LUT_2[37444] = 32'b11111111111111110000110110000111;
assign LUT_2[37445] = 32'b11111111111111101101101110100000;
assign LUT_2[37446] = 32'b11111111111111110111101111000011;
assign LUT_2[37447] = 32'b11111111111111110100100111011100;
assign LUT_2[37448] = 32'b11111111111111101111001001111100;
assign LUT_2[37449] = 32'b11111111111111101100000010010101;
assign LUT_2[37450] = 32'b11111111111111110110000010111000;
assign LUT_2[37451] = 32'b11111111111111110010111011010001;
assign LUT_2[37452] = 32'b11111111111111101011100111100100;
assign LUT_2[37453] = 32'b11111111111111101000011111111101;
assign LUT_2[37454] = 32'b11111111111111110010100000100000;
assign LUT_2[37455] = 32'b11111111111111101111011000111001;
assign LUT_2[37456] = 32'b11111111111111101110111100101001;
assign LUT_2[37457] = 32'b11111111111111101011110101000010;
assign LUT_2[37458] = 32'b11111111111111110101110101100101;
assign LUT_2[37459] = 32'b11111111111111110010101101111110;
assign LUT_2[37460] = 32'b11111111111111101011011010010001;
assign LUT_2[37461] = 32'b11111111111111101000010010101010;
assign LUT_2[37462] = 32'b11111111111111110010010011001101;
assign LUT_2[37463] = 32'b11111111111111101111001011100110;
assign LUT_2[37464] = 32'b11111111111111101001101110000110;
assign LUT_2[37465] = 32'b11111111111111100110100110011111;
assign LUT_2[37466] = 32'b11111111111111110000100111000010;
assign LUT_2[37467] = 32'b11111111111111101101011111011011;
assign LUT_2[37468] = 32'b11111111111111100110001011101110;
assign LUT_2[37469] = 32'b11111111111111100011000100000111;
assign LUT_2[37470] = 32'b11111111111111101101000100101010;
assign LUT_2[37471] = 32'b11111111111111101001111101000011;
assign LUT_2[37472] = 32'b11111111111111110100110100001000;
assign LUT_2[37473] = 32'b11111111111111110001101100100001;
assign LUT_2[37474] = 32'b11111111111111111011101101000100;
assign LUT_2[37475] = 32'b11111111111111111000100101011101;
assign LUT_2[37476] = 32'b11111111111111110001010001110000;
assign LUT_2[37477] = 32'b11111111111111101110001010001001;
assign LUT_2[37478] = 32'b11111111111111111000001010101100;
assign LUT_2[37479] = 32'b11111111111111110101000011000101;
assign LUT_2[37480] = 32'b11111111111111101111100101100101;
assign LUT_2[37481] = 32'b11111111111111101100011101111110;
assign LUT_2[37482] = 32'b11111111111111110110011110100001;
assign LUT_2[37483] = 32'b11111111111111110011010110111010;
assign LUT_2[37484] = 32'b11111111111111101100000011001101;
assign LUT_2[37485] = 32'b11111111111111101000111011100110;
assign LUT_2[37486] = 32'b11111111111111110010111100001001;
assign LUT_2[37487] = 32'b11111111111111101111110100100010;
assign LUT_2[37488] = 32'b11111111111111101111011000010010;
assign LUT_2[37489] = 32'b11111111111111101100010000101011;
assign LUT_2[37490] = 32'b11111111111111110110010001001110;
assign LUT_2[37491] = 32'b11111111111111110011001001100111;
assign LUT_2[37492] = 32'b11111111111111101011110101111010;
assign LUT_2[37493] = 32'b11111111111111101000101110010011;
assign LUT_2[37494] = 32'b11111111111111110010101110110110;
assign LUT_2[37495] = 32'b11111111111111101111100111001111;
assign LUT_2[37496] = 32'b11111111111111101010001001101111;
assign LUT_2[37497] = 32'b11111111111111100111000010001000;
assign LUT_2[37498] = 32'b11111111111111110001000010101011;
assign LUT_2[37499] = 32'b11111111111111101101111011000100;
assign LUT_2[37500] = 32'b11111111111111100110100111010111;
assign LUT_2[37501] = 32'b11111111111111100011011111110000;
assign LUT_2[37502] = 32'b11111111111111101101100000010011;
assign LUT_2[37503] = 32'b11111111111111101010011000101100;
assign LUT_2[37504] = 32'b00000000000000000000100100001011;
assign LUT_2[37505] = 32'b11111111111111111101011100100100;
assign LUT_2[37506] = 32'b00000000000000000111011101000111;
assign LUT_2[37507] = 32'b00000000000000000100010101100000;
assign LUT_2[37508] = 32'b11111111111111111101000001110011;
assign LUT_2[37509] = 32'b11111111111111111001111010001100;
assign LUT_2[37510] = 32'b00000000000000000011111010101111;
assign LUT_2[37511] = 32'b00000000000000000000110011001000;
assign LUT_2[37512] = 32'b11111111111111111011010101101000;
assign LUT_2[37513] = 32'b11111111111111111000001110000001;
assign LUT_2[37514] = 32'b00000000000000000010001110100100;
assign LUT_2[37515] = 32'b11111111111111111111000110111101;
assign LUT_2[37516] = 32'b11111111111111110111110011010000;
assign LUT_2[37517] = 32'b11111111111111110100101011101001;
assign LUT_2[37518] = 32'b11111111111111111110101100001100;
assign LUT_2[37519] = 32'b11111111111111111011100100100101;
assign LUT_2[37520] = 32'b11111111111111111011001000010101;
assign LUT_2[37521] = 32'b11111111111111111000000000101110;
assign LUT_2[37522] = 32'b00000000000000000010000001010001;
assign LUT_2[37523] = 32'b11111111111111111110111001101010;
assign LUT_2[37524] = 32'b11111111111111110111100101111101;
assign LUT_2[37525] = 32'b11111111111111110100011110010110;
assign LUT_2[37526] = 32'b11111111111111111110011110111001;
assign LUT_2[37527] = 32'b11111111111111111011010111010010;
assign LUT_2[37528] = 32'b11111111111111110101111001110010;
assign LUT_2[37529] = 32'b11111111111111110010110010001011;
assign LUT_2[37530] = 32'b11111111111111111100110010101110;
assign LUT_2[37531] = 32'b11111111111111111001101011000111;
assign LUT_2[37532] = 32'b11111111111111110010010111011010;
assign LUT_2[37533] = 32'b11111111111111101111001111110011;
assign LUT_2[37534] = 32'b11111111111111111001010000010110;
assign LUT_2[37535] = 32'b11111111111111110110001000101111;
assign LUT_2[37536] = 32'b00000000000000000000111111110100;
assign LUT_2[37537] = 32'b11111111111111111101111000001101;
assign LUT_2[37538] = 32'b00000000000000000111111000110000;
assign LUT_2[37539] = 32'b00000000000000000100110001001001;
assign LUT_2[37540] = 32'b11111111111111111101011101011100;
assign LUT_2[37541] = 32'b11111111111111111010010101110101;
assign LUT_2[37542] = 32'b00000000000000000100010110011000;
assign LUT_2[37543] = 32'b00000000000000000001001110110001;
assign LUT_2[37544] = 32'b11111111111111111011110001010001;
assign LUT_2[37545] = 32'b11111111111111111000101001101010;
assign LUT_2[37546] = 32'b00000000000000000010101010001101;
assign LUT_2[37547] = 32'b11111111111111111111100010100110;
assign LUT_2[37548] = 32'b11111111111111111000001110111001;
assign LUT_2[37549] = 32'b11111111111111110101000111010010;
assign LUT_2[37550] = 32'b11111111111111111111000111110101;
assign LUT_2[37551] = 32'b11111111111111111100000000001110;
assign LUT_2[37552] = 32'b11111111111111111011100011111110;
assign LUT_2[37553] = 32'b11111111111111111000011100010111;
assign LUT_2[37554] = 32'b00000000000000000010011100111010;
assign LUT_2[37555] = 32'b11111111111111111111010101010011;
assign LUT_2[37556] = 32'b11111111111111111000000001100110;
assign LUT_2[37557] = 32'b11111111111111110100111001111111;
assign LUT_2[37558] = 32'b11111111111111111110111010100010;
assign LUT_2[37559] = 32'b11111111111111111011110010111011;
assign LUT_2[37560] = 32'b11111111111111110110010101011011;
assign LUT_2[37561] = 32'b11111111111111110011001101110100;
assign LUT_2[37562] = 32'b11111111111111111101001110010111;
assign LUT_2[37563] = 32'b11111111111111111010000110110000;
assign LUT_2[37564] = 32'b11111111111111110010110011000011;
assign LUT_2[37565] = 32'b11111111111111101111101011011100;
assign LUT_2[37566] = 32'b11111111111111111001101011111111;
assign LUT_2[37567] = 32'b11111111111111110110100100011000;
assign LUT_2[37568] = 32'b11111111111111111000101100101110;
assign LUT_2[37569] = 32'b11111111111111110101100101000111;
assign LUT_2[37570] = 32'b11111111111111111111100101101010;
assign LUT_2[37571] = 32'b11111111111111111100011110000011;
assign LUT_2[37572] = 32'b11111111111111110101001010010110;
assign LUT_2[37573] = 32'b11111111111111110010000010101111;
assign LUT_2[37574] = 32'b11111111111111111100000011010010;
assign LUT_2[37575] = 32'b11111111111111111000111011101011;
assign LUT_2[37576] = 32'b11111111111111110011011110001011;
assign LUT_2[37577] = 32'b11111111111111110000010110100100;
assign LUT_2[37578] = 32'b11111111111111111010010111000111;
assign LUT_2[37579] = 32'b11111111111111110111001111100000;
assign LUT_2[37580] = 32'b11111111111111101111111011110011;
assign LUT_2[37581] = 32'b11111111111111101100110100001100;
assign LUT_2[37582] = 32'b11111111111111110110110100101111;
assign LUT_2[37583] = 32'b11111111111111110011101101001000;
assign LUT_2[37584] = 32'b11111111111111110011010000111000;
assign LUT_2[37585] = 32'b11111111111111110000001001010001;
assign LUT_2[37586] = 32'b11111111111111111010001001110100;
assign LUT_2[37587] = 32'b11111111111111110111000010001101;
assign LUT_2[37588] = 32'b11111111111111101111101110100000;
assign LUT_2[37589] = 32'b11111111111111101100100110111001;
assign LUT_2[37590] = 32'b11111111111111110110100111011100;
assign LUT_2[37591] = 32'b11111111111111110011011111110101;
assign LUT_2[37592] = 32'b11111111111111101110000010010101;
assign LUT_2[37593] = 32'b11111111111111101010111010101110;
assign LUT_2[37594] = 32'b11111111111111110100111011010001;
assign LUT_2[37595] = 32'b11111111111111110001110011101010;
assign LUT_2[37596] = 32'b11111111111111101010011111111101;
assign LUT_2[37597] = 32'b11111111111111100111011000010110;
assign LUT_2[37598] = 32'b11111111111111110001011000111001;
assign LUT_2[37599] = 32'b11111111111111101110010001010010;
assign LUT_2[37600] = 32'b11111111111111111001001000010111;
assign LUT_2[37601] = 32'b11111111111111110110000000110000;
assign LUT_2[37602] = 32'b00000000000000000000000001010011;
assign LUT_2[37603] = 32'b11111111111111111100111001101100;
assign LUT_2[37604] = 32'b11111111111111110101100101111111;
assign LUT_2[37605] = 32'b11111111111111110010011110011000;
assign LUT_2[37606] = 32'b11111111111111111100011110111011;
assign LUT_2[37607] = 32'b11111111111111111001010111010100;
assign LUT_2[37608] = 32'b11111111111111110011111001110100;
assign LUT_2[37609] = 32'b11111111111111110000110010001101;
assign LUT_2[37610] = 32'b11111111111111111010110010110000;
assign LUT_2[37611] = 32'b11111111111111110111101011001001;
assign LUT_2[37612] = 32'b11111111111111110000010111011100;
assign LUT_2[37613] = 32'b11111111111111101101001111110101;
assign LUT_2[37614] = 32'b11111111111111110111010000011000;
assign LUT_2[37615] = 32'b11111111111111110100001000110001;
assign LUT_2[37616] = 32'b11111111111111110011101100100001;
assign LUT_2[37617] = 32'b11111111111111110000100100111010;
assign LUT_2[37618] = 32'b11111111111111111010100101011101;
assign LUT_2[37619] = 32'b11111111111111110111011101110110;
assign LUT_2[37620] = 32'b11111111111111110000001010001001;
assign LUT_2[37621] = 32'b11111111111111101101000010100010;
assign LUT_2[37622] = 32'b11111111111111110111000011000101;
assign LUT_2[37623] = 32'b11111111111111110011111011011110;
assign LUT_2[37624] = 32'b11111111111111101110011101111110;
assign LUT_2[37625] = 32'b11111111111111101011010110010111;
assign LUT_2[37626] = 32'b11111111111111110101010110111010;
assign LUT_2[37627] = 32'b11111111111111110010001111010011;
assign LUT_2[37628] = 32'b11111111111111101010111011100110;
assign LUT_2[37629] = 32'b11111111111111100111110011111111;
assign LUT_2[37630] = 32'b11111111111111110001110100100010;
assign LUT_2[37631] = 32'b11111111111111101110101100111011;
assign LUT_2[37632] = 32'b00000000000000000000001110100010;
assign LUT_2[37633] = 32'b11111111111111111101000110111011;
assign LUT_2[37634] = 32'b00000000000000000111000111011110;
assign LUT_2[37635] = 32'b00000000000000000011111111110111;
assign LUT_2[37636] = 32'b11111111111111111100101100001010;
assign LUT_2[37637] = 32'b11111111111111111001100100100011;
assign LUT_2[37638] = 32'b00000000000000000011100101000110;
assign LUT_2[37639] = 32'b00000000000000000000011101011111;
assign LUT_2[37640] = 32'b11111111111111111010111111111111;
assign LUT_2[37641] = 32'b11111111111111110111111000011000;
assign LUT_2[37642] = 32'b00000000000000000001111000111011;
assign LUT_2[37643] = 32'b11111111111111111110110001010100;
assign LUT_2[37644] = 32'b11111111111111110111011101100111;
assign LUT_2[37645] = 32'b11111111111111110100010110000000;
assign LUT_2[37646] = 32'b11111111111111111110010110100011;
assign LUT_2[37647] = 32'b11111111111111111011001110111100;
assign LUT_2[37648] = 32'b11111111111111111010110010101100;
assign LUT_2[37649] = 32'b11111111111111110111101011000101;
assign LUT_2[37650] = 32'b00000000000000000001101011101000;
assign LUT_2[37651] = 32'b11111111111111111110100100000001;
assign LUT_2[37652] = 32'b11111111111111110111010000010100;
assign LUT_2[37653] = 32'b11111111111111110100001000101101;
assign LUT_2[37654] = 32'b11111111111111111110001001010000;
assign LUT_2[37655] = 32'b11111111111111111011000001101001;
assign LUT_2[37656] = 32'b11111111111111110101100100001001;
assign LUT_2[37657] = 32'b11111111111111110010011100100010;
assign LUT_2[37658] = 32'b11111111111111111100011101000101;
assign LUT_2[37659] = 32'b11111111111111111001010101011110;
assign LUT_2[37660] = 32'b11111111111111110010000001110001;
assign LUT_2[37661] = 32'b11111111111111101110111010001010;
assign LUT_2[37662] = 32'b11111111111111111000111010101101;
assign LUT_2[37663] = 32'b11111111111111110101110011000110;
assign LUT_2[37664] = 32'b00000000000000000000101010001011;
assign LUT_2[37665] = 32'b11111111111111111101100010100100;
assign LUT_2[37666] = 32'b00000000000000000111100011000111;
assign LUT_2[37667] = 32'b00000000000000000100011011100000;
assign LUT_2[37668] = 32'b11111111111111111101000111110011;
assign LUT_2[37669] = 32'b11111111111111111010000000001100;
assign LUT_2[37670] = 32'b00000000000000000100000000101111;
assign LUT_2[37671] = 32'b00000000000000000000111001001000;
assign LUT_2[37672] = 32'b11111111111111111011011011101000;
assign LUT_2[37673] = 32'b11111111111111111000010100000001;
assign LUT_2[37674] = 32'b00000000000000000010010100100100;
assign LUT_2[37675] = 32'b11111111111111111111001100111101;
assign LUT_2[37676] = 32'b11111111111111110111111001010000;
assign LUT_2[37677] = 32'b11111111111111110100110001101001;
assign LUT_2[37678] = 32'b11111111111111111110110010001100;
assign LUT_2[37679] = 32'b11111111111111111011101010100101;
assign LUT_2[37680] = 32'b11111111111111111011001110010101;
assign LUT_2[37681] = 32'b11111111111111111000000110101110;
assign LUT_2[37682] = 32'b00000000000000000010000111010001;
assign LUT_2[37683] = 32'b11111111111111111110111111101010;
assign LUT_2[37684] = 32'b11111111111111110111101011111101;
assign LUT_2[37685] = 32'b11111111111111110100100100010110;
assign LUT_2[37686] = 32'b11111111111111111110100100111001;
assign LUT_2[37687] = 32'b11111111111111111011011101010010;
assign LUT_2[37688] = 32'b11111111111111110101111111110010;
assign LUT_2[37689] = 32'b11111111111111110010111000001011;
assign LUT_2[37690] = 32'b11111111111111111100111000101110;
assign LUT_2[37691] = 32'b11111111111111111001110001000111;
assign LUT_2[37692] = 32'b11111111111111110010011101011010;
assign LUT_2[37693] = 32'b11111111111111101111010101110011;
assign LUT_2[37694] = 32'b11111111111111111001010110010110;
assign LUT_2[37695] = 32'b11111111111111110110001110101111;
assign LUT_2[37696] = 32'b11111111111111111000010111000101;
assign LUT_2[37697] = 32'b11111111111111110101001111011110;
assign LUT_2[37698] = 32'b11111111111111111111010000000001;
assign LUT_2[37699] = 32'b11111111111111111100001000011010;
assign LUT_2[37700] = 32'b11111111111111110100110100101101;
assign LUT_2[37701] = 32'b11111111111111110001101101000110;
assign LUT_2[37702] = 32'b11111111111111111011101101101001;
assign LUT_2[37703] = 32'b11111111111111111000100110000010;
assign LUT_2[37704] = 32'b11111111111111110011001000100010;
assign LUT_2[37705] = 32'b11111111111111110000000000111011;
assign LUT_2[37706] = 32'b11111111111111111010000001011110;
assign LUT_2[37707] = 32'b11111111111111110110111001110111;
assign LUT_2[37708] = 32'b11111111111111101111100110001010;
assign LUT_2[37709] = 32'b11111111111111101100011110100011;
assign LUT_2[37710] = 32'b11111111111111110110011111000110;
assign LUT_2[37711] = 32'b11111111111111110011010111011111;
assign LUT_2[37712] = 32'b11111111111111110010111011001111;
assign LUT_2[37713] = 32'b11111111111111101111110011101000;
assign LUT_2[37714] = 32'b11111111111111111001110100001011;
assign LUT_2[37715] = 32'b11111111111111110110101100100100;
assign LUT_2[37716] = 32'b11111111111111101111011000110111;
assign LUT_2[37717] = 32'b11111111111111101100010001010000;
assign LUT_2[37718] = 32'b11111111111111110110010001110011;
assign LUT_2[37719] = 32'b11111111111111110011001010001100;
assign LUT_2[37720] = 32'b11111111111111101101101100101100;
assign LUT_2[37721] = 32'b11111111111111101010100101000101;
assign LUT_2[37722] = 32'b11111111111111110100100101101000;
assign LUT_2[37723] = 32'b11111111111111110001011110000001;
assign LUT_2[37724] = 32'b11111111111111101010001010010100;
assign LUT_2[37725] = 32'b11111111111111100111000010101101;
assign LUT_2[37726] = 32'b11111111111111110001000011010000;
assign LUT_2[37727] = 32'b11111111111111101101111011101001;
assign LUT_2[37728] = 32'b11111111111111111000110010101110;
assign LUT_2[37729] = 32'b11111111111111110101101011000111;
assign LUT_2[37730] = 32'b11111111111111111111101011101010;
assign LUT_2[37731] = 32'b11111111111111111100100100000011;
assign LUT_2[37732] = 32'b11111111111111110101010000010110;
assign LUT_2[37733] = 32'b11111111111111110010001000101111;
assign LUT_2[37734] = 32'b11111111111111111100001001010010;
assign LUT_2[37735] = 32'b11111111111111111001000001101011;
assign LUT_2[37736] = 32'b11111111111111110011100100001011;
assign LUT_2[37737] = 32'b11111111111111110000011100100100;
assign LUT_2[37738] = 32'b11111111111111111010011101000111;
assign LUT_2[37739] = 32'b11111111111111110111010101100000;
assign LUT_2[37740] = 32'b11111111111111110000000001110011;
assign LUT_2[37741] = 32'b11111111111111101100111010001100;
assign LUT_2[37742] = 32'b11111111111111110110111010101111;
assign LUT_2[37743] = 32'b11111111111111110011110011001000;
assign LUT_2[37744] = 32'b11111111111111110011010110111000;
assign LUT_2[37745] = 32'b11111111111111110000001111010001;
assign LUT_2[37746] = 32'b11111111111111111010001111110100;
assign LUT_2[37747] = 32'b11111111111111110111001000001101;
assign LUT_2[37748] = 32'b11111111111111101111110100100000;
assign LUT_2[37749] = 32'b11111111111111101100101100111001;
assign LUT_2[37750] = 32'b11111111111111110110101101011100;
assign LUT_2[37751] = 32'b11111111111111110011100101110101;
assign LUT_2[37752] = 32'b11111111111111101110001000010101;
assign LUT_2[37753] = 32'b11111111111111101011000000101110;
assign LUT_2[37754] = 32'b11111111111111110101000001010001;
assign LUT_2[37755] = 32'b11111111111111110001111001101010;
assign LUT_2[37756] = 32'b11111111111111101010100101111101;
assign LUT_2[37757] = 32'b11111111111111100111011110010110;
assign LUT_2[37758] = 32'b11111111111111110001011110111001;
assign LUT_2[37759] = 32'b11111111111111101110010111010010;
assign LUT_2[37760] = 32'b00000000000000000100100010110001;
assign LUT_2[37761] = 32'b00000000000000000001011011001010;
assign LUT_2[37762] = 32'b00000000000000001011011011101101;
assign LUT_2[37763] = 32'b00000000000000001000010100000110;
assign LUT_2[37764] = 32'b00000000000000000001000000011001;
assign LUT_2[37765] = 32'b11111111111111111101111000110010;
assign LUT_2[37766] = 32'b00000000000000000111111001010101;
assign LUT_2[37767] = 32'b00000000000000000100110001101110;
assign LUT_2[37768] = 32'b11111111111111111111010100001110;
assign LUT_2[37769] = 32'b11111111111111111100001100100111;
assign LUT_2[37770] = 32'b00000000000000000110001101001010;
assign LUT_2[37771] = 32'b00000000000000000011000101100011;
assign LUT_2[37772] = 32'b11111111111111111011110001110110;
assign LUT_2[37773] = 32'b11111111111111111000101010001111;
assign LUT_2[37774] = 32'b00000000000000000010101010110010;
assign LUT_2[37775] = 32'b11111111111111111111100011001011;
assign LUT_2[37776] = 32'b11111111111111111111000110111011;
assign LUT_2[37777] = 32'b11111111111111111011111111010100;
assign LUT_2[37778] = 32'b00000000000000000101111111110111;
assign LUT_2[37779] = 32'b00000000000000000010111000010000;
assign LUT_2[37780] = 32'b11111111111111111011100100100011;
assign LUT_2[37781] = 32'b11111111111111111000011100111100;
assign LUT_2[37782] = 32'b00000000000000000010011101011111;
assign LUT_2[37783] = 32'b11111111111111111111010101111000;
assign LUT_2[37784] = 32'b11111111111111111001111000011000;
assign LUT_2[37785] = 32'b11111111111111110110110000110001;
assign LUT_2[37786] = 32'b00000000000000000000110001010100;
assign LUT_2[37787] = 32'b11111111111111111101101001101101;
assign LUT_2[37788] = 32'b11111111111111110110010110000000;
assign LUT_2[37789] = 32'b11111111111111110011001110011001;
assign LUT_2[37790] = 32'b11111111111111111101001110111100;
assign LUT_2[37791] = 32'b11111111111111111010000111010101;
assign LUT_2[37792] = 32'b00000000000000000100111110011010;
assign LUT_2[37793] = 32'b00000000000000000001110110110011;
assign LUT_2[37794] = 32'b00000000000000001011110111010110;
assign LUT_2[37795] = 32'b00000000000000001000101111101111;
assign LUT_2[37796] = 32'b00000000000000000001011100000010;
assign LUT_2[37797] = 32'b11111111111111111110010100011011;
assign LUT_2[37798] = 32'b00000000000000001000010100111110;
assign LUT_2[37799] = 32'b00000000000000000101001101010111;
assign LUT_2[37800] = 32'b11111111111111111111101111110111;
assign LUT_2[37801] = 32'b11111111111111111100101000010000;
assign LUT_2[37802] = 32'b00000000000000000110101000110011;
assign LUT_2[37803] = 32'b00000000000000000011100001001100;
assign LUT_2[37804] = 32'b11111111111111111100001101011111;
assign LUT_2[37805] = 32'b11111111111111111001000101111000;
assign LUT_2[37806] = 32'b00000000000000000011000110011011;
assign LUT_2[37807] = 32'b11111111111111111111111110110100;
assign LUT_2[37808] = 32'b11111111111111111111100010100100;
assign LUT_2[37809] = 32'b11111111111111111100011010111101;
assign LUT_2[37810] = 32'b00000000000000000110011011100000;
assign LUT_2[37811] = 32'b00000000000000000011010011111001;
assign LUT_2[37812] = 32'b11111111111111111100000000001100;
assign LUT_2[37813] = 32'b11111111111111111000111000100101;
assign LUT_2[37814] = 32'b00000000000000000010111001001000;
assign LUT_2[37815] = 32'b11111111111111111111110001100001;
assign LUT_2[37816] = 32'b11111111111111111010010100000001;
assign LUT_2[37817] = 32'b11111111111111110111001100011010;
assign LUT_2[37818] = 32'b00000000000000000001001100111101;
assign LUT_2[37819] = 32'b11111111111111111110000101010110;
assign LUT_2[37820] = 32'b11111111111111110110110001101001;
assign LUT_2[37821] = 32'b11111111111111110011101010000010;
assign LUT_2[37822] = 32'b11111111111111111101101010100101;
assign LUT_2[37823] = 32'b11111111111111111010100010111110;
assign LUT_2[37824] = 32'b11111111111111111100101011010100;
assign LUT_2[37825] = 32'b11111111111111111001100011101101;
assign LUT_2[37826] = 32'b00000000000000000011100100010000;
assign LUT_2[37827] = 32'b00000000000000000000011100101001;
assign LUT_2[37828] = 32'b11111111111111111001001000111100;
assign LUT_2[37829] = 32'b11111111111111110110000001010101;
assign LUT_2[37830] = 32'b00000000000000000000000001111000;
assign LUT_2[37831] = 32'b11111111111111111100111010010001;
assign LUT_2[37832] = 32'b11111111111111110111011100110001;
assign LUT_2[37833] = 32'b11111111111111110100010101001010;
assign LUT_2[37834] = 32'b11111111111111111110010101101101;
assign LUT_2[37835] = 32'b11111111111111111011001110000110;
assign LUT_2[37836] = 32'b11111111111111110011111010011001;
assign LUT_2[37837] = 32'b11111111111111110000110010110010;
assign LUT_2[37838] = 32'b11111111111111111010110011010101;
assign LUT_2[37839] = 32'b11111111111111110111101011101110;
assign LUT_2[37840] = 32'b11111111111111110111001111011110;
assign LUT_2[37841] = 32'b11111111111111110100000111110111;
assign LUT_2[37842] = 32'b11111111111111111110001000011010;
assign LUT_2[37843] = 32'b11111111111111111011000000110011;
assign LUT_2[37844] = 32'b11111111111111110011101101000110;
assign LUT_2[37845] = 32'b11111111111111110000100101011111;
assign LUT_2[37846] = 32'b11111111111111111010100110000010;
assign LUT_2[37847] = 32'b11111111111111110111011110011011;
assign LUT_2[37848] = 32'b11111111111111110010000000111011;
assign LUT_2[37849] = 32'b11111111111111101110111001010100;
assign LUT_2[37850] = 32'b11111111111111111000111001110111;
assign LUT_2[37851] = 32'b11111111111111110101110010010000;
assign LUT_2[37852] = 32'b11111111111111101110011110100011;
assign LUT_2[37853] = 32'b11111111111111101011010110111100;
assign LUT_2[37854] = 32'b11111111111111110101010111011111;
assign LUT_2[37855] = 32'b11111111111111110010001111111000;
assign LUT_2[37856] = 32'b11111111111111111101000110111101;
assign LUT_2[37857] = 32'b11111111111111111001111111010110;
assign LUT_2[37858] = 32'b00000000000000000011111111111001;
assign LUT_2[37859] = 32'b00000000000000000000111000010010;
assign LUT_2[37860] = 32'b11111111111111111001100100100101;
assign LUT_2[37861] = 32'b11111111111111110110011100111110;
assign LUT_2[37862] = 32'b00000000000000000000011101100001;
assign LUT_2[37863] = 32'b11111111111111111101010101111010;
assign LUT_2[37864] = 32'b11111111111111110111111000011010;
assign LUT_2[37865] = 32'b11111111111111110100110000110011;
assign LUT_2[37866] = 32'b11111111111111111110110001010110;
assign LUT_2[37867] = 32'b11111111111111111011101001101111;
assign LUT_2[37868] = 32'b11111111111111110100010110000010;
assign LUT_2[37869] = 32'b11111111111111110001001110011011;
assign LUT_2[37870] = 32'b11111111111111111011001110111110;
assign LUT_2[37871] = 32'b11111111111111111000000111010111;
assign LUT_2[37872] = 32'b11111111111111110111101011000111;
assign LUT_2[37873] = 32'b11111111111111110100100011100000;
assign LUT_2[37874] = 32'b11111111111111111110100100000011;
assign LUT_2[37875] = 32'b11111111111111111011011100011100;
assign LUT_2[37876] = 32'b11111111111111110100001000101111;
assign LUT_2[37877] = 32'b11111111111111110001000001001000;
assign LUT_2[37878] = 32'b11111111111111111011000001101011;
assign LUT_2[37879] = 32'b11111111111111110111111010000100;
assign LUT_2[37880] = 32'b11111111111111110010011100100100;
assign LUT_2[37881] = 32'b11111111111111101111010100111101;
assign LUT_2[37882] = 32'b11111111111111111001010101100000;
assign LUT_2[37883] = 32'b11111111111111110110001101111001;
assign LUT_2[37884] = 32'b11111111111111101110111010001100;
assign LUT_2[37885] = 32'b11111111111111101011110010100101;
assign LUT_2[37886] = 32'b11111111111111110101110011001000;
assign LUT_2[37887] = 32'b11111111111111110010101011100001;
assign LUT_2[37888] = 32'b11111111111111111110001010001111;
assign LUT_2[37889] = 32'b11111111111111111011000010101000;
assign LUT_2[37890] = 32'b00000000000000000101000011001011;
assign LUT_2[37891] = 32'b00000000000000000001111011100100;
assign LUT_2[37892] = 32'b11111111111111111010100111110111;
assign LUT_2[37893] = 32'b11111111111111110111100000010000;
assign LUT_2[37894] = 32'b00000000000000000001100000110011;
assign LUT_2[37895] = 32'b11111111111111111110011001001100;
assign LUT_2[37896] = 32'b11111111111111111000111011101100;
assign LUT_2[37897] = 32'b11111111111111110101110100000101;
assign LUT_2[37898] = 32'b11111111111111111111110100101000;
assign LUT_2[37899] = 32'b11111111111111111100101101000001;
assign LUT_2[37900] = 32'b11111111111111110101011001010100;
assign LUT_2[37901] = 32'b11111111111111110010010001101101;
assign LUT_2[37902] = 32'b11111111111111111100010010010000;
assign LUT_2[37903] = 32'b11111111111111111001001010101001;
assign LUT_2[37904] = 32'b11111111111111111000101110011001;
assign LUT_2[37905] = 32'b11111111111111110101100110110010;
assign LUT_2[37906] = 32'b11111111111111111111100111010101;
assign LUT_2[37907] = 32'b11111111111111111100011111101110;
assign LUT_2[37908] = 32'b11111111111111110101001100000001;
assign LUT_2[37909] = 32'b11111111111111110010000100011010;
assign LUT_2[37910] = 32'b11111111111111111100000100111101;
assign LUT_2[37911] = 32'b11111111111111111000111101010110;
assign LUT_2[37912] = 32'b11111111111111110011011111110110;
assign LUT_2[37913] = 32'b11111111111111110000011000001111;
assign LUT_2[37914] = 32'b11111111111111111010011000110010;
assign LUT_2[37915] = 32'b11111111111111110111010001001011;
assign LUT_2[37916] = 32'b11111111111111101111111101011110;
assign LUT_2[37917] = 32'b11111111111111101100110101110111;
assign LUT_2[37918] = 32'b11111111111111110110110110011010;
assign LUT_2[37919] = 32'b11111111111111110011101110110011;
assign LUT_2[37920] = 32'b11111111111111111110100101111000;
assign LUT_2[37921] = 32'b11111111111111111011011110010001;
assign LUT_2[37922] = 32'b00000000000000000101011110110100;
assign LUT_2[37923] = 32'b00000000000000000010010111001101;
assign LUT_2[37924] = 32'b11111111111111111011000011100000;
assign LUT_2[37925] = 32'b11111111111111110111111011111001;
assign LUT_2[37926] = 32'b00000000000000000001111100011100;
assign LUT_2[37927] = 32'b11111111111111111110110100110101;
assign LUT_2[37928] = 32'b11111111111111111001010111010101;
assign LUT_2[37929] = 32'b11111111111111110110001111101110;
assign LUT_2[37930] = 32'b00000000000000000000010000010001;
assign LUT_2[37931] = 32'b11111111111111111101001000101010;
assign LUT_2[37932] = 32'b11111111111111110101110100111101;
assign LUT_2[37933] = 32'b11111111111111110010101101010110;
assign LUT_2[37934] = 32'b11111111111111111100101101111001;
assign LUT_2[37935] = 32'b11111111111111111001100110010010;
assign LUT_2[37936] = 32'b11111111111111111001001010000010;
assign LUT_2[37937] = 32'b11111111111111110110000010011011;
assign LUT_2[37938] = 32'b00000000000000000000000010111110;
assign LUT_2[37939] = 32'b11111111111111111100111011010111;
assign LUT_2[37940] = 32'b11111111111111110101100111101010;
assign LUT_2[37941] = 32'b11111111111111110010100000000011;
assign LUT_2[37942] = 32'b11111111111111111100100000100110;
assign LUT_2[37943] = 32'b11111111111111111001011000111111;
assign LUT_2[37944] = 32'b11111111111111110011111011011111;
assign LUT_2[37945] = 32'b11111111111111110000110011111000;
assign LUT_2[37946] = 32'b11111111111111111010110100011011;
assign LUT_2[37947] = 32'b11111111111111110111101100110100;
assign LUT_2[37948] = 32'b11111111111111110000011001000111;
assign LUT_2[37949] = 32'b11111111111111101101010001100000;
assign LUT_2[37950] = 32'b11111111111111110111010010000011;
assign LUT_2[37951] = 32'b11111111111111110100001010011100;
assign LUT_2[37952] = 32'b11111111111111110110010010110010;
assign LUT_2[37953] = 32'b11111111111111110011001011001011;
assign LUT_2[37954] = 32'b11111111111111111101001011101110;
assign LUT_2[37955] = 32'b11111111111111111010000100000111;
assign LUT_2[37956] = 32'b11111111111111110010110000011010;
assign LUT_2[37957] = 32'b11111111111111101111101000110011;
assign LUT_2[37958] = 32'b11111111111111111001101001010110;
assign LUT_2[37959] = 32'b11111111111111110110100001101111;
assign LUT_2[37960] = 32'b11111111111111110001000100001111;
assign LUT_2[37961] = 32'b11111111111111101101111100101000;
assign LUT_2[37962] = 32'b11111111111111110111111101001011;
assign LUT_2[37963] = 32'b11111111111111110100110101100100;
assign LUT_2[37964] = 32'b11111111111111101101100001110111;
assign LUT_2[37965] = 32'b11111111111111101010011010010000;
assign LUT_2[37966] = 32'b11111111111111110100011010110011;
assign LUT_2[37967] = 32'b11111111111111110001010011001100;
assign LUT_2[37968] = 32'b11111111111111110000110110111100;
assign LUT_2[37969] = 32'b11111111111111101101101111010101;
assign LUT_2[37970] = 32'b11111111111111110111101111111000;
assign LUT_2[37971] = 32'b11111111111111110100101000010001;
assign LUT_2[37972] = 32'b11111111111111101101010100100100;
assign LUT_2[37973] = 32'b11111111111111101010001100111101;
assign LUT_2[37974] = 32'b11111111111111110100001101100000;
assign LUT_2[37975] = 32'b11111111111111110001000101111001;
assign LUT_2[37976] = 32'b11111111111111101011101000011001;
assign LUT_2[37977] = 32'b11111111111111101000100000110010;
assign LUT_2[37978] = 32'b11111111111111110010100001010101;
assign LUT_2[37979] = 32'b11111111111111101111011001101110;
assign LUT_2[37980] = 32'b11111111111111101000000110000001;
assign LUT_2[37981] = 32'b11111111111111100100111110011010;
assign LUT_2[37982] = 32'b11111111111111101110111110111101;
assign LUT_2[37983] = 32'b11111111111111101011110111010110;
assign LUT_2[37984] = 32'b11111111111111110110101110011011;
assign LUT_2[37985] = 32'b11111111111111110011100110110100;
assign LUT_2[37986] = 32'b11111111111111111101100111010111;
assign LUT_2[37987] = 32'b11111111111111111010011111110000;
assign LUT_2[37988] = 32'b11111111111111110011001100000011;
assign LUT_2[37989] = 32'b11111111111111110000000100011100;
assign LUT_2[37990] = 32'b11111111111111111010000100111111;
assign LUT_2[37991] = 32'b11111111111111110110111101011000;
assign LUT_2[37992] = 32'b11111111111111110001011111111000;
assign LUT_2[37993] = 32'b11111111111111101110011000010001;
assign LUT_2[37994] = 32'b11111111111111111000011000110100;
assign LUT_2[37995] = 32'b11111111111111110101010001001101;
assign LUT_2[37996] = 32'b11111111111111101101111101100000;
assign LUT_2[37997] = 32'b11111111111111101010110101111001;
assign LUT_2[37998] = 32'b11111111111111110100110110011100;
assign LUT_2[37999] = 32'b11111111111111110001101110110101;
assign LUT_2[38000] = 32'b11111111111111110001010010100101;
assign LUT_2[38001] = 32'b11111111111111101110001010111110;
assign LUT_2[38002] = 32'b11111111111111111000001011100001;
assign LUT_2[38003] = 32'b11111111111111110101000011111010;
assign LUT_2[38004] = 32'b11111111111111101101110000001101;
assign LUT_2[38005] = 32'b11111111111111101010101000100110;
assign LUT_2[38006] = 32'b11111111111111110100101001001001;
assign LUT_2[38007] = 32'b11111111111111110001100001100010;
assign LUT_2[38008] = 32'b11111111111111101100000100000010;
assign LUT_2[38009] = 32'b11111111111111101000111100011011;
assign LUT_2[38010] = 32'b11111111111111110010111100111110;
assign LUT_2[38011] = 32'b11111111111111101111110101010111;
assign LUT_2[38012] = 32'b11111111111111101000100001101010;
assign LUT_2[38013] = 32'b11111111111111100101011010000011;
assign LUT_2[38014] = 32'b11111111111111101111011010100110;
assign LUT_2[38015] = 32'b11111111111111101100010010111111;
assign LUT_2[38016] = 32'b00000000000000000010011110011110;
assign LUT_2[38017] = 32'b11111111111111111111010110110111;
assign LUT_2[38018] = 32'b00000000000000001001010111011010;
assign LUT_2[38019] = 32'b00000000000000000110001111110011;
assign LUT_2[38020] = 32'b11111111111111111110111100000110;
assign LUT_2[38021] = 32'b11111111111111111011110100011111;
assign LUT_2[38022] = 32'b00000000000000000101110101000010;
assign LUT_2[38023] = 32'b00000000000000000010101101011011;
assign LUT_2[38024] = 32'b11111111111111111101001111111011;
assign LUT_2[38025] = 32'b11111111111111111010001000010100;
assign LUT_2[38026] = 32'b00000000000000000100001000110111;
assign LUT_2[38027] = 32'b00000000000000000001000001010000;
assign LUT_2[38028] = 32'b11111111111111111001101101100011;
assign LUT_2[38029] = 32'b11111111111111110110100101111100;
assign LUT_2[38030] = 32'b00000000000000000000100110011111;
assign LUT_2[38031] = 32'b11111111111111111101011110111000;
assign LUT_2[38032] = 32'b11111111111111111101000010101000;
assign LUT_2[38033] = 32'b11111111111111111001111011000001;
assign LUT_2[38034] = 32'b00000000000000000011111011100100;
assign LUT_2[38035] = 32'b00000000000000000000110011111101;
assign LUT_2[38036] = 32'b11111111111111111001100000010000;
assign LUT_2[38037] = 32'b11111111111111110110011000101001;
assign LUT_2[38038] = 32'b00000000000000000000011001001100;
assign LUT_2[38039] = 32'b11111111111111111101010001100101;
assign LUT_2[38040] = 32'b11111111111111110111110100000101;
assign LUT_2[38041] = 32'b11111111111111110100101100011110;
assign LUT_2[38042] = 32'b11111111111111111110101101000001;
assign LUT_2[38043] = 32'b11111111111111111011100101011010;
assign LUT_2[38044] = 32'b11111111111111110100010001101101;
assign LUT_2[38045] = 32'b11111111111111110001001010000110;
assign LUT_2[38046] = 32'b11111111111111111011001010101001;
assign LUT_2[38047] = 32'b11111111111111111000000011000010;
assign LUT_2[38048] = 32'b00000000000000000010111010000111;
assign LUT_2[38049] = 32'b11111111111111111111110010100000;
assign LUT_2[38050] = 32'b00000000000000001001110011000011;
assign LUT_2[38051] = 32'b00000000000000000110101011011100;
assign LUT_2[38052] = 32'b11111111111111111111010111101111;
assign LUT_2[38053] = 32'b11111111111111111100010000001000;
assign LUT_2[38054] = 32'b00000000000000000110010000101011;
assign LUT_2[38055] = 32'b00000000000000000011001001000100;
assign LUT_2[38056] = 32'b11111111111111111101101011100100;
assign LUT_2[38057] = 32'b11111111111111111010100011111101;
assign LUT_2[38058] = 32'b00000000000000000100100100100000;
assign LUT_2[38059] = 32'b00000000000000000001011100111001;
assign LUT_2[38060] = 32'b11111111111111111010001001001100;
assign LUT_2[38061] = 32'b11111111111111110111000001100101;
assign LUT_2[38062] = 32'b00000000000000000001000010001000;
assign LUT_2[38063] = 32'b11111111111111111101111010100001;
assign LUT_2[38064] = 32'b11111111111111111101011110010001;
assign LUT_2[38065] = 32'b11111111111111111010010110101010;
assign LUT_2[38066] = 32'b00000000000000000100010111001101;
assign LUT_2[38067] = 32'b00000000000000000001001111100110;
assign LUT_2[38068] = 32'b11111111111111111001111011111001;
assign LUT_2[38069] = 32'b11111111111111110110110100010010;
assign LUT_2[38070] = 32'b00000000000000000000110100110101;
assign LUT_2[38071] = 32'b11111111111111111101101101001110;
assign LUT_2[38072] = 32'b11111111111111111000001111101110;
assign LUT_2[38073] = 32'b11111111111111110101001000000111;
assign LUT_2[38074] = 32'b11111111111111111111001000101010;
assign LUT_2[38075] = 32'b11111111111111111100000001000011;
assign LUT_2[38076] = 32'b11111111111111110100101101010110;
assign LUT_2[38077] = 32'b11111111111111110001100101101111;
assign LUT_2[38078] = 32'b11111111111111111011100110010010;
assign LUT_2[38079] = 32'b11111111111111111000011110101011;
assign LUT_2[38080] = 32'b11111111111111111010100111000001;
assign LUT_2[38081] = 32'b11111111111111110111011111011010;
assign LUT_2[38082] = 32'b00000000000000000001011111111101;
assign LUT_2[38083] = 32'b11111111111111111110011000010110;
assign LUT_2[38084] = 32'b11111111111111110111000100101001;
assign LUT_2[38085] = 32'b11111111111111110011111101000010;
assign LUT_2[38086] = 32'b11111111111111111101111101100101;
assign LUT_2[38087] = 32'b11111111111111111010110101111110;
assign LUT_2[38088] = 32'b11111111111111110101011000011110;
assign LUT_2[38089] = 32'b11111111111111110010010000110111;
assign LUT_2[38090] = 32'b11111111111111111100010001011010;
assign LUT_2[38091] = 32'b11111111111111111001001001110011;
assign LUT_2[38092] = 32'b11111111111111110001110110000110;
assign LUT_2[38093] = 32'b11111111111111101110101110011111;
assign LUT_2[38094] = 32'b11111111111111111000101111000010;
assign LUT_2[38095] = 32'b11111111111111110101100111011011;
assign LUT_2[38096] = 32'b11111111111111110101001011001011;
assign LUT_2[38097] = 32'b11111111111111110010000011100100;
assign LUT_2[38098] = 32'b11111111111111111100000100000111;
assign LUT_2[38099] = 32'b11111111111111111000111100100000;
assign LUT_2[38100] = 32'b11111111111111110001101000110011;
assign LUT_2[38101] = 32'b11111111111111101110100001001100;
assign LUT_2[38102] = 32'b11111111111111111000100001101111;
assign LUT_2[38103] = 32'b11111111111111110101011010001000;
assign LUT_2[38104] = 32'b11111111111111101111111100101000;
assign LUT_2[38105] = 32'b11111111111111101100110101000001;
assign LUT_2[38106] = 32'b11111111111111110110110101100100;
assign LUT_2[38107] = 32'b11111111111111110011101101111101;
assign LUT_2[38108] = 32'b11111111111111101100011010010000;
assign LUT_2[38109] = 32'b11111111111111101001010010101001;
assign LUT_2[38110] = 32'b11111111111111110011010011001100;
assign LUT_2[38111] = 32'b11111111111111110000001011100101;
assign LUT_2[38112] = 32'b11111111111111111011000010101010;
assign LUT_2[38113] = 32'b11111111111111110111111011000011;
assign LUT_2[38114] = 32'b00000000000000000001111011100110;
assign LUT_2[38115] = 32'b11111111111111111110110011111111;
assign LUT_2[38116] = 32'b11111111111111110111100000010010;
assign LUT_2[38117] = 32'b11111111111111110100011000101011;
assign LUT_2[38118] = 32'b11111111111111111110011001001110;
assign LUT_2[38119] = 32'b11111111111111111011010001100111;
assign LUT_2[38120] = 32'b11111111111111110101110100000111;
assign LUT_2[38121] = 32'b11111111111111110010101100100000;
assign LUT_2[38122] = 32'b11111111111111111100101101000011;
assign LUT_2[38123] = 32'b11111111111111111001100101011100;
assign LUT_2[38124] = 32'b11111111111111110010010001101111;
assign LUT_2[38125] = 32'b11111111111111101111001010001000;
assign LUT_2[38126] = 32'b11111111111111111001001010101011;
assign LUT_2[38127] = 32'b11111111111111110110000011000100;
assign LUT_2[38128] = 32'b11111111111111110101100110110100;
assign LUT_2[38129] = 32'b11111111111111110010011111001101;
assign LUT_2[38130] = 32'b11111111111111111100011111110000;
assign LUT_2[38131] = 32'b11111111111111111001011000001001;
assign LUT_2[38132] = 32'b11111111111111110010000100011100;
assign LUT_2[38133] = 32'b11111111111111101110111100110101;
assign LUT_2[38134] = 32'b11111111111111111000111101011000;
assign LUT_2[38135] = 32'b11111111111111110101110101110001;
assign LUT_2[38136] = 32'b11111111111111110000011000010001;
assign LUT_2[38137] = 32'b11111111111111101101010000101010;
assign LUT_2[38138] = 32'b11111111111111110111010001001101;
assign LUT_2[38139] = 32'b11111111111111110100001001100110;
assign LUT_2[38140] = 32'b11111111111111101100110101111001;
assign LUT_2[38141] = 32'b11111111111111101001101110010010;
assign LUT_2[38142] = 32'b11111111111111110011101110110101;
assign LUT_2[38143] = 32'b11111111111111110000100111001110;
assign LUT_2[38144] = 32'b00000000000000000010001000110101;
assign LUT_2[38145] = 32'b11111111111111111111000001001110;
assign LUT_2[38146] = 32'b00000000000000001001000001110001;
assign LUT_2[38147] = 32'b00000000000000000101111010001010;
assign LUT_2[38148] = 32'b11111111111111111110100110011101;
assign LUT_2[38149] = 32'b11111111111111111011011110110110;
assign LUT_2[38150] = 32'b00000000000000000101011111011001;
assign LUT_2[38151] = 32'b00000000000000000010010111110010;
assign LUT_2[38152] = 32'b11111111111111111100111010010010;
assign LUT_2[38153] = 32'b11111111111111111001110010101011;
assign LUT_2[38154] = 32'b00000000000000000011110011001110;
assign LUT_2[38155] = 32'b00000000000000000000101011100111;
assign LUT_2[38156] = 32'b11111111111111111001010111111010;
assign LUT_2[38157] = 32'b11111111111111110110010000010011;
assign LUT_2[38158] = 32'b00000000000000000000010000110110;
assign LUT_2[38159] = 32'b11111111111111111101001001001111;
assign LUT_2[38160] = 32'b11111111111111111100101100111111;
assign LUT_2[38161] = 32'b11111111111111111001100101011000;
assign LUT_2[38162] = 32'b00000000000000000011100101111011;
assign LUT_2[38163] = 32'b00000000000000000000011110010100;
assign LUT_2[38164] = 32'b11111111111111111001001010100111;
assign LUT_2[38165] = 32'b11111111111111110110000011000000;
assign LUT_2[38166] = 32'b00000000000000000000000011100011;
assign LUT_2[38167] = 32'b11111111111111111100111011111100;
assign LUT_2[38168] = 32'b11111111111111110111011110011100;
assign LUT_2[38169] = 32'b11111111111111110100010110110101;
assign LUT_2[38170] = 32'b11111111111111111110010111011000;
assign LUT_2[38171] = 32'b11111111111111111011001111110001;
assign LUT_2[38172] = 32'b11111111111111110011111100000100;
assign LUT_2[38173] = 32'b11111111111111110000110100011101;
assign LUT_2[38174] = 32'b11111111111111111010110101000000;
assign LUT_2[38175] = 32'b11111111111111110111101101011001;
assign LUT_2[38176] = 32'b00000000000000000010100100011110;
assign LUT_2[38177] = 32'b11111111111111111111011100110111;
assign LUT_2[38178] = 32'b00000000000000001001011101011010;
assign LUT_2[38179] = 32'b00000000000000000110010101110011;
assign LUT_2[38180] = 32'b11111111111111111111000010000110;
assign LUT_2[38181] = 32'b11111111111111111011111010011111;
assign LUT_2[38182] = 32'b00000000000000000101111011000010;
assign LUT_2[38183] = 32'b00000000000000000010110011011011;
assign LUT_2[38184] = 32'b11111111111111111101010101111011;
assign LUT_2[38185] = 32'b11111111111111111010001110010100;
assign LUT_2[38186] = 32'b00000000000000000100001110110111;
assign LUT_2[38187] = 32'b00000000000000000001000111010000;
assign LUT_2[38188] = 32'b11111111111111111001110011100011;
assign LUT_2[38189] = 32'b11111111111111110110101011111100;
assign LUT_2[38190] = 32'b00000000000000000000101100011111;
assign LUT_2[38191] = 32'b11111111111111111101100100111000;
assign LUT_2[38192] = 32'b11111111111111111101001000101000;
assign LUT_2[38193] = 32'b11111111111111111010000001000001;
assign LUT_2[38194] = 32'b00000000000000000100000001100100;
assign LUT_2[38195] = 32'b00000000000000000000111001111101;
assign LUT_2[38196] = 32'b11111111111111111001100110010000;
assign LUT_2[38197] = 32'b11111111111111110110011110101001;
assign LUT_2[38198] = 32'b00000000000000000000011111001100;
assign LUT_2[38199] = 32'b11111111111111111101010111100101;
assign LUT_2[38200] = 32'b11111111111111110111111010000101;
assign LUT_2[38201] = 32'b11111111111111110100110010011110;
assign LUT_2[38202] = 32'b11111111111111111110110011000001;
assign LUT_2[38203] = 32'b11111111111111111011101011011010;
assign LUT_2[38204] = 32'b11111111111111110100010111101101;
assign LUT_2[38205] = 32'b11111111111111110001010000000110;
assign LUT_2[38206] = 32'b11111111111111111011010000101001;
assign LUT_2[38207] = 32'b11111111111111111000001001000010;
assign LUT_2[38208] = 32'b11111111111111111010010001011000;
assign LUT_2[38209] = 32'b11111111111111110111001001110001;
assign LUT_2[38210] = 32'b00000000000000000001001010010100;
assign LUT_2[38211] = 32'b11111111111111111110000010101101;
assign LUT_2[38212] = 32'b11111111111111110110101111000000;
assign LUT_2[38213] = 32'b11111111111111110011100111011001;
assign LUT_2[38214] = 32'b11111111111111111101100111111100;
assign LUT_2[38215] = 32'b11111111111111111010100000010101;
assign LUT_2[38216] = 32'b11111111111111110101000010110101;
assign LUT_2[38217] = 32'b11111111111111110001111011001110;
assign LUT_2[38218] = 32'b11111111111111111011111011110001;
assign LUT_2[38219] = 32'b11111111111111111000110100001010;
assign LUT_2[38220] = 32'b11111111111111110001100000011101;
assign LUT_2[38221] = 32'b11111111111111101110011000110110;
assign LUT_2[38222] = 32'b11111111111111111000011001011001;
assign LUT_2[38223] = 32'b11111111111111110101010001110010;
assign LUT_2[38224] = 32'b11111111111111110100110101100010;
assign LUT_2[38225] = 32'b11111111111111110001101101111011;
assign LUT_2[38226] = 32'b11111111111111111011101110011110;
assign LUT_2[38227] = 32'b11111111111111111000100110110111;
assign LUT_2[38228] = 32'b11111111111111110001010011001010;
assign LUT_2[38229] = 32'b11111111111111101110001011100011;
assign LUT_2[38230] = 32'b11111111111111111000001100000110;
assign LUT_2[38231] = 32'b11111111111111110101000100011111;
assign LUT_2[38232] = 32'b11111111111111101111100110111111;
assign LUT_2[38233] = 32'b11111111111111101100011111011000;
assign LUT_2[38234] = 32'b11111111111111110110011111111011;
assign LUT_2[38235] = 32'b11111111111111110011011000010100;
assign LUT_2[38236] = 32'b11111111111111101100000100100111;
assign LUT_2[38237] = 32'b11111111111111101000111101000000;
assign LUT_2[38238] = 32'b11111111111111110010111101100011;
assign LUT_2[38239] = 32'b11111111111111101111110101111100;
assign LUT_2[38240] = 32'b11111111111111111010101101000001;
assign LUT_2[38241] = 32'b11111111111111110111100101011010;
assign LUT_2[38242] = 32'b00000000000000000001100101111101;
assign LUT_2[38243] = 32'b11111111111111111110011110010110;
assign LUT_2[38244] = 32'b11111111111111110111001010101001;
assign LUT_2[38245] = 32'b11111111111111110100000011000010;
assign LUT_2[38246] = 32'b11111111111111111110000011100101;
assign LUT_2[38247] = 32'b11111111111111111010111011111110;
assign LUT_2[38248] = 32'b11111111111111110101011110011110;
assign LUT_2[38249] = 32'b11111111111111110010010110110111;
assign LUT_2[38250] = 32'b11111111111111111100010111011010;
assign LUT_2[38251] = 32'b11111111111111111001001111110011;
assign LUT_2[38252] = 32'b11111111111111110001111100000110;
assign LUT_2[38253] = 32'b11111111111111101110110100011111;
assign LUT_2[38254] = 32'b11111111111111111000110101000010;
assign LUT_2[38255] = 32'b11111111111111110101101101011011;
assign LUT_2[38256] = 32'b11111111111111110101010001001011;
assign LUT_2[38257] = 32'b11111111111111110010001001100100;
assign LUT_2[38258] = 32'b11111111111111111100001010000111;
assign LUT_2[38259] = 32'b11111111111111111001000010100000;
assign LUT_2[38260] = 32'b11111111111111110001101110110011;
assign LUT_2[38261] = 32'b11111111111111101110100111001100;
assign LUT_2[38262] = 32'b11111111111111111000100111101111;
assign LUT_2[38263] = 32'b11111111111111110101100000001000;
assign LUT_2[38264] = 32'b11111111111111110000000010101000;
assign LUT_2[38265] = 32'b11111111111111101100111011000001;
assign LUT_2[38266] = 32'b11111111111111110110111011100100;
assign LUT_2[38267] = 32'b11111111111111110011110011111101;
assign LUT_2[38268] = 32'b11111111111111101100100000010000;
assign LUT_2[38269] = 32'b11111111111111101001011000101001;
assign LUT_2[38270] = 32'b11111111111111110011011001001100;
assign LUT_2[38271] = 32'b11111111111111110000010001100101;
assign LUT_2[38272] = 32'b00000000000000000110011101000100;
assign LUT_2[38273] = 32'b00000000000000000011010101011101;
assign LUT_2[38274] = 32'b00000000000000001101010110000000;
assign LUT_2[38275] = 32'b00000000000000001010001110011001;
assign LUT_2[38276] = 32'b00000000000000000010111010101100;
assign LUT_2[38277] = 32'b11111111111111111111110011000101;
assign LUT_2[38278] = 32'b00000000000000001001110011101000;
assign LUT_2[38279] = 32'b00000000000000000110101100000001;
assign LUT_2[38280] = 32'b00000000000000000001001110100001;
assign LUT_2[38281] = 32'b11111111111111111110000110111010;
assign LUT_2[38282] = 32'b00000000000000001000000111011101;
assign LUT_2[38283] = 32'b00000000000000000100111111110110;
assign LUT_2[38284] = 32'b11111111111111111101101100001001;
assign LUT_2[38285] = 32'b11111111111111111010100100100010;
assign LUT_2[38286] = 32'b00000000000000000100100101000101;
assign LUT_2[38287] = 32'b00000000000000000001011101011110;
assign LUT_2[38288] = 32'b00000000000000000001000001001110;
assign LUT_2[38289] = 32'b11111111111111111101111001100111;
assign LUT_2[38290] = 32'b00000000000000000111111010001010;
assign LUT_2[38291] = 32'b00000000000000000100110010100011;
assign LUT_2[38292] = 32'b11111111111111111101011110110110;
assign LUT_2[38293] = 32'b11111111111111111010010111001111;
assign LUT_2[38294] = 32'b00000000000000000100010111110010;
assign LUT_2[38295] = 32'b00000000000000000001010000001011;
assign LUT_2[38296] = 32'b11111111111111111011110010101011;
assign LUT_2[38297] = 32'b11111111111111111000101011000100;
assign LUT_2[38298] = 32'b00000000000000000010101011100111;
assign LUT_2[38299] = 32'b11111111111111111111100100000000;
assign LUT_2[38300] = 32'b11111111111111111000010000010011;
assign LUT_2[38301] = 32'b11111111111111110101001000101100;
assign LUT_2[38302] = 32'b11111111111111111111001001001111;
assign LUT_2[38303] = 32'b11111111111111111100000001101000;
assign LUT_2[38304] = 32'b00000000000000000110111000101101;
assign LUT_2[38305] = 32'b00000000000000000011110001000110;
assign LUT_2[38306] = 32'b00000000000000001101110001101001;
assign LUT_2[38307] = 32'b00000000000000001010101010000010;
assign LUT_2[38308] = 32'b00000000000000000011010110010101;
assign LUT_2[38309] = 32'b00000000000000000000001110101110;
assign LUT_2[38310] = 32'b00000000000000001010001111010001;
assign LUT_2[38311] = 32'b00000000000000000111000111101010;
assign LUT_2[38312] = 32'b00000000000000000001101010001010;
assign LUT_2[38313] = 32'b11111111111111111110100010100011;
assign LUT_2[38314] = 32'b00000000000000001000100011000110;
assign LUT_2[38315] = 32'b00000000000000000101011011011111;
assign LUT_2[38316] = 32'b11111111111111111110000111110010;
assign LUT_2[38317] = 32'b11111111111111111011000000001011;
assign LUT_2[38318] = 32'b00000000000000000101000000101110;
assign LUT_2[38319] = 32'b00000000000000000001111001000111;
assign LUT_2[38320] = 32'b00000000000000000001011100110111;
assign LUT_2[38321] = 32'b11111111111111111110010101010000;
assign LUT_2[38322] = 32'b00000000000000001000010101110011;
assign LUT_2[38323] = 32'b00000000000000000101001110001100;
assign LUT_2[38324] = 32'b11111111111111111101111010011111;
assign LUT_2[38325] = 32'b11111111111111111010110010111000;
assign LUT_2[38326] = 32'b00000000000000000100110011011011;
assign LUT_2[38327] = 32'b00000000000000000001101011110100;
assign LUT_2[38328] = 32'b11111111111111111100001110010100;
assign LUT_2[38329] = 32'b11111111111111111001000110101101;
assign LUT_2[38330] = 32'b00000000000000000011000111010000;
assign LUT_2[38331] = 32'b11111111111111111111111111101001;
assign LUT_2[38332] = 32'b11111111111111111000101011111100;
assign LUT_2[38333] = 32'b11111111111111110101100100010101;
assign LUT_2[38334] = 32'b11111111111111111111100100111000;
assign LUT_2[38335] = 32'b11111111111111111100011101010001;
assign LUT_2[38336] = 32'b11111111111111111110100101100111;
assign LUT_2[38337] = 32'b11111111111111111011011110000000;
assign LUT_2[38338] = 32'b00000000000000000101011110100011;
assign LUT_2[38339] = 32'b00000000000000000010010110111100;
assign LUT_2[38340] = 32'b11111111111111111011000011001111;
assign LUT_2[38341] = 32'b11111111111111110111111011101000;
assign LUT_2[38342] = 32'b00000000000000000001111100001011;
assign LUT_2[38343] = 32'b11111111111111111110110100100100;
assign LUT_2[38344] = 32'b11111111111111111001010111000100;
assign LUT_2[38345] = 32'b11111111111111110110001111011101;
assign LUT_2[38346] = 32'b00000000000000000000010000000000;
assign LUT_2[38347] = 32'b11111111111111111101001000011001;
assign LUT_2[38348] = 32'b11111111111111110101110100101100;
assign LUT_2[38349] = 32'b11111111111111110010101101000101;
assign LUT_2[38350] = 32'b11111111111111111100101101101000;
assign LUT_2[38351] = 32'b11111111111111111001100110000001;
assign LUT_2[38352] = 32'b11111111111111111001001001110001;
assign LUT_2[38353] = 32'b11111111111111110110000010001010;
assign LUT_2[38354] = 32'b00000000000000000000000010101101;
assign LUT_2[38355] = 32'b11111111111111111100111011000110;
assign LUT_2[38356] = 32'b11111111111111110101100111011001;
assign LUT_2[38357] = 32'b11111111111111110010011111110010;
assign LUT_2[38358] = 32'b11111111111111111100100000010101;
assign LUT_2[38359] = 32'b11111111111111111001011000101110;
assign LUT_2[38360] = 32'b11111111111111110011111011001110;
assign LUT_2[38361] = 32'b11111111111111110000110011100111;
assign LUT_2[38362] = 32'b11111111111111111010110100001010;
assign LUT_2[38363] = 32'b11111111111111110111101100100011;
assign LUT_2[38364] = 32'b11111111111111110000011000110110;
assign LUT_2[38365] = 32'b11111111111111101101010001001111;
assign LUT_2[38366] = 32'b11111111111111110111010001110010;
assign LUT_2[38367] = 32'b11111111111111110100001010001011;
assign LUT_2[38368] = 32'b11111111111111111111000001010000;
assign LUT_2[38369] = 32'b11111111111111111011111001101001;
assign LUT_2[38370] = 32'b00000000000000000101111010001100;
assign LUT_2[38371] = 32'b00000000000000000010110010100101;
assign LUT_2[38372] = 32'b11111111111111111011011110111000;
assign LUT_2[38373] = 32'b11111111111111111000010111010001;
assign LUT_2[38374] = 32'b00000000000000000010010111110100;
assign LUT_2[38375] = 32'b11111111111111111111010000001101;
assign LUT_2[38376] = 32'b11111111111111111001110010101101;
assign LUT_2[38377] = 32'b11111111111111110110101011000110;
assign LUT_2[38378] = 32'b00000000000000000000101011101001;
assign LUT_2[38379] = 32'b11111111111111111101100100000010;
assign LUT_2[38380] = 32'b11111111111111110110010000010101;
assign LUT_2[38381] = 32'b11111111111111110011001000101110;
assign LUT_2[38382] = 32'b11111111111111111101001001010001;
assign LUT_2[38383] = 32'b11111111111111111010000001101010;
assign LUT_2[38384] = 32'b11111111111111111001100101011010;
assign LUT_2[38385] = 32'b11111111111111110110011101110011;
assign LUT_2[38386] = 32'b00000000000000000000011110010110;
assign LUT_2[38387] = 32'b11111111111111111101010110101111;
assign LUT_2[38388] = 32'b11111111111111110110000011000010;
assign LUT_2[38389] = 32'b11111111111111110010111011011011;
assign LUT_2[38390] = 32'b11111111111111111100111011111110;
assign LUT_2[38391] = 32'b11111111111111111001110100010111;
assign LUT_2[38392] = 32'b11111111111111110100010110110111;
assign LUT_2[38393] = 32'b11111111111111110001001111010000;
assign LUT_2[38394] = 32'b11111111111111111011001111110011;
assign LUT_2[38395] = 32'b11111111111111111000001000001100;
assign LUT_2[38396] = 32'b11111111111111110000110100011111;
assign LUT_2[38397] = 32'b11111111111111101101101100111000;
assign LUT_2[38398] = 32'b11111111111111110111101101011011;
assign LUT_2[38399] = 32'b11111111111111110100100101110100;
assign LUT_2[38400] = 32'b00000000000000000010111100000001;
assign LUT_2[38401] = 32'b11111111111111111111110100011010;
assign LUT_2[38402] = 32'b00000000000000001001110100111101;
assign LUT_2[38403] = 32'b00000000000000000110101101010110;
assign LUT_2[38404] = 32'b11111111111111111111011001101001;
assign LUT_2[38405] = 32'b11111111111111111100010010000010;
assign LUT_2[38406] = 32'b00000000000000000110010010100101;
assign LUT_2[38407] = 32'b00000000000000000011001010111110;
assign LUT_2[38408] = 32'b11111111111111111101101101011110;
assign LUT_2[38409] = 32'b11111111111111111010100101110111;
assign LUT_2[38410] = 32'b00000000000000000100100110011010;
assign LUT_2[38411] = 32'b00000000000000000001011110110011;
assign LUT_2[38412] = 32'b11111111111111111010001011000110;
assign LUT_2[38413] = 32'b11111111111111110111000011011111;
assign LUT_2[38414] = 32'b00000000000000000001000100000010;
assign LUT_2[38415] = 32'b11111111111111111101111100011011;
assign LUT_2[38416] = 32'b11111111111111111101100000001011;
assign LUT_2[38417] = 32'b11111111111111111010011000100100;
assign LUT_2[38418] = 32'b00000000000000000100011001000111;
assign LUT_2[38419] = 32'b00000000000000000001010001100000;
assign LUT_2[38420] = 32'b11111111111111111001111101110011;
assign LUT_2[38421] = 32'b11111111111111110110110110001100;
assign LUT_2[38422] = 32'b00000000000000000000110110101111;
assign LUT_2[38423] = 32'b11111111111111111101101111001000;
assign LUT_2[38424] = 32'b11111111111111111000010001101000;
assign LUT_2[38425] = 32'b11111111111111110101001010000001;
assign LUT_2[38426] = 32'b11111111111111111111001010100100;
assign LUT_2[38427] = 32'b11111111111111111100000010111101;
assign LUT_2[38428] = 32'b11111111111111110100101111010000;
assign LUT_2[38429] = 32'b11111111111111110001100111101001;
assign LUT_2[38430] = 32'b11111111111111111011101000001100;
assign LUT_2[38431] = 32'b11111111111111111000100000100101;
assign LUT_2[38432] = 32'b00000000000000000011010111101010;
assign LUT_2[38433] = 32'b00000000000000000000010000000011;
assign LUT_2[38434] = 32'b00000000000000001010010000100110;
assign LUT_2[38435] = 32'b00000000000000000111001000111111;
assign LUT_2[38436] = 32'b11111111111111111111110101010010;
assign LUT_2[38437] = 32'b11111111111111111100101101101011;
assign LUT_2[38438] = 32'b00000000000000000110101110001110;
assign LUT_2[38439] = 32'b00000000000000000011100110100111;
assign LUT_2[38440] = 32'b11111111111111111110001001000111;
assign LUT_2[38441] = 32'b11111111111111111011000001100000;
assign LUT_2[38442] = 32'b00000000000000000101000010000011;
assign LUT_2[38443] = 32'b00000000000000000001111010011100;
assign LUT_2[38444] = 32'b11111111111111111010100110101111;
assign LUT_2[38445] = 32'b11111111111111110111011111001000;
assign LUT_2[38446] = 32'b00000000000000000001011111101011;
assign LUT_2[38447] = 32'b11111111111111111110011000000100;
assign LUT_2[38448] = 32'b11111111111111111101111011110100;
assign LUT_2[38449] = 32'b11111111111111111010110100001101;
assign LUT_2[38450] = 32'b00000000000000000100110100110000;
assign LUT_2[38451] = 32'b00000000000000000001101101001001;
assign LUT_2[38452] = 32'b11111111111111111010011001011100;
assign LUT_2[38453] = 32'b11111111111111110111010001110101;
assign LUT_2[38454] = 32'b00000000000000000001010010011000;
assign LUT_2[38455] = 32'b11111111111111111110001010110001;
assign LUT_2[38456] = 32'b11111111111111111000101101010001;
assign LUT_2[38457] = 32'b11111111111111110101100101101010;
assign LUT_2[38458] = 32'b11111111111111111111100110001101;
assign LUT_2[38459] = 32'b11111111111111111100011110100110;
assign LUT_2[38460] = 32'b11111111111111110101001010111001;
assign LUT_2[38461] = 32'b11111111111111110010000011010010;
assign LUT_2[38462] = 32'b11111111111111111100000011110101;
assign LUT_2[38463] = 32'b11111111111111111000111100001110;
assign LUT_2[38464] = 32'b11111111111111111011000100100100;
assign LUT_2[38465] = 32'b11111111111111110111111100111101;
assign LUT_2[38466] = 32'b00000000000000000001111101100000;
assign LUT_2[38467] = 32'b11111111111111111110110101111001;
assign LUT_2[38468] = 32'b11111111111111110111100010001100;
assign LUT_2[38469] = 32'b11111111111111110100011010100101;
assign LUT_2[38470] = 32'b11111111111111111110011011001000;
assign LUT_2[38471] = 32'b11111111111111111011010011100001;
assign LUT_2[38472] = 32'b11111111111111110101110110000001;
assign LUT_2[38473] = 32'b11111111111111110010101110011010;
assign LUT_2[38474] = 32'b11111111111111111100101110111101;
assign LUT_2[38475] = 32'b11111111111111111001100111010110;
assign LUT_2[38476] = 32'b11111111111111110010010011101001;
assign LUT_2[38477] = 32'b11111111111111101111001100000010;
assign LUT_2[38478] = 32'b11111111111111111001001100100101;
assign LUT_2[38479] = 32'b11111111111111110110000100111110;
assign LUT_2[38480] = 32'b11111111111111110101101000101110;
assign LUT_2[38481] = 32'b11111111111111110010100001000111;
assign LUT_2[38482] = 32'b11111111111111111100100001101010;
assign LUT_2[38483] = 32'b11111111111111111001011010000011;
assign LUT_2[38484] = 32'b11111111111111110010000110010110;
assign LUT_2[38485] = 32'b11111111111111101110111110101111;
assign LUT_2[38486] = 32'b11111111111111111000111111010010;
assign LUT_2[38487] = 32'b11111111111111110101110111101011;
assign LUT_2[38488] = 32'b11111111111111110000011010001011;
assign LUT_2[38489] = 32'b11111111111111101101010010100100;
assign LUT_2[38490] = 32'b11111111111111110111010011000111;
assign LUT_2[38491] = 32'b11111111111111110100001011100000;
assign LUT_2[38492] = 32'b11111111111111101100110111110011;
assign LUT_2[38493] = 32'b11111111111111101001110000001100;
assign LUT_2[38494] = 32'b11111111111111110011110000101111;
assign LUT_2[38495] = 32'b11111111111111110000101001001000;
assign LUT_2[38496] = 32'b11111111111111111011100000001101;
assign LUT_2[38497] = 32'b11111111111111111000011000100110;
assign LUT_2[38498] = 32'b00000000000000000010011001001001;
assign LUT_2[38499] = 32'b11111111111111111111010001100010;
assign LUT_2[38500] = 32'b11111111111111110111111101110101;
assign LUT_2[38501] = 32'b11111111111111110100110110001110;
assign LUT_2[38502] = 32'b11111111111111111110110110110001;
assign LUT_2[38503] = 32'b11111111111111111011101111001010;
assign LUT_2[38504] = 32'b11111111111111110110010001101010;
assign LUT_2[38505] = 32'b11111111111111110011001010000011;
assign LUT_2[38506] = 32'b11111111111111111101001010100110;
assign LUT_2[38507] = 32'b11111111111111111010000010111111;
assign LUT_2[38508] = 32'b11111111111111110010101111010010;
assign LUT_2[38509] = 32'b11111111111111101111100111101011;
assign LUT_2[38510] = 32'b11111111111111111001101000001110;
assign LUT_2[38511] = 32'b11111111111111110110100000100111;
assign LUT_2[38512] = 32'b11111111111111110110000100010111;
assign LUT_2[38513] = 32'b11111111111111110010111100110000;
assign LUT_2[38514] = 32'b11111111111111111100111101010011;
assign LUT_2[38515] = 32'b11111111111111111001110101101100;
assign LUT_2[38516] = 32'b11111111111111110010100001111111;
assign LUT_2[38517] = 32'b11111111111111101111011010011000;
assign LUT_2[38518] = 32'b11111111111111111001011010111011;
assign LUT_2[38519] = 32'b11111111111111110110010011010100;
assign LUT_2[38520] = 32'b11111111111111110000110101110100;
assign LUT_2[38521] = 32'b11111111111111101101101110001101;
assign LUT_2[38522] = 32'b11111111111111110111101110110000;
assign LUT_2[38523] = 32'b11111111111111110100100111001001;
assign LUT_2[38524] = 32'b11111111111111101101010011011100;
assign LUT_2[38525] = 32'b11111111111111101010001011110101;
assign LUT_2[38526] = 32'b11111111111111110100001100011000;
assign LUT_2[38527] = 32'b11111111111111110001000100110001;
assign LUT_2[38528] = 32'b00000000000000000111010000010000;
assign LUT_2[38529] = 32'b00000000000000000100001000101001;
assign LUT_2[38530] = 32'b00000000000000001110001001001100;
assign LUT_2[38531] = 32'b00000000000000001011000001100101;
assign LUT_2[38532] = 32'b00000000000000000011101101111000;
assign LUT_2[38533] = 32'b00000000000000000000100110010001;
assign LUT_2[38534] = 32'b00000000000000001010100110110100;
assign LUT_2[38535] = 32'b00000000000000000111011111001101;
assign LUT_2[38536] = 32'b00000000000000000010000001101101;
assign LUT_2[38537] = 32'b11111111111111111110111010000110;
assign LUT_2[38538] = 32'b00000000000000001000111010101001;
assign LUT_2[38539] = 32'b00000000000000000101110011000010;
assign LUT_2[38540] = 32'b11111111111111111110011111010101;
assign LUT_2[38541] = 32'b11111111111111111011010111101110;
assign LUT_2[38542] = 32'b00000000000000000101011000010001;
assign LUT_2[38543] = 32'b00000000000000000010010000101010;
assign LUT_2[38544] = 32'b00000000000000000001110100011010;
assign LUT_2[38545] = 32'b11111111111111111110101100110011;
assign LUT_2[38546] = 32'b00000000000000001000101101010110;
assign LUT_2[38547] = 32'b00000000000000000101100101101111;
assign LUT_2[38548] = 32'b11111111111111111110010010000010;
assign LUT_2[38549] = 32'b11111111111111111011001010011011;
assign LUT_2[38550] = 32'b00000000000000000101001010111110;
assign LUT_2[38551] = 32'b00000000000000000010000011010111;
assign LUT_2[38552] = 32'b11111111111111111100100101110111;
assign LUT_2[38553] = 32'b11111111111111111001011110010000;
assign LUT_2[38554] = 32'b00000000000000000011011110110011;
assign LUT_2[38555] = 32'b00000000000000000000010111001100;
assign LUT_2[38556] = 32'b11111111111111111001000011011111;
assign LUT_2[38557] = 32'b11111111111111110101111011111000;
assign LUT_2[38558] = 32'b11111111111111111111111100011011;
assign LUT_2[38559] = 32'b11111111111111111100110100110100;
assign LUT_2[38560] = 32'b00000000000000000111101011111001;
assign LUT_2[38561] = 32'b00000000000000000100100100010010;
assign LUT_2[38562] = 32'b00000000000000001110100100110101;
assign LUT_2[38563] = 32'b00000000000000001011011101001110;
assign LUT_2[38564] = 32'b00000000000000000100001001100001;
assign LUT_2[38565] = 32'b00000000000000000001000001111010;
assign LUT_2[38566] = 32'b00000000000000001011000010011101;
assign LUT_2[38567] = 32'b00000000000000000111111010110110;
assign LUT_2[38568] = 32'b00000000000000000010011101010110;
assign LUT_2[38569] = 32'b11111111111111111111010101101111;
assign LUT_2[38570] = 32'b00000000000000001001010110010010;
assign LUT_2[38571] = 32'b00000000000000000110001110101011;
assign LUT_2[38572] = 32'b11111111111111111110111010111110;
assign LUT_2[38573] = 32'b11111111111111111011110011010111;
assign LUT_2[38574] = 32'b00000000000000000101110011111010;
assign LUT_2[38575] = 32'b00000000000000000010101100010011;
assign LUT_2[38576] = 32'b00000000000000000010010000000011;
assign LUT_2[38577] = 32'b11111111111111111111001000011100;
assign LUT_2[38578] = 32'b00000000000000001001001000111111;
assign LUT_2[38579] = 32'b00000000000000000110000001011000;
assign LUT_2[38580] = 32'b11111111111111111110101101101011;
assign LUT_2[38581] = 32'b11111111111111111011100110000100;
assign LUT_2[38582] = 32'b00000000000000000101100110100111;
assign LUT_2[38583] = 32'b00000000000000000010011111000000;
assign LUT_2[38584] = 32'b11111111111111111101000001100000;
assign LUT_2[38585] = 32'b11111111111111111001111001111001;
assign LUT_2[38586] = 32'b00000000000000000011111010011100;
assign LUT_2[38587] = 32'b00000000000000000000110010110101;
assign LUT_2[38588] = 32'b11111111111111111001011111001000;
assign LUT_2[38589] = 32'b11111111111111110110010111100001;
assign LUT_2[38590] = 32'b00000000000000000000011000000100;
assign LUT_2[38591] = 32'b11111111111111111101010000011101;
assign LUT_2[38592] = 32'b11111111111111111111011000110011;
assign LUT_2[38593] = 32'b11111111111111111100010001001100;
assign LUT_2[38594] = 32'b00000000000000000110010001101111;
assign LUT_2[38595] = 32'b00000000000000000011001010001000;
assign LUT_2[38596] = 32'b11111111111111111011110110011011;
assign LUT_2[38597] = 32'b11111111111111111000101110110100;
assign LUT_2[38598] = 32'b00000000000000000010101111010111;
assign LUT_2[38599] = 32'b11111111111111111111100111110000;
assign LUT_2[38600] = 32'b11111111111111111010001010010000;
assign LUT_2[38601] = 32'b11111111111111110111000010101001;
assign LUT_2[38602] = 32'b00000000000000000001000011001100;
assign LUT_2[38603] = 32'b11111111111111111101111011100101;
assign LUT_2[38604] = 32'b11111111111111110110100111111000;
assign LUT_2[38605] = 32'b11111111111111110011100000010001;
assign LUT_2[38606] = 32'b11111111111111111101100000110100;
assign LUT_2[38607] = 32'b11111111111111111010011001001101;
assign LUT_2[38608] = 32'b11111111111111111001111100111101;
assign LUT_2[38609] = 32'b11111111111111110110110101010110;
assign LUT_2[38610] = 32'b00000000000000000000110101111001;
assign LUT_2[38611] = 32'b11111111111111111101101110010010;
assign LUT_2[38612] = 32'b11111111111111110110011010100101;
assign LUT_2[38613] = 32'b11111111111111110011010010111110;
assign LUT_2[38614] = 32'b11111111111111111101010011100001;
assign LUT_2[38615] = 32'b11111111111111111010001011111010;
assign LUT_2[38616] = 32'b11111111111111110100101110011010;
assign LUT_2[38617] = 32'b11111111111111110001100110110011;
assign LUT_2[38618] = 32'b11111111111111111011100111010110;
assign LUT_2[38619] = 32'b11111111111111111000011111101111;
assign LUT_2[38620] = 32'b11111111111111110001001100000010;
assign LUT_2[38621] = 32'b11111111111111101110000100011011;
assign LUT_2[38622] = 32'b11111111111111111000000100111110;
assign LUT_2[38623] = 32'b11111111111111110100111101010111;
assign LUT_2[38624] = 32'b11111111111111111111110100011100;
assign LUT_2[38625] = 32'b11111111111111111100101100110101;
assign LUT_2[38626] = 32'b00000000000000000110101101011000;
assign LUT_2[38627] = 32'b00000000000000000011100101110001;
assign LUT_2[38628] = 32'b11111111111111111100010010000100;
assign LUT_2[38629] = 32'b11111111111111111001001010011101;
assign LUT_2[38630] = 32'b00000000000000000011001011000000;
assign LUT_2[38631] = 32'b00000000000000000000000011011001;
assign LUT_2[38632] = 32'b11111111111111111010100101111001;
assign LUT_2[38633] = 32'b11111111111111110111011110010010;
assign LUT_2[38634] = 32'b00000000000000000001011110110101;
assign LUT_2[38635] = 32'b11111111111111111110010111001110;
assign LUT_2[38636] = 32'b11111111111111110111000011100001;
assign LUT_2[38637] = 32'b11111111111111110011111011111010;
assign LUT_2[38638] = 32'b11111111111111111101111100011101;
assign LUT_2[38639] = 32'b11111111111111111010110100110110;
assign LUT_2[38640] = 32'b11111111111111111010011000100110;
assign LUT_2[38641] = 32'b11111111111111110111010000111111;
assign LUT_2[38642] = 32'b00000000000000000001010001100010;
assign LUT_2[38643] = 32'b11111111111111111110001001111011;
assign LUT_2[38644] = 32'b11111111111111110110110110001110;
assign LUT_2[38645] = 32'b11111111111111110011101110100111;
assign LUT_2[38646] = 32'b11111111111111111101101111001010;
assign LUT_2[38647] = 32'b11111111111111111010100111100011;
assign LUT_2[38648] = 32'b11111111111111110101001010000011;
assign LUT_2[38649] = 32'b11111111111111110010000010011100;
assign LUT_2[38650] = 32'b11111111111111111100000010111111;
assign LUT_2[38651] = 32'b11111111111111111000111011011000;
assign LUT_2[38652] = 32'b11111111111111110001100111101011;
assign LUT_2[38653] = 32'b11111111111111101110100000000100;
assign LUT_2[38654] = 32'b11111111111111111000100000100111;
assign LUT_2[38655] = 32'b11111111111111110101011001000000;
assign LUT_2[38656] = 32'b00000000000000000110111010100111;
assign LUT_2[38657] = 32'b00000000000000000011110011000000;
assign LUT_2[38658] = 32'b00000000000000001101110011100011;
assign LUT_2[38659] = 32'b00000000000000001010101011111100;
assign LUT_2[38660] = 32'b00000000000000000011011000001111;
assign LUT_2[38661] = 32'b00000000000000000000010000101000;
assign LUT_2[38662] = 32'b00000000000000001010010001001011;
assign LUT_2[38663] = 32'b00000000000000000111001001100100;
assign LUT_2[38664] = 32'b00000000000000000001101100000100;
assign LUT_2[38665] = 32'b11111111111111111110100100011101;
assign LUT_2[38666] = 32'b00000000000000001000100101000000;
assign LUT_2[38667] = 32'b00000000000000000101011101011001;
assign LUT_2[38668] = 32'b11111111111111111110001001101100;
assign LUT_2[38669] = 32'b11111111111111111011000010000101;
assign LUT_2[38670] = 32'b00000000000000000101000010101000;
assign LUT_2[38671] = 32'b00000000000000000001111011000001;
assign LUT_2[38672] = 32'b00000000000000000001011110110001;
assign LUT_2[38673] = 32'b11111111111111111110010111001010;
assign LUT_2[38674] = 32'b00000000000000001000010111101101;
assign LUT_2[38675] = 32'b00000000000000000101010000000110;
assign LUT_2[38676] = 32'b11111111111111111101111100011001;
assign LUT_2[38677] = 32'b11111111111111111010110100110010;
assign LUT_2[38678] = 32'b00000000000000000100110101010101;
assign LUT_2[38679] = 32'b00000000000000000001101101101110;
assign LUT_2[38680] = 32'b11111111111111111100010000001110;
assign LUT_2[38681] = 32'b11111111111111111001001000100111;
assign LUT_2[38682] = 32'b00000000000000000011001001001010;
assign LUT_2[38683] = 32'b00000000000000000000000001100011;
assign LUT_2[38684] = 32'b11111111111111111000101101110110;
assign LUT_2[38685] = 32'b11111111111111110101100110001111;
assign LUT_2[38686] = 32'b11111111111111111111100110110010;
assign LUT_2[38687] = 32'b11111111111111111100011111001011;
assign LUT_2[38688] = 32'b00000000000000000111010110010000;
assign LUT_2[38689] = 32'b00000000000000000100001110101001;
assign LUT_2[38690] = 32'b00000000000000001110001111001100;
assign LUT_2[38691] = 32'b00000000000000001011000111100101;
assign LUT_2[38692] = 32'b00000000000000000011110011111000;
assign LUT_2[38693] = 32'b00000000000000000000101100010001;
assign LUT_2[38694] = 32'b00000000000000001010101100110100;
assign LUT_2[38695] = 32'b00000000000000000111100101001101;
assign LUT_2[38696] = 32'b00000000000000000010000111101101;
assign LUT_2[38697] = 32'b11111111111111111111000000000110;
assign LUT_2[38698] = 32'b00000000000000001001000000101001;
assign LUT_2[38699] = 32'b00000000000000000101111001000010;
assign LUT_2[38700] = 32'b11111111111111111110100101010101;
assign LUT_2[38701] = 32'b11111111111111111011011101101110;
assign LUT_2[38702] = 32'b00000000000000000101011110010001;
assign LUT_2[38703] = 32'b00000000000000000010010110101010;
assign LUT_2[38704] = 32'b00000000000000000001111010011010;
assign LUT_2[38705] = 32'b11111111111111111110110010110011;
assign LUT_2[38706] = 32'b00000000000000001000110011010110;
assign LUT_2[38707] = 32'b00000000000000000101101011101111;
assign LUT_2[38708] = 32'b11111111111111111110011000000010;
assign LUT_2[38709] = 32'b11111111111111111011010000011011;
assign LUT_2[38710] = 32'b00000000000000000101010000111110;
assign LUT_2[38711] = 32'b00000000000000000010001001010111;
assign LUT_2[38712] = 32'b11111111111111111100101011110111;
assign LUT_2[38713] = 32'b11111111111111111001100100010000;
assign LUT_2[38714] = 32'b00000000000000000011100100110011;
assign LUT_2[38715] = 32'b00000000000000000000011101001100;
assign LUT_2[38716] = 32'b11111111111111111001001001011111;
assign LUT_2[38717] = 32'b11111111111111110110000001111000;
assign LUT_2[38718] = 32'b00000000000000000000000010011011;
assign LUT_2[38719] = 32'b11111111111111111100111010110100;
assign LUT_2[38720] = 32'b11111111111111111111000011001010;
assign LUT_2[38721] = 32'b11111111111111111011111011100011;
assign LUT_2[38722] = 32'b00000000000000000101111100000110;
assign LUT_2[38723] = 32'b00000000000000000010110100011111;
assign LUT_2[38724] = 32'b11111111111111111011100000110010;
assign LUT_2[38725] = 32'b11111111111111111000011001001011;
assign LUT_2[38726] = 32'b00000000000000000010011001101110;
assign LUT_2[38727] = 32'b11111111111111111111010010000111;
assign LUT_2[38728] = 32'b11111111111111111001110100100111;
assign LUT_2[38729] = 32'b11111111111111110110101101000000;
assign LUT_2[38730] = 32'b00000000000000000000101101100011;
assign LUT_2[38731] = 32'b11111111111111111101100101111100;
assign LUT_2[38732] = 32'b11111111111111110110010010001111;
assign LUT_2[38733] = 32'b11111111111111110011001010101000;
assign LUT_2[38734] = 32'b11111111111111111101001011001011;
assign LUT_2[38735] = 32'b11111111111111111010000011100100;
assign LUT_2[38736] = 32'b11111111111111111001100111010100;
assign LUT_2[38737] = 32'b11111111111111110110011111101101;
assign LUT_2[38738] = 32'b00000000000000000000100000010000;
assign LUT_2[38739] = 32'b11111111111111111101011000101001;
assign LUT_2[38740] = 32'b11111111111111110110000100111100;
assign LUT_2[38741] = 32'b11111111111111110010111101010101;
assign LUT_2[38742] = 32'b11111111111111111100111101111000;
assign LUT_2[38743] = 32'b11111111111111111001110110010001;
assign LUT_2[38744] = 32'b11111111111111110100011000110001;
assign LUT_2[38745] = 32'b11111111111111110001010001001010;
assign LUT_2[38746] = 32'b11111111111111111011010001101101;
assign LUT_2[38747] = 32'b11111111111111111000001010000110;
assign LUT_2[38748] = 32'b11111111111111110000110110011001;
assign LUT_2[38749] = 32'b11111111111111101101101110110010;
assign LUT_2[38750] = 32'b11111111111111110111101111010101;
assign LUT_2[38751] = 32'b11111111111111110100100111101110;
assign LUT_2[38752] = 32'b11111111111111111111011110110011;
assign LUT_2[38753] = 32'b11111111111111111100010111001100;
assign LUT_2[38754] = 32'b00000000000000000110010111101111;
assign LUT_2[38755] = 32'b00000000000000000011010000001000;
assign LUT_2[38756] = 32'b11111111111111111011111100011011;
assign LUT_2[38757] = 32'b11111111111111111000110100110100;
assign LUT_2[38758] = 32'b00000000000000000010110101010111;
assign LUT_2[38759] = 32'b11111111111111111111101101110000;
assign LUT_2[38760] = 32'b11111111111111111010010000010000;
assign LUT_2[38761] = 32'b11111111111111110111001000101001;
assign LUT_2[38762] = 32'b00000000000000000001001001001100;
assign LUT_2[38763] = 32'b11111111111111111110000001100101;
assign LUT_2[38764] = 32'b11111111111111110110101101111000;
assign LUT_2[38765] = 32'b11111111111111110011100110010001;
assign LUT_2[38766] = 32'b11111111111111111101100110110100;
assign LUT_2[38767] = 32'b11111111111111111010011111001101;
assign LUT_2[38768] = 32'b11111111111111111010000010111101;
assign LUT_2[38769] = 32'b11111111111111110110111011010110;
assign LUT_2[38770] = 32'b00000000000000000000111011111001;
assign LUT_2[38771] = 32'b11111111111111111101110100010010;
assign LUT_2[38772] = 32'b11111111111111110110100000100101;
assign LUT_2[38773] = 32'b11111111111111110011011000111110;
assign LUT_2[38774] = 32'b11111111111111111101011001100001;
assign LUT_2[38775] = 32'b11111111111111111010010001111010;
assign LUT_2[38776] = 32'b11111111111111110100110100011010;
assign LUT_2[38777] = 32'b11111111111111110001101100110011;
assign LUT_2[38778] = 32'b11111111111111111011101101010110;
assign LUT_2[38779] = 32'b11111111111111111000100101101111;
assign LUT_2[38780] = 32'b11111111111111110001010010000010;
assign LUT_2[38781] = 32'b11111111111111101110001010011011;
assign LUT_2[38782] = 32'b11111111111111111000001010111110;
assign LUT_2[38783] = 32'b11111111111111110101000011010111;
assign LUT_2[38784] = 32'b00000000000000001011001110110110;
assign LUT_2[38785] = 32'b00000000000000001000000111001111;
assign LUT_2[38786] = 32'b00000000000000010010000111110010;
assign LUT_2[38787] = 32'b00000000000000001111000000001011;
assign LUT_2[38788] = 32'b00000000000000000111101100011110;
assign LUT_2[38789] = 32'b00000000000000000100100100110111;
assign LUT_2[38790] = 32'b00000000000000001110100101011010;
assign LUT_2[38791] = 32'b00000000000000001011011101110011;
assign LUT_2[38792] = 32'b00000000000000000110000000010011;
assign LUT_2[38793] = 32'b00000000000000000010111000101100;
assign LUT_2[38794] = 32'b00000000000000001100111001001111;
assign LUT_2[38795] = 32'b00000000000000001001110001101000;
assign LUT_2[38796] = 32'b00000000000000000010011101111011;
assign LUT_2[38797] = 32'b11111111111111111111010110010100;
assign LUT_2[38798] = 32'b00000000000000001001010110110111;
assign LUT_2[38799] = 32'b00000000000000000110001111010000;
assign LUT_2[38800] = 32'b00000000000000000101110011000000;
assign LUT_2[38801] = 32'b00000000000000000010101011011001;
assign LUT_2[38802] = 32'b00000000000000001100101011111100;
assign LUT_2[38803] = 32'b00000000000000001001100100010101;
assign LUT_2[38804] = 32'b00000000000000000010010000101000;
assign LUT_2[38805] = 32'b11111111111111111111001001000001;
assign LUT_2[38806] = 32'b00000000000000001001001001100100;
assign LUT_2[38807] = 32'b00000000000000000110000001111101;
assign LUT_2[38808] = 32'b00000000000000000000100100011101;
assign LUT_2[38809] = 32'b11111111111111111101011100110110;
assign LUT_2[38810] = 32'b00000000000000000111011101011001;
assign LUT_2[38811] = 32'b00000000000000000100010101110010;
assign LUT_2[38812] = 32'b11111111111111111101000010000101;
assign LUT_2[38813] = 32'b11111111111111111001111010011110;
assign LUT_2[38814] = 32'b00000000000000000011111011000001;
assign LUT_2[38815] = 32'b00000000000000000000110011011010;
assign LUT_2[38816] = 32'b00000000000000001011101010011111;
assign LUT_2[38817] = 32'b00000000000000001000100010111000;
assign LUT_2[38818] = 32'b00000000000000010010100011011011;
assign LUT_2[38819] = 32'b00000000000000001111011011110100;
assign LUT_2[38820] = 32'b00000000000000001000001000000111;
assign LUT_2[38821] = 32'b00000000000000000101000000100000;
assign LUT_2[38822] = 32'b00000000000000001111000001000011;
assign LUT_2[38823] = 32'b00000000000000001011111001011100;
assign LUT_2[38824] = 32'b00000000000000000110011011111100;
assign LUT_2[38825] = 32'b00000000000000000011010100010101;
assign LUT_2[38826] = 32'b00000000000000001101010100111000;
assign LUT_2[38827] = 32'b00000000000000001010001101010001;
assign LUT_2[38828] = 32'b00000000000000000010111001100100;
assign LUT_2[38829] = 32'b11111111111111111111110001111101;
assign LUT_2[38830] = 32'b00000000000000001001110010100000;
assign LUT_2[38831] = 32'b00000000000000000110101010111001;
assign LUT_2[38832] = 32'b00000000000000000110001110101001;
assign LUT_2[38833] = 32'b00000000000000000011000111000010;
assign LUT_2[38834] = 32'b00000000000000001101000111100101;
assign LUT_2[38835] = 32'b00000000000000001001111111111110;
assign LUT_2[38836] = 32'b00000000000000000010101100010001;
assign LUT_2[38837] = 32'b11111111111111111111100100101010;
assign LUT_2[38838] = 32'b00000000000000001001100101001101;
assign LUT_2[38839] = 32'b00000000000000000110011101100110;
assign LUT_2[38840] = 32'b00000000000000000001000000000110;
assign LUT_2[38841] = 32'b11111111111111111101111000011111;
assign LUT_2[38842] = 32'b00000000000000000111111001000010;
assign LUT_2[38843] = 32'b00000000000000000100110001011011;
assign LUT_2[38844] = 32'b11111111111111111101011101101110;
assign LUT_2[38845] = 32'b11111111111111111010010110000111;
assign LUT_2[38846] = 32'b00000000000000000100010110101010;
assign LUT_2[38847] = 32'b00000000000000000001001111000011;
assign LUT_2[38848] = 32'b00000000000000000011010111011001;
assign LUT_2[38849] = 32'b00000000000000000000001111110010;
assign LUT_2[38850] = 32'b00000000000000001010010000010101;
assign LUT_2[38851] = 32'b00000000000000000111001000101110;
assign LUT_2[38852] = 32'b11111111111111111111110101000001;
assign LUT_2[38853] = 32'b11111111111111111100101101011010;
assign LUT_2[38854] = 32'b00000000000000000110101101111101;
assign LUT_2[38855] = 32'b00000000000000000011100110010110;
assign LUT_2[38856] = 32'b11111111111111111110001000110110;
assign LUT_2[38857] = 32'b11111111111111111011000001001111;
assign LUT_2[38858] = 32'b00000000000000000101000001110010;
assign LUT_2[38859] = 32'b00000000000000000001111010001011;
assign LUT_2[38860] = 32'b11111111111111111010100110011110;
assign LUT_2[38861] = 32'b11111111111111110111011110110111;
assign LUT_2[38862] = 32'b00000000000000000001011111011010;
assign LUT_2[38863] = 32'b11111111111111111110010111110011;
assign LUT_2[38864] = 32'b11111111111111111101111011100011;
assign LUT_2[38865] = 32'b11111111111111111010110011111100;
assign LUT_2[38866] = 32'b00000000000000000100110100011111;
assign LUT_2[38867] = 32'b00000000000000000001101100111000;
assign LUT_2[38868] = 32'b11111111111111111010011001001011;
assign LUT_2[38869] = 32'b11111111111111110111010001100100;
assign LUT_2[38870] = 32'b00000000000000000001010010000111;
assign LUT_2[38871] = 32'b11111111111111111110001010100000;
assign LUT_2[38872] = 32'b11111111111111111000101101000000;
assign LUT_2[38873] = 32'b11111111111111110101100101011001;
assign LUT_2[38874] = 32'b11111111111111111111100101111100;
assign LUT_2[38875] = 32'b11111111111111111100011110010101;
assign LUT_2[38876] = 32'b11111111111111110101001010101000;
assign LUT_2[38877] = 32'b11111111111111110010000011000001;
assign LUT_2[38878] = 32'b11111111111111111100000011100100;
assign LUT_2[38879] = 32'b11111111111111111000111011111101;
assign LUT_2[38880] = 32'b00000000000000000011110011000010;
assign LUT_2[38881] = 32'b00000000000000000000101011011011;
assign LUT_2[38882] = 32'b00000000000000001010101011111110;
assign LUT_2[38883] = 32'b00000000000000000111100100010111;
assign LUT_2[38884] = 32'b00000000000000000000010000101010;
assign LUT_2[38885] = 32'b11111111111111111101001001000011;
assign LUT_2[38886] = 32'b00000000000000000111001001100110;
assign LUT_2[38887] = 32'b00000000000000000100000001111111;
assign LUT_2[38888] = 32'b11111111111111111110100100011111;
assign LUT_2[38889] = 32'b11111111111111111011011100111000;
assign LUT_2[38890] = 32'b00000000000000000101011101011011;
assign LUT_2[38891] = 32'b00000000000000000010010101110100;
assign LUT_2[38892] = 32'b11111111111111111011000010000111;
assign LUT_2[38893] = 32'b11111111111111110111111010100000;
assign LUT_2[38894] = 32'b00000000000000000001111011000011;
assign LUT_2[38895] = 32'b11111111111111111110110011011100;
assign LUT_2[38896] = 32'b11111111111111111110010111001100;
assign LUT_2[38897] = 32'b11111111111111111011001111100101;
assign LUT_2[38898] = 32'b00000000000000000101010000001000;
assign LUT_2[38899] = 32'b00000000000000000010001000100001;
assign LUT_2[38900] = 32'b11111111111111111010110100110100;
assign LUT_2[38901] = 32'b11111111111111110111101101001101;
assign LUT_2[38902] = 32'b00000000000000000001101101110000;
assign LUT_2[38903] = 32'b11111111111111111110100110001001;
assign LUT_2[38904] = 32'b11111111111111111001001000101001;
assign LUT_2[38905] = 32'b11111111111111110110000001000010;
assign LUT_2[38906] = 32'b00000000000000000000000001100101;
assign LUT_2[38907] = 32'b11111111111111111100111001111110;
assign LUT_2[38908] = 32'b11111111111111110101100110010001;
assign LUT_2[38909] = 32'b11111111111111110010011110101010;
assign LUT_2[38910] = 32'b11111111111111111100011111001101;
assign LUT_2[38911] = 32'b11111111111111111001010111100110;
assign LUT_2[38912] = 32'b11111111111111110011010100000110;
assign LUT_2[38913] = 32'b11111111111111110000001100011111;
assign LUT_2[38914] = 32'b11111111111111111010001101000010;
assign LUT_2[38915] = 32'b11111111111111110111000101011011;
assign LUT_2[38916] = 32'b11111111111111101111110001101110;
assign LUT_2[38917] = 32'b11111111111111101100101010000111;
assign LUT_2[38918] = 32'b11111111111111110110101010101010;
assign LUT_2[38919] = 32'b11111111111111110011100011000011;
assign LUT_2[38920] = 32'b11111111111111101110000101100011;
assign LUT_2[38921] = 32'b11111111111111101010111101111100;
assign LUT_2[38922] = 32'b11111111111111110100111110011111;
assign LUT_2[38923] = 32'b11111111111111110001110110111000;
assign LUT_2[38924] = 32'b11111111111111101010100011001011;
assign LUT_2[38925] = 32'b11111111111111100111011011100100;
assign LUT_2[38926] = 32'b11111111111111110001011100000111;
assign LUT_2[38927] = 32'b11111111111111101110010100100000;
assign LUT_2[38928] = 32'b11111111111111101101111000010000;
assign LUT_2[38929] = 32'b11111111111111101010110000101001;
assign LUT_2[38930] = 32'b11111111111111110100110001001100;
assign LUT_2[38931] = 32'b11111111111111110001101001100101;
assign LUT_2[38932] = 32'b11111111111111101010010101111000;
assign LUT_2[38933] = 32'b11111111111111100111001110010001;
assign LUT_2[38934] = 32'b11111111111111110001001110110100;
assign LUT_2[38935] = 32'b11111111111111101110000111001101;
assign LUT_2[38936] = 32'b11111111111111101000101001101101;
assign LUT_2[38937] = 32'b11111111111111100101100010000110;
assign LUT_2[38938] = 32'b11111111111111101111100010101001;
assign LUT_2[38939] = 32'b11111111111111101100011011000010;
assign LUT_2[38940] = 32'b11111111111111100101000111010101;
assign LUT_2[38941] = 32'b11111111111111100001111111101110;
assign LUT_2[38942] = 32'b11111111111111101100000000010001;
assign LUT_2[38943] = 32'b11111111111111101000111000101010;
assign LUT_2[38944] = 32'b11111111111111110011101111101111;
assign LUT_2[38945] = 32'b11111111111111110000101000001000;
assign LUT_2[38946] = 32'b11111111111111111010101000101011;
assign LUT_2[38947] = 32'b11111111111111110111100001000100;
assign LUT_2[38948] = 32'b11111111111111110000001101010111;
assign LUT_2[38949] = 32'b11111111111111101101000101110000;
assign LUT_2[38950] = 32'b11111111111111110111000110010011;
assign LUT_2[38951] = 32'b11111111111111110011111110101100;
assign LUT_2[38952] = 32'b11111111111111101110100001001100;
assign LUT_2[38953] = 32'b11111111111111101011011001100101;
assign LUT_2[38954] = 32'b11111111111111110101011010001000;
assign LUT_2[38955] = 32'b11111111111111110010010010100001;
assign LUT_2[38956] = 32'b11111111111111101010111110110100;
assign LUT_2[38957] = 32'b11111111111111100111110111001101;
assign LUT_2[38958] = 32'b11111111111111110001110111110000;
assign LUT_2[38959] = 32'b11111111111111101110110000001001;
assign LUT_2[38960] = 32'b11111111111111101110010011111001;
assign LUT_2[38961] = 32'b11111111111111101011001100010010;
assign LUT_2[38962] = 32'b11111111111111110101001100110101;
assign LUT_2[38963] = 32'b11111111111111110010000101001110;
assign LUT_2[38964] = 32'b11111111111111101010110001100001;
assign LUT_2[38965] = 32'b11111111111111100111101001111010;
assign LUT_2[38966] = 32'b11111111111111110001101010011101;
assign LUT_2[38967] = 32'b11111111111111101110100010110110;
assign LUT_2[38968] = 32'b11111111111111101001000101010110;
assign LUT_2[38969] = 32'b11111111111111100101111101101111;
assign LUT_2[38970] = 32'b11111111111111101111111110010010;
assign LUT_2[38971] = 32'b11111111111111101100110110101011;
assign LUT_2[38972] = 32'b11111111111111100101100010111110;
assign LUT_2[38973] = 32'b11111111111111100010011011010111;
assign LUT_2[38974] = 32'b11111111111111101100011011111010;
assign LUT_2[38975] = 32'b11111111111111101001010100010011;
assign LUT_2[38976] = 32'b11111111111111101011011100101001;
assign LUT_2[38977] = 32'b11111111111111101000010101000010;
assign LUT_2[38978] = 32'b11111111111111110010010101100101;
assign LUT_2[38979] = 32'b11111111111111101111001101111110;
assign LUT_2[38980] = 32'b11111111111111100111111010010001;
assign LUT_2[38981] = 32'b11111111111111100100110010101010;
assign LUT_2[38982] = 32'b11111111111111101110110011001101;
assign LUT_2[38983] = 32'b11111111111111101011101011100110;
assign LUT_2[38984] = 32'b11111111111111100110001110000110;
assign LUT_2[38985] = 32'b11111111111111100011000110011111;
assign LUT_2[38986] = 32'b11111111111111101101000111000010;
assign LUT_2[38987] = 32'b11111111111111101001111111011011;
assign LUT_2[38988] = 32'b11111111111111100010101011101110;
assign LUT_2[38989] = 32'b11111111111111011111100100000111;
assign LUT_2[38990] = 32'b11111111111111101001100100101010;
assign LUT_2[38991] = 32'b11111111111111100110011101000011;
assign LUT_2[38992] = 32'b11111111111111100110000000110011;
assign LUT_2[38993] = 32'b11111111111111100010111001001100;
assign LUT_2[38994] = 32'b11111111111111101100111001101111;
assign LUT_2[38995] = 32'b11111111111111101001110010001000;
assign LUT_2[38996] = 32'b11111111111111100010011110011011;
assign LUT_2[38997] = 32'b11111111111111011111010110110100;
assign LUT_2[38998] = 32'b11111111111111101001010111010111;
assign LUT_2[38999] = 32'b11111111111111100110001111110000;
assign LUT_2[39000] = 32'b11111111111111100000110010010000;
assign LUT_2[39001] = 32'b11111111111111011101101010101001;
assign LUT_2[39002] = 32'b11111111111111100111101011001100;
assign LUT_2[39003] = 32'b11111111111111100100100011100101;
assign LUT_2[39004] = 32'b11111111111111011101001111111000;
assign LUT_2[39005] = 32'b11111111111111011010001000010001;
assign LUT_2[39006] = 32'b11111111111111100100001000110100;
assign LUT_2[39007] = 32'b11111111111111100001000001001101;
assign LUT_2[39008] = 32'b11111111111111101011111000010010;
assign LUT_2[39009] = 32'b11111111111111101000110000101011;
assign LUT_2[39010] = 32'b11111111111111110010110001001110;
assign LUT_2[39011] = 32'b11111111111111101111101001100111;
assign LUT_2[39012] = 32'b11111111111111101000010101111010;
assign LUT_2[39013] = 32'b11111111111111100101001110010011;
assign LUT_2[39014] = 32'b11111111111111101111001110110110;
assign LUT_2[39015] = 32'b11111111111111101100000111001111;
assign LUT_2[39016] = 32'b11111111111111100110101001101111;
assign LUT_2[39017] = 32'b11111111111111100011100010001000;
assign LUT_2[39018] = 32'b11111111111111101101100010101011;
assign LUT_2[39019] = 32'b11111111111111101010011011000100;
assign LUT_2[39020] = 32'b11111111111111100011000111010111;
assign LUT_2[39021] = 32'b11111111111111011111111111110000;
assign LUT_2[39022] = 32'b11111111111111101010000000010011;
assign LUT_2[39023] = 32'b11111111111111100110111000101100;
assign LUT_2[39024] = 32'b11111111111111100110011100011100;
assign LUT_2[39025] = 32'b11111111111111100011010100110101;
assign LUT_2[39026] = 32'b11111111111111101101010101011000;
assign LUT_2[39027] = 32'b11111111111111101010001101110001;
assign LUT_2[39028] = 32'b11111111111111100010111010000100;
assign LUT_2[39029] = 32'b11111111111111011111110010011101;
assign LUT_2[39030] = 32'b11111111111111101001110011000000;
assign LUT_2[39031] = 32'b11111111111111100110101011011001;
assign LUT_2[39032] = 32'b11111111111111100001001101111001;
assign LUT_2[39033] = 32'b11111111111111011110000110010010;
assign LUT_2[39034] = 32'b11111111111111101000000110110101;
assign LUT_2[39035] = 32'b11111111111111100100111111001110;
assign LUT_2[39036] = 32'b11111111111111011101101011100001;
assign LUT_2[39037] = 32'b11111111111111011010100011111010;
assign LUT_2[39038] = 32'b11111111111111100100100100011101;
assign LUT_2[39039] = 32'b11111111111111100001011100110110;
assign LUT_2[39040] = 32'b11111111111111110111101000010101;
assign LUT_2[39041] = 32'b11111111111111110100100000101110;
assign LUT_2[39042] = 32'b11111111111111111110100001010001;
assign LUT_2[39043] = 32'b11111111111111111011011001101010;
assign LUT_2[39044] = 32'b11111111111111110100000101111101;
assign LUT_2[39045] = 32'b11111111111111110000111110010110;
assign LUT_2[39046] = 32'b11111111111111111010111110111001;
assign LUT_2[39047] = 32'b11111111111111110111110111010010;
assign LUT_2[39048] = 32'b11111111111111110010011001110010;
assign LUT_2[39049] = 32'b11111111111111101111010010001011;
assign LUT_2[39050] = 32'b11111111111111111001010010101110;
assign LUT_2[39051] = 32'b11111111111111110110001011000111;
assign LUT_2[39052] = 32'b11111111111111101110110111011010;
assign LUT_2[39053] = 32'b11111111111111101011101111110011;
assign LUT_2[39054] = 32'b11111111111111110101110000010110;
assign LUT_2[39055] = 32'b11111111111111110010101000101111;
assign LUT_2[39056] = 32'b11111111111111110010001100011111;
assign LUT_2[39057] = 32'b11111111111111101111000100111000;
assign LUT_2[39058] = 32'b11111111111111111001000101011011;
assign LUT_2[39059] = 32'b11111111111111110101111101110100;
assign LUT_2[39060] = 32'b11111111111111101110101010000111;
assign LUT_2[39061] = 32'b11111111111111101011100010100000;
assign LUT_2[39062] = 32'b11111111111111110101100011000011;
assign LUT_2[39063] = 32'b11111111111111110010011011011100;
assign LUT_2[39064] = 32'b11111111111111101100111101111100;
assign LUT_2[39065] = 32'b11111111111111101001110110010101;
assign LUT_2[39066] = 32'b11111111111111110011110110111000;
assign LUT_2[39067] = 32'b11111111111111110000101111010001;
assign LUT_2[39068] = 32'b11111111111111101001011011100100;
assign LUT_2[39069] = 32'b11111111111111100110010011111101;
assign LUT_2[39070] = 32'b11111111111111110000010100100000;
assign LUT_2[39071] = 32'b11111111111111101101001100111001;
assign LUT_2[39072] = 32'b11111111111111111000000011111110;
assign LUT_2[39073] = 32'b11111111111111110100111100010111;
assign LUT_2[39074] = 32'b11111111111111111110111100111010;
assign LUT_2[39075] = 32'b11111111111111111011110101010011;
assign LUT_2[39076] = 32'b11111111111111110100100001100110;
assign LUT_2[39077] = 32'b11111111111111110001011001111111;
assign LUT_2[39078] = 32'b11111111111111111011011010100010;
assign LUT_2[39079] = 32'b11111111111111111000010010111011;
assign LUT_2[39080] = 32'b11111111111111110010110101011011;
assign LUT_2[39081] = 32'b11111111111111101111101101110100;
assign LUT_2[39082] = 32'b11111111111111111001101110010111;
assign LUT_2[39083] = 32'b11111111111111110110100110110000;
assign LUT_2[39084] = 32'b11111111111111101111010011000011;
assign LUT_2[39085] = 32'b11111111111111101100001011011100;
assign LUT_2[39086] = 32'b11111111111111110110001011111111;
assign LUT_2[39087] = 32'b11111111111111110011000100011000;
assign LUT_2[39088] = 32'b11111111111111110010101000001000;
assign LUT_2[39089] = 32'b11111111111111101111100000100001;
assign LUT_2[39090] = 32'b11111111111111111001100001000100;
assign LUT_2[39091] = 32'b11111111111111110110011001011101;
assign LUT_2[39092] = 32'b11111111111111101111000101110000;
assign LUT_2[39093] = 32'b11111111111111101011111110001001;
assign LUT_2[39094] = 32'b11111111111111110101111110101100;
assign LUT_2[39095] = 32'b11111111111111110010110111000101;
assign LUT_2[39096] = 32'b11111111111111101101011001100101;
assign LUT_2[39097] = 32'b11111111111111101010010001111110;
assign LUT_2[39098] = 32'b11111111111111110100010010100001;
assign LUT_2[39099] = 32'b11111111111111110001001010111010;
assign LUT_2[39100] = 32'b11111111111111101001110111001101;
assign LUT_2[39101] = 32'b11111111111111100110101111100110;
assign LUT_2[39102] = 32'b11111111111111110000110000001001;
assign LUT_2[39103] = 32'b11111111111111101101101000100010;
assign LUT_2[39104] = 32'b11111111111111101111110000111000;
assign LUT_2[39105] = 32'b11111111111111101100101001010001;
assign LUT_2[39106] = 32'b11111111111111110110101001110100;
assign LUT_2[39107] = 32'b11111111111111110011100010001101;
assign LUT_2[39108] = 32'b11111111111111101100001110100000;
assign LUT_2[39109] = 32'b11111111111111101001000110111001;
assign LUT_2[39110] = 32'b11111111111111110011000111011100;
assign LUT_2[39111] = 32'b11111111111111101111111111110101;
assign LUT_2[39112] = 32'b11111111111111101010100010010101;
assign LUT_2[39113] = 32'b11111111111111100111011010101110;
assign LUT_2[39114] = 32'b11111111111111110001011011010001;
assign LUT_2[39115] = 32'b11111111111111101110010011101010;
assign LUT_2[39116] = 32'b11111111111111100110111111111101;
assign LUT_2[39117] = 32'b11111111111111100011111000010110;
assign LUT_2[39118] = 32'b11111111111111101101111000111001;
assign LUT_2[39119] = 32'b11111111111111101010110001010010;
assign LUT_2[39120] = 32'b11111111111111101010010101000010;
assign LUT_2[39121] = 32'b11111111111111100111001101011011;
assign LUT_2[39122] = 32'b11111111111111110001001101111110;
assign LUT_2[39123] = 32'b11111111111111101110000110010111;
assign LUT_2[39124] = 32'b11111111111111100110110010101010;
assign LUT_2[39125] = 32'b11111111111111100011101011000011;
assign LUT_2[39126] = 32'b11111111111111101101101011100110;
assign LUT_2[39127] = 32'b11111111111111101010100011111111;
assign LUT_2[39128] = 32'b11111111111111100101000110011111;
assign LUT_2[39129] = 32'b11111111111111100001111110111000;
assign LUT_2[39130] = 32'b11111111111111101011111111011011;
assign LUT_2[39131] = 32'b11111111111111101000110111110100;
assign LUT_2[39132] = 32'b11111111111111100001100100000111;
assign LUT_2[39133] = 32'b11111111111111011110011100100000;
assign LUT_2[39134] = 32'b11111111111111101000011101000011;
assign LUT_2[39135] = 32'b11111111111111100101010101011100;
assign LUT_2[39136] = 32'b11111111111111110000001100100001;
assign LUT_2[39137] = 32'b11111111111111101101000100111010;
assign LUT_2[39138] = 32'b11111111111111110111000101011101;
assign LUT_2[39139] = 32'b11111111111111110011111101110110;
assign LUT_2[39140] = 32'b11111111111111101100101010001001;
assign LUT_2[39141] = 32'b11111111111111101001100010100010;
assign LUT_2[39142] = 32'b11111111111111110011100011000101;
assign LUT_2[39143] = 32'b11111111111111110000011011011110;
assign LUT_2[39144] = 32'b11111111111111101010111101111110;
assign LUT_2[39145] = 32'b11111111111111100111110110010111;
assign LUT_2[39146] = 32'b11111111111111110001110110111010;
assign LUT_2[39147] = 32'b11111111111111101110101111010011;
assign LUT_2[39148] = 32'b11111111111111100111011011100110;
assign LUT_2[39149] = 32'b11111111111111100100010011111111;
assign LUT_2[39150] = 32'b11111111111111101110010100100010;
assign LUT_2[39151] = 32'b11111111111111101011001100111011;
assign LUT_2[39152] = 32'b11111111111111101010110000101011;
assign LUT_2[39153] = 32'b11111111111111100111101001000100;
assign LUT_2[39154] = 32'b11111111111111110001101001100111;
assign LUT_2[39155] = 32'b11111111111111101110100010000000;
assign LUT_2[39156] = 32'b11111111111111100111001110010011;
assign LUT_2[39157] = 32'b11111111111111100100000110101100;
assign LUT_2[39158] = 32'b11111111111111101110000111001111;
assign LUT_2[39159] = 32'b11111111111111101010111111101000;
assign LUT_2[39160] = 32'b11111111111111100101100010001000;
assign LUT_2[39161] = 32'b11111111111111100010011010100001;
assign LUT_2[39162] = 32'b11111111111111101100011011000100;
assign LUT_2[39163] = 32'b11111111111111101001010011011101;
assign LUT_2[39164] = 32'b11111111111111100001111111110000;
assign LUT_2[39165] = 32'b11111111111111011110111000001001;
assign LUT_2[39166] = 32'b11111111111111101000111000101100;
assign LUT_2[39167] = 32'b11111111111111100101110001000101;
assign LUT_2[39168] = 32'b11111111111111110111010010101100;
assign LUT_2[39169] = 32'b11111111111111110100001011000101;
assign LUT_2[39170] = 32'b11111111111111111110001011101000;
assign LUT_2[39171] = 32'b11111111111111111011000100000001;
assign LUT_2[39172] = 32'b11111111111111110011110000010100;
assign LUT_2[39173] = 32'b11111111111111110000101000101101;
assign LUT_2[39174] = 32'b11111111111111111010101001010000;
assign LUT_2[39175] = 32'b11111111111111110111100001101001;
assign LUT_2[39176] = 32'b11111111111111110010000100001001;
assign LUT_2[39177] = 32'b11111111111111101110111100100010;
assign LUT_2[39178] = 32'b11111111111111111000111101000101;
assign LUT_2[39179] = 32'b11111111111111110101110101011110;
assign LUT_2[39180] = 32'b11111111111111101110100001110001;
assign LUT_2[39181] = 32'b11111111111111101011011010001010;
assign LUT_2[39182] = 32'b11111111111111110101011010101101;
assign LUT_2[39183] = 32'b11111111111111110010010011000110;
assign LUT_2[39184] = 32'b11111111111111110001110110110110;
assign LUT_2[39185] = 32'b11111111111111101110101111001111;
assign LUT_2[39186] = 32'b11111111111111111000101111110010;
assign LUT_2[39187] = 32'b11111111111111110101101000001011;
assign LUT_2[39188] = 32'b11111111111111101110010100011110;
assign LUT_2[39189] = 32'b11111111111111101011001100110111;
assign LUT_2[39190] = 32'b11111111111111110101001101011010;
assign LUT_2[39191] = 32'b11111111111111110010000101110011;
assign LUT_2[39192] = 32'b11111111111111101100101000010011;
assign LUT_2[39193] = 32'b11111111111111101001100000101100;
assign LUT_2[39194] = 32'b11111111111111110011100001001111;
assign LUT_2[39195] = 32'b11111111111111110000011001101000;
assign LUT_2[39196] = 32'b11111111111111101001000101111011;
assign LUT_2[39197] = 32'b11111111111111100101111110010100;
assign LUT_2[39198] = 32'b11111111111111101111111110110111;
assign LUT_2[39199] = 32'b11111111111111101100110111010000;
assign LUT_2[39200] = 32'b11111111111111110111101110010101;
assign LUT_2[39201] = 32'b11111111111111110100100110101110;
assign LUT_2[39202] = 32'b11111111111111111110100111010001;
assign LUT_2[39203] = 32'b11111111111111111011011111101010;
assign LUT_2[39204] = 32'b11111111111111110100001011111101;
assign LUT_2[39205] = 32'b11111111111111110001000100010110;
assign LUT_2[39206] = 32'b11111111111111111011000100111001;
assign LUT_2[39207] = 32'b11111111111111110111111101010010;
assign LUT_2[39208] = 32'b11111111111111110010011111110010;
assign LUT_2[39209] = 32'b11111111111111101111011000001011;
assign LUT_2[39210] = 32'b11111111111111111001011000101110;
assign LUT_2[39211] = 32'b11111111111111110110010001000111;
assign LUT_2[39212] = 32'b11111111111111101110111101011010;
assign LUT_2[39213] = 32'b11111111111111101011110101110011;
assign LUT_2[39214] = 32'b11111111111111110101110110010110;
assign LUT_2[39215] = 32'b11111111111111110010101110101111;
assign LUT_2[39216] = 32'b11111111111111110010010010011111;
assign LUT_2[39217] = 32'b11111111111111101111001010111000;
assign LUT_2[39218] = 32'b11111111111111111001001011011011;
assign LUT_2[39219] = 32'b11111111111111110110000011110100;
assign LUT_2[39220] = 32'b11111111111111101110110000000111;
assign LUT_2[39221] = 32'b11111111111111101011101000100000;
assign LUT_2[39222] = 32'b11111111111111110101101001000011;
assign LUT_2[39223] = 32'b11111111111111110010100001011100;
assign LUT_2[39224] = 32'b11111111111111101101000011111100;
assign LUT_2[39225] = 32'b11111111111111101001111100010101;
assign LUT_2[39226] = 32'b11111111111111110011111100111000;
assign LUT_2[39227] = 32'b11111111111111110000110101010001;
assign LUT_2[39228] = 32'b11111111111111101001100001100100;
assign LUT_2[39229] = 32'b11111111111111100110011001111101;
assign LUT_2[39230] = 32'b11111111111111110000011010100000;
assign LUT_2[39231] = 32'b11111111111111101101010010111001;
assign LUT_2[39232] = 32'b11111111111111101111011011001111;
assign LUT_2[39233] = 32'b11111111111111101100010011101000;
assign LUT_2[39234] = 32'b11111111111111110110010100001011;
assign LUT_2[39235] = 32'b11111111111111110011001100100100;
assign LUT_2[39236] = 32'b11111111111111101011111000110111;
assign LUT_2[39237] = 32'b11111111111111101000110001010000;
assign LUT_2[39238] = 32'b11111111111111110010110001110011;
assign LUT_2[39239] = 32'b11111111111111101111101010001100;
assign LUT_2[39240] = 32'b11111111111111101010001100101100;
assign LUT_2[39241] = 32'b11111111111111100111000101000101;
assign LUT_2[39242] = 32'b11111111111111110001000101101000;
assign LUT_2[39243] = 32'b11111111111111101101111110000001;
assign LUT_2[39244] = 32'b11111111111111100110101010010100;
assign LUT_2[39245] = 32'b11111111111111100011100010101101;
assign LUT_2[39246] = 32'b11111111111111101101100011010000;
assign LUT_2[39247] = 32'b11111111111111101010011011101001;
assign LUT_2[39248] = 32'b11111111111111101001111111011001;
assign LUT_2[39249] = 32'b11111111111111100110110111110010;
assign LUT_2[39250] = 32'b11111111111111110000111000010101;
assign LUT_2[39251] = 32'b11111111111111101101110000101110;
assign LUT_2[39252] = 32'b11111111111111100110011101000001;
assign LUT_2[39253] = 32'b11111111111111100011010101011010;
assign LUT_2[39254] = 32'b11111111111111101101010101111101;
assign LUT_2[39255] = 32'b11111111111111101010001110010110;
assign LUT_2[39256] = 32'b11111111111111100100110000110110;
assign LUT_2[39257] = 32'b11111111111111100001101001001111;
assign LUT_2[39258] = 32'b11111111111111101011101001110010;
assign LUT_2[39259] = 32'b11111111111111101000100010001011;
assign LUT_2[39260] = 32'b11111111111111100001001110011110;
assign LUT_2[39261] = 32'b11111111111111011110000110110111;
assign LUT_2[39262] = 32'b11111111111111101000000111011010;
assign LUT_2[39263] = 32'b11111111111111100100111111110011;
assign LUT_2[39264] = 32'b11111111111111101111110110111000;
assign LUT_2[39265] = 32'b11111111111111101100101111010001;
assign LUT_2[39266] = 32'b11111111111111110110101111110100;
assign LUT_2[39267] = 32'b11111111111111110011101000001101;
assign LUT_2[39268] = 32'b11111111111111101100010100100000;
assign LUT_2[39269] = 32'b11111111111111101001001100111001;
assign LUT_2[39270] = 32'b11111111111111110011001101011100;
assign LUT_2[39271] = 32'b11111111111111110000000101110101;
assign LUT_2[39272] = 32'b11111111111111101010101000010101;
assign LUT_2[39273] = 32'b11111111111111100111100000101110;
assign LUT_2[39274] = 32'b11111111111111110001100001010001;
assign LUT_2[39275] = 32'b11111111111111101110011001101010;
assign LUT_2[39276] = 32'b11111111111111100111000101111101;
assign LUT_2[39277] = 32'b11111111111111100011111110010110;
assign LUT_2[39278] = 32'b11111111111111101101111110111001;
assign LUT_2[39279] = 32'b11111111111111101010110111010010;
assign LUT_2[39280] = 32'b11111111111111101010011011000010;
assign LUT_2[39281] = 32'b11111111111111100111010011011011;
assign LUT_2[39282] = 32'b11111111111111110001010011111110;
assign LUT_2[39283] = 32'b11111111111111101110001100010111;
assign LUT_2[39284] = 32'b11111111111111100110111000101010;
assign LUT_2[39285] = 32'b11111111111111100011110001000011;
assign LUT_2[39286] = 32'b11111111111111101101110001100110;
assign LUT_2[39287] = 32'b11111111111111101010101001111111;
assign LUT_2[39288] = 32'b11111111111111100101001100011111;
assign LUT_2[39289] = 32'b11111111111111100010000100111000;
assign LUT_2[39290] = 32'b11111111111111101100000101011011;
assign LUT_2[39291] = 32'b11111111111111101000111101110100;
assign LUT_2[39292] = 32'b11111111111111100001101010000111;
assign LUT_2[39293] = 32'b11111111111111011110100010100000;
assign LUT_2[39294] = 32'b11111111111111101000100011000011;
assign LUT_2[39295] = 32'b11111111111111100101011011011100;
assign LUT_2[39296] = 32'b11111111111111111011100110111011;
assign LUT_2[39297] = 32'b11111111111111111000011111010100;
assign LUT_2[39298] = 32'b00000000000000000010011111110111;
assign LUT_2[39299] = 32'b11111111111111111111011000010000;
assign LUT_2[39300] = 32'b11111111111111111000000100100011;
assign LUT_2[39301] = 32'b11111111111111110100111100111100;
assign LUT_2[39302] = 32'b11111111111111111110111101011111;
assign LUT_2[39303] = 32'b11111111111111111011110101111000;
assign LUT_2[39304] = 32'b11111111111111110110011000011000;
assign LUT_2[39305] = 32'b11111111111111110011010000110001;
assign LUT_2[39306] = 32'b11111111111111111101010001010100;
assign LUT_2[39307] = 32'b11111111111111111010001001101101;
assign LUT_2[39308] = 32'b11111111111111110010110110000000;
assign LUT_2[39309] = 32'b11111111111111101111101110011001;
assign LUT_2[39310] = 32'b11111111111111111001101110111100;
assign LUT_2[39311] = 32'b11111111111111110110100111010101;
assign LUT_2[39312] = 32'b11111111111111110110001011000101;
assign LUT_2[39313] = 32'b11111111111111110011000011011110;
assign LUT_2[39314] = 32'b11111111111111111101000100000001;
assign LUT_2[39315] = 32'b11111111111111111001111100011010;
assign LUT_2[39316] = 32'b11111111111111110010101000101101;
assign LUT_2[39317] = 32'b11111111111111101111100001000110;
assign LUT_2[39318] = 32'b11111111111111111001100001101001;
assign LUT_2[39319] = 32'b11111111111111110110011010000010;
assign LUT_2[39320] = 32'b11111111111111110000111100100010;
assign LUT_2[39321] = 32'b11111111111111101101110100111011;
assign LUT_2[39322] = 32'b11111111111111110111110101011110;
assign LUT_2[39323] = 32'b11111111111111110100101101110111;
assign LUT_2[39324] = 32'b11111111111111101101011010001010;
assign LUT_2[39325] = 32'b11111111111111101010010010100011;
assign LUT_2[39326] = 32'b11111111111111110100010011000110;
assign LUT_2[39327] = 32'b11111111111111110001001011011111;
assign LUT_2[39328] = 32'b11111111111111111100000010100100;
assign LUT_2[39329] = 32'b11111111111111111000111010111101;
assign LUT_2[39330] = 32'b00000000000000000010111011100000;
assign LUT_2[39331] = 32'b11111111111111111111110011111001;
assign LUT_2[39332] = 32'b11111111111111111000100000001100;
assign LUT_2[39333] = 32'b11111111111111110101011000100101;
assign LUT_2[39334] = 32'b11111111111111111111011001001000;
assign LUT_2[39335] = 32'b11111111111111111100010001100001;
assign LUT_2[39336] = 32'b11111111111111110110110100000001;
assign LUT_2[39337] = 32'b11111111111111110011101100011010;
assign LUT_2[39338] = 32'b11111111111111111101101100111101;
assign LUT_2[39339] = 32'b11111111111111111010100101010110;
assign LUT_2[39340] = 32'b11111111111111110011010001101001;
assign LUT_2[39341] = 32'b11111111111111110000001010000010;
assign LUT_2[39342] = 32'b11111111111111111010001010100101;
assign LUT_2[39343] = 32'b11111111111111110111000010111110;
assign LUT_2[39344] = 32'b11111111111111110110100110101110;
assign LUT_2[39345] = 32'b11111111111111110011011111000111;
assign LUT_2[39346] = 32'b11111111111111111101011111101010;
assign LUT_2[39347] = 32'b11111111111111111010011000000011;
assign LUT_2[39348] = 32'b11111111111111110011000100010110;
assign LUT_2[39349] = 32'b11111111111111101111111100101111;
assign LUT_2[39350] = 32'b11111111111111111001111101010010;
assign LUT_2[39351] = 32'b11111111111111110110110101101011;
assign LUT_2[39352] = 32'b11111111111111110001011000001011;
assign LUT_2[39353] = 32'b11111111111111101110010000100100;
assign LUT_2[39354] = 32'b11111111111111111000010001000111;
assign LUT_2[39355] = 32'b11111111111111110101001001100000;
assign LUT_2[39356] = 32'b11111111111111101101110101110011;
assign LUT_2[39357] = 32'b11111111111111101010101110001100;
assign LUT_2[39358] = 32'b11111111111111110100101110101111;
assign LUT_2[39359] = 32'b11111111111111110001100111001000;
assign LUT_2[39360] = 32'b11111111111111110011101111011110;
assign LUT_2[39361] = 32'b11111111111111110000100111110111;
assign LUT_2[39362] = 32'b11111111111111111010101000011010;
assign LUT_2[39363] = 32'b11111111111111110111100000110011;
assign LUT_2[39364] = 32'b11111111111111110000001101000110;
assign LUT_2[39365] = 32'b11111111111111101101000101011111;
assign LUT_2[39366] = 32'b11111111111111110111000110000010;
assign LUT_2[39367] = 32'b11111111111111110011111110011011;
assign LUT_2[39368] = 32'b11111111111111101110100000111011;
assign LUT_2[39369] = 32'b11111111111111101011011001010100;
assign LUT_2[39370] = 32'b11111111111111110101011001110111;
assign LUT_2[39371] = 32'b11111111111111110010010010010000;
assign LUT_2[39372] = 32'b11111111111111101010111110100011;
assign LUT_2[39373] = 32'b11111111111111100111110110111100;
assign LUT_2[39374] = 32'b11111111111111110001110111011111;
assign LUT_2[39375] = 32'b11111111111111101110101111111000;
assign LUT_2[39376] = 32'b11111111111111101110010011101000;
assign LUT_2[39377] = 32'b11111111111111101011001100000001;
assign LUT_2[39378] = 32'b11111111111111110101001100100100;
assign LUT_2[39379] = 32'b11111111111111110010000100111101;
assign LUT_2[39380] = 32'b11111111111111101010110001010000;
assign LUT_2[39381] = 32'b11111111111111100111101001101001;
assign LUT_2[39382] = 32'b11111111111111110001101010001100;
assign LUT_2[39383] = 32'b11111111111111101110100010100101;
assign LUT_2[39384] = 32'b11111111111111101001000101000101;
assign LUT_2[39385] = 32'b11111111111111100101111101011110;
assign LUT_2[39386] = 32'b11111111111111101111111110000001;
assign LUT_2[39387] = 32'b11111111111111101100110110011010;
assign LUT_2[39388] = 32'b11111111111111100101100010101101;
assign LUT_2[39389] = 32'b11111111111111100010011011000110;
assign LUT_2[39390] = 32'b11111111111111101100011011101001;
assign LUT_2[39391] = 32'b11111111111111101001010100000010;
assign LUT_2[39392] = 32'b11111111111111110100001011000111;
assign LUT_2[39393] = 32'b11111111111111110001000011100000;
assign LUT_2[39394] = 32'b11111111111111111011000100000011;
assign LUT_2[39395] = 32'b11111111111111110111111100011100;
assign LUT_2[39396] = 32'b11111111111111110000101000101111;
assign LUT_2[39397] = 32'b11111111111111101101100001001000;
assign LUT_2[39398] = 32'b11111111111111110111100001101011;
assign LUT_2[39399] = 32'b11111111111111110100011010000100;
assign LUT_2[39400] = 32'b11111111111111101110111100100100;
assign LUT_2[39401] = 32'b11111111111111101011110100111101;
assign LUT_2[39402] = 32'b11111111111111110101110101100000;
assign LUT_2[39403] = 32'b11111111111111110010101101111001;
assign LUT_2[39404] = 32'b11111111111111101011011010001100;
assign LUT_2[39405] = 32'b11111111111111101000010010100101;
assign LUT_2[39406] = 32'b11111111111111110010010011001000;
assign LUT_2[39407] = 32'b11111111111111101111001011100001;
assign LUT_2[39408] = 32'b11111111111111101110101111010001;
assign LUT_2[39409] = 32'b11111111111111101011100111101010;
assign LUT_2[39410] = 32'b11111111111111110101101000001101;
assign LUT_2[39411] = 32'b11111111111111110010100000100110;
assign LUT_2[39412] = 32'b11111111111111101011001100111001;
assign LUT_2[39413] = 32'b11111111111111101000000101010010;
assign LUT_2[39414] = 32'b11111111111111110010000101110101;
assign LUT_2[39415] = 32'b11111111111111101110111110001110;
assign LUT_2[39416] = 32'b11111111111111101001100000101110;
assign LUT_2[39417] = 32'b11111111111111100110011001000111;
assign LUT_2[39418] = 32'b11111111111111110000011001101010;
assign LUT_2[39419] = 32'b11111111111111101101010010000011;
assign LUT_2[39420] = 32'b11111111111111100101111110010110;
assign LUT_2[39421] = 32'b11111111111111100010110110101111;
assign LUT_2[39422] = 32'b11111111111111101100110111010010;
assign LUT_2[39423] = 32'b11111111111111101001101111101011;
assign LUT_2[39424] = 32'b11111111111111111000000101111000;
assign LUT_2[39425] = 32'b11111111111111110100111110010001;
assign LUT_2[39426] = 32'b11111111111111111110111110110100;
assign LUT_2[39427] = 32'b11111111111111111011110111001101;
assign LUT_2[39428] = 32'b11111111111111110100100011100000;
assign LUT_2[39429] = 32'b11111111111111110001011011111001;
assign LUT_2[39430] = 32'b11111111111111111011011100011100;
assign LUT_2[39431] = 32'b11111111111111111000010100110101;
assign LUT_2[39432] = 32'b11111111111111110010110111010101;
assign LUT_2[39433] = 32'b11111111111111101111101111101110;
assign LUT_2[39434] = 32'b11111111111111111001110000010001;
assign LUT_2[39435] = 32'b11111111111111110110101000101010;
assign LUT_2[39436] = 32'b11111111111111101111010100111101;
assign LUT_2[39437] = 32'b11111111111111101100001101010110;
assign LUT_2[39438] = 32'b11111111111111110110001101111001;
assign LUT_2[39439] = 32'b11111111111111110011000110010010;
assign LUT_2[39440] = 32'b11111111111111110010101010000010;
assign LUT_2[39441] = 32'b11111111111111101111100010011011;
assign LUT_2[39442] = 32'b11111111111111111001100010111110;
assign LUT_2[39443] = 32'b11111111111111110110011011010111;
assign LUT_2[39444] = 32'b11111111111111101111000111101010;
assign LUT_2[39445] = 32'b11111111111111101100000000000011;
assign LUT_2[39446] = 32'b11111111111111110110000000100110;
assign LUT_2[39447] = 32'b11111111111111110010111000111111;
assign LUT_2[39448] = 32'b11111111111111101101011011011111;
assign LUT_2[39449] = 32'b11111111111111101010010011111000;
assign LUT_2[39450] = 32'b11111111111111110100010100011011;
assign LUT_2[39451] = 32'b11111111111111110001001100110100;
assign LUT_2[39452] = 32'b11111111111111101001111001000111;
assign LUT_2[39453] = 32'b11111111111111100110110001100000;
assign LUT_2[39454] = 32'b11111111111111110000110010000011;
assign LUT_2[39455] = 32'b11111111111111101101101010011100;
assign LUT_2[39456] = 32'b11111111111111111000100001100001;
assign LUT_2[39457] = 32'b11111111111111110101011001111010;
assign LUT_2[39458] = 32'b11111111111111111111011010011101;
assign LUT_2[39459] = 32'b11111111111111111100010010110110;
assign LUT_2[39460] = 32'b11111111111111110100111111001001;
assign LUT_2[39461] = 32'b11111111111111110001110111100010;
assign LUT_2[39462] = 32'b11111111111111111011111000000101;
assign LUT_2[39463] = 32'b11111111111111111000110000011110;
assign LUT_2[39464] = 32'b11111111111111110011010010111110;
assign LUT_2[39465] = 32'b11111111111111110000001011010111;
assign LUT_2[39466] = 32'b11111111111111111010001011111010;
assign LUT_2[39467] = 32'b11111111111111110111000100010011;
assign LUT_2[39468] = 32'b11111111111111101111110000100110;
assign LUT_2[39469] = 32'b11111111111111101100101000111111;
assign LUT_2[39470] = 32'b11111111111111110110101001100010;
assign LUT_2[39471] = 32'b11111111111111110011100001111011;
assign LUT_2[39472] = 32'b11111111111111110011000101101011;
assign LUT_2[39473] = 32'b11111111111111101111111110000100;
assign LUT_2[39474] = 32'b11111111111111111001111110100111;
assign LUT_2[39475] = 32'b11111111111111110110110111000000;
assign LUT_2[39476] = 32'b11111111111111101111100011010011;
assign LUT_2[39477] = 32'b11111111111111101100011011101100;
assign LUT_2[39478] = 32'b11111111111111110110011100001111;
assign LUT_2[39479] = 32'b11111111111111110011010100101000;
assign LUT_2[39480] = 32'b11111111111111101101110111001000;
assign LUT_2[39481] = 32'b11111111111111101010101111100001;
assign LUT_2[39482] = 32'b11111111111111110100110000000100;
assign LUT_2[39483] = 32'b11111111111111110001101000011101;
assign LUT_2[39484] = 32'b11111111111111101010010100110000;
assign LUT_2[39485] = 32'b11111111111111100111001101001001;
assign LUT_2[39486] = 32'b11111111111111110001001101101100;
assign LUT_2[39487] = 32'b11111111111111101110000110000101;
assign LUT_2[39488] = 32'b11111111111111110000001110011011;
assign LUT_2[39489] = 32'b11111111111111101101000110110100;
assign LUT_2[39490] = 32'b11111111111111110111000111010111;
assign LUT_2[39491] = 32'b11111111111111110011111111110000;
assign LUT_2[39492] = 32'b11111111111111101100101100000011;
assign LUT_2[39493] = 32'b11111111111111101001100100011100;
assign LUT_2[39494] = 32'b11111111111111110011100100111111;
assign LUT_2[39495] = 32'b11111111111111110000011101011000;
assign LUT_2[39496] = 32'b11111111111111101010111111111000;
assign LUT_2[39497] = 32'b11111111111111100111111000010001;
assign LUT_2[39498] = 32'b11111111111111110001111000110100;
assign LUT_2[39499] = 32'b11111111111111101110110001001101;
assign LUT_2[39500] = 32'b11111111111111100111011101100000;
assign LUT_2[39501] = 32'b11111111111111100100010101111001;
assign LUT_2[39502] = 32'b11111111111111101110010110011100;
assign LUT_2[39503] = 32'b11111111111111101011001110110101;
assign LUT_2[39504] = 32'b11111111111111101010110010100101;
assign LUT_2[39505] = 32'b11111111111111100111101010111110;
assign LUT_2[39506] = 32'b11111111111111110001101011100001;
assign LUT_2[39507] = 32'b11111111111111101110100011111010;
assign LUT_2[39508] = 32'b11111111111111100111010000001101;
assign LUT_2[39509] = 32'b11111111111111100100001000100110;
assign LUT_2[39510] = 32'b11111111111111101110001001001001;
assign LUT_2[39511] = 32'b11111111111111101011000001100010;
assign LUT_2[39512] = 32'b11111111111111100101100100000010;
assign LUT_2[39513] = 32'b11111111111111100010011100011011;
assign LUT_2[39514] = 32'b11111111111111101100011100111110;
assign LUT_2[39515] = 32'b11111111111111101001010101010111;
assign LUT_2[39516] = 32'b11111111111111100010000001101010;
assign LUT_2[39517] = 32'b11111111111111011110111010000011;
assign LUT_2[39518] = 32'b11111111111111101000111010100110;
assign LUT_2[39519] = 32'b11111111111111100101110010111111;
assign LUT_2[39520] = 32'b11111111111111110000101010000100;
assign LUT_2[39521] = 32'b11111111111111101101100010011101;
assign LUT_2[39522] = 32'b11111111111111110111100011000000;
assign LUT_2[39523] = 32'b11111111111111110100011011011001;
assign LUT_2[39524] = 32'b11111111111111101101000111101100;
assign LUT_2[39525] = 32'b11111111111111101010000000000101;
assign LUT_2[39526] = 32'b11111111111111110100000000101000;
assign LUT_2[39527] = 32'b11111111111111110000111001000001;
assign LUT_2[39528] = 32'b11111111111111101011011011100001;
assign LUT_2[39529] = 32'b11111111111111101000010011111010;
assign LUT_2[39530] = 32'b11111111111111110010010100011101;
assign LUT_2[39531] = 32'b11111111111111101111001100110110;
assign LUT_2[39532] = 32'b11111111111111100111111001001001;
assign LUT_2[39533] = 32'b11111111111111100100110001100010;
assign LUT_2[39534] = 32'b11111111111111101110110010000101;
assign LUT_2[39535] = 32'b11111111111111101011101010011110;
assign LUT_2[39536] = 32'b11111111111111101011001110001110;
assign LUT_2[39537] = 32'b11111111111111101000000110100111;
assign LUT_2[39538] = 32'b11111111111111110010000111001010;
assign LUT_2[39539] = 32'b11111111111111101110111111100011;
assign LUT_2[39540] = 32'b11111111111111100111101011110110;
assign LUT_2[39541] = 32'b11111111111111100100100100001111;
assign LUT_2[39542] = 32'b11111111111111101110100100110010;
assign LUT_2[39543] = 32'b11111111111111101011011101001011;
assign LUT_2[39544] = 32'b11111111111111100101111111101011;
assign LUT_2[39545] = 32'b11111111111111100010111000000100;
assign LUT_2[39546] = 32'b11111111111111101100111000100111;
assign LUT_2[39547] = 32'b11111111111111101001110001000000;
assign LUT_2[39548] = 32'b11111111111111100010011101010011;
assign LUT_2[39549] = 32'b11111111111111011111010101101100;
assign LUT_2[39550] = 32'b11111111111111101001010110001111;
assign LUT_2[39551] = 32'b11111111111111100110001110101000;
assign LUT_2[39552] = 32'b11111111111111111100011010000111;
assign LUT_2[39553] = 32'b11111111111111111001010010100000;
assign LUT_2[39554] = 32'b00000000000000000011010011000011;
assign LUT_2[39555] = 32'b00000000000000000000001011011100;
assign LUT_2[39556] = 32'b11111111111111111000110111101111;
assign LUT_2[39557] = 32'b11111111111111110101110000001000;
assign LUT_2[39558] = 32'b11111111111111111111110000101011;
assign LUT_2[39559] = 32'b11111111111111111100101001000100;
assign LUT_2[39560] = 32'b11111111111111110111001011100100;
assign LUT_2[39561] = 32'b11111111111111110100000011111101;
assign LUT_2[39562] = 32'b11111111111111111110000100100000;
assign LUT_2[39563] = 32'b11111111111111111010111100111001;
assign LUT_2[39564] = 32'b11111111111111110011101001001100;
assign LUT_2[39565] = 32'b11111111111111110000100001100101;
assign LUT_2[39566] = 32'b11111111111111111010100010001000;
assign LUT_2[39567] = 32'b11111111111111110111011010100001;
assign LUT_2[39568] = 32'b11111111111111110110111110010001;
assign LUT_2[39569] = 32'b11111111111111110011110110101010;
assign LUT_2[39570] = 32'b11111111111111111101110111001101;
assign LUT_2[39571] = 32'b11111111111111111010101111100110;
assign LUT_2[39572] = 32'b11111111111111110011011011111001;
assign LUT_2[39573] = 32'b11111111111111110000010100010010;
assign LUT_2[39574] = 32'b11111111111111111010010100110101;
assign LUT_2[39575] = 32'b11111111111111110111001101001110;
assign LUT_2[39576] = 32'b11111111111111110001101111101110;
assign LUT_2[39577] = 32'b11111111111111101110101000000111;
assign LUT_2[39578] = 32'b11111111111111111000101000101010;
assign LUT_2[39579] = 32'b11111111111111110101100001000011;
assign LUT_2[39580] = 32'b11111111111111101110001101010110;
assign LUT_2[39581] = 32'b11111111111111101011000101101111;
assign LUT_2[39582] = 32'b11111111111111110101000110010010;
assign LUT_2[39583] = 32'b11111111111111110001111110101011;
assign LUT_2[39584] = 32'b11111111111111111100110101110000;
assign LUT_2[39585] = 32'b11111111111111111001101110001001;
assign LUT_2[39586] = 32'b00000000000000000011101110101100;
assign LUT_2[39587] = 32'b00000000000000000000100111000101;
assign LUT_2[39588] = 32'b11111111111111111001010011011000;
assign LUT_2[39589] = 32'b11111111111111110110001011110001;
assign LUT_2[39590] = 32'b00000000000000000000001100010100;
assign LUT_2[39591] = 32'b11111111111111111101000100101101;
assign LUT_2[39592] = 32'b11111111111111110111100111001101;
assign LUT_2[39593] = 32'b11111111111111110100011111100110;
assign LUT_2[39594] = 32'b11111111111111111110100000001001;
assign LUT_2[39595] = 32'b11111111111111111011011000100010;
assign LUT_2[39596] = 32'b11111111111111110100000100110101;
assign LUT_2[39597] = 32'b11111111111111110000111101001110;
assign LUT_2[39598] = 32'b11111111111111111010111101110001;
assign LUT_2[39599] = 32'b11111111111111110111110110001010;
assign LUT_2[39600] = 32'b11111111111111110111011001111010;
assign LUT_2[39601] = 32'b11111111111111110100010010010011;
assign LUT_2[39602] = 32'b11111111111111111110010010110110;
assign LUT_2[39603] = 32'b11111111111111111011001011001111;
assign LUT_2[39604] = 32'b11111111111111110011110111100010;
assign LUT_2[39605] = 32'b11111111111111110000101111111011;
assign LUT_2[39606] = 32'b11111111111111111010110000011110;
assign LUT_2[39607] = 32'b11111111111111110111101000110111;
assign LUT_2[39608] = 32'b11111111111111110010001011010111;
assign LUT_2[39609] = 32'b11111111111111101111000011110000;
assign LUT_2[39610] = 32'b11111111111111111001000100010011;
assign LUT_2[39611] = 32'b11111111111111110101111100101100;
assign LUT_2[39612] = 32'b11111111111111101110101000111111;
assign LUT_2[39613] = 32'b11111111111111101011100001011000;
assign LUT_2[39614] = 32'b11111111111111110101100001111011;
assign LUT_2[39615] = 32'b11111111111111110010011010010100;
assign LUT_2[39616] = 32'b11111111111111110100100010101010;
assign LUT_2[39617] = 32'b11111111111111110001011011000011;
assign LUT_2[39618] = 32'b11111111111111111011011011100110;
assign LUT_2[39619] = 32'b11111111111111111000010011111111;
assign LUT_2[39620] = 32'b11111111111111110001000000010010;
assign LUT_2[39621] = 32'b11111111111111101101111000101011;
assign LUT_2[39622] = 32'b11111111111111110111111001001110;
assign LUT_2[39623] = 32'b11111111111111110100110001100111;
assign LUT_2[39624] = 32'b11111111111111101111010100000111;
assign LUT_2[39625] = 32'b11111111111111101100001100100000;
assign LUT_2[39626] = 32'b11111111111111110110001101000011;
assign LUT_2[39627] = 32'b11111111111111110011000101011100;
assign LUT_2[39628] = 32'b11111111111111101011110001101111;
assign LUT_2[39629] = 32'b11111111111111101000101010001000;
assign LUT_2[39630] = 32'b11111111111111110010101010101011;
assign LUT_2[39631] = 32'b11111111111111101111100011000100;
assign LUT_2[39632] = 32'b11111111111111101111000110110100;
assign LUT_2[39633] = 32'b11111111111111101011111111001101;
assign LUT_2[39634] = 32'b11111111111111110101111111110000;
assign LUT_2[39635] = 32'b11111111111111110010111000001001;
assign LUT_2[39636] = 32'b11111111111111101011100100011100;
assign LUT_2[39637] = 32'b11111111111111101000011100110101;
assign LUT_2[39638] = 32'b11111111111111110010011101011000;
assign LUT_2[39639] = 32'b11111111111111101111010101110001;
assign LUT_2[39640] = 32'b11111111111111101001111000010001;
assign LUT_2[39641] = 32'b11111111111111100110110000101010;
assign LUT_2[39642] = 32'b11111111111111110000110001001101;
assign LUT_2[39643] = 32'b11111111111111101101101001100110;
assign LUT_2[39644] = 32'b11111111111111100110010101111001;
assign LUT_2[39645] = 32'b11111111111111100011001110010010;
assign LUT_2[39646] = 32'b11111111111111101101001110110101;
assign LUT_2[39647] = 32'b11111111111111101010000111001110;
assign LUT_2[39648] = 32'b11111111111111110100111110010011;
assign LUT_2[39649] = 32'b11111111111111110001110110101100;
assign LUT_2[39650] = 32'b11111111111111111011110111001111;
assign LUT_2[39651] = 32'b11111111111111111000101111101000;
assign LUT_2[39652] = 32'b11111111111111110001011011111011;
assign LUT_2[39653] = 32'b11111111111111101110010100010100;
assign LUT_2[39654] = 32'b11111111111111111000010100110111;
assign LUT_2[39655] = 32'b11111111111111110101001101010000;
assign LUT_2[39656] = 32'b11111111111111101111101111110000;
assign LUT_2[39657] = 32'b11111111111111101100101000001001;
assign LUT_2[39658] = 32'b11111111111111110110101000101100;
assign LUT_2[39659] = 32'b11111111111111110011100001000101;
assign LUT_2[39660] = 32'b11111111111111101100001101011000;
assign LUT_2[39661] = 32'b11111111111111101001000101110001;
assign LUT_2[39662] = 32'b11111111111111110011000110010100;
assign LUT_2[39663] = 32'b11111111111111101111111110101101;
assign LUT_2[39664] = 32'b11111111111111101111100010011101;
assign LUT_2[39665] = 32'b11111111111111101100011010110110;
assign LUT_2[39666] = 32'b11111111111111110110011011011001;
assign LUT_2[39667] = 32'b11111111111111110011010011110010;
assign LUT_2[39668] = 32'b11111111111111101100000000000101;
assign LUT_2[39669] = 32'b11111111111111101000111000011110;
assign LUT_2[39670] = 32'b11111111111111110010111001000001;
assign LUT_2[39671] = 32'b11111111111111101111110001011010;
assign LUT_2[39672] = 32'b11111111111111101010010011111010;
assign LUT_2[39673] = 32'b11111111111111100111001100010011;
assign LUT_2[39674] = 32'b11111111111111110001001100110110;
assign LUT_2[39675] = 32'b11111111111111101110000101001111;
assign LUT_2[39676] = 32'b11111111111111100110110001100010;
assign LUT_2[39677] = 32'b11111111111111100011101001111011;
assign LUT_2[39678] = 32'b11111111111111101101101010011110;
assign LUT_2[39679] = 32'b11111111111111101010100010110111;
assign LUT_2[39680] = 32'b11111111111111111100000100011110;
assign LUT_2[39681] = 32'b11111111111111111000111100110111;
assign LUT_2[39682] = 32'b00000000000000000010111101011010;
assign LUT_2[39683] = 32'b11111111111111111111110101110011;
assign LUT_2[39684] = 32'b11111111111111111000100010000110;
assign LUT_2[39685] = 32'b11111111111111110101011010011111;
assign LUT_2[39686] = 32'b11111111111111111111011011000010;
assign LUT_2[39687] = 32'b11111111111111111100010011011011;
assign LUT_2[39688] = 32'b11111111111111110110110101111011;
assign LUT_2[39689] = 32'b11111111111111110011101110010100;
assign LUT_2[39690] = 32'b11111111111111111101101110110111;
assign LUT_2[39691] = 32'b11111111111111111010100111010000;
assign LUT_2[39692] = 32'b11111111111111110011010011100011;
assign LUT_2[39693] = 32'b11111111111111110000001011111100;
assign LUT_2[39694] = 32'b11111111111111111010001100011111;
assign LUT_2[39695] = 32'b11111111111111110111000100111000;
assign LUT_2[39696] = 32'b11111111111111110110101000101000;
assign LUT_2[39697] = 32'b11111111111111110011100001000001;
assign LUT_2[39698] = 32'b11111111111111111101100001100100;
assign LUT_2[39699] = 32'b11111111111111111010011001111101;
assign LUT_2[39700] = 32'b11111111111111110011000110010000;
assign LUT_2[39701] = 32'b11111111111111101111111110101001;
assign LUT_2[39702] = 32'b11111111111111111001111111001100;
assign LUT_2[39703] = 32'b11111111111111110110110111100101;
assign LUT_2[39704] = 32'b11111111111111110001011010000101;
assign LUT_2[39705] = 32'b11111111111111101110010010011110;
assign LUT_2[39706] = 32'b11111111111111111000010011000001;
assign LUT_2[39707] = 32'b11111111111111110101001011011010;
assign LUT_2[39708] = 32'b11111111111111101101110111101101;
assign LUT_2[39709] = 32'b11111111111111101010110000000110;
assign LUT_2[39710] = 32'b11111111111111110100110000101001;
assign LUT_2[39711] = 32'b11111111111111110001101001000010;
assign LUT_2[39712] = 32'b11111111111111111100100000000111;
assign LUT_2[39713] = 32'b11111111111111111001011000100000;
assign LUT_2[39714] = 32'b00000000000000000011011001000011;
assign LUT_2[39715] = 32'b00000000000000000000010001011100;
assign LUT_2[39716] = 32'b11111111111111111000111101101111;
assign LUT_2[39717] = 32'b11111111111111110101110110001000;
assign LUT_2[39718] = 32'b11111111111111111111110110101011;
assign LUT_2[39719] = 32'b11111111111111111100101111000100;
assign LUT_2[39720] = 32'b11111111111111110111010001100100;
assign LUT_2[39721] = 32'b11111111111111110100001001111101;
assign LUT_2[39722] = 32'b11111111111111111110001010100000;
assign LUT_2[39723] = 32'b11111111111111111011000010111001;
assign LUT_2[39724] = 32'b11111111111111110011101111001100;
assign LUT_2[39725] = 32'b11111111111111110000100111100101;
assign LUT_2[39726] = 32'b11111111111111111010101000001000;
assign LUT_2[39727] = 32'b11111111111111110111100000100001;
assign LUT_2[39728] = 32'b11111111111111110111000100010001;
assign LUT_2[39729] = 32'b11111111111111110011111100101010;
assign LUT_2[39730] = 32'b11111111111111111101111101001101;
assign LUT_2[39731] = 32'b11111111111111111010110101100110;
assign LUT_2[39732] = 32'b11111111111111110011100001111001;
assign LUT_2[39733] = 32'b11111111111111110000011010010010;
assign LUT_2[39734] = 32'b11111111111111111010011010110101;
assign LUT_2[39735] = 32'b11111111111111110111010011001110;
assign LUT_2[39736] = 32'b11111111111111110001110101101110;
assign LUT_2[39737] = 32'b11111111111111101110101110000111;
assign LUT_2[39738] = 32'b11111111111111111000101110101010;
assign LUT_2[39739] = 32'b11111111111111110101100111000011;
assign LUT_2[39740] = 32'b11111111111111101110010011010110;
assign LUT_2[39741] = 32'b11111111111111101011001011101111;
assign LUT_2[39742] = 32'b11111111111111110101001100010010;
assign LUT_2[39743] = 32'b11111111111111110010000100101011;
assign LUT_2[39744] = 32'b11111111111111110100001101000001;
assign LUT_2[39745] = 32'b11111111111111110001000101011010;
assign LUT_2[39746] = 32'b11111111111111111011000101111101;
assign LUT_2[39747] = 32'b11111111111111110111111110010110;
assign LUT_2[39748] = 32'b11111111111111110000101010101001;
assign LUT_2[39749] = 32'b11111111111111101101100011000010;
assign LUT_2[39750] = 32'b11111111111111110111100011100101;
assign LUT_2[39751] = 32'b11111111111111110100011011111110;
assign LUT_2[39752] = 32'b11111111111111101110111110011110;
assign LUT_2[39753] = 32'b11111111111111101011110110110111;
assign LUT_2[39754] = 32'b11111111111111110101110111011010;
assign LUT_2[39755] = 32'b11111111111111110010101111110011;
assign LUT_2[39756] = 32'b11111111111111101011011100000110;
assign LUT_2[39757] = 32'b11111111111111101000010100011111;
assign LUT_2[39758] = 32'b11111111111111110010010101000010;
assign LUT_2[39759] = 32'b11111111111111101111001101011011;
assign LUT_2[39760] = 32'b11111111111111101110110001001011;
assign LUT_2[39761] = 32'b11111111111111101011101001100100;
assign LUT_2[39762] = 32'b11111111111111110101101010000111;
assign LUT_2[39763] = 32'b11111111111111110010100010100000;
assign LUT_2[39764] = 32'b11111111111111101011001110110011;
assign LUT_2[39765] = 32'b11111111111111101000000111001100;
assign LUT_2[39766] = 32'b11111111111111110010000111101111;
assign LUT_2[39767] = 32'b11111111111111101111000000001000;
assign LUT_2[39768] = 32'b11111111111111101001100010101000;
assign LUT_2[39769] = 32'b11111111111111100110011011000001;
assign LUT_2[39770] = 32'b11111111111111110000011011100100;
assign LUT_2[39771] = 32'b11111111111111101101010011111101;
assign LUT_2[39772] = 32'b11111111111111100110000000010000;
assign LUT_2[39773] = 32'b11111111111111100010111000101001;
assign LUT_2[39774] = 32'b11111111111111101100111001001100;
assign LUT_2[39775] = 32'b11111111111111101001110001100101;
assign LUT_2[39776] = 32'b11111111111111110100101000101010;
assign LUT_2[39777] = 32'b11111111111111110001100001000011;
assign LUT_2[39778] = 32'b11111111111111111011100001100110;
assign LUT_2[39779] = 32'b11111111111111111000011001111111;
assign LUT_2[39780] = 32'b11111111111111110001000110010010;
assign LUT_2[39781] = 32'b11111111111111101101111110101011;
assign LUT_2[39782] = 32'b11111111111111110111111111001110;
assign LUT_2[39783] = 32'b11111111111111110100110111100111;
assign LUT_2[39784] = 32'b11111111111111101111011010000111;
assign LUT_2[39785] = 32'b11111111111111101100010010100000;
assign LUT_2[39786] = 32'b11111111111111110110010011000011;
assign LUT_2[39787] = 32'b11111111111111110011001011011100;
assign LUT_2[39788] = 32'b11111111111111101011110111101111;
assign LUT_2[39789] = 32'b11111111111111101000110000001000;
assign LUT_2[39790] = 32'b11111111111111110010110000101011;
assign LUT_2[39791] = 32'b11111111111111101111101001000100;
assign LUT_2[39792] = 32'b11111111111111101111001100110100;
assign LUT_2[39793] = 32'b11111111111111101100000101001101;
assign LUT_2[39794] = 32'b11111111111111110110000101110000;
assign LUT_2[39795] = 32'b11111111111111110010111110001001;
assign LUT_2[39796] = 32'b11111111111111101011101010011100;
assign LUT_2[39797] = 32'b11111111111111101000100010110101;
assign LUT_2[39798] = 32'b11111111111111110010100011011000;
assign LUT_2[39799] = 32'b11111111111111101111011011110001;
assign LUT_2[39800] = 32'b11111111111111101001111110010001;
assign LUT_2[39801] = 32'b11111111111111100110110110101010;
assign LUT_2[39802] = 32'b11111111111111110000110111001101;
assign LUT_2[39803] = 32'b11111111111111101101101111100110;
assign LUT_2[39804] = 32'b11111111111111100110011011111001;
assign LUT_2[39805] = 32'b11111111111111100011010100010010;
assign LUT_2[39806] = 32'b11111111111111101101010100110101;
assign LUT_2[39807] = 32'b11111111111111101010001101001110;
assign LUT_2[39808] = 32'b00000000000000000000011000101101;
assign LUT_2[39809] = 32'b11111111111111111101010001000110;
assign LUT_2[39810] = 32'b00000000000000000111010001101001;
assign LUT_2[39811] = 32'b00000000000000000100001010000010;
assign LUT_2[39812] = 32'b11111111111111111100110110010101;
assign LUT_2[39813] = 32'b11111111111111111001101110101110;
assign LUT_2[39814] = 32'b00000000000000000011101111010001;
assign LUT_2[39815] = 32'b00000000000000000000100111101010;
assign LUT_2[39816] = 32'b11111111111111111011001010001010;
assign LUT_2[39817] = 32'b11111111111111111000000010100011;
assign LUT_2[39818] = 32'b00000000000000000010000011000110;
assign LUT_2[39819] = 32'b11111111111111111110111011011111;
assign LUT_2[39820] = 32'b11111111111111110111100111110010;
assign LUT_2[39821] = 32'b11111111111111110100100000001011;
assign LUT_2[39822] = 32'b11111111111111111110100000101110;
assign LUT_2[39823] = 32'b11111111111111111011011001000111;
assign LUT_2[39824] = 32'b11111111111111111010111100110111;
assign LUT_2[39825] = 32'b11111111111111110111110101010000;
assign LUT_2[39826] = 32'b00000000000000000001110101110011;
assign LUT_2[39827] = 32'b11111111111111111110101110001100;
assign LUT_2[39828] = 32'b11111111111111110111011010011111;
assign LUT_2[39829] = 32'b11111111111111110100010010111000;
assign LUT_2[39830] = 32'b11111111111111111110010011011011;
assign LUT_2[39831] = 32'b11111111111111111011001011110100;
assign LUT_2[39832] = 32'b11111111111111110101101110010100;
assign LUT_2[39833] = 32'b11111111111111110010100110101101;
assign LUT_2[39834] = 32'b11111111111111111100100111010000;
assign LUT_2[39835] = 32'b11111111111111111001011111101001;
assign LUT_2[39836] = 32'b11111111111111110010001011111100;
assign LUT_2[39837] = 32'b11111111111111101111000100010101;
assign LUT_2[39838] = 32'b11111111111111111001000100111000;
assign LUT_2[39839] = 32'b11111111111111110101111101010001;
assign LUT_2[39840] = 32'b00000000000000000000110100010110;
assign LUT_2[39841] = 32'b11111111111111111101101100101111;
assign LUT_2[39842] = 32'b00000000000000000111101101010010;
assign LUT_2[39843] = 32'b00000000000000000100100101101011;
assign LUT_2[39844] = 32'b11111111111111111101010001111110;
assign LUT_2[39845] = 32'b11111111111111111010001010010111;
assign LUT_2[39846] = 32'b00000000000000000100001010111010;
assign LUT_2[39847] = 32'b00000000000000000001000011010011;
assign LUT_2[39848] = 32'b11111111111111111011100101110011;
assign LUT_2[39849] = 32'b11111111111111111000011110001100;
assign LUT_2[39850] = 32'b00000000000000000010011110101111;
assign LUT_2[39851] = 32'b11111111111111111111010111001000;
assign LUT_2[39852] = 32'b11111111111111111000000011011011;
assign LUT_2[39853] = 32'b11111111111111110100111011110100;
assign LUT_2[39854] = 32'b11111111111111111110111100010111;
assign LUT_2[39855] = 32'b11111111111111111011110100110000;
assign LUT_2[39856] = 32'b11111111111111111011011000100000;
assign LUT_2[39857] = 32'b11111111111111111000010000111001;
assign LUT_2[39858] = 32'b00000000000000000010010001011100;
assign LUT_2[39859] = 32'b11111111111111111111001001110101;
assign LUT_2[39860] = 32'b11111111111111110111110110001000;
assign LUT_2[39861] = 32'b11111111111111110100101110100001;
assign LUT_2[39862] = 32'b11111111111111111110101111000100;
assign LUT_2[39863] = 32'b11111111111111111011100111011101;
assign LUT_2[39864] = 32'b11111111111111110110001001111101;
assign LUT_2[39865] = 32'b11111111111111110011000010010110;
assign LUT_2[39866] = 32'b11111111111111111101000010111001;
assign LUT_2[39867] = 32'b11111111111111111001111011010010;
assign LUT_2[39868] = 32'b11111111111111110010100111100101;
assign LUT_2[39869] = 32'b11111111111111101111011111111110;
assign LUT_2[39870] = 32'b11111111111111111001100000100001;
assign LUT_2[39871] = 32'b11111111111111110110011000111010;
assign LUT_2[39872] = 32'b11111111111111111000100001010000;
assign LUT_2[39873] = 32'b11111111111111110101011001101001;
assign LUT_2[39874] = 32'b11111111111111111111011010001100;
assign LUT_2[39875] = 32'b11111111111111111100010010100101;
assign LUT_2[39876] = 32'b11111111111111110100111110111000;
assign LUT_2[39877] = 32'b11111111111111110001110111010001;
assign LUT_2[39878] = 32'b11111111111111111011110111110100;
assign LUT_2[39879] = 32'b11111111111111111000110000001101;
assign LUT_2[39880] = 32'b11111111111111110011010010101101;
assign LUT_2[39881] = 32'b11111111111111110000001011000110;
assign LUT_2[39882] = 32'b11111111111111111010001011101001;
assign LUT_2[39883] = 32'b11111111111111110111000100000010;
assign LUT_2[39884] = 32'b11111111111111101111110000010101;
assign LUT_2[39885] = 32'b11111111111111101100101000101110;
assign LUT_2[39886] = 32'b11111111111111110110101001010001;
assign LUT_2[39887] = 32'b11111111111111110011100001101010;
assign LUT_2[39888] = 32'b11111111111111110011000101011010;
assign LUT_2[39889] = 32'b11111111111111101111111101110011;
assign LUT_2[39890] = 32'b11111111111111111001111110010110;
assign LUT_2[39891] = 32'b11111111111111110110110110101111;
assign LUT_2[39892] = 32'b11111111111111101111100011000010;
assign LUT_2[39893] = 32'b11111111111111101100011011011011;
assign LUT_2[39894] = 32'b11111111111111110110011011111110;
assign LUT_2[39895] = 32'b11111111111111110011010100010111;
assign LUT_2[39896] = 32'b11111111111111101101110110110111;
assign LUT_2[39897] = 32'b11111111111111101010101111010000;
assign LUT_2[39898] = 32'b11111111111111110100101111110011;
assign LUT_2[39899] = 32'b11111111111111110001101000001100;
assign LUT_2[39900] = 32'b11111111111111101010010100011111;
assign LUT_2[39901] = 32'b11111111111111100111001100111000;
assign LUT_2[39902] = 32'b11111111111111110001001101011011;
assign LUT_2[39903] = 32'b11111111111111101110000101110100;
assign LUT_2[39904] = 32'b11111111111111111000111100111001;
assign LUT_2[39905] = 32'b11111111111111110101110101010010;
assign LUT_2[39906] = 32'b11111111111111111111110101110101;
assign LUT_2[39907] = 32'b11111111111111111100101110001110;
assign LUT_2[39908] = 32'b11111111111111110101011010100001;
assign LUT_2[39909] = 32'b11111111111111110010010010111010;
assign LUT_2[39910] = 32'b11111111111111111100010011011101;
assign LUT_2[39911] = 32'b11111111111111111001001011110110;
assign LUT_2[39912] = 32'b11111111111111110011101110010110;
assign LUT_2[39913] = 32'b11111111111111110000100110101111;
assign LUT_2[39914] = 32'b11111111111111111010100111010010;
assign LUT_2[39915] = 32'b11111111111111110111011111101011;
assign LUT_2[39916] = 32'b11111111111111110000001011111110;
assign LUT_2[39917] = 32'b11111111111111101101000100010111;
assign LUT_2[39918] = 32'b11111111111111110111000100111010;
assign LUT_2[39919] = 32'b11111111111111110011111101010011;
assign LUT_2[39920] = 32'b11111111111111110011100001000011;
assign LUT_2[39921] = 32'b11111111111111110000011001011100;
assign LUT_2[39922] = 32'b11111111111111111010011001111111;
assign LUT_2[39923] = 32'b11111111111111110111010010011000;
assign LUT_2[39924] = 32'b11111111111111101111111110101011;
assign LUT_2[39925] = 32'b11111111111111101100110111000100;
assign LUT_2[39926] = 32'b11111111111111110110110111100111;
assign LUT_2[39927] = 32'b11111111111111110011110000000000;
assign LUT_2[39928] = 32'b11111111111111101110010010100000;
assign LUT_2[39929] = 32'b11111111111111101011001010111001;
assign LUT_2[39930] = 32'b11111111111111110101001011011100;
assign LUT_2[39931] = 32'b11111111111111110010000011110101;
assign LUT_2[39932] = 32'b11111111111111101010110000001000;
assign LUT_2[39933] = 32'b11111111111111100111101000100001;
assign LUT_2[39934] = 32'b11111111111111110001101001000100;
assign LUT_2[39935] = 32'b11111111111111101110100001011101;
assign LUT_2[39936] = 32'b11111111111111111010000000001011;
assign LUT_2[39937] = 32'b11111111111111110110111000100100;
assign LUT_2[39938] = 32'b00000000000000000000111001000111;
assign LUT_2[39939] = 32'b11111111111111111101110001100000;
assign LUT_2[39940] = 32'b11111111111111110110011101110011;
assign LUT_2[39941] = 32'b11111111111111110011010110001100;
assign LUT_2[39942] = 32'b11111111111111111101010110101111;
assign LUT_2[39943] = 32'b11111111111111111010001111001000;
assign LUT_2[39944] = 32'b11111111111111110100110001101000;
assign LUT_2[39945] = 32'b11111111111111110001101010000001;
assign LUT_2[39946] = 32'b11111111111111111011101010100100;
assign LUT_2[39947] = 32'b11111111111111111000100010111101;
assign LUT_2[39948] = 32'b11111111111111110001001111010000;
assign LUT_2[39949] = 32'b11111111111111101110000111101001;
assign LUT_2[39950] = 32'b11111111111111111000001000001100;
assign LUT_2[39951] = 32'b11111111111111110101000000100101;
assign LUT_2[39952] = 32'b11111111111111110100100100010101;
assign LUT_2[39953] = 32'b11111111111111110001011100101110;
assign LUT_2[39954] = 32'b11111111111111111011011101010001;
assign LUT_2[39955] = 32'b11111111111111111000010101101010;
assign LUT_2[39956] = 32'b11111111111111110001000001111101;
assign LUT_2[39957] = 32'b11111111111111101101111010010110;
assign LUT_2[39958] = 32'b11111111111111110111111010111001;
assign LUT_2[39959] = 32'b11111111111111110100110011010010;
assign LUT_2[39960] = 32'b11111111111111101111010101110010;
assign LUT_2[39961] = 32'b11111111111111101100001110001011;
assign LUT_2[39962] = 32'b11111111111111110110001110101110;
assign LUT_2[39963] = 32'b11111111111111110011000111000111;
assign LUT_2[39964] = 32'b11111111111111101011110011011010;
assign LUT_2[39965] = 32'b11111111111111101000101011110011;
assign LUT_2[39966] = 32'b11111111111111110010101100010110;
assign LUT_2[39967] = 32'b11111111111111101111100100101111;
assign LUT_2[39968] = 32'b11111111111111111010011011110100;
assign LUT_2[39969] = 32'b11111111111111110111010100001101;
assign LUT_2[39970] = 32'b00000000000000000001010100110000;
assign LUT_2[39971] = 32'b11111111111111111110001101001001;
assign LUT_2[39972] = 32'b11111111111111110110111001011100;
assign LUT_2[39973] = 32'b11111111111111110011110001110101;
assign LUT_2[39974] = 32'b11111111111111111101110010011000;
assign LUT_2[39975] = 32'b11111111111111111010101010110001;
assign LUT_2[39976] = 32'b11111111111111110101001101010001;
assign LUT_2[39977] = 32'b11111111111111110010000101101010;
assign LUT_2[39978] = 32'b11111111111111111100000110001101;
assign LUT_2[39979] = 32'b11111111111111111000111110100110;
assign LUT_2[39980] = 32'b11111111111111110001101010111001;
assign LUT_2[39981] = 32'b11111111111111101110100011010010;
assign LUT_2[39982] = 32'b11111111111111111000100011110101;
assign LUT_2[39983] = 32'b11111111111111110101011100001110;
assign LUT_2[39984] = 32'b11111111111111110100111111111110;
assign LUT_2[39985] = 32'b11111111111111110001111000010111;
assign LUT_2[39986] = 32'b11111111111111111011111000111010;
assign LUT_2[39987] = 32'b11111111111111111000110001010011;
assign LUT_2[39988] = 32'b11111111111111110001011101100110;
assign LUT_2[39989] = 32'b11111111111111101110010101111111;
assign LUT_2[39990] = 32'b11111111111111111000010110100010;
assign LUT_2[39991] = 32'b11111111111111110101001110111011;
assign LUT_2[39992] = 32'b11111111111111101111110001011011;
assign LUT_2[39993] = 32'b11111111111111101100101001110100;
assign LUT_2[39994] = 32'b11111111111111110110101010010111;
assign LUT_2[39995] = 32'b11111111111111110011100010110000;
assign LUT_2[39996] = 32'b11111111111111101100001111000011;
assign LUT_2[39997] = 32'b11111111111111101001000111011100;
assign LUT_2[39998] = 32'b11111111111111110011000111111111;
assign LUT_2[39999] = 32'b11111111111111110000000000011000;
assign LUT_2[40000] = 32'b11111111111111110010001000101110;
assign LUT_2[40001] = 32'b11111111111111101111000001000111;
assign LUT_2[40002] = 32'b11111111111111111001000001101010;
assign LUT_2[40003] = 32'b11111111111111110101111010000011;
assign LUT_2[40004] = 32'b11111111111111101110100110010110;
assign LUT_2[40005] = 32'b11111111111111101011011110101111;
assign LUT_2[40006] = 32'b11111111111111110101011111010010;
assign LUT_2[40007] = 32'b11111111111111110010010111101011;
assign LUT_2[40008] = 32'b11111111111111101100111010001011;
assign LUT_2[40009] = 32'b11111111111111101001110010100100;
assign LUT_2[40010] = 32'b11111111111111110011110011000111;
assign LUT_2[40011] = 32'b11111111111111110000101011100000;
assign LUT_2[40012] = 32'b11111111111111101001010111110011;
assign LUT_2[40013] = 32'b11111111111111100110010000001100;
assign LUT_2[40014] = 32'b11111111111111110000010000101111;
assign LUT_2[40015] = 32'b11111111111111101101001001001000;
assign LUT_2[40016] = 32'b11111111111111101100101100111000;
assign LUT_2[40017] = 32'b11111111111111101001100101010001;
assign LUT_2[40018] = 32'b11111111111111110011100101110100;
assign LUT_2[40019] = 32'b11111111111111110000011110001101;
assign LUT_2[40020] = 32'b11111111111111101001001010100000;
assign LUT_2[40021] = 32'b11111111111111100110000010111001;
assign LUT_2[40022] = 32'b11111111111111110000000011011100;
assign LUT_2[40023] = 32'b11111111111111101100111011110101;
assign LUT_2[40024] = 32'b11111111111111100111011110010101;
assign LUT_2[40025] = 32'b11111111111111100100010110101110;
assign LUT_2[40026] = 32'b11111111111111101110010111010001;
assign LUT_2[40027] = 32'b11111111111111101011001111101010;
assign LUT_2[40028] = 32'b11111111111111100011111011111101;
assign LUT_2[40029] = 32'b11111111111111100000110100010110;
assign LUT_2[40030] = 32'b11111111111111101010110100111001;
assign LUT_2[40031] = 32'b11111111111111100111101101010010;
assign LUT_2[40032] = 32'b11111111111111110010100100010111;
assign LUT_2[40033] = 32'b11111111111111101111011100110000;
assign LUT_2[40034] = 32'b11111111111111111001011101010011;
assign LUT_2[40035] = 32'b11111111111111110110010101101100;
assign LUT_2[40036] = 32'b11111111111111101111000001111111;
assign LUT_2[40037] = 32'b11111111111111101011111010011000;
assign LUT_2[40038] = 32'b11111111111111110101111010111011;
assign LUT_2[40039] = 32'b11111111111111110010110011010100;
assign LUT_2[40040] = 32'b11111111111111101101010101110100;
assign LUT_2[40041] = 32'b11111111111111101010001110001101;
assign LUT_2[40042] = 32'b11111111111111110100001110110000;
assign LUT_2[40043] = 32'b11111111111111110001000111001001;
assign LUT_2[40044] = 32'b11111111111111101001110011011100;
assign LUT_2[40045] = 32'b11111111111111100110101011110101;
assign LUT_2[40046] = 32'b11111111111111110000101100011000;
assign LUT_2[40047] = 32'b11111111111111101101100100110001;
assign LUT_2[40048] = 32'b11111111111111101101001000100001;
assign LUT_2[40049] = 32'b11111111111111101010000000111010;
assign LUT_2[40050] = 32'b11111111111111110100000001011101;
assign LUT_2[40051] = 32'b11111111111111110000111001110110;
assign LUT_2[40052] = 32'b11111111111111101001100110001001;
assign LUT_2[40053] = 32'b11111111111111100110011110100010;
assign LUT_2[40054] = 32'b11111111111111110000011111000101;
assign LUT_2[40055] = 32'b11111111111111101101010111011110;
assign LUT_2[40056] = 32'b11111111111111100111111001111110;
assign LUT_2[40057] = 32'b11111111111111100100110010010111;
assign LUT_2[40058] = 32'b11111111111111101110110010111010;
assign LUT_2[40059] = 32'b11111111111111101011101011010011;
assign LUT_2[40060] = 32'b11111111111111100100010111100110;
assign LUT_2[40061] = 32'b11111111111111100001001111111111;
assign LUT_2[40062] = 32'b11111111111111101011010000100010;
assign LUT_2[40063] = 32'b11111111111111101000001000111011;
assign LUT_2[40064] = 32'b11111111111111111110010100011010;
assign LUT_2[40065] = 32'b11111111111111111011001100110011;
assign LUT_2[40066] = 32'b00000000000000000101001101010110;
assign LUT_2[40067] = 32'b00000000000000000010000101101111;
assign LUT_2[40068] = 32'b11111111111111111010110010000010;
assign LUT_2[40069] = 32'b11111111111111110111101010011011;
assign LUT_2[40070] = 32'b00000000000000000001101010111110;
assign LUT_2[40071] = 32'b11111111111111111110100011010111;
assign LUT_2[40072] = 32'b11111111111111111001000101110111;
assign LUT_2[40073] = 32'b11111111111111110101111110010000;
assign LUT_2[40074] = 32'b11111111111111111111111110110011;
assign LUT_2[40075] = 32'b11111111111111111100110111001100;
assign LUT_2[40076] = 32'b11111111111111110101100011011111;
assign LUT_2[40077] = 32'b11111111111111110010011011111000;
assign LUT_2[40078] = 32'b11111111111111111100011100011011;
assign LUT_2[40079] = 32'b11111111111111111001010100110100;
assign LUT_2[40080] = 32'b11111111111111111000111000100100;
assign LUT_2[40081] = 32'b11111111111111110101110000111101;
assign LUT_2[40082] = 32'b11111111111111111111110001100000;
assign LUT_2[40083] = 32'b11111111111111111100101001111001;
assign LUT_2[40084] = 32'b11111111111111110101010110001100;
assign LUT_2[40085] = 32'b11111111111111110010001110100101;
assign LUT_2[40086] = 32'b11111111111111111100001111001000;
assign LUT_2[40087] = 32'b11111111111111111001000111100001;
assign LUT_2[40088] = 32'b11111111111111110011101010000001;
assign LUT_2[40089] = 32'b11111111111111110000100010011010;
assign LUT_2[40090] = 32'b11111111111111111010100010111101;
assign LUT_2[40091] = 32'b11111111111111110111011011010110;
assign LUT_2[40092] = 32'b11111111111111110000000111101001;
assign LUT_2[40093] = 32'b11111111111111101101000000000010;
assign LUT_2[40094] = 32'b11111111111111110111000000100101;
assign LUT_2[40095] = 32'b11111111111111110011111000111110;
assign LUT_2[40096] = 32'b11111111111111111110110000000011;
assign LUT_2[40097] = 32'b11111111111111111011101000011100;
assign LUT_2[40098] = 32'b00000000000000000101101000111111;
assign LUT_2[40099] = 32'b00000000000000000010100001011000;
assign LUT_2[40100] = 32'b11111111111111111011001101101011;
assign LUT_2[40101] = 32'b11111111111111111000000110000100;
assign LUT_2[40102] = 32'b00000000000000000010000110100111;
assign LUT_2[40103] = 32'b11111111111111111110111111000000;
assign LUT_2[40104] = 32'b11111111111111111001100001100000;
assign LUT_2[40105] = 32'b11111111111111110110011001111001;
assign LUT_2[40106] = 32'b00000000000000000000011010011100;
assign LUT_2[40107] = 32'b11111111111111111101010010110101;
assign LUT_2[40108] = 32'b11111111111111110101111111001000;
assign LUT_2[40109] = 32'b11111111111111110010110111100001;
assign LUT_2[40110] = 32'b11111111111111111100111000000100;
assign LUT_2[40111] = 32'b11111111111111111001110000011101;
assign LUT_2[40112] = 32'b11111111111111111001010100001101;
assign LUT_2[40113] = 32'b11111111111111110110001100100110;
assign LUT_2[40114] = 32'b00000000000000000000001101001001;
assign LUT_2[40115] = 32'b11111111111111111101000101100010;
assign LUT_2[40116] = 32'b11111111111111110101110001110101;
assign LUT_2[40117] = 32'b11111111111111110010101010001110;
assign LUT_2[40118] = 32'b11111111111111111100101010110001;
assign LUT_2[40119] = 32'b11111111111111111001100011001010;
assign LUT_2[40120] = 32'b11111111111111110100000101101010;
assign LUT_2[40121] = 32'b11111111111111110000111110000011;
assign LUT_2[40122] = 32'b11111111111111111010111110100110;
assign LUT_2[40123] = 32'b11111111111111110111110110111111;
assign LUT_2[40124] = 32'b11111111111111110000100011010010;
assign LUT_2[40125] = 32'b11111111111111101101011011101011;
assign LUT_2[40126] = 32'b11111111111111110111011100001110;
assign LUT_2[40127] = 32'b11111111111111110100010100100111;
assign LUT_2[40128] = 32'b11111111111111110110011100111101;
assign LUT_2[40129] = 32'b11111111111111110011010101010110;
assign LUT_2[40130] = 32'b11111111111111111101010101111001;
assign LUT_2[40131] = 32'b11111111111111111010001110010010;
assign LUT_2[40132] = 32'b11111111111111110010111010100101;
assign LUT_2[40133] = 32'b11111111111111101111110010111110;
assign LUT_2[40134] = 32'b11111111111111111001110011100001;
assign LUT_2[40135] = 32'b11111111111111110110101011111010;
assign LUT_2[40136] = 32'b11111111111111110001001110011010;
assign LUT_2[40137] = 32'b11111111111111101110000110110011;
assign LUT_2[40138] = 32'b11111111111111111000000111010110;
assign LUT_2[40139] = 32'b11111111111111110100111111101111;
assign LUT_2[40140] = 32'b11111111111111101101101100000010;
assign LUT_2[40141] = 32'b11111111111111101010100100011011;
assign LUT_2[40142] = 32'b11111111111111110100100100111110;
assign LUT_2[40143] = 32'b11111111111111110001011101010111;
assign LUT_2[40144] = 32'b11111111111111110001000001000111;
assign LUT_2[40145] = 32'b11111111111111101101111001100000;
assign LUT_2[40146] = 32'b11111111111111110111111010000011;
assign LUT_2[40147] = 32'b11111111111111110100110010011100;
assign LUT_2[40148] = 32'b11111111111111101101011110101111;
assign LUT_2[40149] = 32'b11111111111111101010010111001000;
assign LUT_2[40150] = 32'b11111111111111110100010111101011;
assign LUT_2[40151] = 32'b11111111111111110001010000000100;
assign LUT_2[40152] = 32'b11111111111111101011110010100100;
assign LUT_2[40153] = 32'b11111111111111101000101010111101;
assign LUT_2[40154] = 32'b11111111111111110010101011100000;
assign LUT_2[40155] = 32'b11111111111111101111100011111001;
assign LUT_2[40156] = 32'b11111111111111101000010000001100;
assign LUT_2[40157] = 32'b11111111111111100101001000100101;
assign LUT_2[40158] = 32'b11111111111111101111001001001000;
assign LUT_2[40159] = 32'b11111111111111101100000001100001;
assign LUT_2[40160] = 32'b11111111111111110110111000100110;
assign LUT_2[40161] = 32'b11111111111111110011110000111111;
assign LUT_2[40162] = 32'b11111111111111111101110001100010;
assign LUT_2[40163] = 32'b11111111111111111010101001111011;
assign LUT_2[40164] = 32'b11111111111111110011010110001110;
assign LUT_2[40165] = 32'b11111111111111110000001110100111;
assign LUT_2[40166] = 32'b11111111111111111010001111001010;
assign LUT_2[40167] = 32'b11111111111111110111000111100011;
assign LUT_2[40168] = 32'b11111111111111110001101010000011;
assign LUT_2[40169] = 32'b11111111111111101110100010011100;
assign LUT_2[40170] = 32'b11111111111111111000100010111111;
assign LUT_2[40171] = 32'b11111111111111110101011011011000;
assign LUT_2[40172] = 32'b11111111111111101110000111101011;
assign LUT_2[40173] = 32'b11111111111111101011000000000100;
assign LUT_2[40174] = 32'b11111111111111110101000000100111;
assign LUT_2[40175] = 32'b11111111111111110001111001000000;
assign LUT_2[40176] = 32'b11111111111111110001011100110000;
assign LUT_2[40177] = 32'b11111111111111101110010101001001;
assign LUT_2[40178] = 32'b11111111111111111000010101101100;
assign LUT_2[40179] = 32'b11111111111111110101001110000101;
assign LUT_2[40180] = 32'b11111111111111101101111010011000;
assign LUT_2[40181] = 32'b11111111111111101010110010110001;
assign LUT_2[40182] = 32'b11111111111111110100110011010100;
assign LUT_2[40183] = 32'b11111111111111110001101011101101;
assign LUT_2[40184] = 32'b11111111111111101100001110001101;
assign LUT_2[40185] = 32'b11111111111111101001000110100110;
assign LUT_2[40186] = 32'b11111111111111110011000111001001;
assign LUT_2[40187] = 32'b11111111111111101111111111100010;
assign LUT_2[40188] = 32'b11111111111111101000101011110101;
assign LUT_2[40189] = 32'b11111111111111100101100100001110;
assign LUT_2[40190] = 32'b11111111111111101111100100110001;
assign LUT_2[40191] = 32'b11111111111111101100011101001010;
assign LUT_2[40192] = 32'b11111111111111111101111110110001;
assign LUT_2[40193] = 32'b11111111111111111010110111001010;
assign LUT_2[40194] = 32'b00000000000000000100110111101101;
assign LUT_2[40195] = 32'b00000000000000000001110000000110;
assign LUT_2[40196] = 32'b11111111111111111010011100011001;
assign LUT_2[40197] = 32'b11111111111111110111010100110010;
assign LUT_2[40198] = 32'b00000000000000000001010101010101;
assign LUT_2[40199] = 32'b11111111111111111110001101101110;
assign LUT_2[40200] = 32'b11111111111111111000110000001110;
assign LUT_2[40201] = 32'b11111111111111110101101000100111;
assign LUT_2[40202] = 32'b11111111111111111111101001001010;
assign LUT_2[40203] = 32'b11111111111111111100100001100011;
assign LUT_2[40204] = 32'b11111111111111110101001101110110;
assign LUT_2[40205] = 32'b11111111111111110010000110001111;
assign LUT_2[40206] = 32'b11111111111111111100000110110010;
assign LUT_2[40207] = 32'b11111111111111111000111111001011;
assign LUT_2[40208] = 32'b11111111111111111000100010111011;
assign LUT_2[40209] = 32'b11111111111111110101011011010100;
assign LUT_2[40210] = 32'b11111111111111111111011011110111;
assign LUT_2[40211] = 32'b11111111111111111100010100010000;
assign LUT_2[40212] = 32'b11111111111111110101000000100011;
assign LUT_2[40213] = 32'b11111111111111110001111000111100;
assign LUT_2[40214] = 32'b11111111111111111011111001011111;
assign LUT_2[40215] = 32'b11111111111111111000110001111000;
assign LUT_2[40216] = 32'b11111111111111110011010100011000;
assign LUT_2[40217] = 32'b11111111111111110000001100110001;
assign LUT_2[40218] = 32'b11111111111111111010001101010100;
assign LUT_2[40219] = 32'b11111111111111110111000101101101;
assign LUT_2[40220] = 32'b11111111111111101111110010000000;
assign LUT_2[40221] = 32'b11111111111111101100101010011001;
assign LUT_2[40222] = 32'b11111111111111110110101010111100;
assign LUT_2[40223] = 32'b11111111111111110011100011010101;
assign LUT_2[40224] = 32'b11111111111111111110011010011010;
assign LUT_2[40225] = 32'b11111111111111111011010010110011;
assign LUT_2[40226] = 32'b00000000000000000101010011010110;
assign LUT_2[40227] = 32'b00000000000000000010001011101111;
assign LUT_2[40228] = 32'b11111111111111111010111000000010;
assign LUT_2[40229] = 32'b11111111111111110111110000011011;
assign LUT_2[40230] = 32'b00000000000000000001110000111110;
assign LUT_2[40231] = 32'b11111111111111111110101001010111;
assign LUT_2[40232] = 32'b11111111111111111001001011110111;
assign LUT_2[40233] = 32'b11111111111111110110000100010000;
assign LUT_2[40234] = 32'b00000000000000000000000100110011;
assign LUT_2[40235] = 32'b11111111111111111100111101001100;
assign LUT_2[40236] = 32'b11111111111111110101101001011111;
assign LUT_2[40237] = 32'b11111111111111110010100001111000;
assign LUT_2[40238] = 32'b11111111111111111100100010011011;
assign LUT_2[40239] = 32'b11111111111111111001011010110100;
assign LUT_2[40240] = 32'b11111111111111111000111110100100;
assign LUT_2[40241] = 32'b11111111111111110101110110111101;
assign LUT_2[40242] = 32'b11111111111111111111110111100000;
assign LUT_2[40243] = 32'b11111111111111111100101111111001;
assign LUT_2[40244] = 32'b11111111111111110101011100001100;
assign LUT_2[40245] = 32'b11111111111111110010010100100101;
assign LUT_2[40246] = 32'b11111111111111111100010101001000;
assign LUT_2[40247] = 32'b11111111111111111001001101100001;
assign LUT_2[40248] = 32'b11111111111111110011110000000001;
assign LUT_2[40249] = 32'b11111111111111110000101000011010;
assign LUT_2[40250] = 32'b11111111111111111010101000111101;
assign LUT_2[40251] = 32'b11111111111111110111100001010110;
assign LUT_2[40252] = 32'b11111111111111110000001101101001;
assign LUT_2[40253] = 32'b11111111111111101101000110000010;
assign LUT_2[40254] = 32'b11111111111111110111000110100101;
assign LUT_2[40255] = 32'b11111111111111110011111110111110;
assign LUT_2[40256] = 32'b11111111111111110110000111010100;
assign LUT_2[40257] = 32'b11111111111111110010111111101101;
assign LUT_2[40258] = 32'b11111111111111111101000000010000;
assign LUT_2[40259] = 32'b11111111111111111001111000101001;
assign LUT_2[40260] = 32'b11111111111111110010100100111100;
assign LUT_2[40261] = 32'b11111111111111101111011101010101;
assign LUT_2[40262] = 32'b11111111111111111001011101111000;
assign LUT_2[40263] = 32'b11111111111111110110010110010001;
assign LUT_2[40264] = 32'b11111111111111110000111000110001;
assign LUT_2[40265] = 32'b11111111111111101101110001001010;
assign LUT_2[40266] = 32'b11111111111111110111110001101101;
assign LUT_2[40267] = 32'b11111111111111110100101010000110;
assign LUT_2[40268] = 32'b11111111111111101101010110011001;
assign LUT_2[40269] = 32'b11111111111111101010001110110010;
assign LUT_2[40270] = 32'b11111111111111110100001111010101;
assign LUT_2[40271] = 32'b11111111111111110001000111101110;
assign LUT_2[40272] = 32'b11111111111111110000101011011110;
assign LUT_2[40273] = 32'b11111111111111101101100011110111;
assign LUT_2[40274] = 32'b11111111111111110111100100011010;
assign LUT_2[40275] = 32'b11111111111111110100011100110011;
assign LUT_2[40276] = 32'b11111111111111101101001001000110;
assign LUT_2[40277] = 32'b11111111111111101010000001011111;
assign LUT_2[40278] = 32'b11111111111111110100000010000010;
assign LUT_2[40279] = 32'b11111111111111110000111010011011;
assign LUT_2[40280] = 32'b11111111111111101011011100111011;
assign LUT_2[40281] = 32'b11111111111111101000010101010100;
assign LUT_2[40282] = 32'b11111111111111110010010101110111;
assign LUT_2[40283] = 32'b11111111111111101111001110010000;
assign LUT_2[40284] = 32'b11111111111111100111111010100011;
assign LUT_2[40285] = 32'b11111111111111100100110010111100;
assign LUT_2[40286] = 32'b11111111111111101110110011011111;
assign LUT_2[40287] = 32'b11111111111111101011101011111000;
assign LUT_2[40288] = 32'b11111111111111110110100010111101;
assign LUT_2[40289] = 32'b11111111111111110011011011010110;
assign LUT_2[40290] = 32'b11111111111111111101011011111001;
assign LUT_2[40291] = 32'b11111111111111111010010100010010;
assign LUT_2[40292] = 32'b11111111111111110011000000100101;
assign LUT_2[40293] = 32'b11111111111111101111111000111110;
assign LUT_2[40294] = 32'b11111111111111111001111001100001;
assign LUT_2[40295] = 32'b11111111111111110110110001111010;
assign LUT_2[40296] = 32'b11111111111111110001010100011010;
assign LUT_2[40297] = 32'b11111111111111101110001100110011;
assign LUT_2[40298] = 32'b11111111111111111000001101010110;
assign LUT_2[40299] = 32'b11111111111111110101000101101111;
assign LUT_2[40300] = 32'b11111111111111101101110010000010;
assign LUT_2[40301] = 32'b11111111111111101010101010011011;
assign LUT_2[40302] = 32'b11111111111111110100101010111110;
assign LUT_2[40303] = 32'b11111111111111110001100011010111;
assign LUT_2[40304] = 32'b11111111111111110001000111000111;
assign LUT_2[40305] = 32'b11111111111111101101111111100000;
assign LUT_2[40306] = 32'b11111111111111111000000000000011;
assign LUT_2[40307] = 32'b11111111111111110100111000011100;
assign LUT_2[40308] = 32'b11111111111111101101100100101111;
assign LUT_2[40309] = 32'b11111111111111101010011101001000;
assign LUT_2[40310] = 32'b11111111111111110100011101101011;
assign LUT_2[40311] = 32'b11111111111111110001010110000100;
assign LUT_2[40312] = 32'b11111111111111101011111000100100;
assign LUT_2[40313] = 32'b11111111111111101000110000111101;
assign LUT_2[40314] = 32'b11111111111111110010110001100000;
assign LUT_2[40315] = 32'b11111111111111101111101001111001;
assign LUT_2[40316] = 32'b11111111111111101000010110001100;
assign LUT_2[40317] = 32'b11111111111111100101001110100101;
assign LUT_2[40318] = 32'b11111111111111101111001111001000;
assign LUT_2[40319] = 32'b11111111111111101100000111100001;
assign LUT_2[40320] = 32'b00000000000000000010010011000000;
assign LUT_2[40321] = 32'b11111111111111111111001011011001;
assign LUT_2[40322] = 32'b00000000000000001001001011111100;
assign LUT_2[40323] = 32'b00000000000000000110000100010101;
assign LUT_2[40324] = 32'b11111111111111111110110000101000;
assign LUT_2[40325] = 32'b11111111111111111011101001000001;
assign LUT_2[40326] = 32'b00000000000000000101101001100100;
assign LUT_2[40327] = 32'b00000000000000000010100001111101;
assign LUT_2[40328] = 32'b11111111111111111101000100011101;
assign LUT_2[40329] = 32'b11111111111111111001111100110110;
assign LUT_2[40330] = 32'b00000000000000000011111101011001;
assign LUT_2[40331] = 32'b00000000000000000000110101110010;
assign LUT_2[40332] = 32'b11111111111111111001100010000101;
assign LUT_2[40333] = 32'b11111111111111110110011010011110;
assign LUT_2[40334] = 32'b00000000000000000000011011000001;
assign LUT_2[40335] = 32'b11111111111111111101010011011010;
assign LUT_2[40336] = 32'b11111111111111111100110111001010;
assign LUT_2[40337] = 32'b11111111111111111001101111100011;
assign LUT_2[40338] = 32'b00000000000000000011110000000110;
assign LUT_2[40339] = 32'b00000000000000000000101000011111;
assign LUT_2[40340] = 32'b11111111111111111001010100110010;
assign LUT_2[40341] = 32'b11111111111111110110001101001011;
assign LUT_2[40342] = 32'b00000000000000000000001101101110;
assign LUT_2[40343] = 32'b11111111111111111101000110000111;
assign LUT_2[40344] = 32'b11111111111111110111101000100111;
assign LUT_2[40345] = 32'b11111111111111110100100001000000;
assign LUT_2[40346] = 32'b11111111111111111110100001100011;
assign LUT_2[40347] = 32'b11111111111111111011011001111100;
assign LUT_2[40348] = 32'b11111111111111110100000110001111;
assign LUT_2[40349] = 32'b11111111111111110000111110101000;
assign LUT_2[40350] = 32'b11111111111111111010111111001011;
assign LUT_2[40351] = 32'b11111111111111110111110111100100;
assign LUT_2[40352] = 32'b00000000000000000010101110101001;
assign LUT_2[40353] = 32'b11111111111111111111100111000010;
assign LUT_2[40354] = 32'b00000000000000001001100111100101;
assign LUT_2[40355] = 32'b00000000000000000110011111111110;
assign LUT_2[40356] = 32'b11111111111111111111001100010001;
assign LUT_2[40357] = 32'b11111111111111111100000100101010;
assign LUT_2[40358] = 32'b00000000000000000110000101001101;
assign LUT_2[40359] = 32'b00000000000000000010111101100110;
assign LUT_2[40360] = 32'b11111111111111111101100000000110;
assign LUT_2[40361] = 32'b11111111111111111010011000011111;
assign LUT_2[40362] = 32'b00000000000000000100011001000010;
assign LUT_2[40363] = 32'b00000000000000000001010001011011;
assign LUT_2[40364] = 32'b11111111111111111001111101101110;
assign LUT_2[40365] = 32'b11111111111111110110110110000111;
assign LUT_2[40366] = 32'b00000000000000000000110110101010;
assign LUT_2[40367] = 32'b11111111111111111101101111000011;
assign LUT_2[40368] = 32'b11111111111111111101010010110011;
assign LUT_2[40369] = 32'b11111111111111111010001011001100;
assign LUT_2[40370] = 32'b00000000000000000100001011101111;
assign LUT_2[40371] = 32'b00000000000000000001000100001000;
assign LUT_2[40372] = 32'b11111111111111111001110000011011;
assign LUT_2[40373] = 32'b11111111111111110110101000110100;
assign LUT_2[40374] = 32'b00000000000000000000101001010111;
assign LUT_2[40375] = 32'b11111111111111111101100001110000;
assign LUT_2[40376] = 32'b11111111111111111000000100010000;
assign LUT_2[40377] = 32'b11111111111111110100111100101001;
assign LUT_2[40378] = 32'b11111111111111111110111101001100;
assign LUT_2[40379] = 32'b11111111111111111011110101100101;
assign LUT_2[40380] = 32'b11111111111111110100100001111000;
assign LUT_2[40381] = 32'b11111111111111110001011010010001;
assign LUT_2[40382] = 32'b11111111111111111011011010110100;
assign LUT_2[40383] = 32'b11111111111111111000010011001101;
assign LUT_2[40384] = 32'b11111111111111111010011011100011;
assign LUT_2[40385] = 32'b11111111111111110111010011111100;
assign LUT_2[40386] = 32'b00000000000000000001010100011111;
assign LUT_2[40387] = 32'b11111111111111111110001100111000;
assign LUT_2[40388] = 32'b11111111111111110110111001001011;
assign LUT_2[40389] = 32'b11111111111111110011110001100100;
assign LUT_2[40390] = 32'b11111111111111111101110010000111;
assign LUT_2[40391] = 32'b11111111111111111010101010100000;
assign LUT_2[40392] = 32'b11111111111111110101001101000000;
assign LUT_2[40393] = 32'b11111111111111110010000101011001;
assign LUT_2[40394] = 32'b11111111111111111100000101111100;
assign LUT_2[40395] = 32'b11111111111111111000111110010101;
assign LUT_2[40396] = 32'b11111111111111110001101010101000;
assign LUT_2[40397] = 32'b11111111111111101110100011000001;
assign LUT_2[40398] = 32'b11111111111111111000100011100100;
assign LUT_2[40399] = 32'b11111111111111110101011011111101;
assign LUT_2[40400] = 32'b11111111111111110100111111101101;
assign LUT_2[40401] = 32'b11111111111111110001111000000110;
assign LUT_2[40402] = 32'b11111111111111111011111000101001;
assign LUT_2[40403] = 32'b11111111111111111000110001000010;
assign LUT_2[40404] = 32'b11111111111111110001011101010101;
assign LUT_2[40405] = 32'b11111111111111101110010101101110;
assign LUT_2[40406] = 32'b11111111111111111000010110010001;
assign LUT_2[40407] = 32'b11111111111111110101001110101010;
assign LUT_2[40408] = 32'b11111111111111101111110001001010;
assign LUT_2[40409] = 32'b11111111111111101100101001100011;
assign LUT_2[40410] = 32'b11111111111111110110101010000110;
assign LUT_2[40411] = 32'b11111111111111110011100010011111;
assign LUT_2[40412] = 32'b11111111111111101100001110110010;
assign LUT_2[40413] = 32'b11111111111111101001000111001011;
assign LUT_2[40414] = 32'b11111111111111110011000111101110;
assign LUT_2[40415] = 32'b11111111111111110000000000000111;
assign LUT_2[40416] = 32'b11111111111111111010110111001100;
assign LUT_2[40417] = 32'b11111111111111110111101111100101;
assign LUT_2[40418] = 32'b00000000000000000001110000001000;
assign LUT_2[40419] = 32'b11111111111111111110101000100001;
assign LUT_2[40420] = 32'b11111111111111110111010100110100;
assign LUT_2[40421] = 32'b11111111111111110100001101001101;
assign LUT_2[40422] = 32'b11111111111111111110001101110000;
assign LUT_2[40423] = 32'b11111111111111111011000110001001;
assign LUT_2[40424] = 32'b11111111111111110101101000101001;
assign LUT_2[40425] = 32'b11111111111111110010100001000010;
assign LUT_2[40426] = 32'b11111111111111111100100001100101;
assign LUT_2[40427] = 32'b11111111111111111001011001111110;
assign LUT_2[40428] = 32'b11111111111111110010000110010001;
assign LUT_2[40429] = 32'b11111111111111101110111110101010;
assign LUT_2[40430] = 32'b11111111111111111000111111001101;
assign LUT_2[40431] = 32'b11111111111111110101110111100110;
assign LUT_2[40432] = 32'b11111111111111110101011011010110;
assign LUT_2[40433] = 32'b11111111111111110010010011101111;
assign LUT_2[40434] = 32'b11111111111111111100010100010010;
assign LUT_2[40435] = 32'b11111111111111111001001100101011;
assign LUT_2[40436] = 32'b11111111111111110001111000111110;
assign LUT_2[40437] = 32'b11111111111111101110110001010111;
assign LUT_2[40438] = 32'b11111111111111111000110001111010;
assign LUT_2[40439] = 32'b11111111111111110101101010010011;
assign LUT_2[40440] = 32'b11111111111111110000001100110011;
assign LUT_2[40441] = 32'b11111111111111101101000101001100;
assign LUT_2[40442] = 32'b11111111111111110111000101101111;
assign LUT_2[40443] = 32'b11111111111111110011111110001000;
assign LUT_2[40444] = 32'b11111111111111101100101010011011;
assign LUT_2[40445] = 32'b11111111111111101001100010110100;
assign LUT_2[40446] = 32'b11111111111111110011100011010111;
assign LUT_2[40447] = 32'b11111111111111110000011011110000;
assign LUT_2[40448] = 32'b11111111111111111110110001111101;
assign LUT_2[40449] = 32'b11111111111111111011101010010110;
assign LUT_2[40450] = 32'b00000000000000000101101010111001;
assign LUT_2[40451] = 32'b00000000000000000010100011010010;
assign LUT_2[40452] = 32'b11111111111111111011001111100101;
assign LUT_2[40453] = 32'b11111111111111111000000111111110;
assign LUT_2[40454] = 32'b00000000000000000010001000100001;
assign LUT_2[40455] = 32'b11111111111111111111000000111010;
assign LUT_2[40456] = 32'b11111111111111111001100011011010;
assign LUT_2[40457] = 32'b11111111111111110110011011110011;
assign LUT_2[40458] = 32'b00000000000000000000011100010110;
assign LUT_2[40459] = 32'b11111111111111111101010100101111;
assign LUT_2[40460] = 32'b11111111111111110110000001000010;
assign LUT_2[40461] = 32'b11111111111111110010111001011011;
assign LUT_2[40462] = 32'b11111111111111111100111001111110;
assign LUT_2[40463] = 32'b11111111111111111001110010010111;
assign LUT_2[40464] = 32'b11111111111111111001010110000111;
assign LUT_2[40465] = 32'b11111111111111110110001110100000;
assign LUT_2[40466] = 32'b00000000000000000000001111000011;
assign LUT_2[40467] = 32'b11111111111111111101000111011100;
assign LUT_2[40468] = 32'b11111111111111110101110011101111;
assign LUT_2[40469] = 32'b11111111111111110010101100001000;
assign LUT_2[40470] = 32'b11111111111111111100101100101011;
assign LUT_2[40471] = 32'b11111111111111111001100101000100;
assign LUT_2[40472] = 32'b11111111111111110100000111100100;
assign LUT_2[40473] = 32'b11111111111111110000111111111101;
assign LUT_2[40474] = 32'b11111111111111111011000000100000;
assign LUT_2[40475] = 32'b11111111111111110111111000111001;
assign LUT_2[40476] = 32'b11111111111111110000100101001100;
assign LUT_2[40477] = 32'b11111111111111101101011101100101;
assign LUT_2[40478] = 32'b11111111111111110111011110001000;
assign LUT_2[40479] = 32'b11111111111111110100010110100001;
assign LUT_2[40480] = 32'b11111111111111111111001101100110;
assign LUT_2[40481] = 32'b11111111111111111100000101111111;
assign LUT_2[40482] = 32'b00000000000000000110000110100010;
assign LUT_2[40483] = 32'b00000000000000000010111110111011;
assign LUT_2[40484] = 32'b11111111111111111011101011001110;
assign LUT_2[40485] = 32'b11111111111111111000100011100111;
assign LUT_2[40486] = 32'b00000000000000000010100100001010;
assign LUT_2[40487] = 32'b11111111111111111111011100100011;
assign LUT_2[40488] = 32'b11111111111111111001111111000011;
assign LUT_2[40489] = 32'b11111111111111110110110111011100;
assign LUT_2[40490] = 32'b00000000000000000000110111111111;
assign LUT_2[40491] = 32'b11111111111111111101110000011000;
assign LUT_2[40492] = 32'b11111111111111110110011100101011;
assign LUT_2[40493] = 32'b11111111111111110011010101000100;
assign LUT_2[40494] = 32'b11111111111111111101010101100111;
assign LUT_2[40495] = 32'b11111111111111111010001110000000;
assign LUT_2[40496] = 32'b11111111111111111001110001110000;
assign LUT_2[40497] = 32'b11111111111111110110101010001001;
assign LUT_2[40498] = 32'b00000000000000000000101010101100;
assign LUT_2[40499] = 32'b11111111111111111101100011000101;
assign LUT_2[40500] = 32'b11111111111111110110001111011000;
assign LUT_2[40501] = 32'b11111111111111110011000111110001;
assign LUT_2[40502] = 32'b11111111111111111101001000010100;
assign LUT_2[40503] = 32'b11111111111111111010000000101101;
assign LUT_2[40504] = 32'b11111111111111110100100011001101;
assign LUT_2[40505] = 32'b11111111111111110001011011100110;
assign LUT_2[40506] = 32'b11111111111111111011011100001001;
assign LUT_2[40507] = 32'b11111111111111111000010100100010;
assign LUT_2[40508] = 32'b11111111111111110001000000110101;
assign LUT_2[40509] = 32'b11111111111111101101111001001110;
assign LUT_2[40510] = 32'b11111111111111110111111001110001;
assign LUT_2[40511] = 32'b11111111111111110100110010001010;
assign LUT_2[40512] = 32'b11111111111111110110111010100000;
assign LUT_2[40513] = 32'b11111111111111110011110010111001;
assign LUT_2[40514] = 32'b11111111111111111101110011011100;
assign LUT_2[40515] = 32'b11111111111111111010101011110101;
assign LUT_2[40516] = 32'b11111111111111110011011000001000;
assign LUT_2[40517] = 32'b11111111111111110000010000100001;
assign LUT_2[40518] = 32'b11111111111111111010010001000100;
assign LUT_2[40519] = 32'b11111111111111110111001001011101;
assign LUT_2[40520] = 32'b11111111111111110001101011111101;
assign LUT_2[40521] = 32'b11111111111111101110100100010110;
assign LUT_2[40522] = 32'b11111111111111111000100100111001;
assign LUT_2[40523] = 32'b11111111111111110101011101010010;
assign LUT_2[40524] = 32'b11111111111111101110001001100101;
assign LUT_2[40525] = 32'b11111111111111101011000001111110;
assign LUT_2[40526] = 32'b11111111111111110101000010100001;
assign LUT_2[40527] = 32'b11111111111111110001111010111010;
assign LUT_2[40528] = 32'b11111111111111110001011110101010;
assign LUT_2[40529] = 32'b11111111111111101110010111000011;
assign LUT_2[40530] = 32'b11111111111111111000010111100110;
assign LUT_2[40531] = 32'b11111111111111110101001111111111;
assign LUT_2[40532] = 32'b11111111111111101101111100010010;
assign LUT_2[40533] = 32'b11111111111111101010110100101011;
assign LUT_2[40534] = 32'b11111111111111110100110101001110;
assign LUT_2[40535] = 32'b11111111111111110001101101100111;
assign LUT_2[40536] = 32'b11111111111111101100010000000111;
assign LUT_2[40537] = 32'b11111111111111101001001000100000;
assign LUT_2[40538] = 32'b11111111111111110011001001000011;
assign LUT_2[40539] = 32'b11111111111111110000000001011100;
assign LUT_2[40540] = 32'b11111111111111101000101101101111;
assign LUT_2[40541] = 32'b11111111111111100101100110001000;
assign LUT_2[40542] = 32'b11111111111111101111100110101011;
assign LUT_2[40543] = 32'b11111111111111101100011111000100;
assign LUT_2[40544] = 32'b11111111111111110111010110001001;
assign LUT_2[40545] = 32'b11111111111111110100001110100010;
assign LUT_2[40546] = 32'b11111111111111111110001111000101;
assign LUT_2[40547] = 32'b11111111111111111011000111011110;
assign LUT_2[40548] = 32'b11111111111111110011110011110001;
assign LUT_2[40549] = 32'b11111111111111110000101100001010;
assign LUT_2[40550] = 32'b11111111111111111010101100101101;
assign LUT_2[40551] = 32'b11111111111111110111100101000110;
assign LUT_2[40552] = 32'b11111111111111110010000111100110;
assign LUT_2[40553] = 32'b11111111111111101110111111111111;
assign LUT_2[40554] = 32'b11111111111111111001000000100010;
assign LUT_2[40555] = 32'b11111111111111110101111000111011;
assign LUT_2[40556] = 32'b11111111111111101110100101001110;
assign LUT_2[40557] = 32'b11111111111111101011011101100111;
assign LUT_2[40558] = 32'b11111111111111110101011110001010;
assign LUT_2[40559] = 32'b11111111111111110010010110100011;
assign LUT_2[40560] = 32'b11111111111111110001111010010011;
assign LUT_2[40561] = 32'b11111111111111101110110010101100;
assign LUT_2[40562] = 32'b11111111111111111000110011001111;
assign LUT_2[40563] = 32'b11111111111111110101101011101000;
assign LUT_2[40564] = 32'b11111111111111101110010111111011;
assign LUT_2[40565] = 32'b11111111111111101011010000010100;
assign LUT_2[40566] = 32'b11111111111111110101010000110111;
assign LUT_2[40567] = 32'b11111111111111110010001001010000;
assign LUT_2[40568] = 32'b11111111111111101100101011110000;
assign LUT_2[40569] = 32'b11111111111111101001100100001001;
assign LUT_2[40570] = 32'b11111111111111110011100100101100;
assign LUT_2[40571] = 32'b11111111111111110000011101000101;
assign LUT_2[40572] = 32'b11111111111111101001001001011000;
assign LUT_2[40573] = 32'b11111111111111100110000001110001;
assign LUT_2[40574] = 32'b11111111111111110000000010010100;
assign LUT_2[40575] = 32'b11111111111111101100111010101101;
assign LUT_2[40576] = 32'b00000000000000000011000110001100;
assign LUT_2[40577] = 32'b11111111111111111111111110100101;
assign LUT_2[40578] = 32'b00000000000000001001111111001000;
assign LUT_2[40579] = 32'b00000000000000000110110111100001;
assign LUT_2[40580] = 32'b11111111111111111111100011110100;
assign LUT_2[40581] = 32'b11111111111111111100011100001101;
assign LUT_2[40582] = 32'b00000000000000000110011100110000;
assign LUT_2[40583] = 32'b00000000000000000011010101001001;
assign LUT_2[40584] = 32'b11111111111111111101110111101001;
assign LUT_2[40585] = 32'b11111111111111111010110000000010;
assign LUT_2[40586] = 32'b00000000000000000100110000100101;
assign LUT_2[40587] = 32'b00000000000000000001101000111110;
assign LUT_2[40588] = 32'b11111111111111111010010101010001;
assign LUT_2[40589] = 32'b11111111111111110111001101101010;
assign LUT_2[40590] = 32'b00000000000000000001001110001101;
assign LUT_2[40591] = 32'b11111111111111111110000110100110;
assign LUT_2[40592] = 32'b11111111111111111101101010010110;
assign LUT_2[40593] = 32'b11111111111111111010100010101111;
assign LUT_2[40594] = 32'b00000000000000000100100011010010;
assign LUT_2[40595] = 32'b00000000000000000001011011101011;
assign LUT_2[40596] = 32'b11111111111111111010000111111110;
assign LUT_2[40597] = 32'b11111111111111110111000000010111;
assign LUT_2[40598] = 32'b00000000000000000001000000111010;
assign LUT_2[40599] = 32'b11111111111111111101111001010011;
assign LUT_2[40600] = 32'b11111111111111111000011011110011;
assign LUT_2[40601] = 32'b11111111111111110101010100001100;
assign LUT_2[40602] = 32'b11111111111111111111010100101111;
assign LUT_2[40603] = 32'b11111111111111111100001101001000;
assign LUT_2[40604] = 32'b11111111111111110100111001011011;
assign LUT_2[40605] = 32'b11111111111111110001110001110100;
assign LUT_2[40606] = 32'b11111111111111111011110010010111;
assign LUT_2[40607] = 32'b11111111111111111000101010110000;
assign LUT_2[40608] = 32'b00000000000000000011100001110101;
assign LUT_2[40609] = 32'b00000000000000000000011010001110;
assign LUT_2[40610] = 32'b00000000000000001010011010110001;
assign LUT_2[40611] = 32'b00000000000000000111010011001010;
assign LUT_2[40612] = 32'b11111111111111111111111111011101;
assign LUT_2[40613] = 32'b11111111111111111100110111110110;
assign LUT_2[40614] = 32'b00000000000000000110111000011001;
assign LUT_2[40615] = 32'b00000000000000000011110000110010;
assign LUT_2[40616] = 32'b11111111111111111110010011010010;
assign LUT_2[40617] = 32'b11111111111111111011001011101011;
assign LUT_2[40618] = 32'b00000000000000000101001100001110;
assign LUT_2[40619] = 32'b00000000000000000010000100100111;
assign LUT_2[40620] = 32'b11111111111111111010110000111010;
assign LUT_2[40621] = 32'b11111111111111110111101001010011;
assign LUT_2[40622] = 32'b00000000000000000001101001110110;
assign LUT_2[40623] = 32'b11111111111111111110100010001111;
assign LUT_2[40624] = 32'b11111111111111111110000101111111;
assign LUT_2[40625] = 32'b11111111111111111010111110011000;
assign LUT_2[40626] = 32'b00000000000000000100111110111011;
assign LUT_2[40627] = 32'b00000000000000000001110111010100;
assign LUT_2[40628] = 32'b11111111111111111010100011100111;
assign LUT_2[40629] = 32'b11111111111111110111011100000000;
assign LUT_2[40630] = 32'b00000000000000000001011100100011;
assign LUT_2[40631] = 32'b11111111111111111110010100111100;
assign LUT_2[40632] = 32'b11111111111111111000110111011100;
assign LUT_2[40633] = 32'b11111111111111110101101111110101;
assign LUT_2[40634] = 32'b11111111111111111111110000011000;
assign LUT_2[40635] = 32'b11111111111111111100101000110001;
assign LUT_2[40636] = 32'b11111111111111110101010101000100;
assign LUT_2[40637] = 32'b11111111111111110010001101011101;
assign LUT_2[40638] = 32'b11111111111111111100001110000000;
assign LUT_2[40639] = 32'b11111111111111111001000110011001;
assign LUT_2[40640] = 32'b11111111111111111011001110101111;
assign LUT_2[40641] = 32'b11111111111111111000000111001000;
assign LUT_2[40642] = 32'b00000000000000000010000111101011;
assign LUT_2[40643] = 32'b11111111111111111111000000000100;
assign LUT_2[40644] = 32'b11111111111111110111101100010111;
assign LUT_2[40645] = 32'b11111111111111110100100100110000;
assign LUT_2[40646] = 32'b11111111111111111110100101010011;
assign LUT_2[40647] = 32'b11111111111111111011011101101100;
assign LUT_2[40648] = 32'b11111111111111110110000000001100;
assign LUT_2[40649] = 32'b11111111111111110010111000100101;
assign LUT_2[40650] = 32'b11111111111111111100111001001000;
assign LUT_2[40651] = 32'b11111111111111111001110001100001;
assign LUT_2[40652] = 32'b11111111111111110010011101110100;
assign LUT_2[40653] = 32'b11111111111111101111010110001101;
assign LUT_2[40654] = 32'b11111111111111111001010110110000;
assign LUT_2[40655] = 32'b11111111111111110110001111001001;
assign LUT_2[40656] = 32'b11111111111111110101110010111001;
assign LUT_2[40657] = 32'b11111111111111110010101011010010;
assign LUT_2[40658] = 32'b11111111111111111100101011110101;
assign LUT_2[40659] = 32'b11111111111111111001100100001110;
assign LUT_2[40660] = 32'b11111111111111110010010000100001;
assign LUT_2[40661] = 32'b11111111111111101111001000111010;
assign LUT_2[40662] = 32'b11111111111111111001001001011101;
assign LUT_2[40663] = 32'b11111111111111110110000001110110;
assign LUT_2[40664] = 32'b11111111111111110000100100010110;
assign LUT_2[40665] = 32'b11111111111111101101011100101111;
assign LUT_2[40666] = 32'b11111111111111110111011101010010;
assign LUT_2[40667] = 32'b11111111111111110100010101101011;
assign LUT_2[40668] = 32'b11111111111111101101000001111110;
assign LUT_2[40669] = 32'b11111111111111101001111010010111;
assign LUT_2[40670] = 32'b11111111111111110011111010111010;
assign LUT_2[40671] = 32'b11111111111111110000110011010011;
assign LUT_2[40672] = 32'b11111111111111111011101010011000;
assign LUT_2[40673] = 32'b11111111111111111000100010110001;
assign LUT_2[40674] = 32'b00000000000000000010100011010100;
assign LUT_2[40675] = 32'b11111111111111111111011011101101;
assign LUT_2[40676] = 32'b11111111111111111000001000000000;
assign LUT_2[40677] = 32'b11111111111111110101000000011001;
assign LUT_2[40678] = 32'b11111111111111111111000000111100;
assign LUT_2[40679] = 32'b11111111111111111011111001010101;
assign LUT_2[40680] = 32'b11111111111111110110011011110101;
assign LUT_2[40681] = 32'b11111111111111110011010100001110;
assign LUT_2[40682] = 32'b11111111111111111101010100110001;
assign LUT_2[40683] = 32'b11111111111111111010001101001010;
assign LUT_2[40684] = 32'b11111111111111110010111001011101;
assign LUT_2[40685] = 32'b11111111111111101111110001110110;
assign LUT_2[40686] = 32'b11111111111111111001110010011001;
assign LUT_2[40687] = 32'b11111111111111110110101010110010;
assign LUT_2[40688] = 32'b11111111111111110110001110100010;
assign LUT_2[40689] = 32'b11111111111111110011000110111011;
assign LUT_2[40690] = 32'b11111111111111111101000111011110;
assign LUT_2[40691] = 32'b11111111111111111001111111110111;
assign LUT_2[40692] = 32'b11111111111111110010101100001010;
assign LUT_2[40693] = 32'b11111111111111101111100100100011;
assign LUT_2[40694] = 32'b11111111111111111001100101000110;
assign LUT_2[40695] = 32'b11111111111111110110011101011111;
assign LUT_2[40696] = 32'b11111111111111110000111111111111;
assign LUT_2[40697] = 32'b11111111111111101101111000011000;
assign LUT_2[40698] = 32'b11111111111111110111111000111011;
assign LUT_2[40699] = 32'b11111111111111110100110001010100;
assign LUT_2[40700] = 32'b11111111111111101101011101100111;
assign LUT_2[40701] = 32'b11111111111111101010010110000000;
assign LUT_2[40702] = 32'b11111111111111110100010110100011;
assign LUT_2[40703] = 32'b11111111111111110001001110111100;
assign LUT_2[40704] = 32'b00000000000000000010110000100011;
assign LUT_2[40705] = 32'b11111111111111111111101000111100;
assign LUT_2[40706] = 32'b00000000000000001001101001011111;
assign LUT_2[40707] = 32'b00000000000000000110100001111000;
assign LUT_2[40708] = 32'b11111111111111111111001110001011;
assign LUT_2[40709] = 32'b11111111111111111100000110100100;
assign LUT_2[40710] = 32'b00000000000000000110000111000111;
assign LUT_2[40711] = 32'b00000000000000000010111111100000;
assign LUT_2[40712] = 32'b11111111111111111101100010000000;
assign LUT_2[40713] = 32'b11111111111111111010011010011001;
assign LUT_2[40714] = 32'b00000000000000000100011010111100;
assign LUT_2[40715] = 32'b00000000000000000001010011010101;
assign LUT_2[40716] = 32'b11111111111111111001111111101000;
assign LUT_2[40717] = 32'b11111111111111110110111000000001;
assign LUT_2[40718] = 32'b00000000000000000000111000100100;
assign LUT_2[40719] = 32'b11111111111111111101110000111101;
assign LUT_2[40720] = 32'b11111111111111111101010100101101;
assign LUT_2[40721] = 32'b11111111111111111010001101000110;
assign LUT_2[40722] = 32'b00000000000000000100001101101001;
assign LUT_2[40723] = 32'b00000000000000000001000110000010;
assign LUT_2[40724] = 32'b11111111111111111001110010010101;
assign LUT_2[40725] = 32'b11111111111111110110101010101110;
assign LUT_2[40726] = 32'b00000000000000000000101011010001;
assign LUT_2[40727] = 32'b11111111111111111101100011101010;
assign LUT_2[40728] = 32'b11111111111111111000000110001010;
assign LUT_2[40729] = 32'b11111111111111110100111110100011;
assign LUT_2[40730] = 32'b11111111111111111110111111000110;
assign LUT_2[40731] = 32'b11111111111111111011110111011111;
assign LUT_2[40732] = 32'b11111111111111110100100011110010;
assign LUT_2[40733] = 32'b11111111111111110001011100001011;
assign LUT_2[40734] = 32'b11111111111111111011011100101110;
assign LUT_2[40735] = 32'b11111111111111111000010101000111;
assign LUT_2[40736] = 32'b00000000000000000011001100001100;
assign LUT_2[40737] = 32'b00000000000000000000000100100101;
assign LUT_2[40738] = 32'b00000000000000001010000101001000;
assign LUT_2[40739] = 32'b00000000000000000110111101100001;
assign LUT_2[40740] = 32'b11111111111111111111101001110100;
assign LUT_2[40741] = 32'b11111111111111111100100010001101;
assign LUT_2[40742] = 32'b00000000000000000110100010110000;
assign LUT_2[40743] = 32'b00000000000000000011011011001001;
assign LUT_2[40744] = 32'b11111111111111111101111101101001;
assign LUT_2[40745] = 32'b11111111111111111010110110000010;
assign LUT_2[40746] = 32'b00000000000000000100110110100101;
assign LUT_2[40747] = 32'b00000000000000000001101110111110;
assign LUT_2[40748] = 32'b11111111111111111010011011010001;
assign LUT_2[40749] = 32'b11111111111111110111010011101010;
assign LUT_2[40750] = 32'b00000000000000000001010100001101;
assign LUT_2[40751] = 32'b11111111111111111110001100100110;
assign LUT_2[40752] = 32'b11111111111111111101110000010110;
assign LUT_2[40753] = 32'b11111111111111111010101000101111;
assign LUT_2[40754] = 32'b00000000000000000100101001010010;
assign LUT_2[40755] = 32'b00000000000000000001100001101011;
assign LUT_2[40756] = 32'b11111111111111111010001101111110;
assign LUT_2[40757] = 32'b11111111111111110111000110010111;
assign LUT_2[40758] = 32'b00000000000000000001000110111010;
assign LUT_2[40759] = 32'b11111111111111111101111111010011;
assign LUT_2[40760] = 32'b11111111111111111000100001110011;
assign LUT_2[40761] = 32'b11111111111111110101011010001100;
assign LUT_2[40762] = 32'b11111111111111111111011010101111;
assign LUT_2[40763] = 32'b11111111111111111100010011001000;
assign LUT_2[40764] = 32'b11111111111111110100111111011011;
assign LUT_2[40765] = 32'b11111111111111110001110111110100;
assign LUT_2[40766] = 32'b11111111111111111011111000010111;
assign LUT_2[40767] = 32'b11111111111111111000110000110000;
assign LUT_2[40768] = 32'b11111111111111111010111001000110;
assign LUT_2[40769] = 32'b11111111111111110111110001011111;
assign LUT_2[40770] = 32'b00000000000000000001110010000010;
assign LUT_2[40771] = 32'b11111111111111111110101010011011;
assign LUT_2[40772] = 32'b11111111111111110111010110101110;
assign LUT_2[40773] = 32'b11111111111111110100001111000111;
assign LUT_2[40774] = 32'b11111111111111111110001111101010;
assign LUT_2[40775] = 32'b11111111111111111011001000000011;
assign LUT_2[40776] = 32'b11111111111111110101101010100011;
assign LUT_2[40777] = 32'b11111111111111110010100010111100;
assign LUT_2[40778] = 32'b11111111111111111100100011011111;
assign LUT_2[40779] = 32'b11111111111111111001011011111000;
assign LUT_2[40780] = 32'b11111111111111110010001000001011;
assign LUT_2[40781] = 32'b11111111111111101111000000100100;
assign LUT_2[40782] = 32'b11111111111111111001000001000111;
assign LUT_2[40783] = 32'b11111111111111110101111001100000;
assign LUT_2[40784] = 32'b11111111111111110101011101010000;
assign LUT_2[40785] = 32'b11111111111111110010010101101001;
assign LUT_2[40786] = 32'b11111111111111111100010110001100;
assign LUT_2[40787] = 32'b11111111111111111001001110100101;
assign LUT_2[40788] = 32'b11111111111111110001111010111000;
assign LUT_2[40789] = 32'b11111111111111101110110011010001;
assign LUT_2[40790] = 32'b11111111111111111000110011110100;
assign LUT_2[40791] = 32'b11111111111111110101101100001101;
assign LUT_2[40792] = 32'b11111111111111110000001110101101;
assign LUT_2[40793] = 32'b11111111111111101101000111000110;
assign LUT_2[40794] = 32'b11111111111111110111000111101001;
assign LUT_2[40795] = 32'b11111111111111110100000000000010;
assign LUT_2[40796] = 32'b11111111111111101100101100010101;
assign LUT_2[40797] = 32'b11111111111111101001100100101110;
assign LUT_2[40798] = 32'b11111111111111110011100101010001;
assign LUT_2[40799] = 32'b11111111111111110000011101101010;
assign LUT_2[40800] = 32'b11111111111111111011010100101111;
assign LUT_2[40801] = 32'b11111111111111111000001101001000;
assign LUT_2[40802] = 32'b00000000000000000010001101101011;
assign LUT_2[40803] = 32'b11111111111111111111000110000100;
assign LUT_2[40804] = 32'b11111111111111110111110010010111;
assign LUT_2[40805] = 32'b11111111111111110100101010110000;
assign LUT_2[40806] = 32'b11111111111111111110101011010011;
assign LUT_2[40807] = 32'b11111111111111111011100011101100;
assign LUT_2[40808] = 32'b11111111111111110110000110001100;
assign LUT_2[40809] = 32'b11111111111111110010111110100101;
assign LUT_2[40810] = 32'b11111111111111111100111111001000;
assign LUT_2[40811] = 32'b11111111111111111001110111100001;
assign LUT_2[40812] = 32'b11111111111111110010100011110100;
assign LUT_2[40813] = 32'b11111111111111101111011100001101;
assign LUT_2[40814] = 32'b11111111111111111001011100110000;
assign LUT_2[40815] = 32'b11111111111111110110010101001001;
assign LUT_2[40816] = 32'b11111111111111110101111000111001;
assign LUT_2[40817] = 32'b11111111111111110010110001010010;
assign LUT_2[40818] = 32'b11111111111111111100110001110101;
assign LUT_2[40819] = 32'b11111111111111111001101010001110;
assign LUT_2[40820] = 32'b11111111111111110010010110100001;
assign LUT_2[40821] = 32'b11111111111111101111001110111010;
assign LUT_2[40822] = 32'b11111111111111111001001111011101;
assign LUT_2[40823] = 32'b11111111111111110110000111110110;
assign LUT_2[40824] = 32'b11111111111111110000101010010110;
assign LUT_2[40825] = 32'b11111111111111101101100010101111;
assign LUT_2[40826] = 32'b11111111111111110111100011010010;
assign LUT_2[40827] = 32'b11111111111111110100011011101011;
assign LUT_2[40828] = 32'b11111111111111101101000111111110;
assign LUT_2[40829] = 32'b11111111111111101010000000010111;
assign LUT_2[40830] = 32'b11111111111111110100000000111010;
assign LUT_2[40831] = 32'b11111111111111110000111001010011;
assign LUT_2[40832] = 32'b00000000000000000111000100110010;
assign LUT_2[40833] = 32'b00000000000000000011111101001011;
assign LUT_2[40834] = 32'b00000000000000001101111101101110;
assign LUT_2[40835] = 32'b00000000000000001010110110000111;
assign LUT_2[40836] = 32'b00000000000000000011100010011010;
assign LUT_2[40837] = 32'b00000000000000000000011010110011;
assign LUT_2[40838] = 32'b00000000000000001010011011010110;
assign LUT_2[40839] = 32'b00000000000000000111010011101111;
assign LUT_2[40840] = 32'b00000000000000000001110110001111;
assign LUT_2[40841] = 32'b11111111111111111110101110101000;
assign LUT_2[40842] = 32'b00000000000000001000101111001011;
assign LUT_2[40843] = 32'b00000000000000000101100111100100;
assign LUT_2[40844] = 32'b11111111111111111110010011110111;
assign LUT_2[40845] = 32'b11111111111111111011001100010000;
assign LUT_2[40846] = 32'b00000000000000000101001100110011;
assign LUT_2[40847] = 32'b00000000000000000010000101001100;
assign LUT_2[40848] = 32'b00000000000000000001101000111100;
assign LUT_2[40849] = 32'b11111111111111111110100001010101;
assign LUT_2[40850] = 32'b00000000000000001000100001111000;
assign LUT_2[40851] = 32'b00000000000000000101011010010001;
assign LUT_2[40852] = 32'b11111111111111111110000110100100;
assign LUT_2[40853] = 32'b11111111111111111010111110111101;
assign LUT_2[40854] = 32'b00000000000000000100111111100000;
assign LUT_2[40855] = 32'b00000000000000000001110111111001;
assign LUT_2[40856] = 32'b11111111111111111100011010011001;
assign LUT_2[40857] = 32'b11111111111111111001010010110010;
assign LUT_2[40858] = 32'b00000000000000000011010011010101;
assign LUT_2[40859] = 32'b00000000000000000000001011101110;
assign LUT_2[40860] = 32'b11111111111111111000111000000001;
assign LUT_2[40861] = 32'b11111111111111110101110000011010;
assign LUT_2[40862] = 32'b11111111111111111111110000111101;
assign LUT_2[40863] = 32'b11111111111111111100101001010110;
assign LUT_2[40864] = 32'b00000000000000000111100000011011;
assign LUT_2[40865] = 32'b00000000000000000100011000110100;
assign LUT_2[40866] = 32'b00000000000000001110011001010111;
assign LUT_2[40867] = 32'b00000000000000001011010001110000;
assign LUT_2[40868] = 32'b00000000000000000011111110000011;
assign LUT_2[40869] = 32'b00000000000000000000110110011100;
assign LUT_2[40870] = 32'b00000000000000001010110110111111;
assign LUT_2[40871] = 32'b00000000000000000111101111011000;
assign LUT_2[40872] = 32'b00000000000000000010010001111000;
assign LUT_2[40873] = 32'b11111111111111111111001010010001;
assign LUT_2[40874] = 32'b00000000000000001001001010110100;
assign LUT_2[40875] = 32'b00000000000000000110000011001101;
assign LUT_2[40876] = 32'b11111111111111111110101111100000;
assign LUT_2[40877] = 32'b11111111111111111011100111111001;
assign LUT_2[40878] = 32'b00000000000000000101101000011100;
assign LUT_2[40879] = 32'b00000000000000000010100000110101;
assign LUT_2[40880] = 32'b00000000000000000010000100100101;
assign LUT_2[40881] = 32'b11111111111111111110111100111110;
assign LUT_2[40882] = 32'b00000000000000001000111101100001;
assign LUT_2[40883] = 32'b00000000000000000101110101111010;
assign LUT_2[40884] = 32'b11111111111111111110100010001101;
assign LUT_2[40885] = 32'b11111111111111111011011010100110;
assign LUT_2[40886] = 32'b00000000000000000101011011001001;
assign LUT_2[40887] = 32'b00000000000000000010010011100010;
assign LUT_2[40888] = 32'b11111111111111111100110110000010;
assign LUT_2[40889] = 32'b11111111111111111001101110011011;
assign LUT_2[40890] = 32'b00000000000000000011101110111110;
assign LUT_2[40891] = 32'b00000000000000000000100111010111;
assign LUT_2[40892] = 32'b11111111111111111001010011101010;
assign LUT_2[40893] = 32'b11111111111111110110001100000011;
assign LUT_2[40894] = 32'b00000000000000000000001100100110;
assign LUT_2[40895] = 32'b11111111111111111101000100111111;
assign LUT_2[40896] = 32'b11111111111111111111001101010101;
assign LUT_2[40897] = 32'b11111111111111111100000101101110;
assign LUT_2[40898] = 32'b00000000000000000110000110010001;
assign LUT_2[40899] = 32'b00000000000000000010111110101010;
assign LUT_2[40900] = 32'b11111111111111111011101010111101;
assign LUT_2[40901] = 32'b11111111111111111000100011010110;
assign LUT_2[40902] = 32'b00000000000000000010100011111001;
assign LUT_2[40903] = 32'b11111111111111111111011100010010;
assign LUT_2[40904] = 32'b11111111111111111001111110110010;
assign LUT_2[40905] = 32'b11111111111111110110110111001011;
assign LUT_2[40906] = 32'b00000000000000000000110111101110;
assign LUT_2[40907] = 32'b11111111111111111101110000000111;
assign LUT_2[40908] = 32'b11111111111111110110011100011010;
assign LUT_2[40909] = 32'b11111111111111110011010100110011;
assign LUT_2[40910] = 32'b11111111111111111101010101010110;
assign LUT_2[40911] = 32'b11111111111111111010001101101111;
assign LUT_2[40912] = 32'b11111111111111111001110001011111;
assign LUT_2[40913] = 32'b11111111111111110110101001111000;
assign LUT_2[40914] = 32'b00000000000000000000101010011011;
assign LUT_2[40915] = 32'b11111111111111111101100010110100;
assign LUT_2[40916] = 32'b11111111111111110110001111000111;
assign LUT_2[40917] = 32'b11111111111111110011000111100000;
assign LUT_2[40918] = 32'b11111111111111111101001000000011;
assign LUT_2[40919] = 32'b11111111111111111010000000011100;
assign LUT_2[40920] = 32'b11111111111111110100100010111100;
assign LUT_2[40921] = 32'b11111111111111110001011011010101;
assign LUT_2[40922] = 32'b11111111111111111011011011111000;
assign LUT_2[40923] = 32'b11111111111111111000010100010001;
assign LUT_2[40924] = 32'b11111111111111110001000000100100;
assign LUT_2[40925] = 32'b11111111111111101101111000111101;
assign LUT_2[40926] = 32'b11111111111111110111111001100000;
assign LUT_2[40927] = 32'b11111111111111110100110001111001;
assign LUT_2[40928] = 32'b11111111111111111111101000111110;
assign LUT_2[40929] = 32'b11111111111111111100100001010111;
assign LUT_2[40930] = 32'b00000000000000000110100001111010;
assign LUT_2[40931] = 32'b00000000000000000011011010010011;
assign LUT_2[40932] = 32'b11111111111111111100000110100110;
assign LUT_2[40933] = 32'b11111111111111111000111110111111;
assign LUT_2[40934] = 32'b00000000000000000010111111100010;
assign LUT_2[40935] = 32'b11111111111111111111110111111011;
assign LUT_2[40936] = 32'b11111111111111111010011010011011;
assign LUT_2[40937] = 32'b11111111111111110111010010110100;
assign LUT_2[40938] = 32'b00000000000000000001010011010111;
assign LUT_2[40939] = 32'b11111111111111111110001011110000;
assign LUT_2[40940] = 32'b11111111111111110110111000000011;
assign LUT_2[40941] = 32'b11111111111111110011110000011100;
assign LUT_2[40942] = 32'b11111111111111111101110000111111;
assign LUT_2[40943] = 32'b11111111111111111010101001011000;
assign LUT_2[40944] = 32'b11111111111111111010001101001000;
assign LUT_2[40945] = 32'b11111111111111110111000101100001;
assign LUT_2[40946] = 32'b00000000000000000001000110000100;
assign LUT_2[40947] = 32'b11111111111111111101111110011101;
assign LUT_2[40948] = 32'b11111111111111110110101010110000;
assign LUT_2[40949] = 32'b11111111111111110011100011001001;
assign LUT_2[40950] = 32'b11111111111111111101100011101100;
assign LUT_2[40951] = 32'b11111111111111111010011100000101;
assign LUT_2[40952] = 32'b11111111111111110100111110100101;
assign LUT_2[40953] = 32'b11111111111111110001110110111110;
assign LUT_2[40954] = 32'b11111111111111111011110111100001;
assign LUT_2[40955] = 32'b11111111111111111000101111111010;
assign LUT_2[40956] = 32'b11111111111111110001011100001101;
assign LUT_2[40957] = 32'b11111111111111101110010100100110;
assign LUT_2[40958] = 32'b11111111111111111000010101001001;
assign LUT_2[40959] = 32'b11111111111111110101001101100010;
assign LUT_2[40960] = 32'b11111111111111110001101111111101;
assign LUT_2[40961] = 32'b11111111111111101110101000010110;
assign LUT_2[40962] = 32'b11111111111111111000101000111001;
assign LUT_2[40963] = 32'b11111111111111110101100001010010;
assign LUT_2[40964] = 32'b11111111111111101110001101100101;
assign LUT_2[40965] = 32'b11111111111111101011000101111110;
assign LUT_2[40966] = 32'b11111111111111110101000110100001;
assign LUT_2[40967] = 32'b11111111111111110001111110111010;
assign LUT_2[40968] = 32'b11111111111111101100100001011010;
assign LUT_2[40969] = 32'b11111111111111101001011001110011;
assign LUT_2[40970] = 32'b11111111111111110011011010010110;
assign LUT_2[40971] = 32'b11111111111111110000010010101111;
assign LUT_2[40972] = 32'b11111111111111101000111111000010;
assign LUT_2[40973] = 32'b11111111111111100101110111011011;
assign LUT_2[40974] = 32'b11111111111111101111110111111110;
assign LUT_2[40975] = 32'b11111111111111101100110000010111;
assign LUT_2[40976] = 32'b11111111111111101100010100000111;
assign LUT_2[40977] = 32'b11111111111111101001001100100000;
assign LUT_2[40978] = 32'b11111111111111110011001101000011;
assign LUT_2[40979] = 32'b11111111111111110000000101011100;
assign LUT_2[40980] = 32'b11111111111111101000110001101111;
assign LUT_2[40981] = 32'b11111111111111100101101010001000;
assign LUT_2[40982] = 32'b11111111111111101111101010101011;
assign LUT_2[40983] = 32'b11111111111111101100100011000100;
assign LUT_2[40984] = 32'b11111111111111100111000101100100;
assign LUT_2[40985] = 32'b11111111111111100011111101111101;
assign LUT_2[40986] = 32'b11111111111111101101111110100000;
assign LUT_2[40987] = 32'b11111111111111101010110110111001;
assign LUT_2[40988] = 32'b11111111111111100011100011001100;
assign LUT_2[40989] = 32'b11111111111111100000011011100101;
assign LUT_2[40990] = 32'b11111111111111101010011100001000;
assign LUT_2[40991] = 32'b11111111111111100111010100100001;
assign LUT_2[40992] = 32'b11111111111111110010001011100110;
assign LUT_2[40993] = 32'b11111111111111101111000011111111;
assign LUT_2[40994] = 32'b11111111111111111001000100100010;
assign LUT_2[40995] = 32'b11111111111111110101111100111011;
assign LUT_2[40996] = 32'b11111111111111101110101001001110;
assign LUT_2[40997] = 32'b11111111111111101011100001100111;
assign LUT_2[40998] = 32'b11111111111111110101100010001010;
assign LUT_2[40999] = 32'b11111111111111110010011010100011;
assign LUT_2[41000] = 32'b11111111111111101100111101000011;
assign LUT_2[41001] = 32'b11111111111111101001110101011100;
assign LUT_2[41002] = 32'b11111111111111110011110101111111;
assign LUT_2[41003] = 32'b11111111111111110000101110011000;
assign LUT_2[41004] = 32'b11111111111111101001011010101011;
assign LUT_2[41005] = 32'b11111111111111100110010011000100;
assign LUT_2[41006] = 32'b11111111111111110000010011100111;
assign LUT_2[41007] = 32'b11111111111111101101001100000000;
assign LUT_2[41008] = 32'b11111111111111101100101111110000;
assign LUT_2[41009] = 32'b11111111111111101001101000001001;
assign LUT_2[41010] = 32'b11111111111111110011101000101100;
assign LUT_2[41011] = 32'b11111111111111110000100001000101;
assign LUT_2[41012] = 32'b11111111111111101001001101011000;
assign LUT_2[41013] = 32'b11111111111111100110000101110001;
assign LUT_2[41014] = 32'b11111111111111110000000110010100;
assign LUT_2[41015] = 32'b11111111111111101100111110101101;
assign LUT_2[41016] = 32'b11111111111111100111100001001101;
assign LUT_2[41017] = 32'b11111111111111100100011001100110;
assign LUT_2[41018] = 32'b11111111111111101110011010001001;
assign LUT_2[41019] = 32'b11111111111111101011010010100010;
assign LUT_2[41020] = 32'b11111111111111100011111110110101;
assign LUT_2[41021] = 32'b11111111111111100000110111001110;
assign LUT_2[41022] = 32'b11111111111111101010110111110001;
assign LUT_2[41023] = 32'b11111111111111100111110000001010;
assign LUT_2[41024] = 32'b11111111111111101001111000100000;
assign LUT_2[41025] = 32'b11111111111111100110110000111001;
assign LUT_2[41026] = 32'b11111111111111110000110001011100;
assign LUT_2[41027] = 32'b11111111111111101101101001110101;
assign LUT_2[41028] = 32'b11111111111111100110010110001000;
assign LUT_2[41029] = 32'b11111111111111100011001110100001;
assign LUT_2[41030] = 32'b11111111111111101101001111000100;
assign LUT_2[41031] = 32'b11111111111111101010000111011101;
assign LUT_2[41032] = 32'b11111111111111100100101001111101;
assign LUT_2[41033] = 32'b11111111111111100001100010010110;
assign LUT_2[41034] = 32'b11111111111111101011100010111001;
assign LUT_2[41035] = 32'b11111111111111101000011011010010;
assign LUT_2[41036] = 32'b11111111111111100001000111100101;
assign LUT_2[41037] = 32'b11111111111111011101111111111110;
assign LUT_2[41038] = 32'b11111111111111101000000000100001;
assign LUT_2[41039] = 32'b11111111111111100100111000111010;
assign LUT_2[41040] = 32'b11111111111111100100011100101010;
assign LUT_2[41041] = 32'b11111111111111100001010101000011;
assign LUT_2[41042] = 32'b11111111111111101011010101100110;
assign LUT_2[41043] = 32'b11111111111111101000001101111111;
assign LUT_2[41044] = 32'b11111111111111100000111010010010;
assign LUT_2[41045] = 32'b11111111111111011101110010101011;
assign LUT_2[41046] = 32'b11111111111111100111110011001110;
assign LUT_2[41047] = 32'b11111111111111100100101011100111;
assign LUT_2[41048] = 32'b11111111111111011111001110000111;
assign LUT_2[41049] = 32'b11111111111111011100000110100000;
assign LUT_2[41050] = 32'b11111111111111100110000111000011;
assign LUT_2[41051] = 32'b11111111111111100010111111011100;
assign LUT_2[41052] = 32'b11111111111111011011101011101111;
assign LUT_2[41053] = 32'b11111111111111011000100100001000;
assign LUT_2[41054] = 32'b11111111111111100010100100101011;
assign LUT_2[41055] = 32'b11111111111111011111011101000100;
assign LUT_2[41056] = 32'b11111111111111101010010100001001;
assign LUT_2[41057] = 32'b11111111111111100111001100100010;
assign LUT_2[41058] = 32'b11111111111111110001001101000101;
assign LUT_2[41059] = 32'b11111111111111101110000101011110;
assign LUT_2[41060] = 32'b11111111111111100110110001110001;
assign LUT_2[41061] = 32'b11111111111111100011101010001010;
assign LUT_2[41062] = 32'b11111111111111101101101010101101;
assign LUT_2[41063] = 32'b11111111111111101010100011000110;
assign LUT_2[41064] = 32'b11111111111111100101000101100110;
assign LUT_2[41065] = 32'b11111111111111100001111101111111;
assign LUT_2[41066] = 32'b11111111111111101011111110100010;
assign LUT_2[41067] = 32'b11111111111111101000110110111011;
assign LUT_2[41068] = 32'b11111111111111100001100011001110;
assign LUT_2[41069] = 32'b11111111111111011110011011100111;
assign LUT_2[41070] = 32'b11111111111111101000011100001010;
assign LUT_2[41071] = 32'b11111111111111100101010100100011;
assign LUT_2[41072] = 32'b11111111111111100100111000010011;
assign LUT_2[41073] = 32'b11111111111111100001110000101100;
assign LUT_2[41074] = 32'b11111111111111101011110001001111;
assign LUT_2[41075] = 32'b11111111111111101000101001101000;
assign LUT_2[41076] = 32'b11111111111111100001010101111011;
assign LUT_2[41077] = 32'b11111111111111011110001110010100;
assign LUT_2[41078] = 32'b11111111111111101000001110110111;
assign LUT_2[41079] = 32'b11111111111111100101000111010000;
assign LUT_2[41080] = 32'b11111111111111011111101001110000;
assign LUT_2[41081] = 32'b11111111111111011100100010001001;
assign LUT_2[41082] = 32'b11111111111111100110100010101100;
assign LUT_2[41083] = 32'b11111111111111100011011011000101;
assign LUT_2[41084] = 32'b11111111111111011100000111011000;
assign LUT_2[41085] = 32'b11111111111111011000111111110001;
assign LUT_2[41086] = 32'b11111111111111100011000000010100;
assign LUT_2[41087] = 32'b11111111111111011111111000101101;
assign LUT_2[41088] = 32'b11111111111111110110000100001100;
assign LUT_2[41089] = 32'b11111111111111110010111100100101;
assign LUT_2[41090] = 32'b11111111111111111100111101001000;
assign LUT_2[41091] = 32'b11111111111111111001110101100001;
assign LUT_2[41092] = 32'b11111111111111110010100001110100;
assign LUT_2[41093] = 32'b11111111111111101111011010001101;
assign LUT_2[41094] = 32'b11111111111111111001011010110000;
assign LUT_2[41095] = 32'b11111111111111110110010011001001;
assign LUT_2[41096] = 32'b11111111111111110000110101101001;
assign LUT_2[41097] = 32'b11111111111111101101101110000010;
assign LUT_2[41098] = 32'b11111111111111110111101110100101;
assign LUT_2[41099] = 32'b11111111111111110100100110111110;
assign LUT_2[41100] = 32'b11111111111111101101010011010001;
assign LUT_2[41101] = 32'b11111111111111101010001011101010;
assign LUT_2[41102] = 32'b11111111111111110100001100001101;
assign LUT_2[41103] = 32'b11111111111111110001000100100110;
assign LUT_2[41104] = 32'b11111111111111110000101000010110;
assign LUT_2[41105] = 32'b11111111111111101101100000101111;
assign LUT_2[41106] = 32'b11111111111111110111100001010010;
assign LUT_2[41107] = 32'b11111111111111110100011001101011;
assign LUT_2[41108] = 32'b11111111111111101101000101111110;
assign LUT_2[41109] = 32'b11111111111111101001111110010111;
assign LUT_2[41110] = 32'b11111111111111110011111110111010;
assign LUT_2[41111] = 32'b11111111111111110000110111010011;
assign LUT_2[41112] = 32'b11111111111111101011011001110011;
assign LUT_2[41113] = 32'b11111111111111101000010010001100;
assign LUT_2[41114] = 32'b11111111111111110010010010101111;
assign LUT_2[41115] = 32'b11111111111111101111001011001000;
assign LUT_2[41116] = 32'b11111111111111100111110111011011;
assign LUT_2[41117] = 32'b11111111111111100100101111110100;
assign LUT_2[41118] = 32'b11111111111111101110110000010111;
assign LUT_2[41119] = 32'b11111111111111101011101000110000;
assign LUT_2[41120] = 32'b11111111111111110110011111110101;
assign LUT_2[41121] = 32'b11111111111111110011011000001110;
assign LUT_2[41122] = 32'b11111111111111111101011000110001;
assign LUT_2[41123] = 32'b11111111111111111010010001001010;
assign LUT_2[41124] = 32'b11111111111111110010111101011101;
assign LUT_2[41125] = 32'b11111111111111101111110101110110;
assign LUT_2[41126] = 32'b11111111111111111001110110011001;
assign LUT_2[41127] = 32'b11111111111111110110101110110010;
assign LUT_2[41128] = 32'b11111111111111110001010001010010;
assign LUT_2[41129] = 32'b11111111111111101110001001101011;
assign LUT_2[41130] = 32'b11111111111111111000001010001110;
assign LUT_2[41131] = 32'b11111111111111110101000010100111;
assign LUT_2[41132] = 32'b11111111111111101101101110111010;
assign LUT_2[41133] = 32'b11111111111111101010100111010011;
assign LUT_2[41134] = 32'b11111111111111110100100111110110;
assign LUT_2[41135] = 32'b11111111111111110001100000001111;
assign LUT_2[41136] = 32'b11111111111111110001000011111111;
assign LUT_2[41137] = 32'b11111111111111101101111100011000;
assign LUT_2[41138] = 32'b11111111111111110111111100111011;
assign LUT_2[41139] = 32'b11111111111111110100110101010100;
assign LUT_2[41140] = 32'b11111111111111101101100001100111;
assign LUT_2[41141] = 32'b11111111111111101010011010000000;
assign LUT_2[41142] = 32'b11111111111111110100011010100011;
assign LUT_2[41143] = 32'b11111111111111110001010010111100;
assign LUT_2[41144] = 32'b11111111111111101011110101011100;
assign LUT_2[41145] = 32'b11111111111111101000101101110101;
assign LUT_2[41146] = 32'b11111111111111110010101110011000;
assign LUT_2[41147] = 32'b11111111111111101111100110110001;
assign LUT_2[41148] = 32'b11111111111111101000010011000100;
assign LUT_2[41149] = 32'b11111111111111100101001011011101;
assign LUT_2[41150] = 32'b11111111111111101111001100000000;
assign LUT_2[41151] = 32'b11111111111111101100000100011001;
assign LUT_2[41152] = 32'b11111111111111101110001100101111;
assign LUT_2[41153] = 32'b11111111111111101011000101001000;
assign LUT_2[41154] = 32'b11111111111111110101000101101011;
assign LUT_2[41155] = 32'b11111111111111110001111110000100;
assign LUT_2[41156] = 32'b11111111111111101010101010010111;
assign LUT_2[41157] = 32'b11111111111111100111100010110000;
assign LUT_2[41158] = 32'b11111111111111110001100011010011;
assign LUT_2[41159] = 32'b11111111111111101110011011101100;
assign LUT_2[41160] = 32'b11111111111111101000111110001100;
assign LUT_2[41161] = 32'b11111111111111100101110110100101;
assign LUT_2[41162] = 32'b11111111111111101111110111001000;
assign LUT_2[41163] = 32'b11111111111111101100101111100001;
assign LUT_2[41164] = 32'b11111111111111100101011011110100;
assign LUT_2[41165] = 32'b11111111111111100010010100001101;
assign LUT_2[41166] = 32'b11111111111111101100010100110000;
assign LUT_2[41167] = 32'b11111111111111101001001101001001;
assign LUT_2[41168] = 32'b11111111111111101000110000111001;
assign LUT_2[41169] = 32'b11111111111111100101101001010010;
assign LUT_2[41170] = 32'b11111111111111101111101001110101;
assign LUT_2[41171] = 32'b11111111111111101100100010001110;
assign LUT_2[41172] = 32'b11111111111111100101001110100001;
assign LUT_2[41173] = 32'b11111111111111100010000110111010;
assign LUT_2[41174] = 32'b11111111111111101100000111011101;
assign LUT_2[41175] = 32'b11111111111111101000111111110110;
assign LUT_2[41176] = 32'b11111111111111100011100010010110;
assign LUT_2[41177] = 32'b11111111111111100000011010101111;
assign LUT_2[41178] = 32'b11111111111111101010011011010010;
assign LUT_2[41179] = 32'b11111111111111100111010011101011;
assign LUT_2[41180] = 32'b11111111111111011111111111111110;
assign LUT_2[41181] = 32'b11111111111111011100111000010111;
assign LUT_2[41182] = 32'b11111111111111100110111000111010;
assign LUT_2[41183] = 32'b11111111111111100011110001010011;
assign LUT_2[41184] = 32'b11111111111111101110101000011000;
assign LUT_2[41185] = 32'b11111111111111101011100000110001;
assign LUT_2[41186] = 32'b11111111111111110101100001010100;
assign LUT_2[41187] = 32'b11111111111111110010011001101101;
assign LUT_2[41188] = 32'b11111111111111101011000110000000;
assign LUT_2[41189] = 32'b11111111111111100111111110011001;
assign LUT_2[41190] = 32'b11111111111111110001111110111100;
assign LUT_2[41191] = 32'b11111111111111101110110111010101;
assign LUT_2[41192] = 32'b11111111111111101001011001110101;
assign LUT_2[41193] = 32'b11111111111111100110010010001110;
assign LUT_2[41194] = 32'b11111111111111110000010010110001;
assign LUT_2[41195] = 32'b11111111111111101101001011001010;
assign LUT_2[41196] = 32'b11111111111111100101110111011101;
assign LUT_2[41197] = 32'b11111111111111100010101111110110;
assign LUT_2[41198] = 32'b11111111111111101100110000011001;
assign LUT_2[41199] = 32'b11111111111111101001101000110010;
assign LUT_2[41200] = 32'b11111111111111101001001100100010;
assign LUT_2[41201] = 32'b11111111111111100110000100111011;
assign LUT_2[41202] = 32'b11111111111111110000000101011110;
assign LUT_2[41203] = 32'b11111111111111101100111101110111;
assign LUT_2[41204] = 32'b11111111111111100101101010001010;
assign LUT_2[41205] = 32'b11111111111111100010100010100011;
assign LUT_2[41206] = 32'b11111111111111101100100011000110;
assign LUT_2[41207] = 32'b11111111111111101001011011011111;
assign LUT_2[41208] = 32'b11111111111111100011111101111111;
assign LUT_2[41209] = 32'b11111111111111100000110110011000;
assign LUT_2[41210] = 32'b11111111111111101010110110111011;
assign LUT_2[41211] = 32'b11111111111111100111101111010100;
assign LUT_2[41212] = 32'b11111111111111100000011011100111;
assign LUT_2[41213] = 32'b11111111111111011101010100000000;
assign LUT_2[41214] = 32'b11111111111111100111010100100011;
assign LUT_2[41215] = 32'b11111111111111100100001100111100;
assign LUT_2[41216] = 32'b11111111111111110101101110100011;
assign LUT_2[41217] = 32'b11111111111111110010100110111100;
assign LUT_2[41218] = 32'b11111111111111111100100111011111;
assign LUT_2[41219] = 32'b11111111111111111001011111111000;
assign LUT_2[41220] = 32'b11111111111111110010001100001011;
assign LUT_2[41221] = 32'b11111111111111101111000100100100;
assign LUT_2[41222] = 32'b11111111111111111001000101000111;
assign LUT_2[41223] = 32'b11111111111111110101111101100000;
assign LUT_2[41224] = 32'b11111111111111110000100000000000;
assign LUT_2[41225] = 32'b11111111111111101101011000011001;
assign LUT_2[41226] = 32'b11111111111111110111011000111100;
assign LUT_2[41227] = 32'b11111111111111110100010001010101;
assign LUT_2[41228] = 32'b11111111111111101100111101101000;
assign LUT_2[41229] = 32'b11111111111111101001110110000001;
assign LUT_2[41230] = 32'b11111111111111110011110110100100;
assign LUT_2[41231] = 32'b11111111111111110000101110111101;
assign LUT_2[41232] = 32'b11111111111111110000010010101101;
assign LUT_2[41233] = 32'b11111111111111101101001011000110;
assign LUT_2[41234] = 32'b11111111111111110111001011101001;
assign LUT_2[41235] = 32'b11111111111111110100000100000010;
assign LUT_2[41236] = 32'b11111111111111101100110000010101;
assign LUT_2[41237] = 32'b11111111111111101001101000101110;
assign LUT_2[41238] = 32'b11111111111111110011101001010001;
assign LUT_2[41239] = 32'b11111111111111110000100001101010;
assign LUT_2[41240] = 32'b11111111111111101011000100001010;
assign LUT_2[41241] = 32'b11111111111111100111111100100011;
assign LUT_2[41242] = 32'b11111111111111110001111101000110;
assign LUT_2[41243] = 32'b11111111111111101110110101011111;
assign LUT_2[41244] = 32'b11111111111111100111100001110010;
assign LUT_2[41245] = 32'b11111111111111100100011010001011;
assign LUT_2[41246] = 32'b11111111111111101110011010101110;
assign LUT_2[41247] = 32'b11111111111111101011010011000111;
assign LUT_2[41248] = 32'b11111111111111110110001010001100;
assign LUT_2[41249] = 32'b11111111111111110011000010100101;
assign LUT_2[41250] = 32'b11111111111111111101000011001000;
assign LUT_2[41251] = 32'b11111111111111111001111011100001;
assign LUT_2[41252] = 32'b11111111111111110010100111110100;
assign LUT_2[41253] = 32'b11111111111111101111100000001101;
assign LUT_2[41254] = 32'b11111111111111111001100000110000;
assign LUT_2[41255] = 32'b11111111111111110110011001001001;
assign LUT_2[41256] = 32'b11111111111111110000111011101001;
assign LUT_2[41257] = 32'b11111111111111101101110100000010;
assign LUT_2[41258] = 32'b11111111111111110111110100100101;
assign LUT_2[41259] = 32'b11111111111111110100101100111110;
assign LUT_2[41260] = 32'b11111111111111101101011001010001;
assign LUT_2[41261] = 32'b11111111111111101010010001101010;
assign LUT_2[41262] = 32'b11111111111111110100010010001101;
assign LUT_2[41263] = 32'b11111111111111110001001010100110;
assign LUT_2[41264] = 32'b11111111111111110000101110010110;
assign LUT_2[41265] = 32'b11111111111111101101100110101111;
assign LUT_2[41266] = 32'b11111111111111110111100111010010;
assign LUT_2[41267] = 32'b11111111111111110100011111101011;
assign LUT_2[41268] = 32'b11111111111111101101001011111110;
assign LUT_2[41269] = 32'b11111111111111101010000100010111;
assign LUT_2[41270] = 32'b11111111111111110100000100111010;
assign LUT_2[41271] = 32'b11111111111111110000111101010011;
assign LUT_2[41272] = 32'b11111111111111101011011111110011;
assign LUT_2[41273] = 32'b11111111111111101000011000001100;
assign LUT_2[41274] = 32'b11111111111111110010011000101111;
assign LUT_2[41275] = 32'b11111111111111101111010001001000;
assign LUT_2[41276] = 32'b11111111111111100111111101011011;
assign LUT_2[41277] = 32'b11111111111111100100110101110100;
assign LUT_2[41278] = 32'b11111111111111101110110110010111;
assign LUT_2[41279] = 32'b11111111111111101011101110110000;
assign LUT_2[41280] = 32'b11111111111111101101110111000110;
assign LUT_2[41281] = 32'b11111111111111101010101111011111;
assign LUT_2[41282] = 32'b11111111111111110100110000000010;
assign LUT_2[41283] = 32'b11111111111111110001101000011011;
assign LUT_2[41284] = 32'b11111111111111101010010100101110;
assign LUT_2[41285] = 32'b11111111111111100111001101000111;
assign LUT_2[41286] = 32'b11111111111111110001001101101010;
assign LUT_2[41287] = 32'b11111111111111101110000110000011;
assign LUT_2[41288] = 32'b11111111111111101000101000100011;
assign LUT_2[41289] = 32'b11111111111111100101100000111100;
assign LUT_2[41290] = 32'b11111111111111101111100001011111;
assign LUT_2[41291] = 32'b11111111111111101100011001111000;
assign LUT_2[41292] = 32'b11111111111111100101000110001011;
assign LUT_2[41293] = 32'b11111111111111100001111110100100;
assign LUT_2[41294] = 32'b11111111111111101011111111000111;
assign LUT_2[41295] = 32'b11111111111111101000110111100000;
assign LUT_2[41296] = 32'b11111111111111101000011011010000;
assign LUT_2[41297] = 32'b11111111111111100101010011101001;
assign LUT_2[41298] = 32'b11111111111111101111010100001100;
assign LUT_2[41299] = 32'b11111111111111101100001100100101;
assign LUT_2[41300] = 32'b11111111111111100100111000111000;
assign LUT_2[41301] = 32'b11111111111111100001110001010001;
assign LUT_2[41302] = 32'b11111111111111101011110001110100;
assign LUT_2[41303] = 32'b11111111111111101000101010001101;
assign LUT_2[41304] = 32'b11111111111111100011001100101101;
assign LUT_2[41305] = 32'b11111111111111100000000101000110;
assign LUT_2[41306] = 32'b11111111111111101010000101101001;
assign LUT_2[41307] = 32'b11111111111111100110111110000010;
assign LUT_2[41308] = 32'b11111111111111011111101010010101;
assign LUT_2[41309] = 32'b11111111111111011100100010101110;
assign LUT_2[41310] = 32'b11111111111111100110100011010001;
assign LUT_2[41311] = 32'b11111111111111100011011011101010;
assign LUT_2[41312] = 32'b11111111111111101110010010101111;
assign LUT_2[41313] = 32'b11111111111111101011001011001000;
assign LUT_2[41314] = 32'b11111111111111110101001011101011;
assign LUT_2[41315] = 32'b11111111111111110010000100000100;
assign LUT_2[41316] = 32'b11111111111111101010110000010111;
assign LUT_2[41317] = 32'b11111111111111100111101000110000;
assign LUT_2[41318] = 32'b11111111111111110001101001010011;
assign LUT_2[41319] = 32'b11111111111111101110100001101100;
assign LUT_2[41320] = 32'b11111111111111101001000100001100;
assign LUT_2[41321] = 32'b11111111111111100101111100100101;
assign LUT_2[41322] = 32'b11111111111111101111111101001000;
assign LUT_2[41323] = 32'b11111111111111101100110101100001;
assign LUT_2[41324] = 32'b11111111111111100101100001110100;
assign LUT_2[41325] = 32'b11111111111111100010011010001101;
assign LUT_2[41326] = 32'b11111111111111101100011010110000;
assign LUT_2[41327] = 32'b11111111111111101001010011001001;
assign LUT_2[41328] = 32'b11111111111111101000110110111001;
assign LUT_2[41329] = 32'b11111111111111100101101111010010;
assign LUT_2[41330] = 32'b11111111111111101111101111110101;
assign LUT_2[41331] = 32'b11111111111111101100101000001110;
assign LUT_2[41332] = 32'b11111111111111100101010100100001;
assign LUT_2[41333] = 32'b11111111111111100010001100111010;
assign LUT_2[41334] = 32'b11111111111111101100001101011101;
assign LUT_2[41335] = 32'b11111111111111101001000101110110;
assign LUT_2[41336] = 32'b11111111111111100011101000010110;
assign LUT_2[41337] = 32'b11111111111111100000100000101111;
assign LUT_2[41338] = 32'b11111111111111101010100001010010;
assign LUT_2[41339] = 32'b11111111111111100111011001101011;
assign LUT_2[41340] = 32'b11111111111111100000000101111110;
assign LUT_2[41341] = 32'b11111111111111011100111110010111;
assign LUT_2[41342] = 32'b11111111111111100110111110111010;
assign LUT_2[41343] = 32'b11111111111111100011110111010011;
assign LUT_2[41344] = 32'b11111111111111111010000010110010;
assign LUT_2[41345] = 32'b11111111111111110110111011001011;
assign LUT_2[41346] = 32'b00000000000000000000111011101110;
assign LUT_2[41347] = 32'b11111111111111111101110100000111;
assign LUT_2[41348] = 32'b11111111111111110110100000011010;
assign LUT_2[41349] = 32'b11111111111111110011011000110011;
assign LUT_2[41350] = 32'b11111111111111111101011001010110;
assign LUT_2[41351] = 32'b11111111111111111010010001101111;
assign LUT_2[41352] = 32'b11111111111111110100110100001111;
assign LUT_2[41353] = 32'b11111111111111110001101100101000;
assign LUT_2[41354] = 32'b11111111111111111011101101001011;
assign LUT_2[41355] = 32'b11111111111111111000100101100100;
assign LUT_2[41356] = 32'b11111111111111110001010001110111;
assign LUT_2[41357] = 32'b11111111111111101110001010010000;
assign LUT_2[41358] = 32'b11111111111111111000001010110011;
assign LUT_2[41359] = 32'b11111111111111110101000011001100;
assign LUT_2[41360] = 32'b11111111111111110100100110111100;
assign LUT_2[41361] = 32'b11111111111111110001011111010101;
assign LUT_2[41362] = 32'b11111111111111111011011111111000;
assign LUT_2[41363] = 32'b11111111111111111000011000010001;
assign LUT_2[41364] = 32'b11111111111111110001000100100100;
assign LUT_2[41365] = 32'b11111111111111101101111100111101;
assign LUT_2[41366] = 32'b11111111111111110111111101100000;
assign LUT_2[41367] = 32'b11111111111111110100110101111001;
assign LUT_2[41368] = 32'b11111111111111101111011000011001;
assign LUT_2[41369] = 32'b11111111111111101100010000110010;
assign LUT_2[41370] = 32'b11111111111111110110010001010101;
assign LUT_2[41371] = 32'b11111111111111110011001001101110;
assign LUT_2[41372] = 32'b11111111111111101011110110000001;
assign LUT_2[41373] = 32'b11111111111111101000101110011010;
assign LUT_2[41374] = 32'b11111111111111110010101110111101;
assign LUT_2[41375] = 32'b11111111111111101111100111010110;
assign LUT_2[41376] = 32'b11111111111111111010011110011011;
assign LUT_2[41377] = 32'b11111111111111110111010110110100;
assign LUT_2[41378] = 32'b00000000000000000001010111010111;
assign LUT_2[41379] = 32'b11111111111111111110001111110000;
assign LUT_2[41380] = 32'b11111111111111110110111100000011;
assign LUT_2[41381] = 32'b11111111111111110011110100011100;
assign LUT_2[41382] = 32'b11111111111111111101110100111111;
assign LUT_2[41383] = 32'b11111111111111111010101101011000;
assign LUT_2[41384] = 32'b11111111111111110101001111111000;
assign LUT_2[41385] = 32'b11111111111111110010001000010001;
assign LUT_2[41386] = 32'b11111111111111111100001000110100;
assign LUT_2[41387] = 32'b11111111111111111001000001001101;
assign LUT_2[41388] = 32'b11111111111111110001101101100000;
assign LUT_2[41389] = 32'b11111111111111101110100101111001;
assign LUT_2[41390] = 32'b11111111111111111000100110011100;
assign LUT_2[41391] = 32'b11111111111111110101011110110101;
assign LUT_2[41392] = 32'b11111111111111110101000010100101;
assign LUT_2[41393] = 32'b11111111111111110001111010111110;
assign LUT_2[41394] = 32'b11111111111111111011111011100001;
assign LUT_2[41395] = 32'b11111111111111111000110011111010;
assign LUT_2[41396] = 32'b11111111111111110001100000001101;
assign LUT_2[41397] = 32'b11111111111111101110011000100110;
assign LUT_2[41398] = 32'b11111111111111111000011001001001;
assign LUT_2[41399] = 32'b11111111111111110101010001100010;
assign LUT_2[41400] = 32'b11111111111111101111110100000010;
assign LUT_2[41401] = 32'b11111111111111101100101100011011;
assign LUT_2[41402] = 32'b11111111111111110110101100111110;
assign LUT_2[41403] = 32'b11111111111111110011100101010111;
assign LUT_2[41404] = 32'b11111111111111101100010001101010;
assign LUT_2[41405] = 32'b11111111111111101001001010000011;
assign LUT_2[41406] = 32'b11111111111111110011001010100110;
assign LUT_2[41407] = 32'b11111111111111110000000010111111;
assign LUT_2[41408] = 32'b11111111111111110010001011010101;
assign LUT_2[41409] = 32'b11111111111111101111000011101110;
assign LUT_2[41410] = 32'b11111111111111111001000100010001;
assign LUT_2[41411] = 32'b11111111111111110101111100101010;
assign LUT_2[41412] = 32'b11111111111111101110101000111101;
assign LUT_2[41413] = 32'b11111111111111101011100001010110;
assign LUT_2[41414] = 32'b11111111111111110101100001111001;
assign LUT_2[41415] = 32'b11111111111111110010011010010010;
assign LUT_2[41416] = 32'b11111111111111101100111100110010;
assign LUT_2[41417] = 32'b11111111111111101001110101001011;
assign LUT_2[41418] = 32'b11111111111111110011110101101110;
assign LUT_2[41419] = 32'b11111111111111110000101110000111;
assign LUT_2[41420] = 32'b11111111111111101001011010011010;
assign LUT_2[41421] = 32'b11111111111111100110010010110011;
assign LUT_2[41422] = 32'b11111111111111110000010011010110;
assign LUT_2[41423] = 32'b11111111111111101101001011101111;
assign LUT_2[41424] = 32'b11111111111111101100101111011111;
assign LUT_2[41425] = 32'b11111111111111101001100111111000;
assign LUT_2[41426] = 32'b11111111111111110011101000011011;
assign LUT_2[41427] = 32'b11111111111111110000100000110100;
assign LUT_2[41428] = 32'b11111111111111101001001101000111;
assign LUT_2[41429] = 32'b11111111111111100110000101100000;
assign LUT_2[41430] = 32'b11111111111111110000000110000011;
assign LUT_2[41431] = 32'b11111111111111101100111110011100;
assign LUT_2[41432] = 32'b11111111111111100111100000111100;
assign LUT_2[41433] = 32'b11111111111111100100011001010101;
assign LUT_2[41434] = 32'b11111111111111101110011001111000;
assign LUT_2[41435] = 32'b11111111111111101011010010010001;
assign LUT_2[41436] = 32'b11111111111111100011111110100100;
assign LUT_2[41437] = 32'b11111111111111100000110110111101;
assign LUT_2[41438] = 32'b11111111111111101010110111100000;
assign LUT_2[41439] = 32'b11111111111111100111101111111001;
assign LUT_2[41440] = 32'b11111111111111110010100110111110;
assign LUT_2[41441] = 32'b11111111111111101111011111010111;
assign LUT_2[41442] = 32'b11111111111111111001011111111010;
assign LUT_2[41443] = 32'b11111111111111110110011000010011;
assign LUT_2[41444] = 32'b11111111111111101111000100100110;
assign LUT_2[41445] = 32'b11111111111111101011111100111111;
assign LUT_2[41446] = 32'b11111111111111110101111101100010;
assign LUT_2[41447] = 32'b11111111111111110010110101111011;
assign LUT_2[41448] = 32'b11111111111111101101011000011011;
assign LUT_2[41449] = 32'b11111111111111101010010000110100;
assign LUT_2[41450] = 32'b11111111111111110100010001010111;
assign LUT_2[41451] = 32'b11111111111111110001001001110000;
assign LUT_2[41452] = 32'b11111111111111101001110110000011;
assign LUT_2[41453] = 32'b11111111111111100110101110011100;
assign LUT_2[41454] = 32'b11111111111111110000101110111111;
assign LUT_2[41455] = 32'b11111111111111101101100111011000;
assign LUT_2[41456] = 32'b11111111111111101101001011001000;
assign LUT_2[41457] = 32'b11111111111111101010000011100001;
assign LUT_2[41458] = 32'b11111111111111110100000100000100;
assign LUT_2[41459] = 32'b11111111111111110000111100011101;
assign LUT_2[41460] = 32'b11111111111111101001101000110000;
assign LUT_2[41461] = 32'b11111111111111100110100001001001;
assign LUT_2[41462] = 32'b11111111111111110000100001101100;
assign LUT_2[41463] = 32'b11111111111111101101011010000101;
assign LUT_2[41464] = 32'b11111111111111100111111100100101;
assign LUT_2[41465] = 32'b11111111111111100100110100111110;
assign LUT_2[41466] = 32'b11111111111111101110110101100001;
assign LUT_2[41467] = 32'b11111111111111101011101101111010;
assign LUT_2[41468] = 32'b11111111111111100100011010001101;
assign LUT_2[41469] = 32'b11111111111111100001010010100110;
assign LUT_2[41470] = 32'b11111111111111101011010011001001;
assign LUT_2[41471] = 32'b11111111111111101000001011100010;
assign LUT_2[41472] = 32'b11111111111111110110100001101111;
assign LUT_2[41473] = 32'b11111111111111110011011010001000;
assign LUT_2[41474] = 32'b11111111111111111101011010101011;
assign LUT_2[41475] = 32'b11111111111111111010010011000100;
assign LUT_2[41476] = 32'b11111111111111110010111111010111;
assign LUT_2[41477] = 32'b11111111111111101111110111110000;
assign LUT_2[41478] = 32'b11111111111111111001111000010011;
assign LUT_2[41479] = 32'b11111111111111110110110000101100;
assign LUT_2[41480] = 32'b11111111111111110001010011001100;
assign LUT_2[41481] = 32'b11111111111111101110001011100101;
assign LUT_2[41482] = 32'b11111111111111111000001100001000;
assign LUT_2[41483] = 32'b11111111111111110101000100100001;
assign LUT_2[41484] = 32'b11111111111111101101110000110100;
assign LUT_2[41485] = 32'b11111111111111101010101001001101;
assign LUT_2[41486] = 32'b11111111111111110100101001110000;
assign LUT_2[41487] = 32'b11111111111111110001100010001001;
assign LUT_2[41488] = 32'b11111111111111110001000101111001;
assign LUT_2[41489] = 32'b11111111111111101101111110010010;
assign LUT_2[41490] = 32'b11111111111111110111111110110101;
assign LUT_2[41491] = 32'b11111111111111110100110111001110;
assign LUT_2[41492] = 32'b11111111111111101101100011100001;
assign LUT_2[41493] = 32'b11111111111111101010011011111010;
assign LUT_2[41494] = 32'b11111111111111110100011100011101;
assign LUT_2[41495] = 32'b11111111111111110001010100110110;
assign LUT_2[41496] = 32'b11111111111111101011110111010110;
assign LUT_2[41497] = 32'b11111111111111101000101111101111;
assign LUT_2[41498] = 32'b11111111111111110010110000010010;
assign LUT_2[41499] = 32'b11111111111111101111101000101011;
assign LUT_2[41500] = 32'b11111111111111101000010100111110;
assign LUT_2[41501] = 32'b11111111111111100101001101010111;
assign LUT_2[41502] = 32'b11111111111111101111001101111010;
assign LUT_2[41503] = 32'b11111111111111101100000110010011;
assign LUT_2[41504] = 32'b11111111111111110110111101011000;
assign LUT_2[41505] = 32'b11111111111111110011110101110001;
assign LUT_2[41506] = 32'b11111111111111111101110110010100;
assign LUT_2[41507] = 32'b11111111111111111010101110101101;
assign LUT_2[41508] = 32'b11111111111111110011011011000000;
assign LUT_2[41509] = 32'b11111111111111110000010011011001;
assign LUT_2[41510] = 32'b11111111111111111010010011111100;
assign LUT_2[41511] = 32'b11111111111111110111001100010101;
assign LUT_2[41512] = 32'b11111111111111110001101110110101;
assign LUT_2[41513] = 32'b11111111111111101110100111001110;
assign LUT_2[41514] = 32'b11111111111111111000100111110001;
assign LUT_2[41515] = 32'b11111111111111110101100000001010;
assign LUT_2[41516] = 32'b11111111111111101110001100011101;
assign LUT_2[41517] = 32'b11111111111111101011000100110110;
assign LUT_2[41518] = 32'b11111111111111110101000101011001;
assign LUT_2[41519] = 32'b11111111111111110001111101110010;
assign LUT_2[41520] = 32'b11111111111111110001100001100010;
assign LUT_2[41521] = 32'b11111111111111101110011001111011;
assign LUT_2[41522] = 32'b11111111111111111000011010011110;
assign LUT_2[41523] = 32'b11111111111111110101010010110111;
assign LUT_2[41524] = 32'b11111111111111101101111111001010;
assign LUT_2[41525] = 32'b11111111111111101010110111100011;
assign LUT_2[41526] = 32'b11111111111111110100111000000110;
assign LUT_2[41527] = 32'b11111111111111110001110000011111;
assign LUT_2[41528] = 32'b11111111111111101100010010111111;
assign LUT_2[41529] = 32'b11111111111111101001001011011000;
assign LUT_2[41530] = 32'b11111111111111110011001011111011;
assign LUT_2[41531] = 32'b11111111111111110000000100010100;
assign LUT_2[41532] = 32'b11111111111111101000110000100111;
assign LUT_2[41533] = 32'b11111111111111100101101001000000;
assign LUT_2[41534] = 32'b11111111111111101111101001100011;
assign LUT_2[41535] = 32'b11111111111111101100100001111100;
assign LUT_2[41536] = 32'b11111111111111101110101010010010;
assign LUT_2[41537] = 32'b11111111111111101011100010101011;
assign LUT_2[41538] = 32'b11111111111111110101100011001110;
assign LUT_2[41539] = 32'b11111111111111110010011011100111;
assign LUT_2[41540] = 32'b11111111111111101011000111111010;
assign LUT_2[41541] = 32'b11111111111111101000000000010011;
assign LUT_2[41542] = 32'b11111111111111110010000000110110;
assign LUT_2[41543] = 32'b11111111111111101110111001001111;
assign LUT_2[41544] = 32'b11111111111111101001011011101111;
assign LUT_2[41545] = 32'b11111111111111100110010100001000;
assign LUT_2[41546] = 32'b11111111111111110000010100101011;
assign LUT_2[41547] = 32'b11111111111111101101001101000100;
assign LUT_2[41548] = 32'b11111111111111100101111001010111;
assign LUT_2[41549] = 32'b11111111111111100010110001110000;
assign LUT_2[41550] = 32'b11111111111111101100110010010011;
assign LUT_2[41551] = 32'b11111111111111101001101010101100;
assign LUT_2[41552] = 32'b11111111111111101001001110011100;
assign LUT_2[41553] = 32'b11111111111111100110000110110101;
assign LUT_2[41554] = 32'b11111111111111110000000111011000;
assign LUT_2[41555] = 32'b11111111111111101100111111110001;
assign LUT_2[41556] = 32'b11111111111111100101101100000100;
assign LUT_2[41557] = 32'b11111111111111100010100100011101;
assign LUT_2[41558] = 32'b11111111111111101100100101000000;
assign LUT_2[41559] = 32'b11111111111111101001011101011001;
assign LUT_2[41560] = 32'b11111111111111100011111111111001;
assign LUT_2[41561] = 32'b11111111111111100000111000010010;
assign LUT_2[41562] = 32'b11111111111111101010111000110101;
assign LUT_2[41563] = 32'b11111111111111100111110001001110;
assign LUT_2[41564] = 32'b11111111111111100000011101100001;
assign LUT_2[41565] = 32'b11111111111111011101010101111010;
assign LUT_2[41566] = 32'b11111111111111100111010110011101;
assign LUT_2[41567] = 32'b11111111111111100100001110110110;
assign LUT_2[41568] = 32'b11111111111111101111000101111011;
assign LUT_2[41569] = 32'b11111111111111101011111110010100;
assign LUT_2[41570] = 32'b11111111111111110101111110110111;
assign LUT_2[41571] = 32'b11111111111111110010110111010000;
assign LUT_2[41572] = 32'b11111111111111101011100011100011;
assign LUT_2[41573] = 32'b11111111111111101000011011111100;
assign LUT_2[41574] = 32'b11111111111111110010011100011111;
assign LUT_2[41575] = 32'b11111111111111101111010100111000;
assign LUT_2[41576] = 32'b11111111111111101001110111011000;
assign LUT_2[41577] = 32'b11111111111111100110101111110001;
assign LUT_2[41578] = 32'b11111111111111110000110000010100;
assign LUT_2[41579] = 32'b11111111111111101101101000101101;
assign LUT_2[41580] = 32'b11111111111111100110010101000000;
assign LUT_2[41581] = 32'b11111111111111100011001101011001;
assign LUT_2[41582] = 32'b11111111111111101101001101111100;
assign LUT_2[41583] = 32'b11111111111111101010000110010101;
assign LUT_2[41584] = 32'b11111111111111101001101010000101;
assign LUT_2[41585] = 32'b11111111111111100110100010011110;
assign LUT_2[41586] = 32'b11111111111111110000100011000001;
assign LUT_2[41587] = 32'b11111111111111101101011011011010;
assign LUT_2[41588] = 32'b11111111111111100110000111101101;
assign LUT_2[41589] = 32'b11111111111111100011000000000110;
assign LUT_2[41590] = 32'b11111111111111101101000000101001;
assign LUT_2[41591] = 32'b11111111111111101001111001000010;
assign LUT_2[41592] = 32'b11111111111111100100011011100010;
assign LUT_2[41593] = 32'b11111111111111100001010011111011;
assign LUT_2[41594] = 32'b11111111111111101011010100011110;
assign LUT_2[41595] = 32'b11111111111111101000001100110111;
assign LUT_2[41596] = 32'b11111111111111100000111001001010;
assign LUT_2[41597] = 32'b11111111111111011101110001100011;
assign LUT_2[41598] = 32'b11111111111111100111110010000110;
assign LUT_2[41599] = 32'b11111111111111100100101010011111;
assign LUT_2[41600] = 32'b11111111111111111010110101111110;
assign LUT_2[41601] = 32'b11111111111111110111101110010111;
assign LUT_2[41602] = 32'b00000000000000000001101110111010;
assign LUT_2[41603] = 32'b11111111111111111110100111010011;
assign LUT_2[41604] = 32'b11111111111111110111010011100110;
assign LUT_2[41605] = 32'b11111111111111110100001011111111;
assign LUT_2[41606] = 32'b11111111111111111110001100100010;
assign LUT_2[41607] = 32'b11111111111111111011000100111011;
assign LUT_2[41608] = 32'b11111111111111110101100111011011;
assign LUT_2[41609] = 32'b11111111111111110010011111110100;
assign LUT_2[41610] = 32'b11111111111111111100100000010111;
assign LUT_2[41611] = 32'b11111111111111111001011000110000;
assign LUT_2[41612] = 32'b11111111111111110010000101000011;
assign LUT_2[41613] = 32'b11111111111111101110111101011100;
assign LUT_2[41614] = 32'b11111111111111111000111101111111;
assign LUT_2[41615] = 32'b11111111111111110101110110011000;
assign LUT_2[41616] = 32'b11111111111111110101011010001000;
assign LUT_2[41617] = 32'b11111111111111110010010010100001;
assign LUT_2[41618] = 32'b11111111111111111100010011000100;
assign LUT_2[41619] = 32'b11111111111111111001001011011101;
assign LUT_2[41620] = 32'b11111111111111110001110111110000;
assign LUT_2[41621] = 32'b11111111111111101110110000001001;
assign LUT_2[41622] = 32'b11111111111111111000110000101100;
assign LUT_2[41623] = 32'b11111111111111110101101001000101;
assign LUT_2[41624] = 32'b11111111111111110000001011100101;
assign LUT_2[41625] = 32'b11111111111111101101000011111110;
assign LUT_2[41626] = 32'b11111111111111110111000100100001;
assign LUT_2[41627] = 32'b11111111111111110011111100111010;
assign LUT_2[41628] = 32'b11111111111111101100101001001101;
assign LUT_2[41629] = 32'b11111111111111101001100001100110;
assign LUT_2[41630] = 32'b11111111111111110011100010001001;
assign LUT_2[41631] = 32'b11111111111111110000011010100010;
assign LUT_2[41632] = 32'b11111111111111111011010001100111;
assign LUT_2[41633] = 32'b11111111111111111000001010000000;
assign LUT_2[41634] = 32'b00000000000000000010001010100011;
assign LUT_2[41635] = 32'b11111111111111111111000010111100;
assign LUT_2[41636] = 32'b11111111111111110111101111001111;
assign LUT_2[41637] = 32'b11111111111111110100100111101000;
assign LUT_2[41638] = 32'b11111111111111111110101000001011;
assign LUT_2[41639] = 32'b11111111111111111011100000100100;
assign LUT_2[41640] = 32'b11111111111111110110000011000100;
assign LUT_2[41641] = 32'b11111111111111110010111011011101;
assign LUT_2[41642] = 32'b11111111111111111100111100000000;
assign LUT_2[41643] = 32'b11111111111111111001110100011001;
assign LUT_2[41644] = 32'b11111111111111110010100000101100;
assign LUT_2[41645] = 32'b11111111111111101111011001000101;
assign LUT_2[41646] = 32'b11111111111111111001011001101000;
assign LUT_2[41647] = 32'b11111111111111110110010010000001;
assign LUT_2[41648] = 32'b11111111111111110101110101110001;
assign LUT_2[41649] = 32'b11111111111111110010101110001010;
assign LUT_2[41650] = 32'b11111111111111111100101110101101;
assign LUT_2[41651] = 32'b11111111111111111001100111000110;
assign LUT_2[41652] = 32'b11111111111111110010010011011001;
assign LUT_2[41653] = 32'b11111111111111101111001011110010;
assign LUT_2[41654] = 32'b11111111111111111001001100010101;
assign LUT_2[41655] = 32'b11111111111111110110000100101110;
assign LUT_2[41656] = 32'b11111111111111110000100111001110;
assign LUT_2[41657] = 32'b11111111111111101101011111100111;
assign LUT_2[41658] = 32'b11111111111111110111100000001010;
assign LUT_2[41659] = 32'b11111111111111110100011000100011;
assign LUT_2[41660] = 32'b11111111111111101101000100110110;
assign LUT_2[41661] = 32'b11111111111111101001111101001111;
assign LUT_2[41662] = 32'b11111111111111110011111101110010;
assign LUT_2[41663] = 32'b11111111111111110000110110001011;
assign LUT_2[41664] = 32'b11111111111111110010111110100001;
assign LUT_2[41665] = 32'b11111111111111101111110110111010;
assign LUT_2[41666] = 32'b11111111111111111001110111011101;
assign LUT_2[41667] = 32'b11111111111111110110101111110110;
assign LUT_2[41668] = 32'b11111111111111101111011100001001;
assign LUT_2[41669] = 32'b11111111111111101100010100100010;
assign LUT_2[41670] = 32'b11111111111111110110010101000101;
assign LUT_2[41671] = 32'b11111111111111110011001101011110;
assign LUT_2[41672] = 32'b11111111111111101101101111111110;
assign LUT_2[41673] = 32'b11111111111111101010101000010111;
assign LUT_2[41674] = 32'b11111111111111110100101000111010;
assign LUT_2[41675] = 32'b11111111111111110001100001010011;
assign LUT_2[41676] = 32'b11111111111111101010001101100110;
assign LUT_2[41677] = 32'b11111111111111100111000101111111;
assign LUT_2[41678] = 32'b11111111111111110001000110100010;
assign LUT_2[41679] = 32'b11111111111111101101111110111011;
assign LUT_2[41680] = 32'b11111111111111101101100010101011;
assign LUT_2[41681] = 32'b11111111111111101010011011000100;
assign LUT_2[41682] = 32'b11111111111111110100011011100111;
assign LUT_2[41683] = 32'b11111111111111110001010100000000;
assign LUT_2[41684] = 32'b11111111111111101010000000010011;
assign LUT_2[41685] = 32'b11111111111111100110111000101100;
assign LUT_2[41686] = 32'b11111111111111110000111001001111;
assign LUT_2[41687] = 32'b11111111111111101101110001101000;
assign LUT_2[41688] = 32'b11111111111111101000010100001000;
assign LUT_2[41689] = 32'b11111111111111100101001100100001;
assign LUT_2[41690] = 32'b11111111111111101111001101000100;
assign LUT_2[41691] = 32'b11111111111111101100000101011101;
assign LUT_2[41692] = 32'b11111111111111100100110001110000;
assign LUT_2[41693] = 32'b11111111111111100001101010001001;
assign LUT_2[41694] = 32'b11111111111111101011101010101100;
assign LUT_2[41695] = 32'b11111111111111101000100011000101;
assign LUT_2[41696] = 32'b11111111111111110011011010001010;
assign LUT_2[41697] = 32'b11111111111111110000010010100011;
assign LUT_2[41698] = 32'b11111111111111111010010011000110;
assign LUT_2[41699] = 32'b11111111111111110111001011011111;
assign LUT_2[41700] = 32'b11111111111111101111110111110010;
assign LUT_2[41701] = 32'b11111111111111101100110000001011;
assign LUT_2[41702] = 32'b11111111111111110110110000101110;
assign LUT_2[41703] = 32'b11111111111111110011101001000111;
assign LUT_2[41704] = 32'b11111111111111101110001011100111;
assign LUT_2[41705] = 32'b11111111111111101011000100000000;
assign LUT_2[41706] = 32'b11111111111111110101000100100011;
assign LUT_2[41707] = 32'b11111111111111110001111100111100;
assign LUT_2[41708] = 32'b11111111111111101010101001001111;
assign LUT_2[41709] = 32'b11111111111111100111100001101000;
assign LUT_2[41710] = 32'b11111111111111110001100010001011;
assign LUT_2[41711] = 32'b11111111111111101110011010100100;
assign LUT_2[41712] = 32'b11111111111111101101111110010100;
assign LUT_2[41713] = 32'b11111111111111101010110110101101;
assign LUT_2[41714] = 32'b11111111111111110100110111010000;
assign LUT_2[41715] = 32'b11111111111111110001101111101001;
assign LUT_2[41716] = 32'b11111111111111101010011011111100;
assign LUT_2[41717] = 32'b11111111111111100111010100010101;
assign LUT_2[41718] = 32'b11111111111111110001010100111000;
assign LUT_2[41719] = 32'b11111111111111101110001101010001;
assign LUT_2[41720] = 32'b11111111111111101000101111110001;
assign LUT_2[41721] = 32'b11111111111111100101101000001010;
assign LUT_2[41722] = 32'b11111111111111101111101000101101;
assign LUT_2[41723] = 32'b11111111111111101100100001000110;
assign LUT_2[41724] = 32'b11111111111111100101001101011001;
assign LUT_2[41725] = 32'b11111111111111100010000101110010;
assign LUT_2[41726] = 32'b11111111111111101100000110010101;
assign LUT_2[41727] = 32'b11111111111111101000111110101110;
assign LUT_2[41728] = 32'b11111111111111111010100000010101;
assign LUT_2[41729] = 32'b11111111111111110111011000101110;
assign LUT_2[41730] = 32'b00000000000000000001011001010001;
assign LUT_2[41731] = 32'b11111111111111111110010001101010;
assign LUT_2[41732] = 32'b11111111111111110110111101111101;
assign LUT_2[41733] = 32'b11111111111111110011110110010110;
assign LUT_2[41734] = 32'b11111111111111111101110110111001;
assign LUT_2[41735] = 32'b11111111111111111010101111010010;
assign LUT_2[41736] = 32'b11111111111111110101010001110010;
assign LUT_2[41737] = 32'b11111111111111110010001010001011;
assign LUT_2[41738] = 32'b11111111111111111100001010101110;
assign LUT_2[41739] = 32'b11111111111111111001000011000111;
assign LUT_2[41740] = 32'b11111111111111110001101111011010;
assign LUT_2[41741] = 32'b11111111111111101110100111110011;
assign LUT_2[41742] = 32'b11111111111111111000101000010110;
assign LUT_2[41743] = 32'b11111111111111110101100000101111;
assign LUT_2[41744] = 32'b11111111111111110101000100011111;
assign LUT_2[41745] = 32'b11111111111111110001111100111000;
assign LUT_2[41746] = 32'b11111111111111111011111101011011;
assign LUT_2[41747] = 32'b11111111111111111000110101110100;
assign LUT_2[41748] = 32'b11111111111111110001100010000111;
assign LUT_2[41749] = 32'b11111111111111101110011010100000;
assign LUT_2[41750] = 32'b11111111111111111000011011000011;
assign LUT_2[41751] = 32'b11111111111111110101010011011100;
assign LUT_2[41752] = 32'b11111111111111101111110101111100;
assign LUT_2[41753] = 32'b11111111111111101100101110010101;
assign LUT_2[41754] = 32'b11111111111111110110101110111000;
assign LUT_2[41755] = 32'b11111111111111110011100111010001;
assign LUT_2[41756] = 32'b11111111111111101100010011100100;
assign LUT_2[41757] = 32'b11111111111111101001001011111101;
assign LUT_2[41758] = 32'b11111111111111110011001100100000;
assign LUT_2[41759] = 32'b11111111111111110000000100111001;
assign LUT_2[41760] = 32'b11111111111111111010111011111110;
assign LUT_2[41761] = 32'b11111111111111110111110100010111;
assign LUT_2[41762] = 32'b00000000000000000001110100111010;
assign LUT_2[41763] = 32'b11111111111111111110101101010011;
assign LUT_2[41764] = 32'b11111111111111110111011001100110;
assign LUT_2[41765] = 32'b11111111111111110100010001111111;
assign LUT_2[41766] = 32'b11111111111111111110010010100010;
assign LUT_2[41767] = 32'b11111111111111111011001010111011;
assign LUT_2[41768] = 32'b11111111111111110101101101011011;
assign LUT_2[41769] = 32'b11111111111111110010100101110100;
assign LUT_2[41770] = 32'b11111111111111111100100110010111;
assign LUT_2[41771] = 32'b11111111111111111001011110110000;
assign LUT_2[41772] = 32'b11111111111111110010001011000011;
assign LUT_2[41773] = 32'b11111111111111101111000011011100;
assign LUT_2[41774] = 32'b11111111111111111001000011111111;
assign LUT_2[41775] = 32'b11111111111111110101111100011000;
assign LUT_2[41776] = 32'b11111111111111110101100000001000;
assign LUT_2[41777] = 32'b11111111111111110010011000100001;
assign LUT_2[41778] = 32'b11111111111111111100011001000100;
assign LUT_2[41779] = 32'b11111111111111111001010001011101;
assign LUT_2[41780] = 32'b11111111111111110001111101110000;
assign LUT_2[41781] = 32'b11111111111111101110110110001001;
assign LUT_2[41782] = 32'b11111111111111111000110110101100;
assign LUT_2[41783] = 32'b11111111111111110101101111000101;
assign LUT_2[41784] = 32'b11111111111111110000010001100101;
assign LUT_2[41785] = 32'b11111111111111101101001001111110;
assign LUT_2[41786] = 32'b11111111111111110111001010100001;
assign LUT_2[41787] = 32'b11111111111111110100000010111010;
assign LUT_2[41788] = 32'b11111111111111101100101111001101;
assign LUT_2[41789] = 32'b11111111111111101001100111100110;
assign LUT_2[41790] = 32'b11111111111111110011101000001001;
assign LUT_2[41791] = 32'b11111111111111110000100000100010;
assign LUT_2[41792] = 32'b11111111111111110010101000111000;
assign LUT_2[41793] = 32'b11111111111111101111100001010001;
assign LUT_2[41794] = 32'b11111111111111111001100001110100;
assign LUT_2[41795] = 32'b11111111111111110110011010001101;
assign LUT_2[41796] = 32'b11111111111111101111000110100000;
assign LUT_2[41797] = 32'b11111111111111101011111110111001;
assign LUT_2[41798] = 32'b11111111111111110101111111011100;
assign LUT_2[41799] = 32'b11111111111111110010110111110101;
assign LUT_2[41800] = 32'b11111111111111101101011010010101;
assign LUT_2[41801] = 32'b11111111111111101010010010101110;
assign LUT_2[41802] = 32'b11111111111111110100010011010001;
assign LUT_2[41803] = 32'b11111111111111110001001011101010;
assign LUT_2[41804] = 32'b11111111111111101001110111111101;
assign LUT_2[41805] = 32'b11111111111111100110110000010110;
assign LUT_2[41806] = 32'b11111111111111110000110000111001;
assign LUT_2[41807] = 32'b11111111111111101101101001010010;
assign LUT_2[41808] = 32'b11111111111111101101001101000010;
assign LUT_2[41809] = 32'b11111111111111101010000101011011;
assign LUT_2[41810] = 32'b11111111111111110100000101111110;
assign LUT_2[41811] = 32'b11111111111111110000111110010111;
assign LUT_2[41812] = 32'b11111111111111101001101010101010;
assign LUT_2[41813] = 32'b11111111111111100110100011000011;
assign LUT_2[41814] = 32'b11111111111111110000100011100110;
assign LUT_2[41815] = 32'b11111111111111101101011011111111;
assign LUT_2[41816] = 32'b11111111111111100111111110011111;
assign LUT_2[41817] = 32'b11111111111111100100110110111000;
assign LUT_2[41818] = 32'b11111111111111101110110111011011;
assign LUT_2[41819] = 32'b11111111111111101011101111110100;
assign LUT_2[41820] = 32'b11111111111111100100011100000111;
assign LUT_2[41821] = 32'b11111111111111100001010100100000;
assign LUT_2[41822] = 32'b11111111111111101011010101000011;
assign LUT_2[41823] = 32'b11111111111111101000001101011100;
assign LUT_2[41824] = 32'b11111111111111110011000100100001;
assign LUT_2[41825] = 32'b11111111111111101111111100111010;
assign LUT_2[41826] = 32'b11111111111111111001111101011101;
assign LUT_2[41827] = 32'b11111111111111110110110101110110;
assign LUT_2[41828] = 32'b11111111111111101111100010001001;
assign LUT_2[41829] = 32'b11111111111111101100011010100010;
assign LUT_2[41830] = 32'b11111111111111110110011011000101;
assign LUT_2[41831] = 32'b11111111111111110011010011011110;
assign LUT_2[41832] = 32'b11111111111111101101110101111110;
assign LUT_2[41833] = 32'b11111111111111101010101110010111;
assign LUT_2[41834] = 32'b11111111111111110100101110111010;
assign LUT_2[41835] = 32'b11111111111111110001100111010011;
assign LUT_2[41836] = 32'b11111111111111101010010011100110;
assign LUT_2[41837] = 32'b11111111111111100111001011111111;
assign LUT_2[41838] = 32'b11111111111111110001001100100010;
assign LUT_2[41839] = 32'b11111111111111101110000100111011;
assign LUT_2[41840] = 32'b11111111111111101101101000101011;
assign LUT_2[41841] = 32'b11111111111111101010100001000100;
assign LUT_2[41842] = 32'b11111111111111110100100001100111;
assign LUT_2[41843] = 32'b11111111111111110001011010000000;
assign LUT_2[41844] = 32'b11111111111111101010000110010011;
assign LUT_2[41845] = 32'b11111111111111100110111110101100;
assign LUT_2[41846] = 32'b11111111111111110000111111001111;
assign LUT_2[41847] = 32'b11111111111111101101110111101000;
assign LUT_2[41848] = 32'b11111111111111101000011010001000;
assign LUT_2[41849] = 32'b11111111111111100101010010100001;
assign LUT_2[41850] = 32'b11111111111111101111010011000100;
assign LUT_2[41851] = 32'b11111111111111101100001011011101;
assign LUT_2[41852] = 32'b11111111111111100100110111110000;
assign LUT_2[41853] = 32'b11111111111111100001110000001001;
assign LUT_2[41854] = 32'b11111111111111101011110000101100;
assign LUT_2[41855] = 32'b11111111111111101000101001000101;
assign LUT_2[41856] = 32'b11111111111111111110110100100100;
assign LUT_2[41857] = 32'b11111111111111111011101100111101;
assign LUT_2[41858] = 32'b00000000000000000101101101100000;
assign LUT_2[41859] = 32'b00000000000000000010100101111001;
assign LUT_2[41860] = 32'b11111111111111111011010010001100;
assign LUT_2[41861] = 32'b11111111111111111000001010100101;
assign LUT_2[41862] = 32'b00000000000000000010001011001000;
assign LUT_2[41863] = 32'b11111111111111111111000011100001;
assign LUT_2[41864] = 32'b11111111111111111001100110000001;
assign LUT_2[41865] = 32'b11111111111111110110011110011010;
assign LUT_2[41866] = 32'b00000000000000000000011110111101;
assign LUT_2[41867] = 32'b11111111111111111101010111010110;
assign LUT_2[41868] = 32'b11111111111111110110000011101001;
assign LUT_2[41869] = 32'b11111111111111110010111100000010;
assign LUT_2[41870] = 32'b11111111111111111100111100100101;
assign LUT_2[41871] = 32'b11111111111111111001110100111110;
assign LUT_2[41872] = 32'b11111111111111111001011000101110;
assign LUT_2[41873] = 32'b11111111111111110110010001000111;
assign LUT_2[41874] = 32'b00000000000000000000010001101010;
assign LUT_2[41875] = 32'b11111111111111111101001010000011;
assign LUT_2[41876] = 32'b11111111111111110101110110010110;
assign LUT_2[41877] = 32'b11111111111111110010101110101111;
assign LUT_2[41878] = 32'b11111111111111111100101111010010;
assign LUT_2[41879] = 32'b11111111111111111001100111101011;
assign LUT_2[41880] = 32'b11111111111111110100001010001011;
assign LUT_2[41881] = 32'b11111111111111110001000010100100;
assign LUT_2[41882] = 32'b11111111111111111011000011000111;
assign LUT_2[41883] = 32'b11111111111111110111111011100000;
assign LUT_2[41884] = 32'b11111111111111110000100111110011;
assign LUT_2[41885] = 32'b11111111111111101101100000001100;
assign LUT_2[41886] = 32'b11111111111111110111100000101111;
assign LUT_2[41887] = 32'b11111111111111110100011001001000;
assign LUT_2[41888] = 32'b11111111111111111111010000001101;
assign LUT_2[41889] = 32'b11111111111111111100001000100110;
assign LUT_2[41890] = 32'b00000000000000000110001001001001;
assign LUT_2[41891] = 32'b00000000000000000011000001100010;
assign LUT_2[41892] = 32'b11111111111111111011101101110101;
assign LUT_2[41893] = 32'b11111111111111111000100110001110;
assign LUT_2[41894] = 32'b00000000000000000010100110110001;
assign LUT_2[41895] = 32'b11111111111111111111011111001010;
assign LUT_2[41896] = 32'b11111111111111111010000001101010;
assign LUT_2[41897] = 32'b11111111111111110110111010000011;
assign LUT_2[41898] = 32'b00000000000000000000111010100110;
assign LUT_2[41899] = 32'b11111111111111111101110010111111;
assign LUT_2[41900] = 32'b11111111111111110110011111010010;
assign LUT_2[41901] = 32'b11111111111111110011010111101011;
assign LUT_2[41902] = 32'b11111111111111111101011000001110;
assign LUT_2[41903] = 32'b11111111111111111010010000100111;
assign LUT_2[41904] = 32'b11111111111111111001110100010111;
assign LUT_2[41905] = 32'b11111111111111110110101100110000;
assign LUT_2[41906] = 32'b00000000000000000000101101010011;
assign LUT_2[41907] = 32'b11111111111111111101100101101100;
assign LUT_2[41908] = 32'b11111111111111110110010001111111;
assign LUT_2[41909] = 32'b11111111111111110011001010011000;
assign LUT_2[41910] = 32'b11111111111111111101001010111011;
assign LUT_2[41911] = 32'b11111111111111111010000011010100;
assign LUT_2[41912] = 32'b11111111111111110100100101110100;
assign LUT_2[41913] = 32'b11111111111111110001011110001101;
assign LUT_2[41914] = 32'b11111111111111111011011110110000;
assign LUT_2[41915] = 32'b11111111111111111000010111001001;
assign LUT_2[41916] = 32'b11111111111111110001000011011100;
assign LUT_2[41917] = 32'b11111111111111101101111011110101;
assign LUT_2[41918] = 32'b11111111111111110111111100011000;
assign LUT_2[41919] = 32'b11111111111111110100110100110001;
assign LUT_2[41920] = 32'b11111111111111110110111101000111;
assign LUT_2[41921] = 32'b11111111111111110011110101100000;
assign LUT_2[41922] = 32'b11111111111111111101110110000011;
assign LUT_2[41923] = 32'b11111111111111111010101110011100;
assign LUT_2[41924] = 32'b11111111111111110011011010101111;
assign LUT_2[41925] = 32'b11111111111111110000010011001000;
assign LUT_2[41926] = 32'b11111111111111111010010011101011;
assign LUT_2[41927] = 32'b11111111111111110111001100000100;
assign LUT_2[41928] = 32'b11111111111111110001101110100100;
assign LUT_2[41929] = 32'b11111111111111101110100110111101;
assign LUT_2[41930] = 32'b11111111111111111000100111100000;
assign LUT_2[41931] = 32'b11111111111111110101011111111001;
assign LUT_2[41932] = 32'b11111111111111101110001100001100;
assign LUT_2[41933] = 32'b11111111111111101011000100100101;
assign LUT_2[41934] = 32'b11111111111111110101000101001000;
assign LUT_2[41935] = 32'b11111111111111110001111101100001;
assign LUT_2[41936] = 32'b11111111111111110001100001010001;
assign LUT_2[41937] = 32'b11111111111111101110011001101010;
assign LUT_2[41938] = 32'b11111111111111111000011010001101;
assign LUT_2[41939] = 32'b11111111111111110101010010100110;
assign LUT_2[41940] = 32'b11111111111111101101111110111001;
assign LUT_2[41941] = 32'b11111111111111101010110111010010;
assign LUT_2[41942] = 32'b11111111111111110100110111110101;
assign LUT_2[41943] = 32'b11111111111111110001110000001110;
assign LUT_2[41944] = 32'b11111111111111101100010010101110;
assign LUT_2[41945] = 32'b11111111111111101001001011000111;
assign LUT_2[41946] = 32'b11111111111111110011001011101010;
assign LUT_2[41947] = 32'b11111111111111110000000100000011;
assign LUT_2[41948] = 32'b11111111111111101000110000010110;
assign LUT_2[41949] = 32'b11111111111111100101101000101111;
assign LUT_2[41950] = 32'b11111111111111101111101001010010;
assign LUT_2[41951] = 32'b11111111111111101100100001101011;
assign LUT_2[41952] = 32'b11111111111111110111011000110000;
assign LUT_2[41953] = 32'b11111111111111110100010001001001;
assign LUT_2[41954] = 32'b11111111111111111110010001101100;
assign LUT_2[41955] = 32'b11111111111111111011001010000101;
assign LUT_2[41956] = 32'b11111111111111110011110110011000;
assign LUT_2[41957] = 32'b11111111111111110000101110110001;
assign LUT_2[41958] = 32'b11111111111111111010101111010100;
assign LUT_2[41959] = 32'b11111111111111110111100111101101;
assign LUT_2[41960] = 32'b11111111111111110010001010001101;
assign LUT_2[41961] = 32'b11111111111111101111000010100110;
assign LUT_2[41962] = 32'b11111111111111111001000011001001;
assign LUT_2[41963] = 32'b11111111111111110101111011100010;
assign LUT_2[41964] = 32'b11111111111111101110100111110101;
assign LUT_2[41965] = 32'b11111111111111101011100000001110;
assign LUT_2[41966] = 32'b11111111111111110101100000110001;
assign LUT_2[41967] = 32'b11111111111111110010011001001010;
assign LUT_2[41968] = 32'b11111111111111110001111100111010;
assign LUT_2[41969] = 32'b11111111111111101110110101010011;
assign LUT_2[41970] = 32'b11111111111111111000110101110110;
assign LUT_2[41971] = 32'b11111111111111110101101110001111;
assign LUT_2[41972] = 32'b11111111111111101110011010100010;
assign LUT_2[41973] = 32'b11111111111111101011010010111011;
assign LUT_2[41974] = 32'b11111111111111110101010011011110;
assign LUT_2[41975] = 32'b11111111111111110010001011110111;
assign LUT_2[41976] = 32'b11111111111111101100101110010111;
assign LUT_2[41977] = 32'b11111111111111101001100110110000;
assign LUT_2[41978] = 32'b11111111111111110011100111010011;
assign LUT_2[41979] = 32'b11111111111111110000011111101100;
assign LUT_2[41980] = 32'b11111111111111101001001011111111;
assign LUT_2[41981] = 32'b11111111111111100110000100011000;
assign LUT_2[41982] = 32'b11111111111111110000000100111011;
assign LUT_2[41983] = 32'b11111111111111101100111101010100;
assign LUT_2[41984] = 32'b11111111111111111000011100000010;
assign LUT_2[41985] = 32'b11111111111111110101010100011011;
assign LUT_2[41986] = 32'b11111111111111111111010100111110;
assign LUT_2[41987] = 32'b11111111111111111100001101010111;
assign LUT_2[41988] = 32'b11111111111111110100111001101010;
assign LUT_2[41989] = 32'b11111111111111110001110010000011;
assign LUT_2[41990] = 32'b11111111111111111011110010100110;
assign LUT_2[41991] = 32'b11111111111111111000101010111111;
assign LUT_2[41992] = 32'b11111111111111110011001101011111;
assign LUT_2[41993] = 32'b11111111111111110000000101111000;
assign LUT_2[41994] = 32'b11111111111111111010000110011011;
assign LUT_2[41995] = 32'b11111111111111110110111110110100;
assign LUT_2[41996] = 32'b11111111111111101111101011000111;
assign LUT_2[41997] = 32'b11111111111111101100100011100000;
assign LUT_2[41998] = 32'b11111111111111110110100100000011;
assign LUT_2[41999] = 32'b11111111111111110011011100011100;
assign LUT_2[42000] = 32'b11111111111111110011000000001100;
assign LUT_2[42001] = 32'b11111111111111101111111000100101;
assign LUT_2[42002] = 32'b11111111111111111001111001001000;
assign LUT_2[42003] = 32'b11111111111111110110110001100001;
assign LUT_2[42004] = 32'b11111111111111101111011101110100;
assign LUT_2[42005] = 32'b11111111111111101100010110001101;
assign LUT_2[42006] = 32'b11111111111111110110010110110000;
assign LUT_2[42007] = 32'b11111111111111110011001111001001;
assign LUT_2[42008] = 32'b11111111111111101101110001101001;
assign LUT_2[42009] = 32'b11111111111111101010101010000010;
assign LUT_2[42010] = 32'b11111111111111110100101010100101;
assign LUT_2[42011] = 32'b11111111111111110001100010111110;
assign LUT_2[42012] = 32'b11111111111111101010001111010001;
assign LUT_2[42013] = 32'b11111111111111100111000111101010;
assign LUT_2[42014] = 32'b11111111111111110001001000001101;
assign LUT_2[42015] = 32'b11111111111111101110000000100110;
assign LUT_2[42016] = 32'b11111111111111111000110111101011;
assign LUT_2[42017] = 32'b11111111111111110101110000000100;
assign LUT_2[42018] = 32'b11111111111111111111110000100111;
assign LUT_2[42019] = 32'b11111111111111111100101001000000;
assign LUT_2[42020] = 32'b11111111111111110101010101010011;
assign LUT_2[42021] = 32'b11111111111111110010001101101100;
assign LUT_2[42022] = 32'b11111111111111111100001110001111;
assign LUT_2[42023] = 32'b11111111111111111001000110101000;
assign LUT_2[42024] = 32'b11111111111111110011101001001000;
assign LUT_2[42025] = 32'b11111111111111110000100001100001;
assign LUT_2[42026] = 32'b11111111111111111010100010000100;
assign LUT_2[42027] = 32'b11111111111111110111011010011101;
assign LUT_2[42028] = 32'b11111111111111110000000110110000;
assign LUT_2[42029] = 32'b11111111111111101100111111001001;
assign LUT_2[42030] = 32'b11111111111111110110111111101100;
assign LUT_2[42031] = 32'b11111111111111110011111000000101;
assign LUT_2[42032] = 32'b11111111111111110011011011110101;
assign LUT_2[42033] = 32'b11111111111111110000010100001110;
assign LUT_2[42034] = 32'b11111111111111111010010100110001;
assign LUT_2[42035] = 32'b11111111111111110111001101001010;
assign LUT_2[42036] = 32'b11111111111111101111111001011101;
assign LUT_2[42037] = 32'b11111111111111101100110001110110;
assign LUT_2[42038] = 32'b11111111111111110110110010011001;
assign LUT_2[42039] = 32'b11111111111111110011101010110010;
assign LUT_2[42040] = 32'b11111111111111101110001101010010;
assign LUT_2[42041] = 32'b11111111111111101011000101101011;
assign LUT_2[42042] = 32'b11111111111111110101000110001110;
assign LUT_2[42043] = 32'b11111111111111110001111110100111;
assign LUT_2[42044] = 32'b11111111111111101010101010111010;
assign LUT_2[42045] = 32'b11111111111111100111100011010011;
assign LUT_2[42046] = 32'b11111111111111110001100011110110;
assign LUT_2[42047] = 32'b11111111111111101110011100001111;
assign LUT_2[42048] = 32'b11111111111111110000100100100101;
assign LUT_2[42049] = 32'b11111111111111101101011100111110;
assign LUT_2[42050] = 32'b11111111111111110111011101100001;
assign LUT_2[42051] = 32'b11111111111111110100010101111010;
assign LUT_2[42052] = 32'b11111111111111101101000010001101;
assign LUT_2[42053] = 32'b11111111111111101001111010100110;
assign LUT_2[42054] = 32'b11111111111111110011111011001001;
assign LUT_2[42055] = 32'b11111111111111110000110011100010;
assign LUT_2[42056] = 32'b11111111111111101011010110000010;
assign LUT_2[42057] = 32'b11111111111111101000001110011011;
assign LUT_2[42058] = 32'b11111111111111110010001110111110;
assign LUT_2[42059] = 32'b11111111111111101111000111010111;
assign LUT_2[42060] = 32'b11111111111111100111110011101010;
assign LUT_2[42061] = 32'b11111111111111100100101100000011;
assign LUT_2[42062] = 32'b11111111111111101110101100100110;
assign LUT_2[42063] = 32'b11111111111111101011100100111111;
assign LUT_2[42064] = 32'b11111111111111101011001000101111;
assign LUT_2[42065] = 32'b11111111111111101000000001001000;
assign LUT_2[42066] = 32'b11111111111111110010000001101011;
assign LUT_2[42067] = 32'b11111111111111101110111010000100;
assign LUT_2[42068] = 32'b11111111111111100111100110010111;
assign LUT_2[42069] = 32'b11111111111111100100011110110000;
assign LUT_2[42070] = 32'b11111111111111101110011111010011;
assign LUT_2[42071] = 32'b11111111111111101011010111101100;
assign LUT_2[42072] = 32'b11111111111111100101111010001100;
assign LUT_2[42073] = 32'b11111111111111100010110010100101;
assign LUT_2[42074] = 32'b11111111111111101100110011001000;
assign LUT_2[42075] = 32'b11111111111111101001101011100001;
assign LUT_2[42076] = 32'b11111111111111100010010111110100;
assign LUT_2[42077] = 32'b11111111111111011111010000001101;
assign LUT_2[42078] = 32'b11111111111111101001010000110000;
assign LUT_2[42079] = 32'b11111111111111100110001001001001;
assign LUT_2[42080] = 32'b11111111111111110001000000001110;
assign LUT_2[42081] = 32'b11111111111111101101111000100111;
assign LUT_2[42082] = 32'b11111111111111110111111001001010;
assign LUT_2[42083] = 32'b11111111111111110100110001100011;
assign LUT_2[42084] = 32'b11111111111111101101011101110110;
assign LUT_2[42085] = 32'b11111111111111101010010110001111;
assign LUT_2[42086] = 32'b11111111111111110100010110110010;
assign LUT_2[42087] = 32'b11111111111111110001001111001011;
assign LUT_2[42088] = 32'b11111111111111101011110001101011;
assign LUT_2[42089] = 32'b11111111111111101000101010000100;
assign LUT_2[42090] = 32'b11111111111111110010101010100111;
assign LUT_2[42091] = 32'b11111111111111101111100011000000;
assign LUT_2[42092] = 32'b11111111111111101000001111010011;
assign LUT_2[42093] = 32'b11111111111111100101000111101100;
assign LUT_2[42094] = 32'b11111111111111101111001000001111;
assign LUT_2[42095] = 32'b11111111111111101100000000101000;
assign LUT_2[42096] = 32'b11111111111111101011100100011000;
assign LUT_2[42097] = 32'b11111111111111101000011100110001;
assign LUT_2[42098] = 32'b11111111111111110010011101010100;
assign LUT_2[42099] = 32'b11111111111111101111010101101101;
assign LUT_2[42100] = 32'b11111111111111101000000010000000;
assign LUT_2[42101] = 32'b11111111111111100100111010011001;
assign LUT_2[42102] = 32'b11111111111111101110111010111100;
assign LUT_2[42103] = 32'b11111111111111101011110011010101;
assign LUT_2[42104] = 32'b11111111111111100110010101110101;
assign LUT_2[42105] = 32'b11111111111111100011001110001110;
assign LUT_2[42106] = 32'b11111111111111101101001110110001;
assign LUT_2[42107] = 32'b11111111111111101010000111001010;
assign LUT_2[42108] = 32'b11111111111111100010110011011101;
assign LUT_2[42109] = 32'b11111111111111011111101011110110;
assign LUT_2[42110] = 32'b11111111111111101001101100011001;
assign LUT_2[42111] = 32'b11111111111111100110100100110010;
assign LUT_2[42112] = 32'b11111111111111111100110000010001;
assign LUT_2[42113] = 32'b11111111111111111001101000101010;
assign LUT_2[42114] = 32'b00000000000000000011101001001101;
assign LUT_2[42115] = 32'b00000000000000000000100001100110;
assign LUT_2[42116] = 32'b11111111111111111001001101111001;
assign LUT_2[42117] = 32'b11111111111111110110000110010010;
assign LUT_2[42118] = 32'b00000000000000000000000110110101;
assign LUT_2[42119] = 32'b11111111111111111100111111001110;
assign LUT_2[42120] = 32'b11111111111111110111100001101110;
assign LUT_2[42121] = 32'b11111111111111110100011010000111;
assign LUT_2[42122] = 32'b11111111111111111110011010101010;
assign LUT_2[42123] = 32'b11111111111111111011010011000011;
assign LUT_2[42124] = 32'b11111111111111110011111111010110;
assign LUT_2[42125] = 32'b11111111111111110000110111101111;
assign LUT_2[42126] = 32'b11111111111111111010111000010010;
assign LUT_2[42127] = 32'b11111111111111110111110000101011;
assign LUT_2[42128] = 32'b11111111111111110111010100011011;
assign LUT_2[42129] = 32'b11111111111111110100001100110100;
assign LUT_2[42130] = 32'b11111111111111111110001101010111;
assign LUT_2[42131] = 32'b11111111111111111011000101110000;
assign LUT_2[42132] = 32'b11111111111111110011110010000011;
assign LUT_2[42133] = 32'b11111111111111110000101010011100;
assign LUT_2[42134] = 32'b11111111111111111010101010111111;
assign LUT_2[42135] = 32'b11111111111111110111100011011000;
assign LUT_2[42136] = 32'b11111111111111110010000101111000;
assign LUT_2[42137] = 32'b11111111111111101110111110010001;
assign LUT_2[42138] = 32'b11111111111111111000111110110100;
assign LUT_2[42139] = 32'b11111111111111110101110111001101;
assign LUT_2[42140] = 32'b11111111111111101110100011100000;
assign LUT_2[42141] = 32'b11111111111111101011011011111001;
assign LUT_2[42142] = 32'b11111111111111110101011100011100;
assign LUT_2[42143] = 32'b11111111111111110010010100110101;
assign LUT_2[42144] = 32'b11111111111111111101001011111010;
assign LUT_2[42145] = 32'b11111111111111111010000100010011;
assign LUT_2[42146] = 32'b00000000000000000100000100110110;
assign LUT_2[42147] = 32'b00000000000000000000111101001111;
assign LUT_2[42148] = 32'b11111111111111111001101001100010;
assign LUT_2[42149] = 32'b11111111111111110110100001111011;
assign LUT_2[42150] = 32'b00000000000000000000100010011110;
assign LUT_2[42151] = 32'b11111111111111111101011010110111;
assign LUT_2[42152] = 32'b11111111111111110111111101010111;
assign LUT_2[42153] = 32'b11111111111111110100110101110000;
assign LUT_2[42154] = 32'b11111111111111111110110110010011;
assign LUT_2[42155] = 32'b11111111111111111011101110101100;
assign LUT_2[42156] = 32'b11111111111111110100011010111111;
assign LUT_2[42157] = 32'b11111111111111110001010011011000;
assign LUT_2[42158] = 32'b11111111111111111011010011111011;
assign LUT_2[42159] = 32'b11111111111111111000001100010100;
assign LUT_2[42160] = 32'b11111111111111110111110000000100;
assign LUT_2[42161] = 32'b11111111111111110100101000011101;
assign LUT_2[42162] = 32'b11111111111111111110101001000000;
assign LUT_2[42163] = 32'b11111111111111111011100001011001;
assign LUT_2[42164] = 32'b11111111111111110100001101101100;
assign LUT_2[42165] = 32'b11111111111111110001000110000101;
assign LUT_2[42166] = 32'b11111111111111111011000110101000;
assign LUT_2[42167] = 32'b11111111111111110111111111000001;
assign LUT_2[42168] = 32'b11111111111111110010100001100001;
assign LUT_2[42169] = 32'b11111111111111101111011001111010;
assign LUT_2[42170] = 32'b11111111111111111001011010011101;
assign LUT_2[42171] = 32'b11111111111111110110010010110110;
assign LUT_2[42172] = 32'b11111111111111101110111111001001;
assign LUT_2[42173] = 32'b11111111111111101011110111100010;
assign LUT_2[42174] = 32'b11111111111111110101111000000101;
assign LUT_2[42175] = 32'b11111111111111110010110000011110;
assign LUT_2[42176] = 32'b11111111111111110100111000110100;
assign LUT_2[42177] = 32'b11111111111111110001110001001101;
assign LUT_2[42178] = 32'b11111111111111111011110001110000;
assign LUT_2[42179] = 32'b11111111111111111000101010001001;
assign LUT_2[42180] = 32'b11111111111111110001010110011100;
assign LUT_2[42181] = 32'b11111111111111101110001110110101;
assign LUT_2[42182] = 32'b11111111111111111000001111011000;
assign LUT_2[42183] = 32'b11111111111111110101000111110001;
assign LUT_2[42184] = 32'b11111111111111101111101010010001;
assign LUT_2[42185] = 32'b11111111111111101100100010101010;
assign LUT_2[42186] = 32'b11111111111111110110100011001101;
assign LUT_2[42187] = 32'b11111111111111110011011011100110;
assign LUT_2[42188] = 32'b11111111111111101100000111111001;
assign LUT_2[42189] = 32'b11111111111111101001000000010010;
assign LUT_2[42190] = 32'b11111111111111110011000000110101;
assign LUT_2[42191] = 32'b11111111111111101111111001001110;
assign LUT_2[42192] = 32'b11111111111111101111011100111110;
assign LUT_2[42193] = 32'b11111111111111101100010101010111;
assign LUT_2[42194] = 32'b11111111111111110110010101111010;
assign LUT_2[42195] = 32'b11111111111111110011001110010011;
assign LUT_2[42196] = 32'b11111111111111101011111010100110;
assign LUT_2[42197] = 32'b11111111111111101000110010111111;
assign LUT_2[42198] = 32'b11111111111111110010110011100010;
assign LUT_2[42199] = 32'b11111111111111101111101011111011;
assign LUT_2[42200] = 32'b11111111111111101010001110011011;
assign LUT_2[42201] = 32'b11111111111111100111000110110100;
assign LUT_2[42202] = 32'b11111111111111110001000111010111;
assign LUT_2[42203] = 32'b11111111111111101101111111110000;
assign LUT_2[42204] = 32'b11111111111111100110101100000011;
assign LUT_2[42205] = 32'b11111111111111100011100100011100;
assign LUT_2[42206] = 32'b11111111111111101101100100111111;
assign LUT_2[42207] = 32'b11111111111111101010011101011000;
assign LUT_2[42208] = 32'b11111111111111110101010100011101;
assign LUT_2[42209] = 32'b11111111111111110010001100110110;
assign LUT_2[42210] = 32'b11111111111111111100001101011001;
assign LUT_2[42211] = 32'b11111111111111111001000101110010;
assign LUT_2[42212] = 32'b11111111111111110001110010000101;
assign LUT_2[42213] = 32'b11111111111111101110101010011110;
assign LUT_2[42214] = 32'b11111111111111111000101011000001;
assign LUT_2[42215] = 32'b11111111111111110101100011011010;
assign LUT_2[42216] = 32'b11111111111111110000000101111010;
assign LUT_2[42217] = 32'b11111111111111101100111110010011;
assign LUT_2[42218] = 32'b11111111111111110110111110110110;
assign LUT_2[42219] = 32'b11111111111111110011110111001111;
assign LUT_2[42220] = 32'b11111111111111101100100011100010;
assign LUT_2[42221] = 32'b11111111111111101001011011111011;
assign LUT_2[42222] = 32'b11111111111111110011011100011110;
assign LUT_2[42223] = 32'b11111111111111110000010100110111;
assign LUT_2[42224] = 32'b11111111111111101111111000100111;
assign LUT_2[42225] = 32'b11111111111111101100110001000000;
assign LUT_2[42226] = 32'b11111111111111110110110001100011;
assign LUT_2[42227] = 32'b11111111111111110011101001111100;
assign LUT_2[42228] = 32'b11111111111111101100010110001111;
assign LUT_2[42229] = 32'b11111111111111101001001110101000;
assign LUT_2[42230] = 32'b11111111111111110011001111001011;
assign LUT_2[42231] = 32'b11111111111111110000000111100100;
assign LUT_2[42232] = 32'b11111111111111101010101010000100;
assign LUT_2[42233] = 32'b11111111111111100111100010011101;
assign LUT_2[42234] = 32'b11111111111111110001100011000000;
assign LUT_2[42235] = 32'b11111111111111101110011011011001;
assign LUT_2[42236] = 32'b11111111111111100111000111101100;
assign LUT_2[42237] = 32'b11111111111111100100000000000101;
assign LUT_2[42238] = 32'b11111111111111101110000000101000;
assign LUT_2[42239] = 32'b11111111111111101010111001000001;
assign LUT_2[42240] = 32'b11111111111111111100011010101000;
assign LUT_2[42241] = 32'b11111111111111111001010011000001;
assign LUT_2[42242] = 32'b00000000000000000011010011100100;
assign LUT_2[42243] = 32'b00000000000000000000001011111101;
assign LUT_2[42244] = 32'b11111111111111111000111000010000;
assign LUT_2[42245] = 32'b11111111111111110101110000101001;
assign LUT_2[42246] = 32'b11111111111111111111110001001100;
assign LUT_2[42247] = 32'b11111111111111111100101001100101;
assign LUT_2[42248] = 32'b11111111111111110111001100000101;
assign LUT_2[42249] = 32'b11111111111111110100000100011110;
assign LUT_2[42250] = 32'b11111111111111111110000101000001;
assign LUT_2[42251] = 32'b11111111111111111010111101011010;
assign LUT_2[42252] = 32'b11111111111111110011101001101101;
assign LUT_2[42253] = 32'b11111111111111110000100010000110;
assign LUT_2[42254] = 32'b11111111111111111010100010101001;
assign LUT_2[42255] = 32'b11111111111111110111011011000010;
assign LUT_2[42256] = 32'b11111111111111110110111110110010;
assign LUT_2[42257] = 32'b11111111111111110011110111001011;
assign LUT_2[42258] = 32'b11111111111111111101110111101110;
assign LUT_2[42259] = 32'b11111111111111111010110000000111;
assign LUT_2[42260] = 32'b11111111111111110011011100011010;
assign LUT_2[42261] = 32'b11111111111111110000010100110011;
assign LUT_2[42262] = 32'b11111111111111111010010101010110;
assign LUT_2[42263] = 32'b11111111111111110111001101101111;
assign LUT_2[42264] = 32'b11111111111111110001110000001111;
assign LUT_2[42265] = 32'b11111111111111101110101000101000;
assign LUT_2[42266] = 32'b11111111111111111000101001001011;
assign LUT_2[42267] = 32'b11111111111111110101100001100100;
assign LUT_2[42268] = 32'b11111111111111101110001101110111;
assign LUT_2[42269] = 32'b11111111111111101011000110010000;
assign LUT_2[42270] = 32'b11111111111111110101000110110011;
assign LUT_2[42271] = 32'b11111111111111110001111111001100;
assign LUT_2[42272] = 32'b11111111111111111100110110010001;
assign LUT_2[42273] = 32'b11111111111111111001101110101010;
assign LUT_2[42274] = 32'b00000000000000000011101111001101;
assign LUT_2[42275] = 32'b00000000000000000000100111100110;
assign LUT_2[42276] = 32'b11111111111111111001010011111001;
assign LUT_2[42277] = 32'b11111111111111110110001100010010;
assign LUT_2[42278] = 32'b00000000000000000000001100110101;
assign LUT_2[42279] = 32'b11111111111111111101000101001110;
assign LUT_2[42280] = 32'b11111111111111110111100111101110;
assign LUT_2[42281] = 32'b11111111111111110100100000000111;
assign LUT_2[42282] = 32'b11111111111111111110100000101010;
assign LUT_2[42283] = 32'b11111111111111111011011001000011;
assign LUT_2[42284] = 32'b11111111111111110100000101010110;
assign LUT_2[42285] = 32'b11111111111111110000111101101111;
assign LUT_2[42286] = 32'b11111111111111111010111110010010;
assign LUT_2[42287] = 32'b11111111111111110111110110101011;
assign LUT_2[42288] = 32'b11111111111111110111011010011011;
assign LUT_2[42289] = 32'b11111111111111110100010010110100;
assign LUT_2[42290] = 32'b11111111111111111110010011010111;
assign LUT_2[42291] = 32'b11111111111111111011001011110000;
assign LUT_2[42292] = 32'b11111111111111110011111000000011;
assign LUT_2[42293] = 32'b11111111111111110000110000011100;
assign LUT_2[42294] = 32'b11111111111111111010110000111111;
assign LUT_2[42295] = 32'b11111111111111110111101001011000;
assign LUT_2[42296] = 32'b11111111111111110010001011111000;
assign LUT_2[42297] = 32'b11111111111111101111000100010001;
assign LUT_2[42298] = 32'b11111111111111111001000100110100;
assign LUT_2[42299] = 32'b11111111111111110101111101001101;
assign LUT_2[42300] = 32'b11111111111111101110101001100000;
assign LUT_2[42301] = 32'b11111111111111101011100001111001;
assign LUT_2[42302] = 32'b11111111111111110101100010011100;
assign LUT_2[42303] = 32'b11111111111111110010011010110101;
assign LUT_2[42304] = 32'b11111111111111110100100011001011;
assign LUT_2[42305] = 32'b11111111111111110001011011100100;
assign LUT_2[42306] = 32'b11111111111111111011011100000111;
assign LUT_2[42307] = 32'b11111111111111111000010100100000;
assign LUT_2[42308] = 32'b11111111111111110001000000110011;
assign LUT_2[42309] = 32'b11111111111111101101111001001100;
assign LUT_2[42310] = 32'b11111111111111110111111001101111;
assign LUT_2[42311] = 32'b11111111111111110100110010001000;
assign LUT_2[42312] = 32'b11111111111111101111010100101000;
assign LUT_2[42313] = 32'b11111111111111101100001101000001;
assign LUT_2[42314] = 32'b11111111111111110110001101100100;
assign LUT_2[42315] = 32'b11111111111111110011000101111101;
assign LUT_2[42316] = 32'b11111111111111101011110010010000;
assign LUT_2[42317] = 32'b11111111111111101000101010101001;
assign LUT_2[42318] = 32'b11111111111111110010101011001100;
assign LUT_2[42319] = 32'b11111111111111101111100011100101;
assign LUT_2[42320] = 32'b11111111111111101111000111010101;
assign LUT_2[42321] = 32'b11111111111111101011111111101110;
assign LUT_2[42322] = 32'b11111111111111110110000000010001;
assign LUT_2[42323] = 32'b11111111111111110010111000101010;
assign LUT_2[42324] = 32'b11111111111111101011100100111101;
assign LUT_2[42325] = 32'b11111111111111101000011101010110;
assign LUT_2[42326] = 32'b11111111111111110010011101111001;
assign LUT_2[42327] = 32'b11111111111111101111010110010010;
assign LUT_2[42328] = 32'b11111111111111101001111000110010;
assign LUT_2[42329] = 32'b11111111111111100110110001001011;
assign LUT_2[42330] = 32'b11111111111111110000110001101110;
assign LUT_2[42331] = 32'b11111111111111101101101010000111;
assign LUT_2[42332] = 32'b11111111111111100110010110011010;
assign LUT_2[42333] = 32'b11111111111111100011001110110011;
assign LUT_2[42334] = 32'b11111111111111101101001111010110;
assign LUT_2[42335] = 32'b11111111111111101010000111101111;
assign LUT_2[42336] = 32'b11111111111111110100111110110100;
assign LUT_2[42337] = 32'b11111111111111110001110111001101;
assign LUT_2[42338] = 32'b11111111111111111011110111110000;
assign LUT_2[42339] = 32'b11111111111111111000110000001001;
assign LUT_2[42340] = 32'b11111111111111110001011100011100;
assign LUT_2[42341] = 32'b11111111111111101110010100110101;
assign LUT_2[42342] = 32'b11111111111111111000010101011000;
assign LUT_2[42343] = 32'b11111111111111110101001101110001;
assign LUT_2[42344] = 32'b11111111111111101111110000010001;
assign LUT_2[42345] = 32'b11111111111111101100101000101010;
assign LUT_2[42346] = 32'b11111111111111110110101001001101;
assign LUT_2[42347] = 32'b11111111111111110011100001100110;
assign LUT_2[42348] = 32'b11111111111111101100001101111001;
assign LUT_2[42349] = 32'b11111111111111101001000110010010;
assign LUT_2[42350] = 32'b11111111111111110011000110110101;
assign LUT_2[42351] = 32'b11111111111111101111111111001110;
assign LUT_2[42352] = 32'b11111111111111101111100010111110;
assign LUT_2[42353] = 32'b11111111111111101100011011010111;
assign LUT_2[42354] = 32'b11111111111111110110011011111010;
assign LUT_2[42355] = 32'b11111111111111110011010100010011;
assign LUT_2[42356] = 32'b11111111111111101100000000100110;
assign LUT_2[42357] = 32'b11111111111111101000111000111111;
assign LUT_2[42358] = 32'b11111111111111110010111001100010;
assign LUT_2[42359] = 32'b11111111111111101111110001111011;
assign LUT_2[42360] = 32'b11111111111111101010010100011011;
assign LUT_2[42361] = 32'b11111111111111100111001100110100;
assign LUT_2[42362] = 32'b11111111111111110001001101010111;
assign LUT_2[42363] = 32'b11111111111111101110000101110000;
assign LUT_2[42364] = 32'b11111111111111100110110010000011;
assign LUT_2[42365] = 32'b11111111111111100011101010011100;
assign LUT_2[42366] = 32'b11111111111111101101101010111111;
assign LUT_2[42367] = 32'b11111111111111101010100011011000;
assign LUT_2[42368] = 32'b00000000000000000000101110110111;
assign LUT_2[42369] = 32'b11111111111111111101100111010000;
assign LUT_2[42370] = 32'b00000000000000000111100111110011;
assign LUT_2[42371] = 32'b00000000000000000100100000001100;
assign LUT_2[42372] = 32'b11111111111111111101001100011111;
assign LUT_2[42373] = 32'b11111111111111111010000100111000;
assign LUT_2[42374] = 32'b00000000000000000100000101011011;
assign LUT_2[42375] = 32'b00000000000000000000111101110100;
assign LUT_2[42376] = 32'b11111111111111111011100000010100;
assign LUT_2[42377] = 32'b11111111111111111000011000101101;
assign LUT_2[42378] = 32'b00000000000000000010011001010000;
assign LUT_2[42379] = 32'b11111111111111111111010001101001;
assign LUT_2[42380] = 32'b11111111111111110111111101111100;
assign LUT_2[42381] = 32'b11111111111111110100110110010101;
assign LUT_2[42382] = 32'b11111111111111111110110110111000;
assign LUT_2[42383] = 32'b11111111111111111011101111010001;
assign LUT_2[42384] = 32'b11111111111111111011010011000001;
assign LUT_2[42385] = 32'b11111111111111111000001011011010;
assign LUT_2[42386] = 32'b00000000000000000010001011111101;
assign LUT_2[42387] = 32'b11111111111111111111000100010110;
assign LUT_2[42388] = 32'b11111111111111110111110000101001;
assign LUT_2[42389] = 32'b11111111111111110100101001000010;
assign LUT_2[42390] = 32'b11111111111111111110101001100101;
assign LUT_2[42391] = 32'b11111111111111111011100001111110;
assign LUT_2[42392] = 32'b11111111111111110110000100011110;
assign LUT_2[42393] = 32'b11111111111111110010111100110111;
assign LUT_2[42394] = 32'b11111111111111111100111101011010;
assign LUT_2[42395] = 32'b11111111111111111001110101110011;
assign LUT_2[42396] = 32'b11111111111111110010100010000110;
assign LUT_2[42397] = 32'b11111111111111101111011010011111;
assign LUT_2[42398] = 32'b11111111111111111001011011000010;
assign LUT_2[42399] = 32'b11111111111111110110010011011011;
assign LUT_2[42400] = 32'b00000000000000000001001010100000;
assign LUT_2[42401] = 32'b11111111111111111110000010111001;
assign LUT_2[42402] = 32'b00000000000000001000000011011100;
assign LUT_2[42403] = 32'b00000000000000000100111011110101;
assign LUT_2[42404] = 32'b11111111111111111101101000001000;
assign LUT_2[42405] = 32'b11111111111111111010100000100001;
assign LUT_2[42406] = 32'b00000000000000000100100001000100;
assign LUT_2[42407] = 32'b00000000000000000001011001011101;
assign LUT_2[42408] = 32'b11111111111111111011111011111101;
assign LUT_2[42409] = 32'b11111111111111111000110100010110;
assign LUT_2[42410] = 32'b00000000000000000010110100111001;
assign LUT_2[42411] = 32'b11111111111111111111101101010010;
assign LUT_2[42412] = 32'b11111111111111111000011001100101;
assign LUT_2[42413] = 32'b11111111111111110101010001111110;
assign LUT_2[42414] = 32'b11111111111111111111010010100001;
assign LUT_2[42415] = 32'b11111111111111111100001010111010;
assign LUT_2[42416] = 32'b11111111111111111011101110101010;
assign LUT_2[42417] = 32'b11111111111111111000100111000011;
assign LUT_2[42418] = 32'b00000000000000000010100111100110;
assign LUT_2[42419] = 32'b11111111111111111111011111111111;
assign LUT_2[42420] = 32'b11111111111111111000001100010010;
assign LUT_2[42421] = 32'b11111111111111110101000100101011;
assign LUT_2[42422] = 32'b11111111111111111111000101001110;
assign LUT_2[42423] = 32'b11111111111111111011111101100111;
assign LUT_2[42424] = 32'b11111111111111110110100000000111;
assign LUT_2[42425] = 32'b11111111111111110011011000100000;
assign LUT_2[42426] = 32'b11111111111111111101011001000011;
assign LUT_2[42427] = 32'b11111111111111111010010001011100;
assign LUT_2[42428] = 32'b11111111111111110010111101101111;
assign LUT_2[42429] = 32'b11111111111111101111110110001000;
assign LUT_2[42430] = 32'b11111111111111111001110110101011;
assign LUT_2[42431] = 32'b11111111111111110110101111000100;
assign LUT_2[42432] = 32'b11111111111111111000110111011010;
assign LUT_2[42433] = 32'b11111111111111110101101111110011;
assign LUT_2[42434] = 32'b11111111111111111111110000010110;
assign LUT_2[42435] = 32'b11111111111111111100101000101111;
assign LUT_2[42436] = 32'b11111111111111110101010101000010;
assign LUT_2[42437] = 32'b11111111111111110010001101011011;
assign LUT_2[42438] = 32'b11111111111111111100001101111110;
assign LUT_2[42439] = 32'b11111111111111111001000110010111;
assign LUT_2[42440] = 32'b11111111111111110011101000110111;
assign LUT_2[42441] = 32'b11111111111111110000100001010000;
assign LUT_2[42442] = 32'b11111111111111111010100001110011;
assign LUT_2[42443] = 32'b11111111111111110111011010001100;
assign LUT_2[42444] = 32'b11111111111111110000000110011111;
assign LUT_2[42445] = 32'b11111111111111101100111110111000;
assign LUT_2[42446] = 32'b11111111111111110110111111011011;
assign LUT_2[42447] = 32'b11111111111111110011110111110100;
assign LUT_2[42448] = 32'b11111111111111110011011011100100;
assign LUT_2[42449] = 32'b11111111111111110000010011111101;
assign LUT_2[42450] = 32'b11111111111111111010010100100000;
assign LUT_2[42451] = 32'b11111111111111110111001100111001;
assign LUT_2[42452] = 32'b11111111111111101111111001001100;
assign LUT_2[42453] = 32'b11111111111111101100110001100101;
assign LUT_2[42454] = 32'b11111111111111110110110010001000;
assign LUT_2[42455] = 32'b11111111111111110011101010100001;
assign LUT_2[42456] = 32'b11111111111111101110001101000001;
assign LUT_2[42457] = 32'b11111111111111101011000101011010;
assign LUT_2[42458] = 32'b11111111111111110101000101111101;
assign LUT_2[42459] = 32'b11111111111111110001111110010110;
assign LUT_2[42460] = 32'b11111111111111101010101010101001;
assign LUT_2[42461] = 32'b11111111111111100111100011000010;
assign LUT_2[42462] = 32'b11111111111111110001100011100101;
assign LUT_2[42463] = 32'b11111111111111101110011011111110;
assign LUT_2[42464] = 32'b11111111111111111001010011000011;
assign LUT_2[42465] = 32'b11111111111111110110001011011100;
assign LUT_2[42466] = 32'b00000000000000000000001011111111;
assign LUT_2[42467] = 32'b11111111111111111101000100011000;
assign LUT_2[42468] = 32'b11111111111111110101110000101011;
assign LUT_2[42469] = 32'b11111111111111110010101001000100;
assign LUT_2[42470] = 32'b11111111111111111100101001100111;
assign LUT_2[42471] = 32'b11111111111111111001100010000000;
assign LUT_2[42472] = 32'b11111111111111110100000100100000;
assign LUT_2[42473] = 32'b11111111111111110000111100111001;
assign LUT_2[42474] = 32'b11111111111111111010111101011100;
assign LUT_2[42475] = 32'b11111111111111110111110101110101;
assign LUT_2[42476] = 32'b11111111111111110000100010001000;
assign LUT_2[42477] = 32'b11111111111111101101011010100001;
assign LUT_2[42478] = 32'b11111111111111110111011011000100;
assign LUT_2[42479] = 32'b11111111111111110100010011011101;
assign LUT_2[42480] = 32'b11111111111111110011110111001101;
assign LUT_2[42481] = 32'b11111111111111110000101111100110;
assign LUT_2[42482] = 32'b11111111111111111010110000001001;
assign LUT_2[42483] = 32'b11111111111111110111101000100010;
assign LUT_2[42484] = 32'b11111111111111110000010100110101;
assign LUT_2[42485] = 32'b11111111111111101101001101001110;
assign LUT_2[42486] = 32'b11111111111111110111001101110001;
assign LUT_2[42487] = 32'b11111111111111110100000110001010;
assign LUT_2[42488] = 32'b11111111111111101110101000101010;
assign LUT_2[42489] = 32'b11111111111111101011100001000011;
assign LUT_2[42490] = 32'b11111111111111110101100001100110;
assign LUT_2[42491] = 32'b11111111111111110010011001111111;
assign LUT_2[42492] = 32'b11111111111111101011000110010010;
assign LUT_2[42493] = 32'b11111111111111100111111110101011;
assign LUT_2[42494] = 32'b11111111111111110001111111001110;
assign LUT_2[42495] = 32'b11111111111111101110110111100111;
assign LUT_2[42496] = 32'b11111111111111111101001101110100;
assign LUT_2[42497] = 32'b11111111111111111010000110001101;
assign LUT_2[42498] = 32'b00000000000000000100000110110000;
assign LUT_2[42499] = 32'b00000000000000000000111111001001;
assign LUT_2[42500] = 32'b11111111111111111001101011011100;
assign LUT_2[42501] = 32'b11111111111111110110100011110101;
assign LUT_2[42502] = 32'b00000000000000000000100100011000;
assign LUT_2[42503] = 32'b11111111111111111101011100110001;
assign LUT_2[42504] = 32'b11111111111111110111111111010001;
assign LUT_2[42505] = 32'b11111111111111110100110111101010;
assign LUT_2[42506] = 32'b11111111111111111110111000001101;
assign LUT_2[42507] = 32'b11111111111111111011110000100110;
assign LUT_2[42508] = 32'b11111111111111110100011100111001;
assign LUT_2[42509] = 32'b11111111111111110001010101010010;
assign LUT_2[42510] = 32'b11111111111111111011010101110101;
assign LUT_2[42511] = 32'b11111111111111111000001110001110;
assign LUT_2[42512] = 32'b11111111111111110111110001111110;
assign LUT_2[42513] = 32'b11111111111111110100101010010111;
assign LUT_2[42514] = 32'b11111111111111111110101010111010;
assign LUT_2[42515] = 32'b11111111111111111011100011010011;
assign LUT_2[42516] = 32'b11111111111111110100001111100110;
assign LUT_2[42517] = 32'b11111111111111110001000111111111;
assign LUT_2[42518] = 32'b11111111111111111011001000100010;
assign LUT_2[42519] = 32'b11111111111111111000000000111011;
assign LUT_2[42520] = 32'b11111111111111110010100011011011;
assign LUT_2[42521] = 32'b11111111111111101111011011110100;
assign LUT_2[42522] = 32'b11111111111111111001011100010111;
assign LUT_2[42523] = 32'b11111111111111110110010100110000;
assign LUT_2[42524] = 32'b11111111111111101111000001000011;
assign LUT_2[42525] = 32'b11111111111111101011111001011100;
assign LUT_2[42526] = 32'b11111111111111110101111001111111;
assign LUT_2[42527] = 32'b11111111111111110010110010011000;
assign LUT_2[42528] = 32'b11111111111111111101101001011101;
assign LUT_2[42529] = 32'b11111111111111111010100001110110;
assign LUT_2[42530] = 32'b00000000000000000100100010011001;
assign LUT_2[42531] = 32'b00000000000000000001011010110010;
assign LUT_2[42532] = 32'b11111111111111111010000111000101;
assign LUT_2[42533] = 32'b11111111111111110110111111011110;
assign LUT_2[42534] = 32'b00000000000000000001000000000001;
assign LUT_2[42535] = 32'b11111111111111111101111000011010;
assign LUT_2[42536] = 32'b11111111111111111000011010111010;
assign LUT_2[42537] = 32'b11111111111111110101010011010011;
assign LUT_2[42538] = 32'b11111111111111111111010011110110;
assign LUT_2[42539] = 32'b11111111111111111100001100001111;
assign LUT_2[42540] = 32'b11111111111111110100111000100010;
assign LUT_2[42541] = 32'b11111111111111110001110000111011;
assign LUT_2[42542] = 32'b11111111111111111011110001011110;
assign LUT_2[42543] = 32'b11111111111111111000101001110111;
assign LUT_2[42544] = 32'b11111111111111111000001101100111;
assign LUT_2[42545] = 32'b11111111111111110101000110000000;
assign LUT_2[42546] = 32'b11111111111111111111000110100011;
assign LUT_2[42547] = 32'b11111111111111111011111110111100;
assign LUT_2[42548] = 32'b11111111111111110100101011001111;
assign LUT_2[42549] = 32'b11111111111111110001100011101000;
assign LUT_2[42550] = 32'b11111111111111111011100100001011;
assign LUT_2[42551] = 32'b11111111111111111000011100100100;
assign LUT_2[42552] = 32'b11111111111111110010111111000100;
assign LUT_2[42553] = 32'b11111111111111101111110111011101;
assign LUT_2[42554] = 32'b11111111111111111001111000000000;
assign LUT_2[42555] = 32'b11111111111111110110110000011001;
assign LUT_2[42556] = 32'b11111111111111101111011100101100;
assign LUT_2[42557] = 32'b11111111111111101100010101000101;
assign LUT_2[42558] = 32'b11111111111111110110010101101000;
assign LUT_2[42559] = 32'b11111111111111110011001110000001;
assign LUT_2[42560] = 32'b11111111111111110101010110010111;
assign LUT_2[42561] = 32'b11111111111111110010001110110000;
assign LUT_2[42562] = 32'b11111111111111111100001111010011;
assign LUT_2[42563] = 32'b11111111111111111001000111101100;
assign LUT_2[42564] = 32'b11111111111111110001110011111111;
assign LUT_2[42565] = 32'b11111111111111101110101100011000;
assign LUT_2[42566] = 32'b11111111111111111000101100111011;
assign LUT_2[42567] = 32'b11111111111111110101100101010100;
assign LUT_2[42568] = 32'b11111111111111110000000111110100;
assign LUT_2[42569] = 32'b11111111111111101101000000001101;
assign LUT_2[42570] = 32'b11111111111111110111000000110000;
assign LUT_2[42571] = 32'b11111111111111110011111001001001;
assign LUT_2[42572] = 32'b11111111111111101100100101011100;
assign LUT_2[42573] = 32'b11111111111111101001011101110101;
assign LUT_2[42574] = 32'b11111111111111110011011110011000;
assign LUT_2[42575] = 32'b11111111111111110000010110110001;
assign LUT_2[42576] = 32'b11111111111111101111111010100001;
assign LUT_2[42577] = 32'b11111111111111101100110010111010;
assign LUT_2[42578] = 32'b11111111111111110110110011011101;
assign LUT_2[42579] = 32'b11111111111111110011101011110110;
assign LUT_2[42580] = 32'b11111111111111101100011000001001;
assign LUT_2[42581] = 32'b11111111111111101001010000100010;
assign LUT_2[42582] = 32'b11111111111111110011010001000101;
assign LUT_2[42583] = 32'b11111111111111110000001001011110;
assign LUT_2[42584] = 32'b11111111111111101010101011111110;
assign LUT_2[42585] = 32'b11111111111111100111100100010111;
assign LUT_2[42586] = 32'b11111111111111110001100100111010;
assign LUT_2[42587] = 32'b11111111111111101110011101010011;
assign LUT_2[42588] = 32'b11111111111111100111001001100110;
assign LUT_2[42589] = 32'b11111111111111100100000001111111;
assign LUT_2[42590] = 32'b11111111111111101110000010100010;
assign LUT_2[42591] = 32'b11111111111111101010111010111011;
assign LUT_2[42592] = 32'b11111111111111110101110010000000;
assign LUT_2[42593] = 32'b11111111111111110010101010011001;
assign LUT_2[42594] = 32'b11111111111111111100101010111100;
assign LUT_2[42595] = 32'b11111111111111111001100011010101;
assign LUT_2[42596] = 32'b11111111111111110010001111101000;
assign LUT_2[42597] = 32'b11111111111111101111001000000001;
assign LUT_2[42598] = 32'b11111111111111111001001000100100;
assign LUT_2[42599] = 32'b11111111111111110110000000111101;
assign LUT_2[42600] = 32'b11111111111111110000100011011101;
assign LUT_2[42601] = 32'b11111111111111101101011011110110;
assign LUT_2[42602] = 32'b11111111111111110111011100011001;
assign LUT_2[42603] = 32'b11111111111111110100010100110010;
assign LUT_2[42604] = 32'b11111111111111101101000001000101;
assign LUT_2[42605] = 32'b11111111111111101001111001011110;
assign LUT_2[42606] = 32'b11111111111111110011111010000001;
assign LUT_2[42607] = 32'b11111111111111110000110010011010;
assign LUT_2[42608] = 32'b11111111111111110000010110001010;
assign LUT_2[42609] = 32'b11111111111111101101001110100011;
assign LUT_2[42610] = 32'b11111111111111110111001111000110;
assign LUT_2[42611] = 32'b11111111111111110100000111011111;
assign LUT_2[42612] = 32'b11111111111111101100110011110010;
assign LUT_2[42613] = 32'b11111111111111101001101100001011;
assign LUT_2[42614] = 32'b11111111111111110011101100101110;
assign LUT_2[42615] = 32'b11111111111111110000100101000111;
assign LUT_2[42616] = 32'b11111111111111101011000111100111;
assign LUT_2[42617] = 32'b11111111111111101000000000000000;
assign LUT_2[42618] = 32'b11111111111111110010000000100011;
assign LUT_2[42619] = 32'b11111111111111101110111000111100;
assign LUT_2[42620] = 32'b11111111111111100111100101001111;
assign LUT_2[42621] = 32'b11111111111111100100011101101000;
assign LUT_2[42622] = 32'b11111111111111101110011110001011;
assign LUT_2[42623] = 32'b11111111111111101011010110100100;
assign LUT_2[42624] = 32'b00000000000000000001100010000011;
assign LUT_2[42625] = 32'b11111111111111111110011010011100;
assign LUT_2[42626] = 32'b00000000000000001000011010111111;
assign LUT_2[42627] = 32'b00000000000000000101010011011000;
assign LUT_2[42628] = 32'b11111111111111111101111111101011;
assign LUT_2[42629] = 32'b11111111111111111010111000000100;
assign LUT_2[42630] = 32'b00000000000000000100111000100111;
assign LUT_2[42631] = 32'b00000000000000000001110001000000;
assign LUT_2[42632] = 32'b11111111111111111100010011100000;
assign LUT_2[42633] = 32'b11111111111111111001001011111001;
assign LUT_2[42634] = 32'b00000000000000000011001100011100;
assign LUT_2[42635] = 32'b00000000000000000000000100110101;
assign LUT_2[42636] = 32'b11111111111111111000110001001000;
assign LUT_2[42637] = 32'b11111111111111110101101001100001;
assign LUT_2[42638] = 32'b11111111111111111111101010000100;
assign LUT_2[42639] = 32'b11111111111111111100100010011101;
assign LUT_2[42640] = 32'b11111111111111111100000110001101;
assign LUT_2[42641] = 32'b11111111111111111000111110100110;
assign LUT_2[42642] = 32'b00000000000000000010111111001001;
assign LUT_2[42643] = 32'b11111111111111111111110111100010;
assign LUT_2[42644] = 32'b11111111111111111000100011110101;
assign LUT_2[42645] = 32'b11111111111111110101011100001110;
assign LUT_2[42646] = 32'b11111111111111111111011100110001;
assign LUT_2[42647] = 32'b11111111111111111100010101001010;
assign LUT_2[42648] = 32'b11111111111111110110110111101010;
assign LUT_2[42649] = 32'b11111111111111110011110000000011;
assign LUT_2[42650] = 32'b11111111111111111101110000100110;
assign LUT_2[42651] = 32'b11111111111111111010101000111111;
assign LUT_2[42652] = 32'b11111111111111110011010101010010;
assign LUT_2[42653] = 32'b11111111111111110000001101101011;
assign LUT_2[42654] = 32'b11111111111111111010001110001110;
assign LUT_2[42655] = 32'b11111111111111110111000110100111;
assign LUT_2[42656] = 32'b00000000000000000001111101101100;
assign LUT_2[42657] = 32'b11111111111111111110110110000101;
assign LUT_2[42658] = 32'b00000000000000001000110110101000;
assign LUT_2[42659] = 32'b00000000000000000101101111000001;
assign LUT_2[42660] = 32'b11111111111111111110011011010100;
assign LUT_2[42661] = 32'b11111111111111111011010011101101;
assign LUT_2[42662] = 32'b00000000000000000101010100010000;
assign LUT_2[42663] = 32'b00000000000000000010001100101001;
assign LUT_2[42664] = 32'b11111111111111111100101111001001;
assign LUT_2[42665] = 32'b11111111111111111001100111100010;
assign LUT_2[42666] = 32'b00000000000000000011101000000101;
assign LUT_2[42667] = 32'b00000000000000000000100000011110;
assign LUT_2[42668] = 32'b11111111111111111001001100110001;
assign LUT_2[42669] = 32'b11111111111111110110000101001010;
assign LUT_2[42670] = 32'b00000000000000000000000101101101;
assign LUT_2[42671] = 32'b11111111111111111100111110000110;
assign LUT_2[42672] = 32'b11111111111111111100100001110110;
assign LUT_2[42673] = 32'b11111111111111111001011010001111;
assign LUT_2[42674] = 32'b00000000000000000011011010110010;
assign LUT_2[42675] = 32'b00000000000000000000010011001011;
assign LUT_2[42676] = 32'b11111111111111111000111111011110;
assign LUT_2[42677] = 32'b11111111111111110101110111110111;
assign LUT_2[42678] = 32'b11111111111111111111111000011010;
assign LUT_2[42679] = 32'b11111111111111111100110000110011;
assign LUT_2[42680] = 32'b11111111111111110111010011010011;
assign LUT_2[42681] = 32'b11111111111111110100001011101100;
assign LUT_2[42682] = 32'b11111111111111111110001100001111;
assign LUT_2[42683] = 32'b11111111111111111011000100101000;
assign LUT_2[42684] = 32'b11111111111111110011110000111011;
assign LUT_2[42685] = 32'b11111111111111110000101001010100;
assign LUT_2[42686] = 32'b11111111111111111010101001110111;
assign LUT_2[42687] = 32'b11111111111111110111100010010000;
assign LUT_2[42688] = 32'b11111111111111111001101010100110;
assign LUT_2[42689] = 32'b11111111111111110110100010111111;
assign LUT_2[42690] = 32'b00000000000000000000100011100010;
assign LUT_2[42691] = 32'b11111111111111111101011011111011;
assign LUT_2[42692] = 32'b11111111111111110110001000001110;
assign LUT_2[42693] = 32'b11111111111111110011000000100111;
assign LUT_2[42694] = 32'b11111111111111111101000001001010;
assign LUT_2[42695] = 32'b11111111111111111001111001100011;
assign LUT_2[42696] = 32'b11111111111111110100011100000011;
assign LUT_2[42697] = 32'b11111111111111110001010100011100;
assign LUT_2[42698] = 32'b11111111111111111011010100111111;
assign LUT_2[42699] = 32'b11111111111111111000001101011000;
assign LUT_2[42700] = 32'b11111111111111110000111001101011;
assign LUT_2[42701] = 32'b11111111111111101101110010000100;
assign LUT_2[42702] = 32'b11111111111111110111110010100111;
assign LUT_2[42703] = 32'b11111111111111110100101011000000;
assign LUT_2[42704] = 32'b11111111111111110100001110110000;
assign LUT_2[42705] = 32'b11111111111111110001000111001001;
assign LUT_2[42706] = 32'b11111111111111111011000111101100;
assign LUT_2[42707] = 32'b11111111111111111000000000000101;
assign LUT_2[42708] = 32'b11111111111111110000101100011000;
assign LUT_2[42709] = 32'b11111111111111101101100100110001;
assign LUT_2[42710] = 32'b11111111111111110111100101010100;
assign LUT_2[42711] = 32'b11111111111111110100011101101101;
assign LUT_2[42712] = 32'b11111111111111101111000000001101;
assign LUT_2[42713] = 32'b11111111111111101011111000100110;
assign LUT_2[42714] = 32'b11111111111111110101111001001001;
assign LUT_2[42715] = 32'b11111111111111110010110001100010;
assign LUT_2[42716] = 32'b11111111111111101011011101110101;
assign LUT_2[42717] = 32'b11111111111111101000010110001110;
assign LUT_2[42718] = 32'b11111111111111110010010110110001;
assign LUT_2[42719] = 32'b11111111111111101111001111001010;
assign LUT_2[42720] = 32'b11111111111111111010000110001111;
assign LUT_2[42721] = 32'b11111111111111110110111110101000;
assign LUT_2[42722] = 32'b00000000000000000000111111001011;
assign LUT_2[42723] = 32'b11111111111111111101110111100100;
assign LUT_2[42724] = 32'b11111111111111110110100011110111;
assign LUT_2[42725] = 32'b11111111111111110011011100010000;
assign LUT_2[42726] = 32'b11111111111111111101011100110011;
assign LUT_2[42727] = 32'b11111111111111111010010101001100;
assign LUT_2[42728] = 32'b11111111111111110100110111101100;
assign LUT_2[42729] = 32'b11111111111111110001110000000101;
assign LUT_2[42730] = 32'b11111111111111111011110000101000;
assign LUT_2[42731] = 32'b11111111111111111000101001000001;
assign LUT_2[42732] = 32'b11111111111111110001010101010100;
assign LUT_2[42733] = 32'b11111111111111101110001101101101;
assign LUT_2[42734] = 32'b11111111111111111000001110010000;
assign LUT_2[42735] = 32'b11111111111111110101000110101001;
assign LUT_2[42736] = 32'b11111111111111110100101010011001;
assign LUT_2[42737] = 32'b11111111111111110001100010110010;
assign LUT_2[42738] = 32'b11111111111111111011100011010101;
assign LUT_2[42739] = 32'b11111111111111111000011011101110;
assign LUT_2[42740] = 32'b11111111111111110001001000000001;
assign LUT_2[42741] = 32'b11111111111111101110000000011010;
assign LUT_2[42742] = 32'b11111111111111111000000000111101;
assign LUT_2[42743] = 32'b11111111111111110100111001010110;
assign LUT_2[42744] = 32'b11111111111111101111011011110110;
assign LUT_2[42745] = 32'b11111111111111101100010100001111;
assign LUT_2[42746] = 32'b11111111111111110110010100110010;
assign LUT_2[42747] = 32'b11111111111111110011001101001011;
assign LUT_2[42748] = 32'b11111111111111101011111001011110;
assign LUT_2[42749] = 32'b11111111111111101000110001110111;
assign LUT_2[42750] = 32'b11111111111111110010110010011010;
assign LUT_2[42751] = 32'b11111111111111101111101010110011;
assign LUT_2[42752] = 32'b00000000000000000001001100011010;
assign LUT_2[42753] = 32'b11111111111111111110000100110011;
assign LUT_2[42754] = 32'b00000000000000001000000101010110;
assign LUT_2[42755] = 32'b00000000000000000100111101101111;
assign LUT_2[42756] = 32'b11111111111111111101101010000010;
assign LUT_2[42757] = 32'b11111111111111111010100010011011;
assign LUT_2[42758] = 32'b00000000000000000100100010111110;
assign LUT_2[42759] = 32'b00000000000000000001011011010111;
assign LUT_2[42760] = 32'b11111111111111111011111101110111;
assign LUT_2[42761] = 32'b11111111111111111000110110010000;
assign LUT_2[42762] = 32'b00000000000000000010110110110011;
assign LUT_2[42763] = 32'b11111111111111111111101111001100;
assign LUT_2[42764] = 32'b11111111111111111000011011011111;
assign LUT_2[42765] = 32'b11111111111111110101010011111000;
assign LUT_2[42766] = 32'b11111111111111111111010100011011;
assign LUT_2[42767] = 32'b11111111111111111100001100110100;
assign LUT_2[42768] = 32'b11111111111111111011110000100100;
assign LUT_2[42769] = 32'b11111111111111111000101000111101;
assign LUT_2[42770] = 32'b00000000000000000010101001100000;
assign LUT_2[42771] = 32'b11111111111111111111100001111001;
assign LUT_2[42772] = 32'b11111111111111111000001110001100;
assign LUT_2[42773] = 32'b11111111111111110101000110100101;
assign LUT_2[42774] = 32'b11111111111111111111000111001000;
assign LUT_2[42775] = 32'b11111111111111111011111111100001;
assign LUT_2[42776] = 32'b11111111111111110110100010000001;
assign LUT_2[42777] = 32'b11111111111111110011011010011010;
assign LUT_2[42778] = 32'b11111111111111111101011010111101;
assign LUT_2[42779] = 32'b11111111111111111010010011010110;
assign LUT_2[42780] = 32'b11111111111111110010111111101001;
assign LUT_2[42781] = 32'b11111111111111101111111000000010;
assign LUT_2[42782] = 32'b11111111111111111001111000100101;
assign LUT_2[42783] = 32'b11111111111111110110110000111110;
assign LUT_2[42784] = 32'b00000000000000000001101000000011;
assign LUT_2[42785] = 32'b11111111111111111110100000011100;
assign LUT_2[42786] = 32'b00000000000000001000100000111111;
assign LUT_2[42787] = 32'b00000000000000000101011001011000;
assign LUT_2[42788] = 32'b11111111111111111110000101101011;
assign LUT_2[42789] = 32'b11111111111111111010111110000100;
assign LUT_2[42790] = 32'b00000000000000000100111110100111;
assign LUT_2[42791] = 32'b00000000000000000001110111000000;
assign LUT_2[42792] = 32'b11111111111111111100011001100000;
assign LUT_2[42793] = 32'b11111111111111111001010001111001;
assign LUT_2[42794] = 32'b00000000000000000011010010011100;
assign LUT_2[42795] = 32'b00000000000000000000001010110101;
assign LUT_2[42796] = 32'b11111111111111111000110111001000;
assign LUT_2[42797] = 32'b11111111111111110101101111100001;
assign LUT_2[42798] = 32'b11111111111111111111110000000100;
assign LUT_2[42799] = 32'b11111111111111111100101000011101;
assign LUT_2[42800] = 32'b11111111111111111100001100001101;
assign LUT_2[42801] = 32'b11111111111111111001000100100110;
assign LUT_2[42802] = 32'b00000000000000000011000101001001;
assign LUT_2[42803] = 32'b11111111111111111111111101100010;
assign LUT_2[42804] = 32'b11111111111111111000101001110101;
assign LUT_2[42805] = 32'b11111111111111110101100010001110;
assign LUT_2[42806] = 32'b11111111111111111111100010110001;
assign LUT_2[42807] = 32'b11111111111111111100011011001010;
assign LUT_2[42808] = 32'b11111111111111110110111101101010;
assign LUT_2[42809] = 32'b11111111111111110011110110000011;
assign LUT_2[42810] = 32'b11111111111111111101110110100110;
assign LUT_2[42811] = 32'b11111111111111111010101110111111;
assign LUT_2[42812] = 32'b11111111111111110011011011010010;
assign LUT_2[42813] = 32'b11111111111111110000010011101011;
assign LUT_2[42814] = 32'b11111111111111111010010100001110;
assign LUT_2[42815] = 32'b11111111111111110111001100100111;
assign LUT_2[42816] = 32'b11111111111111111001010100111101;
assign LUT_2[42817] = 32'b11111111111111110110001101010110;
assign LUT_2[42818] = 32'b00000000000000000000001101111001;
assign LUT_2[42819] = 32'b11111111111111111101000110010010;
assign LUT_2[42820] = 32'b11111111111111110101110010100101;
assign LUT_2[42821] = 32'b11111111111111110010101010111110;
assign LUT_2[42822] = 32'b11111111111111111100101011100001;
assign LUT_2[42823] = 32'b11111111111111111001100011111010;
assign LUT_2[42824] = 32'b11111111111111110100000110011010;
assign LUT_2[42825] = 32'b11111111111111110000111110110011;
assign LUT_2[42826] = 32'b11111111111111111010111111010110;
assign LUT_2[42827] = 32'b11111111111111110111110111101111;
assign LUT_2[42828] = 32'b11111111111111110000100100000010;
assign LUT_2[42829] = 32'b11111111111111101101011100011011;
assign LUT_2[42830] = 32'b11111111111111110111011100111110;
assign LUT_2[42831] = 32'b11111111111111110100010101010111;
assign LUT_2[42832] = 32'b11111111111111110011111001000111;
assign LUT_2[42833] = 32'b11111111111111110000110001100000;
assign LUT_2[42834] = 32'b11111111111111111010110010000011;
assign LUT_2[42835] = 32'b11111111111111110111101010011100;
assign LUT_2[42836] = 32'b11111111111111110000010110101111;
assign LUT_2[42837] = 32'b11111111111111101101001111001000;
assign LUT_2[42838] = 32'b11111111111111110111001111101011;
assign LUT_2[42839] = 32'b11111111111111110100001000000100;
assign LUT_2[42840] = 32'b11111111111111101110101010100100;
assign LUT_2[42841] = 32'b11111111111111101011100010111101;
assign LUT_2[42842] = 32'b11111111111111110101100011100000;
assign LUT_2[42843] = 32'b11111111111111110010011011111001;
assign LUT_2[42844] = 32'b11111111111111101011001000001100;
assign LUT_2[42845] = 32'b11111111111111101000000000100101;
assign LUT_2[42846] = 32'b11111111111111110010000001001000;
assign LUT_2[42847] = 32'b11111111111111101110111001100001;
assign LUT_2[42848] = 32'b11111111111111111001110000100110;
assign LUT_2[42849] = 32'b11111111111111110110101000111111;
assign LUT_2[42850] = 32'b00000000000000000000101001100010;
assign LUT_2[42851] = 32'b11111111111111111101100001111011;
assign LUT_2[42852] = 32'b11111111111111110110001110001110;
assign LUT_2[42853] = 32'b11111111111111110011000110100111;
assign LUT_2[42854] = 32'b11111111111111111101000111001010;
assign LUT_2[42855] = 32'b11111111111111111001111111100011;
assign LUT_2[42856] = 32'b11111111111111110100100010000011;
assign LUT_2[42857] = 32'b11111111111111110001011010011100;
assign LUT_2[42858] = 32'b11111111111111111011011010111111;
assign LUT_2[42859] = 32'b11111111111111111000010011011000;
assign LUT_2[42860] = 32'b11111111111111110000111111101011;
assign LUT_2[42861] = 32'b11111111111111101101111000000100;
assign LUT_2[42862] = 32'b11111111111111110111111000100111;
assign LUT_2[42863] = 32'b11111111111111110100110001000000;
assign LUT_2[42864] = 32'b11111111111111110100010100110000;
assign LUT_2[42865] = 32'b11111111111111110001001101001001;
assign LUT_2[42866] = 32'b11111111111111111011001101101100;
assign LUT_2[42867] = 32'b11111111111111111000000110000101;
assign LUT_2[42868] = 32'b11111111111111110000110010011000;
assign LUT_2[42869] = 32'b11111111111111101101101010110001;
assign LUT_2[42870] = 32'b11111111111111110111101011010100;
assign LUT_2[42871] = 32'b11111111111111110100100011101101;
assign LUT_2[42872] = 32'b11111111111111101111000110001101;
assign LUT_2[42873] = 32'b11111111111111101011111110100110;
assign LUT_2[42874] = 32'b11111111111111110101111111001001;
assign LUT_2[42875] = 32'b11111111111111110010110111100010;
assign LUT_2[42876] = 32'b11111111111111101011100011110101;
assign LUT_2[42877] = 32'b11111111111111101000011100001110;
assign LUT_2[42878] = 32'b11111111111111110010011100110001;
assign LUT_2[42879] = 32'b11111111111111101111010101001010;
assign LUT_2[42880] = 32'b00000000000000000101100000101001;
assign LUT_2[42881] = 32'b00000000000000000010011001000010;
assign LUT_2[42882] = 32'b00000000000000001100011001100101;
assign LUT_2[42883] = 32'b00000000000000001001010001111110;
assign LUT_2[42884] = 32'b00000000000000000001111110010001;
assign LUT_2[42885] = 32'b11111111111111111110110110101010;
assign LUT_2[42886] = 32'b00000000000000001000110111001101;
assign LUT_2[42887] = 32'b00000000000000000101101111100110;
assign LUT_2[42888] = 32'b00000000000000000000010010000110;
assign LUT_2[42889] = 32'b11111111111111111101001010011111;
assign LUT_2[42890] = 32'b00000000000000000111001011000010;
assign LUT_2[42891] = 32'b00000000000000000100000011011011;
assign LUT_2[42892] = 32'b11111111111111111100101111101110;
assign LUT_2[42893] = 32'b11111111111111111001101000000111;
assign LUT_2[42894] = 32'b00000000000000000011101000101010;
assign LUT_2[42895] = 32'b00000000000000000000100001000011;
assign LUT_2[42896] = 32'b00000000000000000000000100110011;
assign LUT_2[42897] = 32'b11111111111111111100111101001100;
assign LUT_2[42898] = 32'b00000000000000000110111101101111;
assign LUT_2[42899] = 32'b00000000000000000011110110001000;
assign LUT_2[42900] = 32'b11111111111111111100100010011011;
assign LUT_2[42901] = 32'b11111111111111111001011010110100;
assign LUT_2[42902] = 32'b00000000000000000011011011010111;
assign LUT_2[42903] = 32'b00000000000000000000010011110000;
assign LUT_2[42904] = 32'b11111111111111111010110110010000;
assign LUT_2[42905] = 32'b11111111111111110111101110101001;
assign LUT_2[42906] = 32'b00000000000000000001101111001100;
assign LUT_2[42907] = 32'b11111111111111111110100111100101;
assign LUT_2[42908] = 32'b11111111111111110111010011111000;
assign LUT_2[42909] = 32'b11111111111111110100001100010001;
assign LUT_2[42910] = 32'b11111111111111111110001100110100;
assign LUT_2[42911] = 32'b11111111111111111011000101001101;
assign LUT_2[42912] = 32'b00000000000000000101111100010010;
assign LUT_2[42913] = 32'b00000000000000000010110100101011;
assign LUT_2[42914] = 32'b00000000000000001100110101001110;
assign LUT_2[42915] = 32'b00000000000000001001101101100111;
assign LUT_2[42916] = 32'b00000000000000000010011001111010;
assign LUT_2[42917] = 32'b11111111111111111111010010010011;
assign LUT_2[42918] = 32'b00000000000000001001010010110110;
assign LUT_2[42919] = 32'b00000000000000000110001011001111;
assign LUT_2[42920] = 32'b00000000000000000000101101101111;
assign LUT_2[42921] = 32'b11111111111111111101100110001000;
assign LUT_2[42922] = 32'b00000000000000000111100110101011;
assign LUT_2[42923] = 32'b00000000000000000100011111000100;
assign LUT_2[42924] = 32'b11111111111111111101001011010111;
assign LUT_2[42925] = 32'b11111111111111111010000011110000;
assign LUT_2[42926] = 32'b00000000000000000100000100010011;
assign LUT_2[42927] = 32'b00000000000000000000111100101100;
assign LUT_2[42928] = 32'b00000000000000000000100000011100;
assign LUT_2[42929] = 32'b11111111111111111101011000110101;
assign LUT_2[42930] = 32'b00000000000000000111011001011000;
assign LUT_2[42931] = 32'b00000000000000000100010001110001;
assign LUT_2[42932] = 32'b11111111111111111100111110000100;
assign LUT_2[42933] = 32'b11111111111111111001110110011101;
assign LUT_2[42934] = 32'b00000000000000000011110111000000;
assign LUT_2[42935] = 32'b00000000000000000000101111011001;
assign LUT_2[42936] = 32'b11111111111111111011010001111001;
assign LUT_2[42937] = 32'b11111111111111111000001010010010;
assign LUT_2[42938] = 32'b00000000000000000010001010110101;
assign LUT_2[42939] = 32'b11111111111111111111000011001110;
assign LUT_2[42940] = 32'b11111111111111110111101111100001;
assign LUT_2[42941] = 32'b11111111111111110100100111111010;
assign LUT_2[42942] = 32'b11111111111111111110101000011101;
assign LUT_2[42943] = 32'b11111111111111111011100000110110;
assign LUT_2[42944] = 32'b11111111111111111101101001001100;
assign LUT_2[42945] = 32'b11111111111111111010100001100101;
assign LUT_2[42946] = 32'b00000000000000000100100010001000;
assign LUT_2[42947] = 32'b00000000000000000001011010100001;
assign LUT_2[42948] = 32'b11111111111111111010000110110100;
assign LUT_2[42949] = 32'b11111111111111110110111111001101;
assign LUT_2[42950] = 32'b00000000000000000000111111110000;
assign LUT_2[42951] = 32'b11111111111111111101111000001001;
assign LUT_2[42952] = 32'b11111111111111111000011010101001;
assign LUT_2[42953] = 32'b11111111111111110101010011000010;
assign LUT_2[42954] = 32'b11111111111111111111010011100101;
assign LUT_2[42955] = 32'b11111111111111111100001011111110;
assign LUT_2[42956] = 32'b11111111111111110100111000010001;
assign LUT_2[42957] = 32'b11111111111111110001110000101010;
assign LUT_2[42958] = 32'b11111111111111111011110001001101;
assign LUT_2[42959] = 32'b11111111111111111000101001100110;
assign LUT_2[42960] = 32'b11111111111111111000001101010110;
assign LUT_2[42961] = 32'b11111111111111110101000101101111;
assign LUT_2[42962] = 32'b11111111111111111111000110010010;
assign LUT_2[42963] = 32'b11111111111111111011111110101011;
assign LUT_2[42964] = 32'b11111111111111110100101010111110;
assign LUT_2[42965] = 32'b11111111111111110001100011010111;
assign LUT_2[42966] = 32'b11111111111111111011100011111010;
assign LUT_2[42967] = 32'b11111111111111111000011100010011;
assign LUT_2[42968] = 32'b11111111111111110010111110110011;
assign LUT_2[42969] = 32'b11111111111111101111110111001100;
assign LUT_2[42970] = 32'b11111111111111111001110111101111;
assign LUT_2[42971] = 32'b11111111111111110110110000001000;
assign LUT_2[42972] = 32'b11111111111111101111011100011011;
assign LUT_2[42973] = 32'b11111111111111101100010100110100;
assign LUT_2[42974] = 32'b11111111111111110110010101010111;
assign LUT_2[42975] = 32'b11111111111111110011001101110000;
assign LUT_2[42976] = 32'b11111111111111111110000100110101;
assign LUT_2[42977] = 32'b11111111111111111010111101001110;
assign LUT_2[42978] = 32'b00000000000000000100111101110001;
assign LUT_2[42979] = 32'b00000000000000000001110110001010;
assign LUT_2[42980] = 32'b11111111111111111010100010011101;
assign LUT_2[42981] = 32'b11111111111111110111011010110110;
assign LUT_2[42982] = 32'b00000000000000000001011011011001;
assign LUT_2[42983] = 32'b11111111111111111110010011110010;
assign LUT_2[42984] = 32'b11111111111111111000110110010010;
assign LUT_2[42985] = 32'b11111111111111110101101110101011;
assign LUT_2[42986] = 32'b11111111111111111111101111001110;
assign LUT_2[42987] = 32'b11111111111111111100100111100111;
assign LUT_2[42988] = 32'b11111111111111110101010011111010;
assign LUT_2[42989] = 32'b11111111111111110010001100010011;
assign LUT_2[42990] = 32'b11111111111111111100001100110110;
assign LUT_2[42991] = 32'b11111111111111111001000101001111;
assign LUT_2[42992] = 32'b11111111111111111000101000111111;
assign LUT_2[42993] = 32'b11111111111111110101100001011000;
assign LUT_2[42994] = 32'b11111111111111111111100001111011;
assign LUT_2[42995] = 32'b11111111111111111100011010010100;
assign LUT_2[42996] = 32'b11111111111111110101000110100111;
assign LUT_2[42997] = 32'b11111111111111110001111111000000;
assign LUT_2[42998] = 32'b11111111111111111011111111100011;
assign LUT_2[42999] = 32'b11111111111111111000110111111100;
assign LUT_2[43000] = 32'b11111111111111110011011010011100;
assign LUT_2[43001] = 32'b11111111111111110000010010110101;
assign LUT_2[43002] = 32'b11111111111111111010010011011000;
assign LUT_2[43003] = 32'b11111111111111110111001011110001;
assign LUT_2[43004] = 32'b11111111111111101111111000000100;
assign LUT_2[43005] = 32'b11111111111111101100110000011101;
assign LUT_2[43006] = 32'b11111111111111110110110001000000;
assign LUT_2[43007] = 32'b11111111111111110011101001011001;
assign LUT_2[43008] = 32'b11111111111111101101100101111001;
assign LUT_2[43009] = 32'b11111111111111101010011110010010;
assign LUT_2[43010] = 32'b11111111111111110100011110110101;
assign LUT_2[43011] = 32'b11111111111111110001010111001110;
assign LUT_2[43012] = 32'b11111111111111101010000011100001;
assign LUT_2[43013] = 32'b11111111111111100110111011111010;
assign LUT_2[43014] = 32'b11111111111111110000111100011101;
assign LUT_2[43015] = 32'b11111111111111101101110100110110;
assign LUT_2[43016] = 32'b11111111111111101000010111010110;
assign LUT_2[43017] = 32'b11111111111111100101001111101111;
assign LUT_2[43018] = 32'b11111111111111101111010000010010;
assign LUT_2[43019] = 32'b11111111111111101100001000101011;
assign LUT_2[43020] = 32'b11111111111111100100110100111110;
assign LUT_2[43021] = 32'b11111111111111100001101101010111;
assign LUT_2[43022] = 32'b11111111111111101011101101111010;
assign LUT_2[43023] = 32'b11111111111111101000100110010011;
assign LUT_2[43024] = 32'b11111111111111101000001010000011;
assign LUT_2[43025] = 32'b11111111111111100101000010011100;
assign LUT_2[43026] = 32'b11111111111111101111000010111111;
assign LUT_2[43027] = 32'b11111111111111101011111011011000;
assign LUT_2[43028] = 32'b11111111111111100100100111101011;
assign LUT_2[43029] = 32'b11111111111111100001100000000100;
assign LUT_2[43030] = 32'b11111111111111101011100000100111;
assign LUT_2[43031] = 32'b11111111111111101000011001000000;
assign LUT_2[43032] = 32'b11111111111111100010111011100000;
assign LUT_2[43033] = 32'b11111111111111011111110011111001;
assign LUT_2[43034] = 32'b11111111111111101001110100011100;
assign LUT_2[43035] = 32'b11111111111111100110101100110101;
assign LUT_2[43036] = 32'b11111111111111011111011001001000;
assign LUT_2[43037] = 32'b11111111111111011100010001100001;
assign LUT_2[43038] = 32'b11111111111111100110010010000100;
assign LUT_2[43039] = 32'b11111111111111100011001010011101;
assign LUT_2[43040] = 32'b11111111111111101110000001100010;
assign LUT_2[43041] = 32'b11111111111111101010111001111011;
assign LUT_2[43042] = 32'b11111111111111110100111010011110;
assign LUT_2[43043] = 32'b11111111111111110001110010110111;
assign LUT_2[43044] = 32'b11111111111111101010011111001010;
assign LUT_2[43045] = 32'b11111111111111100111010111100011;
assign LUT_2[43046] = 32'b11111111111111110001011000000110;
assign LUT_2[43047] = 32'b11111111111111101110010000011111;
assign LUT_2[43048] = 32'b11111111111111101000110010111111;
assign LUT_2[43049] = 32'b11111111111111100101101011011000;
assign LUT_2[43050] = 32'b11111111111111101111101011111011;
assign LUT_2[43051] = 32'b11111111111111101100100100010100;
assign LUT_2[43052] = 32'b11111111111111100101010000100111;
assign LUT_2[43053] = 32'b11111111111111100010001001000000;
assign LUT_2[43054] = 32'b11111111111111101100001001100011;
assign LUT_2[43055] = 32'b11111111111111101001000001111100;
assign LUT_2[43056] = 32'b11111111111111101000100101101100;
assign LUT_2[43057] = 32'b11111111111111100101011110000101;
assign LUT_2[43058] = 32'b11111111111111101111011110101000;
assign LUT_2[43059] = 32'b11111111111111101100010111000001;
assign LUT_2[43060] = 32'b11111111111111100101000011010100;
assign LUT_2[43061] = 32'b11111111111111100001111011101101;
assign LUT_2[43062] = 32'b11111111111111101011111100010000;
assign LUT_2[43063] = 32'b11111111111111101000110100101001;
assign LUT_2[43064] = 32'b11111111111111100011010111001001;
assign LUT_2[43065] = 32'b11111111111111100000001111100010;
assign LUT_2[43066] = 32'b11111111111111101010010000000101;
assign LUT_2[43067] = 32'b11111111111111100111001000011110;
assign LUT_2[43068] = 32'b11111111111111011111110100110001;
assign LUT_2[43069] = 32'b11111111111111011100101101001010;
assign LUT_2[43070] = 32'b11111111111111100110101101101101;
assign LUT_2[43071] = 32'b11111111111111100011100110000110;
assign LUT_2[43072] = 32'b11111111111111100101101110011100;
assign LUT_2[43073] = 32'b11111111111111100010100110110101;
assign LUT_2[43074] = 32'b11111111111111101100100111011000;
assign LUT_2[43075] = 32'b11111111111111101001011111110001;
assign LUT_2[43076] = 32'b11111111111111100010001100000100;
assign LUT_2[43077] = 32'b11111111111111011111000100011101;
assign LUT_2[43078] = 32'b11111111111111101001000101000000;
assign LUT_2[43079] = 32'b11111111111111100101111101011001;
assign LUT_2[43080] = 32'b11111111111111100000011111111001;
assign LUT_2[43081] = 32'b11111111111111011101011000010010;
assign LUT_2[43082] = 32'b11111111111111100111011000110101;
assign LUT_2[43083] = 32'b11111111111111100100010001001110;
assign LUT_2[43084] = 32'b11111111111111011100111101100001;
assign LUT_2[43085] = 32'b11111111111111011001110101111010;
assign LUT_2[43086] = 32'b11111111111111100011110110011101;
assign LUT_2[43087] = 32'b11111111111111100000101110110110;
assign LUT_2[43088] = 32'b11111111111111100000010010100110;
assign LUT_2[43089] = 32'b11111111111111011101001010111111;
assign LUT_2[43090] = 32'b11111111111111100111001011100010;
assign LUT_2[43091] = 32'b11111111111111100100000011111011;
assign LUT_2[43092] = 32'b11111111111111011100110000001110;
assign LUT_2[43093] = 32'b11111111111111011001101000100111;
assign LUT_2[43094] = 32'b11111111111111100011101001001010;
assign LUT_2[43095] = 32'b11111111111111100000100001100011;
assign LUT_2[43096] = 32'b11111111111111011011000100000011;
assign LUT_2[43097] = 32'b11111111111111010111111100011100;
assign LUT_2[43098] = 32'b11111111111111100001111100111111;
assign LUT_2[43099] = 32'b11111111111111011110110101011000;
assign LUT_2[43100] = 32'b11111111111111010111100001101011;
assign LUT_2[43101] = 32'b11111111111111010100011010000100;
assign LUT_2[43102] = 32'b11111111111111011110011010100111;
assign LUT_2[43103] = 32'b11111111111111011011010011000000;
assign LUT_2[43104] = 32'b11111111111111100110001010000101;
assign LUT_2[43105] = 32'b11111111111111100011000010011110;
assign LUT_2[43106] = 32'b11111111111111101101000011000001;
assign LUT_2[43107] = 32'b11111111111111101001111011011010;
assign LUT_2[43108] = 32'b11111111111111100010100111101101;
assign LUT_2[43109] = 32'b11111111111111011111100000000110;
assign LUT_2[43110] = 32'b11111111111111101001100000101001;
assign LUT_2[43111] = 32'b11111111111111100110011001000010;
assign LUT_2[43112] = 32'b11111111111111100000111011100010;
assign LUT_2[43113] = 32'b11111111111111011101110011111011;
assign LUT_2[43114] = 32'b11111111111111100111110100011110;
assign LUT_2[43115] = 32'b11111111111111100100101100110111;
assign LUT_2[43116] = 32'b11111111111111011101011001001010;
assign LUT_2[43117] = 32'b11111111111111011010010001100011;
assign LUT_2[43118] = 32'b11111111111111100100010010000110;
assign LUT_2[43119] = 32'b11111111111111100001001010011111;
assign LUT_2[43120] = 32'b11111111111111100000101110001111;
assign LUT_2[43121] = 32'b11111111111111011101100110101000;
assign LUT_2[43122] = 32'b11111111111111100111100111001011;
assign LUT_2[43123] = 32'b11111111111111100100011111100100;
assign LUT_2[43124] = 32'b11111111111111011101001011110111;
assign LUT_2[43125] = 32'b11111111111111011010000100010000;
assign LUT_2[43126] = 32'b11111111111111100100000100110011;
assign LUT_2[43127] = 32'b11111111111111100000111101001100;
assign LUT_2[43128] = 32'b11111111111111011011011111101100;
assign LUT_2[43129] = 32'b11111111111111011000011000000101;
assign LUT_2[43130] = 32'b11111111111111100010011000101000;
assign LUT_2[43131] = 32'b11111111111111011111010001000001;
assign LUT_2[43132] = 32'b11111111111111010111111101010100;
assign LUT_2[43133] = 32'b11111111111111010100110101101101;
assign LUT_2[43134] = 32'b11111111111111011110110110010000;
assign LUT_2[43135] = 32'b11111111111111011011101110101001;
assign LUT_2[43136] = 32'b11111111111111110001111010001000;
assign LUT_2[43137] = 32'b11111111111111101110110010100001;
assign LUT_2[43138] = 32'b11111111111111111000110011000100;
assign LUT_2[43139] = 32'b11111111111111110101101011011101;
assign LUT_2[43140] = 32'b11111111111111101110010111110000;
assign LUT_2[43141] = 32'b11111111111111101011010000001001;
assign LUT_2[43142] = 32'b11111111111111110101010000101100;
assign LUT_2[43143] = 32'b11111111111111110010001001000101;
assign LUT_2[43144] = 32'b11111111111111101100101011100101;
assign LUT_2[43145] = 32'b11111111111111101001100011111110;
assign LUT_2[43146] = 32'b11111111111111110011100100100001;
assign LUT_2[43147] = 32'b11111111111111110000011100111010;
assign LUT_2[43148] = 32'b11111111111111101001001001001101;
assign LUT_2[43149] = 32'b11111111111111100110000001100110;
assign LUT_2[43150] = 32'b11111111111111110000000010001001;
assign LUT_2[43151] = 32'b11111111111111101100111010100010;
assign LUT_2[43152] = 32'b11111111111111101100011110010010;
assign LUT_2[43153] = 32'b11111111111111101001010110101011;
assign LUT_2[43154] = 32'b11111111111111110011010111001110;
assign LUT_2[43155] = 32'b11111111111111110000001111100111;
assign LUT_2[43156] = 32'b11111111111111101000111011111010;
assign LUT_2[43157] = 32'b11111111111111100101110100010011;
assign LUT_2[43158] = 32'b11111111111111101111110100110110;
assign LUT_2[43159] = 32'b11111111111111101100101101001111;
assign LUT_2[43160] = 32'b11111111111111100111001111101111;
assign LUT_2[43161] = 32'b11111111111111100100001000001000;
assign LUT_2[43162] = 32'b11111111111111101110001000101011;
assign LUT_2[43163] = 32'b11111111111111101011000001000100;
assign LUT_2[43164] = 32'b11111111111111100011101101010111;
assign LUT_2[43165] = 32'b11111111111111100000100101110000;
assign LUT_2[43166] = 32'b11111111111111101010100110010011;
assign LUT_2[43167] = 32'b11111111111111100111011110101100;
assign LUT_2[43168] = 32'b11111111111111110010010101110001;
assign LUT_2[43169] = 32'b11111111111111101111001110001010;
assign LUT_2[43170] = 32'b11111111111111111001001110101101;
assign LUT_2[43171] = 32'b11111111111111110110000111000110;
assign LUT_2[43172] = 32'b11111111111111101110110011011001;
assign LUT_2[43173] = 32'b11111111111111101011101011110010;
assign LUT_2[43174] = 32'b11111111111111110101101100010101;
assign LUT_2[43175] = 32'b11111111111111110010100100101110;
assign LUT_2[43176] = 32'b11111111111111101101000111001110;
assign LUT_2[43177] = 32'b11111111111111101001111111100111;
assign LUT_2[43178] = 32'b11111111111111110100000000001010;
assign LUT_2[43179] = 32'b11111111111111110000111000100011;
assign LUT_2[43180] = 32'b11111111111111101001100100110110;
assign LUT_2[43181] = 32'b11111111111111100110011101001111;
assign LUT_2[43182] = 32'b11111111111111110000011101110010;
assign LUT_2[43183] = 32'b11111111111111101101010110001011;
assign LUT_2[43184] = 32'b11111111111111101100111001111011;
assign LUT_2[43185] = 32'b11111111111111101001110010010100;
assign LUT_2[43186] = 32'b11111111111111110011110010110111;
assign LUT_2[43187] = 32'b11111111111111110000101011010000;
assign LUT_2[43188] = 32'b11111111111111101001010111100011;
assign LUT_2[43189] = 32'b11111111111111100110001111111100;
assign LUT_2[43190] = 32'b11111111111111110000010000011111;
assign LUT_2[43191] = 32'b11111111111111101101001000111000;
assign LUT_2[43192] = 32'b11111111111111100111101011011000;
assign LUT_2[43193] = 32'b11111111111111100100100011110001;
assign LUT_2[43194] = 32'b11111111111111101110100100010100;
assign LUT_2[43195] = 32'b11111111111111101011011100101101;
assign LUT_2[43196] = 32'b11111111111111100100001001000000;
assign LUT_2[43197] = 32'b11111111111111100001000001011001;
assign LUT_2[43198] = 32'b11111111111111101011000001111100;
assign LUT_2[43199] = 32'b11111111111111100111111010010101;
assign LUT_2[43200] = 32'b11111111111111101010000010101011;
assign LUT_2[43201] = 32'b11111111111111100110111011000100;
assign LUT_2[43202] = 32'b11111111111111110000111011100111;
assign LUT_2[43203] = 32'b11111111111111101101110100000000;
assign LUT_2[43204] = 32'b11111111111111100110100000010011;
assign LUT_2[43205] = 32'b11111111111111100011011000101100;
assign LUT_2[43206] = 32'b11111111111111101101011001001111;
assign LUT_2[43207] = 32'b11111111111111101010010001101000;
assign LUT_2[43208] = 32'b11111111111111100100110100001000;
assign LUT_2[43209] = 32'b11111111111111100001101100100001;
assign LUT_2[43210] = 32'b11111111111111101011101101000100;
assign LUT_2[43211] = 32'b11111111111111101000100101011101;
assign LUT_2[43212] = 32'b11111111111111100001010001110000;
assign LUT_2[43213] = 32'b11111111111111011110001010001001;
assign LUT_2[43214] = 32'b11111111111111101000001010101100;
assign LUT_2[43215] = 32'b11111111111111100101000011000101;
assign LUT_2[43216] = 32'b11111111111111100100100110110101;
assign LUT_2[43217] = 32'b11111111111111100001011111001110;
assign LUT_2[43218] = 32'b11111111111111101011011111110001;
assign LUT_2[43219] = 32'b11111111111111101000011000001010;
assign LUT_2[43220] = 32'b11111111111111100001000100011101;
assign LUT_2[43221] = 32'b11111111111111011101111100110110;
assign LUT_2[43222] = 32'b11111111111111100111111101011001;
assign LUT_2[43223] = 32'b11111111111111100100110101110010;
assign LUT_2[43224] = 32'b11111111111111011111011000010010;
assign LUT_2[43225] = 32'b11111111111111011100010000101011;
assign LUT_2[43226] = 32'b11111111111111100110010001001110;
assign LUT_2[43227] = 32'b11111111111111100011001001100111;
assign LUT_2[43228] = 32'b11111111111111011011110101111010;
assign LUT_2[43229] = 32'b11111111111111011000101110010011;
assign LUT_2[43230] = 32'b11111111111111100010101110110110;
assign LUT_2[43231] = 32'b11111111111111011111100111001111;
assign LUT_2[43232] = 32'b11111111111111101010011110010100;
assign LUT_2[43233] = 32'b11111111111111100111010110101101;
assign LUT_2[43234] = 32'b11111111111111110001010111010000;
assign LUT_2[43235] = 32'b11111111111111101110001111101001;
assign LUT_2[43236] = 32'b11111111111111100110111011111100;
assign LUT_2[43237] = 32'b11111111111111100011110100010101;
assign LUT_2[43238] = 32'b11111111111111101101110100111000;
assign LUT_2[43239] = 32'b11111111111111101010101101010001;
assign LUT_2[43240] = 32'b11111111111111100101001111110001;
assign LUT_2[43241] = 32'b11111111111111100010001000001010;
assign LUT_2[43242] = 32'b11111111111111101100001000101101;
assign LUT_2[43243] = 32'b11111111111111101001000001000110;
assign LUT_2[43244] = 32'b11111111111111100001101101011001;
assign LUT_2[43245] = 32'b11111111111111011110100101110010;
assign LUT_2[43246] = 32'b11111111111111101000100110010101;
assign LUT_2[43247] = 32'b11111111111111100101011110101110;
assign LUT_2[43248] = 32'b11111111111111100101000010011110;
assign LUT_2[43249] = 32'b11111111111111100001111010110111;
assign LUT_2[43250] = 32'b11111111111111101011111011011010;
assign LUT_2[43251] = 32'b11111111111111101000110011110011;
assign LUT_2[43252] = 32'b11111111111111100001100000000110;
assign LUT_2[43253] = 32'b11111111111111011110011000011111;
assign LUT_2[43254] = 32'b11111111111111101000011001000010;
assign LUT_2[43255] = 32'b11111111111111100101010001011011;
assign LUT_2[43256] = 32'b11111111111111011111110011111011;
assign LUT_2[43257] = 32'b11111111111111011100101100010100;
assign LUT_2[43258] = 32'b11111111111111100110101100110111;
assign LUT_2[43259] = 32'b11111111111111100011100101010000;
assign LUT_2[43260] = 32'b11111111111111011100010001100011;
assign LUT_2[43261] = 32'b11111111111111011001001001111100;
assign LUT_2[43262] = 32'b11111111111111100011001010011111;
assign LUT_2[43263] = 32'b11111111111111100000000010111000;
assign LUT_2[43264] = 32'b11111111111111110001100100011111;
assign LUT_2[43265] = 32'b11111111111111101110011100111000;
assign LUT_2[43266] = 32'b11111111111111111000011101011011;
assign LUT_2[43267] = 32'b11111111111111110101010101110100;
assign LUT_2[43268] = 32'b11111111111111101110000010000111;
assign LUT_2[43269] = 32'b11111111111111101010111010100000;
assign LUT_2[43270] = 32'b11111111111111110100111011000011;
assign LUT_2[43271] = 32'b11111111111111110001110011011100;
assign LUT_2[43272] = 32'b11111111111111101100010101111100;
assign LUT_2[43273] = 32'b11111111111111101001001110010101;
assign LUT_2[43274] = 32'b11111111111111110011001110111000;
assign LUT_2[43275] = 32'b11111111111111110000000111010001;
assign LUT_2[43276] = 32'b11111111111111101000110011100100;
assign LUT_2[43277] = 32'b11111111111111100101101011111101;
assign LUT_2[43278] = 32'b11111111111111101111101100100000;
assign LUT_2[43279] = 32'b11111111111111101100100100111001;
assign LUT_2[43280] = 32'b11111111111111101100001000101001;
assign LUT_2[43281] = 32'b11111111111111101001000001000010;
assign LUT_2[43282] = 32'b11111111111111110011000001100101;
assign LUT_2[43283] = 32'b11111111111111101111111001111110;
assign LUT_2[43284] = 32'b11111111111111101000100110010001;
assign LUT_2[43285] = 32'b11111111111111100101011110101010;
assign LUT_2[43286] = 32'b11111111111111101111011111001101;
assign LUT_2[43287] = 32'b11111111111111101100010111100110;
assign LUT_2[43288] = 32'b11111111111111100110111010000110;
assign LUT_2[43289] = 32'b11111111111111100011110010011111;
assign LUT_2[43290] = 32'b11111111111111101101110011000010;
assign LUT_2[43291] = 32'b11111111111111101010101011011011;
assign LUT_2[43292] = 32'b11111111111111100011010111101110;
assign LUT_2[43293] = 32'b11111111111111100000010000000111;
assign LUT_2[43294] = 32'b11111111111111101010010000101010;
assign LUT_2[43295] = 32'b11111111111111100111001001000011;
assign LUT_2[43296] = 32'b11111111111111110010000000001000;
assign LUT_2[43297] = 32'b11111111111111101110111000100001;
assign LUT_2[43298] = 32'b11111111111111111000111001000100;
assign LUT_2[43299] = 32'b11111111111111110101110001011101;
assign LUT_2[43300] = 32'b11111111111111101110011101110000;
assign LUT_2[43301] = 32'b11111111111111101011010110001001;
assign LUT_2[43302] = 32'b11111111111111110101010110101100;
assign LUT_2[43303] = 32'b11111111111111110010001111000101;
assign LUT_2[43304] = 32'b11111111111111101100110001100101;
assign LUT_2[43305] = 32'b11111111111111101001101001111110;
assign LUT_2[43306] = 32'b11111111111111110011101010100001;
assign LUT_2[43307] = 32'b11111111111111110000100010111010;
assign LUT_2[43308] = 32'b11111111111111101001001111001101;
assign LUT_2[43309] = 32'b11111111111111100110000111100110;
assign LUT_2[43310] = 32'b11111111111111110000001000001001;
assign LUT_2[43311] = 32'b11111111111111101101000000100010;
assign LUT_2[43312] = 32'b11111111111111101100100100010010;
assign LUT_2[43313] = 32'b11111111111111101001011100101011;
assign LUT_2[43314] = 32'b11111111111111110011011101001110;
assign LUT_2[43315] = 32'b11111111111111110000010101100111;
assign LUT_2[43316] = 32'b11111111111111101001000001111010;
assign LUT_2[43317] = 32'b11111111111111100101111010010011;
assign LUT_2[43318] = 32'b11111111111111101111111010110110;
assign LUT_2[43319] = 32'b11111111111111101100110011001111;
assign LUT_2[43320] = 32'b11111111111111100111010101101111;
assign LUT_2[43321] = 32'b11111111111111100100001110001000;
assign LUT_2[43322] = 32'b11111111111111101110001110101011;
assign LUT_2[43323] = 32'b11111111111111101011000111000100;
assign LUT_2[43324] = 32'b11111111111111100011110011010111;
assign LUT_2[43325] = 32'b11111111111111100000101011110000;
assign LUT_2[43326] = 32'b11111111111111101010101100010011;
assign LUT_2[43327] = 32'b11111111111111100111100100101100;
assign LUT_2[43328] = 32'b11111111111111101001101101000010;
assign LUT_2[43329] = 32'b11111111111111100110100101011011;
assign LUT_2[43330] = 32'b11111111111111110000100101111110;
assign LUT_2[43331] = 32'b11111111111111101101011110010111;
assign LUT_2[43332] = 32'b11111111111111100110001010101010;
assign LUT_2[43333] = 32'b11111111111111100011000011000011;
assign LUT_2[43334] = 32'b11111111111111101101000011100110;
assign LUT_2[43335] = 32'b11111111111111101001111011111111;
assign LUT_2[43336] = 32'b11111111111111100100011110011111;
assign LUT_2[43337] = 32'b11111111111111100001010110111000;
assign LUT_2[43338] = 32'b11111111111111101011010111011011;
assign LUT_2[43339] = 32'b11111111111111101000001111110100;
assign LUT_2[43340] = 32'b11111111111111100000111100000111;
assign LUT_2[43341] = 32'b11111111111111011101110100100000;
assign LUT_2[43342] = 32'b11111111111111100111110101000011;
assign LUT_2[43343] = 32'b11111111111111100100101101011100;
assign LUT_2[43344] = 32'b11111111111111100100010001001100;
assign LUT_2[43345] = 32'b11111111111111100001001001100101;
assign LUT_2[43346] = 32'b11111111111111101011001010001000;
assign LUT_2[43347] = 32'b11111111111111101000000010100001;
assign LUT_2[43348] = 32'b11111111111111100000101110110100;
assign LUT_2[43349] = 32'b11111111111111011101100111001101;
assign LUT_2[43350] = 32'b11111111111111100111100111110000;
assign LUT_2[43351] = 32'b11111111111111100100100000001001;
assign LUT_2[43352] = 32'b11111111111111011111000010101001;
assign LUT_2[43353] = 32'b11111111111111011011111011000010;
assign LUT_2[43354] = 32'b11111111111111100101111011100101;
assign LUT_2[43355] = 32'b11111111111111100010110011111110;
assign LUT_2[43356] = 32'b11111111111111011011100000010001;
assign LUT_2[43357] = 32'b11111111111111011000011000101010;
assign LUT_2[43358] = 32'b11111111111111100010011001001101;
assign LUT_2[43359] = 32'b11111111111111011111010001100110;
assign LUT_2[43360] = 32'b11111111111111101010001000101011;
assign LUT_2[43361] = 32'b11111111111111100111000001000100;
assign LUT_2[43362] = 32'b11111111111111110001000001100111;
assign LUT_2[43363] = 32'b11111111111111101101111010000000;
assign LUT_2[43364] = 32'b11111111111111100110100110010011;
assign LUT_2[43365] = 32'b11111111111111100011011110101100;
assign LUT_2[43366] = 32'b11111111111111101101011111001111;
assign LUT_2[43367] = 32'b11111111111111101010010111101000;
assign LUT_2[43368] = 32'b11111111111111100100111010001000;
assign LUT_2[43369] = 32'b11111111111111100001110010100001;
assign LUT_2[43370] = 32'b11111111111111101011110011000100;
assign LUT_2[43371] = 32'b11111111111111101000101011011101;
assign LUT_2[43372] = 32'b11111111111111100001010111110000;
assign LUT_2[43373] = 32'b11111111111111011110010000001001;
assign LUT_2[43374] = 32'b11111111111111101000010000101100;
assign LUT_2[43375] = 32'b11111111111111100101001001000101;
assign LUT_2[43376] = 32'b11111111111111100100101100110101;
assign LUT_2[43377] = 32'b11111111111111100001100101001110;
assign LUT_2[43378] = 32'b11111111111111101011100101110001;
assign LUT_2[43379] = 32'b11111111111111101000011110001010;
assign LUT_2[43380] = 32'b11111111111111100001001010011101;
assign LUT_2[43381] = 32'b11111111111111011110000010110110;
assign LUT_2[43382] = 32'b11111111111111101000000011011001;
assign LUT_2[43383] = 32'b11111111111111100100111011110010;
assign LUT_2[43384] = 32'b11111111111111011111011110010010;
assign LUT_2[43385] = 32'b11111111111111011100010110101011;
assign LUT_2[43386] = 32'b11111111111111100110010111001110;
assign LUT_2[43387] = 32'b11111111111111100011001111100111;
assign LUT_2[43388] = 32'b11111111111111011011111011111010;
assign LUT_2[43389] = 32'b11111111111111011000110100010011;
assign LUT_2[43390] = 32'b11111111111111100010110100110110;
assign LUT_2[43391] = 32'b11111111111111011111101101001111;
assign LUT_2[43392] = 32'b11111111111111110101111000101110;
assign LUT_2[43393] = 32'b11111111111111110010110001000111;
assign LUT_2[43394] = 32'b11111111111111111100110001101010;
assign LUT_2[43395] = 32'b11111111111111111001101010000011;
assign LUT_2[43396] = 32'b11111111111111110010010110010110;
assign LUT_2[43397] = 32'b11111111111111101111001110101111;
assign LUT_2[43398] = 32'b11111111111111111001001111010010;
assign LUT_2[43399] = 32'b11111111111111110110000111101011;
assign LUT_2[43400] = 32'b11111111111111110000101010001011;
assign LUT_2[43401] = 32'b11111111111111101101100010100100;
assign LUT_2[43402] = 32'b11111111111111110111100011000111;
assign LUT_2[43403] = 32'b11111111111111110100011011100000;
assign LUT_2[43404] = 32'b11111111111111101101000111110011;
assign LUT_2[43405] = 32'b11111111111111101010000000001100;
assign LUT_2[43406] = 32'b11111111111111110100000000101111;
assign LUT_2[43407] = 32'b11111111111111110000111001001000;
assign LUT_2[43408] = 32'b11111111111111110000011100111000;
assign LUT_2[43409] = 32'b11111111111111101101010101010001;
assign LUT_2[43410] = 32'b11111111111111110111010101110100;
assign LUT_2[43411] = 32'b11111111111111110100001110001101;
assign LUT_2[43412] = 32'b11111111111111101100111010100000;
assign LUT_2[43413] = 32'b11111111111111101001110010111001;
assign LUT_2[43414] = 32'b11111111111111110011110011011100;
assign LUT_2[43415] = 32'b11111111111111110000101011110101;
assign LUT_2[43416] = 32'b11111111111111101011001110010101;
assign LUT_2[43417] = 32'b11111111111111101000000110101110;
assign LUT_2[43418] = 32'b11111111111111110010000111010001;
assign LUT_2[43419] = 32'b11111111111111101110111111101010;
assign LUT_2[43420] = 32'b11111111111111100111101011111101;
assign LUT_2[43421] = 32'b11111111111111100100100100010110;
assign LUT_2[43422] = 32'b11111111111111101110100100111001;
assign LUT_2[43423] = 32'b11111111111111101011011101010010;
assign LUT_2[43424] = 32'b11111111111111110110010100010111;
assign LUT_2[43425] = 32'b11111111111111110011001100110000;
assign LUT_2[43426] = 32'b11111111111111111101001101010011;
assign LUT_2[43427] = 32'b11111111111111111010000101101100;
assign LUT_2[43428] = 32'b11111111111111110010110001111111;
assign LUT_2[43429] = 32'b11111111111111101111101010011000;
assign LUT_2[43430] = 32'b11111111111111111001101010111011;
assign LUT_2[43431] = 32'b11111111111111110110100011010100;
assign LUT_2[43432] = 32'b11111111111111110001000101110100;
assign LUT_2[43433] = 32'b11111111111111101101111110001101;
assign LUT_2[43434] = 32'b11111111111111110111111110110000;
assign LUT_2[43435] = 32'b11111111111111110100110111001001;
assign LUT_2[43436] = 32'b11111111111111101101100011011100;
assign LUT_2[43437] = 32'b11111111111111101010011011110101;
assign LUT_2[43438] = 32'b11111111111111110100011100011000;
assign LUT_2[43439] = 32'b11111111111111110001010100110001;
assign LUT_2[43440] = 32'b11111111111111110000111000100001;
assign LUT_2[43441] = 32'b11111111111111101101110000111010;
assign LUT_2[43442] = 32'b11111111111111110111110001011101;
assign LUT_2[43443] = 32'b11111111111111110100101001110110;
assign LUT_2[43444] = 32'b11111111111111101101010110001001;
assign LUT_2[43445] = 32'b11111111111111101010001110100010;
assign LUT_2[43446] = 32'b11111111111111110100001111000101;
assign LUT_2[43447] = 32'b11111111111111110001000111011110;
assign LUT_2[43448] = 32'b11111111111111101011101001111110;
assign LUT_2[43449] = 32'b11111111111111101000100010010111;
assign LUT_2[43450] = 32'b11111111111111110010100010111010;
assign LUT_2[43451] = 32'b11111111111111101111011011010011;
assign LUT_2[43452] = 32'b11111111111111101000000111100110;
assign LUT_2[43453] = 32'b11111111111111100100111111111111;
assign LUT_2[43454] = 32'b11111111111111101111000000100010;
assign LUT_2[43455] = 32'b11111111111111101011111000111011;
assign LUT_2[43456] = 32'b11111111111111101110000001010001;
assign LUT_2[43457] = 32'b11111111111111101010111001101010;
assign LUT_2[43458] = 32'b11111111111111110100111010001101;
assign LUT_2[43459] = 32'b11111111111111110001110010100110;
assign LUT_2[43460] = 32'b11111111111111101010011110111001;
assign LUT_2[43461] = 32'b11111111111111100111010111010010;
assign LUT_2[43462] = 32'b11111111111111110001010111110101;
assign LUT_2[43463] = 32'b11111111111111101110010000001110;
assign LUT_2[43464] = 32'b11111111111111101000110010101110;
assign LUT_2[43465] = 32'b11111111111111100101101011000111;
assign LUT_2[43466] = 32'b11111111111111101111101011101010;
assign LUT_2[43467] = 32'b11111111111111101100100100000011;
assign LUT_2[43468] = 32'b11111111111111100101010000010110;
assign LUT_2[43469] = 32'b11111111111111100010001000101111;
assign LUT_2[43470] = 32'b11111111111111101100001001010010;
assign LUT_2[43471] = 32'b11111111111111101001000001101011;
assign LUT_2[43472] = 32'b11111111111111101000100101011011;
assign LUT_2[43473] = 32'b11111111111111100101011101110100;
assign LUT_2[43474] = 32'b11111111111111101111011110010111;
assign LUT_2[43475] = 32'b11111111111111101100010110110000;
assign LUT_2[43476] = 32'b11111111111111100101000011000011;
assign LUT_2[43477] = 32'b11111111111111100001111011011100;
assign LUT_2[43478] = 32'b11111111111111101011111011111111;
assign LUT_2[43479] = 32'b11111111111111101000110100011000;
assign LUT_2[43480] = 32'b11111111111111100011010110111000;
assign LUT_2[43481] = 32'b11111111111111100000001111010001;
assign LUT_2[43482] = 32'b11111111111111101010001111110100;
assign LUT_2[43483] = 32'b11111111111111100111001000001101;
assign LUT_2[43484] = 32'b11111111111111011111110100100000;
assign LUT_2[43485] = 32'b11111111111111011100101100111001;
assign LUT_2[43486] = 32'b11111111111111100110101101011100;
assign LUT_2[43487] = 32'b11111111111111100011100101110101;
assign LUT_2[43488] = 32'b11111111111111101110011100111010;
assign LUT_2[43489] = 32'b11111111111111101011010101010011;
assign LUT_2[43490] = 32'b11111111111111110101010101110110;
assign LUT_2[43491] = 32'b11111111111111110010001110001111;
assign LUT_2[43492] = 32'b11111111111111101010111010100010;
assign LUT_2[43493] = 32'b11111111111111100111110010111011;
assign LUT_2[43494] = 32'b11111111111111110001110011011110;
assign LUT_2[43495] = 32'b11111111111111101110101011110111;
assign LUT_2[43496] = 32'b11111111111111101001001110010111;
assign LUT_2[43497] = 32'b11111111111111100110000110110000;
assign LUT_2[43498] = 32'b11111111111111110000000111010011;
assign LUT_2[43499] = 32'b11111111111111101100111111101100;
assign LUT_2[43500] = 32'b11111111111111100101101011111111;
assign LUT_2[43501] = 32'b11111111111111100010100100011000;
assign LUT_2[43502] = 32'b11111111111111101100100100111011;
assign LUT_2[43503] = 32'b11111111111111101001011101010100;
assign LUT_2[43504] = 32'b11111111111111101001000001000100;
assign LUT_2[43505] = 32'b11111111111111100101111001011101;
assign LUT_2[43506] = 32'b11111111111111101111111010000000;
assign LUT_2[43507] = 32'b11111111111111101100110010011001;
assign LUT_2[43508] = 32'b11111111111111100101011110101100;
assign LUT_2[43509] = 32'b11111111111111100010010111000101;
assign LUT_2[43510] = 32'b11111111111111101100010111101000;
assign LUT_2[43511] = 32'b11111111111111101001010000000001;
assign LUT_2[43512] = 32'b11111111111111100011110010100001;
assign LUT_2[43513] = 32'b11111111111111100000101010111010;
assign LUT_2[43514] = 32'b11111111111111101010101011011101;
assign LUT_2[43515] = 32'b11111111111111100111100011110110;
assign LUT_2[43516] = 32'b11111111111111100000010000001001;
assign LUT_2[43517] = 32'b11111111111111011101001000100010;
assign LUT_2[43518] = 32'b11111111111111100111001001000101;
assign LUT_2[43519] = 32'b11111111111111100100000001011110;
assign LUT_2[43520] = 32'b11111111111111110010010111101011;
assign LUT_2[43521] = 32'b11111111111111101111010000000100;
assign LUT_2[43522] = 32'b11111111111111111001010000100111;
assign LUT_2[43523] = 32'b11111111111111110110001001000000;
assign LUT_2[43524] = 32'b11111111111111101110110101010011;
assign LUT_2[43525] = 32'b11111111111111101011101101101100;
assign LUT_2[43526] = 32'b11111111111111110101101110001111;
assign LUT_2[43527] = 32'b11111111111111110010100110101000;
assign LUT_2[43528] = 32'b11111111111111101101001001001000;
assign LUT_2[43529] = 32'b11111111111111101010000001100001;
assign LUT_2[43530] = 32'b11111111111111110100000010000100;
assign LUT_2[43531] = 32'b11111111111111110000111010011101;
assign LUT_2[43532] = 32'b11111111111111101001100110110000;
assign LUT_2[43533] = 32'b11111111111111100110011111001001;
assign LUT_2[43534] = 32'b11111111111111110000011111101100;
assign LUT_2[43535] = 32'b11111111111111101101011000000101;
assign LUT_2[43536] = 32'b11111111111111101100111011110101;
assign LUT_2[43537] = 32'b11111111111111101001110100001110;
assign LUT_2[43538] = 32'b11111111111111110011110100110001;
assign LUT_2[43539] = 32'b11111111111111110000101101001010;
assign LUT_2[43540] = 32'b11111111111111101001011001011101;
assign LUT_2[43541] = 32'b11111111111111100110010001110110;
assign LUT_2[43542] = 32'b11111111111111110000010010011001;
assign LUT_2[43543] = 32'b11111111111111101101001010110010;
assign LUT_2[43544] = 32'b11111111111111100111101101010010;
assign LUT_2[43545] = 32'b11111111111111100100100101101011;
assign LUT_2[43546] = 32'b11111111111111101110100110001110;
assign LUT_2[43547] = 32'b11111111111111101011011110100111;
assign LUT_2[43548] = 32'b11111111111111100100001010111010;
assign LUT_2[43549] = 32'b11111111111111100001000011010011;
assign LUT_2[43550] = 32'b11111111111111101011000011110110;
assign LUT_2[43551] = 32'b11111111111111100111111100001111;
assign LUT_2[43552] = 32'b11111111111111110010110011010100;
assign LUT_2[43553] = 32'b11111111111111101111101011101101;
assign LUT_2[43554] = 32'b11111111111111111001101100010000;
assign LUT_2[43555] = 32'b11111111111111110110100100101001;
assign LUT_2[43556] = 32'b11111111111111101111010000111100;
assign LUT_2[43557] = 32'b11111111111111101100001001010101;
assign LUT_2[43558] = 32'b11111111111111110110001001111000;
assign LUT_2[43559] = 32'b11111111111111110011000010010001;
assign LUT_2[43560] = 32'b11111111111111101101100100110001;
assign LUT_2[43561] = 32'b11111111111111101010011101001010;
assign LUT_2[43562] = 32'b11111111111111110100011101101101;
assign LUT_2[43563] = 32'b11111111111111110001010110000110;
assign LUT_2[43564] = 32'b11111111111111101010000010011001;
assign LUT_2[43565] = 32'b11111111111111100110111010110010;
assign LUT_2[43566] = 32'b11111111111111110000111011010101;
assign LUT_2[43567] = 32'b11111111111111101101110011101110;
assign LUT_2[43568] = 32'b11111111111111101101010111011110;
assign LUT_2[43569] = 32'b11111111111111101010001111110111;
assign LUT_2[43570] = 32'b11111111111111110100010000011010;
assign LUT_2[43571] = 32'b11111111111111110001001000110011;
assign LUT_2[43572] = 32'b11111111111111101001110101000110;
assign LUT_2[43573] = 32'b11111111111111100110101101011111;
assign LUT_2[43574] = 32'b11111111111111110000101110000010;
assign LUT_2[43575] = 32'b11111111111111101101100110011011;
assign LUT_2[43576] = 32'b11111111111111101000001000111011;
assign LUT_2[43577] = 32'b11111111111111100101000001010100;
assign LUT_2[43578] = 32'b11111111111111101111000001110111;
assign LUT_2[43579] = 32'b11111111111111101011111010010000;
assign LUT_2[43580] = 32'b11111111111111100100100110100011;
assign LUT_2[43581] = 32'b11111111111111100001011110111100;
assign LUT_2[43582] = 32'b11111111111111101011011111011111;
assign LUT_2[43583] = 32'b11111111111111101000010111111000;
assign LUT_2[43584] = 32'b11111111111111101010100000001110;
assign LUT_2[43585] = 32'b11111111111111100111011000100111;
assign LUT_2[43586] = 32'b11111111111111110001011001001010;
assign LUT_2[43587] = 32'b11111111111111101110010001100011;
assign LUT_2[43588] = 32'b11111111111111100110111101110110;
assign LUT_2[43589] = 32'b11111111111111100011110110001111;
assign LUT_2[43590] = 32'b11111111111111101101110110110010;
assign LUT_2[43591] = 32'b11111111111111101010101111001011;
assign LUT_2[43592] = 32'b11111111111111100101010001101011;
assign LUT_2[43593] = 32'b11111111111111100010001010000100;
assign LUT_2[43594] = 32'b11111111111111101100001010100111;
assign LUT_2[43595] = 32'b11111111111111101001000011000000;
assign LUT_2[43596] = 32'b11111111111111100001101111010011;
assign LUT_2[43597] = 32'b11111111111111011110100111101100;
assign LUT_2[43598] = 32'b11111111111111101000101000001111;
assign LUT_2[43599] = 32'b11111111111111100101100000101000;
assign LUT_2[43600] = 32'b11111111111111100101000100011000;
assign LUT_2[43601] = 32'b11111111111111100001111100110001;
assign LUT_2[43602] = 32'b11111111111111101011111101010100;
assign LUT_2[43603] = 32'b11111111111111101000110101101101;
assign LUT_2[43604] = 32'b11111111111111100001100010000000;
assign LUT_2[43605] = 32'b11111111111111011110011010011001;
assign LUT_2[43606] = 32'b11111111111111101000011010111100;
assign LUT_2[43607] = 32'b11111111111111100101010011010101;
assign LUT_2[43608] = 32'b11111111111111011111110101110101;
assign LUT_2[43609] = 32'b11111111111111011100101110001110;
assign LUT_2[43610] = 32'b11111111111111100110101110110001;
assign LUT_2[43611] = 32'b11111111111111100011100111001010;
assign LUT_2[43612] = 32'b11111111111111011100010011011101;
assign LUT_2[43613] = 32'b11111111111111011001001011110110;
assign LUT_2[43614] = 32'b11111111111111100011001100011001;
assign LUT_2[43615] = 32'b11111111111111100000000100110010;
assign LUT_2[43616] = 32'b11111111111111101010111011110111;
assign LUT_2[43617] = 32'b11111111111111100111110100010000;
assign LUT_2[43618] = 32'b11111111111111110001110100110011;
assign LUT_2[43619] = 32'b11111111111111101110101101001100;
assign LUT_2[43620] = 32'b11111111111111100111011001011111;
assign LUT_2[43621] = 32'b11111111111111100100010001111000;
assign LUT_2[43622] = 32'b11111111111111101110010010011011;
assign LUT_2[43623] = 32'b11111111111111101011001010110100;
assign LUT_2[43624] = 32'b11111111111111100101101101010100;
assign LUT_2[43625] = 32'b11111111111111100010100101101101;
assign LUT_2[43626] = 32'b11111111111111101100100110010000;
assign LUT_2[43627] = 32'b11111111111111101001011110101001;
assign LUT_2[43628] = 32'b11111111111111100010001010111100;
assign LUT_2[43629] = 32'b11111111111111011111000011010101;
assign LUT_2[43630] = 32'b11111111111111101001000011111000;
assign LUT_2[43631] = 32'b11111111111111100101111100010001;
assign LUT_2[43632] = 32'b11111111111111100101100000000001;
assign LUT_2[43633] = 32'b11111111111111100010011000011010;
assign LUT_2[43634] = 32'b11111111111111101100011000111101;
assign LUT_2[43635] = 32'b11111111111111101001010001010110;
assign LUT_2[43636] = 32'b11111111111111100001111101101001;
assign LUT_2[43637] = 32'b11111111111111011110110110000010;
assign LUT_2[43638] = 32'b11111111111111101000110110100101;
assign LUT_2[43639] = 32'b11111111111111100101101110111110;
assign LUT_2[43640] = 32'b11111111111111100000010001011110;
assign LUT_2[43641] = 32'b11111111111111011101001001110111;
assign LUT_2[43642] = 32'b11111111111111100111001010011010;
assign LUT_2[43643] = 32'b11111111111111100100000010110011;
assign LUT_2[43644] = 32'b11111111111111011100101111000110;
assign LUT_2[43645] = 32'b11111111111111011001100111011111;
assign LUT_2[43646] = 32'b11111111111111100011101000000010;
assign LUT_2[43647] = 32'b11111111111111100000100000011011;
assign LUT_2[43648] = 32'b11111111111111110110101011111010;
assign LUT_2[43649] = 32'b11111111111111110011100100010011;
assign LUT_2[43650] = 32'b11111111111111111101100100110110;
assign LUT_2[43651] = 32'b11111111111111111010011101001111;
assign LUT_2[43652] = 32'b11111111111111110011001001100010;
assign LUT_2[43653] = 32'b11111111111111110000000001111011;
assign LUT_2[43654] = 32'b11111111111111111010000010011110;
assign LUT_2[43655] = 32'b11111111111111110110111010110111;
assign LUT_2[43656] = 32'b11111111111111110001011101010111;
assign LUT_2[43657] = 32'b11111111111111101110010101110000;
assign LUT_2[43658] = 32'b11111111111111111000010110010011;
assign LUT_2[43659] = 32'b11111111111111110101001110101100;
assign LUT_2[43660] = 32'b11111111111111101101111010111111;
assign LUT_2[43661] = 32'b11111111111111101010110011011000;
assign LUT_2[43662] = 32'b11111111111111110100110011111011;
assign LUT_2[43663] = 32'b11111111111111110001101100010100;
assign LUT_2[43664] = 32'b11111111111111110001010000000100;
assign LUT_2[43665] = 32'b11111111111111101110001000011101;
assign LUT_2[43666] = 32'b11111111111111111000001001000000;
assign LUT_2[43667] = 32'b11111111111111110101000001011001;
assign LUT_2[43668] = 32'b11111111111111101101101101101100;
assign LUT_2[43669] = 32'b11111111111111101010100110000101;
assign LUT_2[43670] = 32'b11111111111111110100100110101000;
assign LUT_2[43671] = 32'b11111111111111110001011111000001;
assign LUT_2[43672] = 32'b11111111111111101100000001100001;
assign LUT_2[43673] = 32'b11111111111111101000111001111010;
assign LUT_2[43674] = 32'b11111111111111110010111010011101;
assign LUT_2[43675] = 32'b11111111111111101111110010110110;
assign LUT_2[43676] = 32'b11111111111111101000011111001001;
assign LUT_2[43677] = 32'b11111111111111100101010111100010;
assign LUT_2[43678] = 32'b11111111111111101111011000000101;
assign LUT_2[43679] = 32'b11111111111111101100010000011110;
assign LUT_2[43680] = 32'b11111111111111110111000111100011;
assign LUT_2[43681] = 32'b11111111111111110011111111111100;
assign LUT_2[43682] = 32'b11111111111111111110000000011111;
assign LUT_2[43683] = 32'b11111111111111111010111000111000;
assign LUT_2[43684] = 32'b11111111111111110011100101001011;
assign LUT_2[43685] = 32'b11111111111111110000011101100100;
assign LUT_2[43686] = 32'b11111111111111111010011110000111;
assign LUT_2[43687] = 32'b11111111111111110111010110100000;
assign LUT_2[43688] = 32'b11111111111111110001111001000000;
assign LUT_2[43689] = 32'b11111111111111101110110001011001;
assign LUT_2[43690] = 32'b11111111111111111000110001111100;
assign LUT_2[43691] = 32'b11111111111111110101101010010101;
assign LUT_2[43692] = 32'b11111111111111101110010110101000;
assign LUT_2[43693] = 32'b11111111111111101011001111000001;
assign LUT_2[43694] = 32'b11111111111111110101001111100100;
assign LUT_2[43695] = 32'b11111111111111110010000111111101;
assign LUT_2[43696] = 32'b11111111111111110001101011101101;
assign LUT_2[43697] = 32'b11111111111111101110100100000110;
assign LUT_2[43698] = 32'b11111111111111111000100100101001;
assign LUT_2[43699] = 32'b11111111111111110101011101000010;
assign LUT_2[43700] = 32'b11111111111111101110001001010101;
assign LUT_2[43701] = 32'b11111111111111101011000001101110;
assign LUT_2[43702] = 32'b11111111111111110101000010010001;
assign LUT_2[43703] = 32'b11111111111111110001111010101010;
assign LUT_2[43704] = 32'b11111111111111101100011101001010;
assign LUT_2[43705] = 32'b11111111111111101001010101100011;
assign LUT_2[43706] = 32'b11111111111111110011010110000110;
assign LUT_2[43707] = 32'b11111111111111110000001110011111;
assign LUT_2[43708] = 32'b11111111111111101000111010110010;
assign LUT_2[43709] = 32'b11111111111111100101110011001011;
assign LUT_2[43710] = 32'b11111111111111101111110011101110;
assign LUT_2[43711] = 32'b11111111111111101100101100000111;
assign LUT_2[43712] = 32'b11111111111111101110110100011101;
assign LUT_2[43713] = 32'b11111111111111101011101100110110;
assign LUT_2[43714] = 32'b11111111111111110101101101011001;
assign LUT_2[43715] = 32'b11111111111111110010100101110010;
assign LUT_2[43716] = 32'b11111111111111101011010010000101;
assign LUT_2[43717] = 32'b11111111111111101000001010011110;
assign LUT_2[43718] = 32'b11111111111111110010001011000001;
assign LUT_2[43719] = 32'b11111111111111101111000011011010;
assign LUT_2[43720] = 32'b11111111111111101001100101111010;
assign LUT_2[43721] = 32'b11111111111111100110011110010011;
assign LUT_2[43722] = 32'b11111111111111110000011110110110;
assign LUT_2[43723] = 32'b11111111111111101101010111001111;
assign LUT_2[43724] = 32'b11111111111111100110000011100010;
assign LUT_2[43725] = 32'b11111111111111100010111011111011;
assign LUT_2[43726] = 32'b11111111111111101100111100011110;
assign LUT_2[43727] = 32'b11111111111111101001110100110111;
assign LUT_2[43728] = 32'b11111111111111101001011000100111;
assign LUT_2[43729] = 32'b11111111111111100110010001000000;
assign LUT_2[43730] = 32'b11111111111111110000010001100011;
assign LUT_2[43731] = 32'b11111111111111101101001001111100;
assign LUT_2[43732] = 32'b11111111111111100101110110001111;
assign LUT_2[43733] = 32'b11111111111111100010101110101000;
assign LUT_2[43734] = 32'b11111111111111101100101111001011;
assign LUT_2[43735] = 32'b11111111111111101001100111100100;
assign LUT_2[43736] = 32'b11111111111111100100001010000100;
assign LUT_2[43737] = 32'b11111111111111100001000010011101;
assign LUT_2[43738] = 32'b11111111111111101011000011000000;
assign LUT_2[43739] = 32'b11111111111111100111111011011001;
assign LUT_2[43740] = 32'b11111111111111100000100111101100;
assign LUT_2[43741] = 32'b11111111111111011101100000000101;
assign LUT_2[43742] = 32'b11111111111111100111100000101000;
assign LUT_2[43743] = 32'b11111111111111100100011001000001;
assign LUT_2[43744] = 32'b11111111111111101111010000000110;
assign LUT_2[43745] = 32'b11111111111111101100001000011111;
assign LUT_2[43746] = 32'b11111111111111110110001001000010;
assign LUT_2[43747] = 32'b11111111111111110011000001011011;
assign LUT_2[43748] = 32'b11111111111111101011101101101110;
assign LUT_2[43749] = 32'b11111111111111101000100110000111;
assign LUT_2[43750] = 32'b11111111111111110010100110101010;
assign LUT_2[43751] = 32'b11111111111111101111011111000011;
assign LUT_2[43752] = 32'b11111111111111101010000001100011;
assign LUT_2[43753] = 32'b11111111111111100110111001111100;
assign LUT_2[43754] = 32'b11111111111111110000111010011111;
assign LUT_2[43755] = 32'b11111111111111101101110010111000;
assign LUT_2[43756] = 32'b11111111111111100110011111001011;
assign LUT_2[43757] = 32'b11111111111111100011010111100100;
assign LUT_2[43758] = 32'b11111111111111101101011000000111;
assign LUT_2[43759] = 32'b11111111111111101010010000100000;
assign LUT_2[43760] = 32'b11111111111111101001110100010000;
assign LUT_2[43761] = 32'b11111111111111100110101100101001;
assign LUT_2[43762] = 32'b11111111111111110000101101001100;
assign LUT_2[43763] = 32'b11111111111111101101100101100101;
assign LUT_2[43764] = 32'b11111111111111100110010001111000;
assign LUT_2[43765] = 32'b11111111111111100011001010010001;
assign LUT_2[43766] = 32'b11111111111111101101001010110100;
assign LUT_2[43767] = 32'b11111111111111101010000011001101;
assign LUT_2[43768] = 32'b11111111111111100100100101101101;
assign LUT_2[43769] = 32'b11111111111111100001011110000110;
assign LUT_2[43770] = 32'b11111111111111101011011110101001;
assign LUT_2[43771] = 32'b11111111111111101000010111000010;
assign LUT_2[43772] = 32'b11111111111111100001000011010101;
assign LUT_2[43773] = 32'b11111111111111011101111011101110;
assign LUT_2[43774] = 32'b11111111111111100111111100010001;
assign LUT_2[43775] = 32'b11111111111111100100110100101010;
assign LUT_2[43776] = 32'b11111111111111110110010110010001;
assign LUT_2[43777] = 32'b11111111111111110011001110101010;
assign LUT_2[43778] = 32'b11111111111111111101001111001101;
assign LUT_2[43779] = 32'b11111111111111111010000111100110;
assign LUT_2[43780] = 32'b11111111111111110010110011111001;
assign LUT_2[43781] = 32'b11111111111111101111101100010010;
assign LUT_2[43782] = 32'b11111111111111111001101100110101;
assign LUT_2[43783] = 32'b11111111111111110110100101001110;
assign LUT_2[43784] = 32'b11111111111111110001000111101110;
assign LUT_2[43785] = 32'b11111111111111101110000000000111;
assign LUT_2[43786] = 32'b11111111111111111000000000101010;
assign LUT_2[43787] = 32'b11111111111111110100111001000011;
assign LUT_2[43788] = 32'b11111111111111101101100101010110;
assign LUT_2[43789] = 32'b11111111111111101010011101101111;
assign LUT_2[43790] = 32'b11111111111111110100011110010010;
assign LUT_2[43791] = 32'b11111111111111110001010110101011;
assign LUT_2[43792] = 32'b11111111111111110000111010011011;
assign LUT_2[43793] = 32'b11111111111111101101110010110100;
assign LUT_2[43794] = 32'b11111111111111110111110011010111;
assign LUT_2[43795] = 32'b11111111111111110100101011110000;
assign LUT_2[43796] = 32'b11111111111111101101011000000011;
assign LUT_2[43797] = 32'b11111111111111101010010000011100;
assign LUT_2[43798] = 32'b11111111111111110100010000111111;
assign LUT_2[43799] = 32'b11111111111111110001001001011000;
assign LUT_2[43800] = 32'b11111111111111101011101011111000;
assign LUT_2[43801] = 32'b11111111111111101000100100010001;
assign LUT_2[43802] = 32'b11111111111111110010100100110100;
assign LUT_2[43803] = 32'b11111111111111101111011101001101;
assign LUT_2[43804] = 32'b11111111111111101000001001100000;
assign LUT_2[43805] = 32'b11111111111111100101000001111001;
assign LUT_2[43806] = 32'b11111111111111101111000010011100;
assign LUT_2[43807] = 32'b11111111111111101011111010110101;
assign LUT_2[43808] = 32'b11111111111111110110110001111010;
assign LUT_2[43809] = 32'b11111111111111110011101010010011;
assign LUT_2[43810] = 32'b11111111111111111101101010110110;
assign LUT_2[43811] = 32'b11111111111111111010100011001111;
assign LUT_2[43812] = 32'b11111111111111110011001111100010;
assign LUT_2[43813] = 32'b11111111111111110000000111111011;
assign LUT_2[43814] = 32'b11111111111111111010001000011110;
assign LUT_2[43815] = 32'b11111111111111110111000000110111;
assign LUT_2[43816] = 32'b11111111111111110001100011010111;
assign LUT_2[43817] = 32'b11111111111111101110011011110000;
assign LUT_2[43818] = 32'b11111111111111111000011100010011;
assign LUT_2[43819] = 32'b11111111111111110101010100101100;
assign LUT_2[43820] = 32'b11111111111111101110000000111111;
assign LUT_2[43821] = 32'b11111111111111101010111001011000;
assign LUT_2[43822] = 32'b11111111111111110100111001111011;
assign LUT_2[43823] = 32'b11111111111111110001110010010100;
assign LUT_2[43824] = 32'b11111111111111110001010110000100;
assign LUT_2[43825] = 32'b11111111111111101110001110011101;
assign LUT_2[43826] = 32'b11111111111111111000001111000000;
assign LUT_2[43827] = 32'b11111111111111110101000111011001;
assign LUT_2[43828] = 32'b11111111111111101101110011101100;
assign LUT_2[43829] = 32'b11111111111111101010101100000101;
assign LUT_2[43830] = 32'b11111111111111110100101100101000;
assign LUT_2[43831] = 32'b11111111111111110001100101000001;
assign LUT_2[43832] = 32'b11111111111111101100000111100001;
assign LUT_2[43833] = 32'b11111111111111101000111111111010;
assign LUT_2[43834] = 32'b11111111111111110011000000011101;
assign LUT_2[43835] = 32'b11111111111111101111111000110110;
assign LUT_2[43836] = 32'b11111111111111101000100101001001;
assign LUT_2[43837] = 32'b11111111111111100101011101100010;
assign LUT_2[43838] = 32'b11111111111111101111011110000101;
assign LUT_2[43839] = 32'b11111111111111101100010110011110;
assign LUT_2[43840] = 32'b11111111111111101110011110110100;
assign LUT_2[43841] = 32'b11111111111111101011010111001101;
assign LUT_2[43842] = 32'b11111111111111110101010111110000;
assign LUT_2[43843] = 32'b11111111111111110010010000001001;
assign LUT_2[43844] = 32'b11111111111111101010111100011100;
assign LUT_2[43845] = 32'b11111111111111100111110100110101;
assign LUT_2[43846] = 32'b11111111111111110001110101011000;
assign LUT_2[43847] = 32'b11111111111111101110101101110001;
assign LUT_2[43848] = 32'b11111111111111101001010000010001;
assign LUT_2[43849] = 32'b11111111111111100110001000101010;
assign LUT_2[43850] = 32'b11111111111111110000001001001101;
assign LUT_2[43851] = 32'b11111111111111101101000001100110;
assign LUT_2[43852] = 32'b11111111111111100101101101111001;
assign LUT_2[43853] = 32'b11111111111111100010100110010010;
assign LUT_2[43854] = 32'b11111111111111101100100110110101;
assign LUT_2[43855] = 32'b11111111111111101001011111001110;
assign LUT_2[43856] = 32'b11111111111111101001000010111110;
assign LUT_2[43857] = 32'b11111111111111100101111011010111;
assign LUT_2[43858] = 32'b11111111111111101111111011111010;
assign LUT_2[43859] = 32'b11111111111111101100110100010011;
assign LUT_2[43860] = 32'b11111111111111100101100000100110;
assign LUT_2[43861] = 32'b11111111111111100010011000111111;
assign LUT_2[43862] = 32'b11111111111111101100011001100010;
assign LUT_2[43863] = 32'b11111111111111101001010001111011;
assign LUT_2[43864] = 32'b11111111111111100011110100011011;
assign LUT_2[43865] = 32'b11111111111111100000101100110100;
assign LUT_2[43866] = 32'b11111111111111101010101101010111;
assign LUT_2[43867] = 32'b11111111111111100111100101110000;
assign LUT_2[43868] = 32'b11111111111111100000010010000011;
assign LUT_2[43869] = 32'b11111111111111011101001010011100;
assign LUT_2[43870] = 32'b11111111111111100111001010111111;
assign LUT_2[43871] = 32'b11111111111111100100000011011000;
assign LUT_2[43872] = 32'b11111111111111101110111010011101;
assign LUT_2[43873] = 32'b11111111111111101011110010110110;
assign LUT_2[43874] = 32'b11111111111111110101110011011001;
assign LUT_2[43875] = 32'b11111111111111110010101011110010;
assign LUT_2[43876] = 32'b11111111111111101011011000000101;
assign LUT_2[43877] = 32'b11111111111111101000010000011110;
assign LUT_2[43878] = 32'b11111111111111110010010001000001;
assign LUT_2[43879] = 32'b11111111111111101111001001011010;
assign LUT_2[43880] = 32'b11111111111111101001101011111010;
assign LUT_2[43881] = 32'b11111111111111100110100100010011;
assign LUT_2[43882] = 32'b11111111111111110000100100110110;
assign LUT_2[43883] = 32'b11111111111111101101011101001111;
assign LUT_2[43884] = 32'b11111111111111100110001001100010;
assign LUT_2[43885] = 32'b11111111111111100011000001111011;
assign LUT_2[43886] = 32'b11111111111111101101000010011110;
assign LUT_2[43887] = 32'b11111111111111101001111010110111;
assign LUT_2[43888] = 32'b11111111111111101001011110100111;
assign LUT_2[43889] = 32'b11111111111111100110010111000000;
assign LUT_2[43890] = 32'b11111111111111110000010111100011;
assign LUT_2[43891] = 32'b11111111111111101101001111111100;
assign LUT_2[43892] = 32'b11111111111111100101111100001111;
assign LUT_2[43893] = 32'b11111111111111100010110100101000;
assign LUT_2[43894] = 32'b11111111111111101100110101001011;
assign LUT_2[43895] = 32'b11111111111111101001101101100100;
assign LUT_2[43896] = 32'b11111111111111100100010000000100;
assign LUT_2[43897] = 32'b11111111111111100001001000011101;
assign LUT_2[43898] = 32'b11111111111111101011001001000000;
assign LUT_2[43899] = 32'b11111111111111101000000001011001;
assign LUT_2[43900] = 32'b11111111111111100000101101101100;
assign LUT_2[43901] = 32'b11111111111111011101100110000101;
assign LUT_2[43902] = 32'b11111111111111100111100110101000;
assign LUT_2[43903] = 32'b11111111111111100100011111000001;
assign LUT_2[43904] = 32'b11111111111111111010101010100000;
assign LUT_2[43905] = 32'b11111111111111110111100010111001;
assign LUT_2[43906] = 32'b00000000000000000001100011011100;
assign LUT_2[43907] = 32'b11111111111111111110011011110101;
assign LUT_2[43908] = 32'b11111111111111110111001000001000;
assign LUT_2[43909] = 32'b11111111111111110100000000100001;
assign LUT_2[43910] = 32'b11111111111111111110000001000100;
assign LUT_2[43911] = 32'b11111111111111111010111001011101;
assign LUT_2[43912] = 32'b11111111111111110101011011111101;
assign LUT_2[43913] = 32'b11111111111111110010010100010110;
assign LUT_2[43914] = 32'b11111111111111111100010100111001;
assign LUT_2[43915] = 32'b11111111111111111001001101010010;
assign LUT_2[43916] = 32'b11111111111111110001111001100101;
assign LUT_2[43917] = 32'b11111111111111101110110001111110;
assign LUT_2[43918] = 32'b11111111111111111000110010100001;
assign LUT_2[43919] = 32'b11111111111111110101101010111010;
assign LUT_2[43920] = 32'b11111111111111110101001110101010;
assign LUT_2[43921] = 32'b11111111111111110010000111000011;
assign LUT_2[43922] = 32'b11111111111111111100000111100110;
assign LUT_2[43923] = 32'b11111111111111111000111111111111;
assign LUT_2[43924] = 32'b11111111111111110001101100010010;
assign LUT_2[43925] = 32'b11111111111111101110100100101011;
assign LUT_2[43926] = 32'b11111111111111111000100101001110;
assign LUT_2[43927] = 32'b11111111111111110101011101100111;
assign LUT_2[43928] = 32'b11111111111111110000000000000111;
assign LUT_2[43929] = 32'b11111111111111101100111000100000;
assign LUT_2[43930] = 32'b11111111111111110110111001000011;
assign LUT_2[43931] = 32'b11111111111111110011110001011100;
assign LUT_2[43932] = 32'b11111111111111101100011101101111;
assign LUT_2[43933] = 32'b11111111111111101001010110001000;
assign LUT_2[43934] = 32'b11111111111111110011010110101011;
assign LUT_2[43935] = 32'b11111111111111110000001111000100;
assign LUT_2[43936] = 32'b11111111111111111011000110001001;
assign LUT_2[43937] = 32'b11111111111111110111111110100010;
assign LUT_2[43938] = 32'b00000000000000000001111111000101;
assign LUT_2[43939] = 32'b11111111111111111110110111011110;
assign LUT_2[43940] = 32'b11111111111111110111100011110001;
assign LUT_2[43941] = 32'b11111111111111110100011100001010;
assign LUT_2[43942] = 32'b11111111111111111110011100101101;
assign LUT_2[43943] = 32'b11111111111111111011010101000110;
assign LUT_2[43944] = 32'b11111111111111110101110111100110;
assign LUT_2[43945] = 32'b11111111111111110010101111111111;
assign LUT_2[43946] = 32'b11111111111111111100110000100010;
assign LUT_2[43947] = 32'b11111111111111111001101000111011;
assign LUT_2[43948] = 32'b11111111111111110010010101001110;
assign LUT_2[43949] = 32'b11111111111111101111001101100111;
assign LUT_2[43950] = 32'b11111111111111111001001110001010;
assign LUT_2[43951] = 32'b11111111111111110110000110100011;
assign LUT_2[43952] = 32'b11111111111111110101101010010011;
assign LUT_2[43953] = 32'b11111111111111110010100010101100;
assign LUT_2[43954] = 32'b11111111111111111100100011001111;
assign LUT_2[43955] = 32'b11111111111111111001011011101000;
assign LUT_2[43956] = 32'b11111111111111110010000111111011;
assign LUT_2[43957] = 32'b11111111111111101111000000010100;
assign LUT_2[43958] = 32'b11111111111111111001000000110111;
assign LUT_2[43959] = 32'b11111111111111110101111001010000;
assign LUT_2[43960] = 32'b11111111111111110000011011110000;
assign LUT_2[43961] = 32'b11111111111111101101010100001001;
assign LUT_2[43962] = 32'b11111111111111110111010100101100;
assign LUT_2[43963] = 32'b11111111111111110100001101000101;
assign LUT_2[43964] = 32'b11111111111111101100111001011000;
assign LUT_2[43965] = 32'b11111111111111101001110001110001;
assign LUT_2[43966] = 32'b11111111111111110011110010010100;
assign LUT_2[43967] = 32'b11111111111111110000101010101101;
assign LUT_2[43968] = 32'b11111111111111110010110011000011;
assign LUT_2[43969] = 32'b11111111111111101111101011011100;
assign LUT_2[43970] = 32'b11111111111111111001101011111111;
assign LUT_2[43971] = 32'b11111111111111110110100100011000;
assign LUT_2[43972] = 32'b11111111111111101111010000101011;
assign LUT_2[43973] = 32'b11111111111111101100001001000100;
assign LUT_2[43974] = 32'b11111111111111110110001001100111;
assign LUT_2[43975] = 32'b11111111111111110011000010000000;
assign LUT_2[43976] = 32'b11111111111111101101100100100000;
assign LUT_2[43977] = 32'b11111111111111101010011100111001;
assign LUT_2[43978] = 32'b11111111111111110100011101011100;
assign LUT_2[43979] = 32'b11111111111111110001010101110101;
assign LUT_2[43980] = 32'b11111111111111101010000010001000;
assign LUT_2[43981] = 32'b11111111111111100110111010100001;
assign LUT_2[43982] = 32'b11111111111111110000111011000100;
assign LUT_2[43983] = 32'b11111111111111101101110011011101;
assign LUT_2[43984] = 32'b11111111111111101101010111001101;
assign LUT_2[43985] = 32'b11111111111111101010001111100110;
assign LUT_2[43986] = 32'b11111111111111110100010000001001;
assign LUT_2[43987] = 32'b11111111111111110001001000100010;
assign LUT_2[43988] = 32'b11111111111111101001110100110101;
assign LUT_2[43989] = 32'b11111111111111100110101101001110;
assign LUT_2[43990] = 32'b11111111111111110000101101110001;
assign LUT_2[43991] = 32'b11111111111111101101100110001010;
assign LUT_2[43992] = 32'b11111111111111101000001000101010;
assign LUT_2[43993] = 32'b11111111111111100101000001000011;
assign LUT_2[43994] = 32'b11111111111111101111000001100110;
assign LUT_2[43995] = 32'b11111111111111101011111001111111;
assign LUT_2[43996] = 32'b11111111111111100100100110010010;
assign LUT_2[43997] = 32'b11111111111111100001011110101011;
assign LUT_2[43998] = 32'b11111111111111101011011111001110;
assign LUT_2[43999] = 32'b11111111111111101000010111100111;
assign LUT_2[44000] = 32'b11111111111111110011001110101100;
assign LUT_2[44001] = 32'b11111111111111110000000111000101;
assign LUT_2[44002] = 32'b11111111111111111010000111101000;
assign LUT_2[44003] = 32'b11111111111111110111000000000001;
assign LUT_2[44004] = 32'b11111111111111101111101100010100;
assign LUT_2[44005] = 32'b11111111111111101100100100101101;
assign LUT_2[44006] = 32'b11111111111111110110100101010000;
assign LUT_2[44007] = 32'b11111111111111110011011101101001;
assign LUT_2[44008] = 32'b11111111111111101110000000001001;
assign LUT_2[44009] = 32'b11111111111111101010111000100010;
assign LUT_2[44010] = 32'b11111111111111110100111001000101;
assign LUT_2[44011] = 32'b11111111111111110001110001011110;
assign LUT_2[44012] = 32'b11111111111111101010011101110001;
assign LUT_2[44013] = 32'b11111111111111100111010110001010;
assign LUT_2[44014] = 32'b11111111111111110001010110101101;
assign LUT_2[44015] = 32'b11111111111111101110001111000110;
assign LUT_2[44016] = 32'b11111111111111101101110010110110;
assign LUT_2[44017] = 32'b11111111111111101010101011001111;
assign LUT_2[44018] = 32'b11111111111111110100101011110010;
assign LUT_2[44019] = 32'b11111111111111110001100100001011;
assign LUT_2[44020] = 32'b11111111111111101010010000011110;
assign LUT_2[44021] = 32'b11111111111111100111001000110111;
assign LUT_2[44022] = 32'b11111111111111110001001001011010;
assign LUT_2[44023] = 32'b11111111111111101110000001110011;
assign LUT_2[44024] = 32'b11111111111111101000100100010011;
assign LUT_2[44025] = 32'b11111111111111100101011100101100;
assign LUT_2[44026] = 32'b11111111111111101111011101001111;
assign LUT_2[44027] = 32'b11111111111111101100010101101000;
assign LUT_2[44028] = 32'b11111111111111100101000001111011;
assign LUT_2[44029] = 32'b11111111111111100001111010010100;
assign LUT_2[44030] = 32'b11111111111111101011111010110111;
assign LUT_2[44031] = 32'b11111111111111101000110011010000;
assign LUT_2[44032] = 32'b11111111111111110100010001111110;
assign LUT_2[44033] = 32'b11111111111111110001001010010111;
assign LUT_2[44034] = 32'b11111111111111111011001010111010;
assign LUT_2[44035] = 32'b11111111111111111000000011010011;
assign LUT_2[44036] = 32'b11111111111111110000101111100110;
assign LUT_2[44037] = 32'b11111111111111101101100111111111;
assign LUT_2[44038] = 32'b11111111111111110111101000100010;
assign LUT_2[44039] = 32'b11111111111111110100100000111011;
assign LUT_2[44040] = 32'b11111111111111101111000011011011;
assign LUT_2[44041] = 32'b11111111111111101011111011110100;
assign LUT_2[44042] = 32'b11111111111111110101111100010111;
assign LUT_2[44043] = 32'b11111111111111110010110100110000;
assign LUT_2[44044] = 32'b11111111111111101011100001000011;
assign LUT_2[44045] = 32'b11111111111111101000011001011100;
assign LUT_2[44046] = 32'b11111111111111110010011001111111;
assign LUT_2[44047] = 32'b11111111111111101111010010011000;
assign LUT_2[44048] = 32'b11111111111111101110110110001000;
assign LUT_2[44049] = 32'b11111111111111101011101110100001;
assign LUT_2[44050] = 32'b11111111111111110101101111000100;
assign LUT_2[44051] = 32'b11111111111111110010100111011101;
assign LUT_2[44052] = 32'b11111111111111101011010011110000;
assign LUT_2[44053] = 32'b11111111111111101000001100001001;
assign LUT_2[44054] = 32'b11111111111111110010001100101100;
assign LUT_2[44055] = 32'b11111111111111101111000101000101;
assign LUT_2[44056] = 32'b11111111111111101001100111100101;
assign LUT_2[44057] = 32'b11111111111111100110011111111110;
assign LUT_2[44058] = 32'b11111111111111110000100000100001;
assign LUT_2[44059] = 32'b11111111111111101101011000111010;
assign LUT_2[44060] = 32'b11111111111111100110000101001101;
assign LUT_2[44061] = 32'b11111111111111100010111101100110;
assign LUT_2[44062] = 32'b11111111111111101100111110001001;
assign LUT_2[44063] = 32'b11111111111111101001110110100010;
assign LUT_2[44064] = 32'b11111111111111110100101101100111;
assign LUT_2[44065] = 32'b11111111111111110001100110000000;
assign LUT_2[44066] = 32'b11111111111111111011100110100011;
assign LUT_2[44067] = 32'b11111111111111111000011110111100;
assign LUT_2[44068] = 32'b11111111111111110001001011001111;
assign LUT_2[44069] = 32'b11111111111111101110000011101000;
assign LUT_2[44070] = 32'b11111111111111111000000100001011;
assign LUT_2[44071] = 32'b11111111111111110100111100100100;
assign LUT_2[44072] = 32'b11111111111111101111011111000100;
assign LUT_2[44073] = 32'b11111111111111101100010111011101;
assign LUT_2[44074] = 32'b11111111111111110110011000000000;
assign LUT_2[44075] = 32'b11111111111111110011010000011001;
assign LUT_2[44076] = 32'b11111111111111101011111100101100;
assign LUT_2[44077] = 32'b11111111111111101000110101000101;
assign LUT_2[44078] = 32'b11111111111111110010110101101000;
assign LUT_2[44079] = 32'b11111111111111101111101110000001;
assign LUT_2[44080] = 32'b11111111111111101111010001110001;
assign LUT_2[44081] = 32'b11111111111111101100001010001010;
assign LUT_2[44082] = 32'b11111111111111110110001010101101;
assign LUT_2[44083] = 32'b11111111111111110011000011000110;
assign LUT_2[44084] = 32'b11111111111111101011101111011001;
assign LUT_2[44085] = 32'b11111111111111101000100111110010;
assign LUT_2[44086] = 32'b11111111111111110010101000010101;
assign LUT_2[44087] = 32'b11111111111111101111100000101110;
assign LUT_2[44088] = 32'b11111111111111101010000011001110;
assign LUT_2[44089] = 32'b11111111111111100110111011100111;
assign LUT_2[44090] = 32'b11111111111111110000111100001010;
assign LUT_2[44091] = 32'b11111111111111101101110100100011;
assign LUT_2[44092] = 32'b11111111111111100110100000110110;
assign LUT_2[44093] = 32'b11111111111111100011011001001111;
assign LUT_2[44094] = 32'b11111111111111101101011001110010;
assign LUT_2[44095] = 32'b11111111111111101010010010001011;
assign LUT_2[44096] = 32'b11111111111111101100011010100001;
assign LUT_2[44097] = 32'b11111111111111101001010010111010;
assign LUT_2[44098] = 32'b11111111111111110011010011011101;
assign LUT_2[44099] = 32'b11111111111111110000001011110110;
assign LUT_2[44100] = 32'b11111111111111101000111000001001;
assign LUT_2[44101] = 32'b11111111111111100101110000100010;
assign LUT_2[44102] = 32'b11111111111111101111110001000101;
assign LUT_2[44103] = 32'b11111111111111101100101001011110;
assign LUT_2[44104] = 32'b11111111111111100111001011111110;
assign LUT_2[44105] = 32'b11111111111111100100000100010111;
assign LUT_2[44106] = 32'b11111111111111101110000100111010;
assign LUT_2[44107] = 32'b11111111111111101010111101010011;
assign LUT_2[44108] = 32'b11111111111111100011101001100110;
assign LUT_2[44109] = 32'b11111111111111100000100001111111;
assign LUT_2[44110] = 32'b11111111111111101010100010100010;
assign LUT_2[44111] = 32'b11111111111111100111011010111011;
assign LUT_2[44112] = 32'b11111111111111100110111110101011;
assign LUT_2[44113] = 32'b11111111111111100011110111000100;
assign LUT_2[44114] = 32'b11111111111111101101110111100111;
assign LUT_2[44115] = 32'b11111111111111101010110000000000;
assign LUT_2[44116] = 32'b11111111111111100011011100010011;
assign LUT_2[44117] = 32'b11111111111111100000010100101100;
assign LUT_2[44118] = 32'b11111111111111101010010101001111;
assign LUT_2[44119] = 32'b11111111111111100111001101101000;
assign LUT_2[44120] = 32'b11111111111111100001110000001000;
assign LUT_2[44121] = 32'b11111111111111011110101000100001;
assign LUT_2[44122] = 32'b11111111111111101000101001000100;
assign LUT_2[44123] = 32'b11111111111111100101100001011101;
assign LUT_2[44124] = 32'b11111111111111011110001101110000;
assign LUT_2[44125] = 32'b11111111111111011011000110001001;
assign LUT_2[44126] = 32'b11111111111111100101000110101100;
assign LUT_2[44127] = 32'b11111111111111100001111111000101;
assign LUT_2[44128] = 32'b11111111111111101100110110001010;
assign LUT_2[44129] = 32'b11111111111111101001101110100011;
assign LUT_2[44130] = 32'b11111111111111110011101111000110;
assign LUT_2[44131] = 32'b11111111111111110000100111011111;
assign LUT_2[44132] = 32'b11111111111111101001010011110010;
assign LUT_2[44133] = 32'b11111111111111100110001100001011;
assign LUT_2[44134] = 32'b11111111111111110000001100101110;
assign LUT_2[44135] = 32'b11111111111111101101000101000111;
assign LUT_2[44136] = 32'b11111111111111100111100111100111;
assign LUT_2[44137] = 32'b11111111111111100100100000000000;
assign LUT_2[44138] = 32'b11111111111111101110100000100011;
assign LUT_2[44139] = 32'b11111111111111101011011000111100;
assign LUT_2[44140] = 32'b11111111111111100100000101001111;
assign LUT_2[44141] = 32'b11111111111111100000111101101000;
assign LUT_2[44142] = 32'b11111111111111101010111110001011;
assign LUT_2[44143] = 32'b11111111111111100111110110100100;
assign LUT_2[44144] = 32'b11111111111111100111011010010100;
assign LUT_2[44145] = 32'b11111111111111100100010010101101;
assign LUT_2[44146] = 32'b11111111111111101110010011010000;
assign LUT_2[44147] = 32'b11111111111111101011001011101001;
assign LUT_2[44148] = 32'b11111111111111100011110111111100;
assign LUT_2[44149] = 32'b11111111111111100000110000010101;
assign LUT_2[44150] = 32'b11111111111111101010110000111000;
assign LUT_2[44151] = 32'b11111111111111100111101001010001;
assign LUT_2[44152] = 32'b11111111111111100010001011110001;
assign LUT_2[44153] = 32'b11111111111111011111000100001010;
assign LUT_2[44154] = 32'b11111111111111101001000100101101;
assign LUT_2[44155] = 32'b11111111111111100101111101000110;
assign LUT_2[44156] = 32'b11111111111111011110101001011001;
assign LUT_2[44157] = 32'b11111111111111011011100001110010;
assign LUT_2[44158] = 32'b11111111111111100101100010010101;
assign LUT_2[44159] = 32'b11111111111111100010011010101110;
assign LUT_2[44160] = 32'b11111111111111111000100110001101;
assign LUT_2[44161] = 32'b11111111111111110101011110100110;
assign LUT_2[44162] = 32'b11111111111111111111011111001001;
assign LUT_2[44163] = 32'b11111111111111111100010111100010;
assign LUT_2[44164] = 32'b11111111111111110101000011110101;
assign LUT_2[44165] = 32'b11111111111111110001111100001110;
assign LUT_2[44166] = 32'b11111111111111111011111100110001;
assign LUT_2[44167] = 32'b11111111111111111000110101001010;
assign LUT_2[44168] = 32'b11111111111111110011010111101010;
assign LUT_2[44169] = 32'b11111111111111110000010000000011;
assign LUT_2[44170] = 32'b11111111111111111010010000100110;
assign LUT_2[44171] = 32'b11111111111111110111001000111111;
assign LUT_2[44172] = 32'b11111111111111101111110101010010;
assign LUT_2[44173] = 32'b11111111111111101100101101101011;
assign LUT_2[44174] = 32'b11111111111111110110101110001110;
assign LUT_2[44175] = 32'b11111111111111110011100110100111;
assign LUT_2[44176] = 32'b11111111111111110011001010010111;
assign LUT_2[44177] = 32'b11111111111111110000000010110000;
assign LUT_2[44178] = 32'b11111111111111111010000011010011;
assign LUT_2[44179] = 32'b11111111111111110110111011101100;
assign LUT_2[44180] = 32'b11111111111111101111100111111111;
assign LUT_2[44181] = 32'b11111111111111101100100000011000;
assign LUT_2[44182] = 32'b11111111111111110110100000111011;
assign LUT_2[44183] = 32'b11111111111111110011011001010100;
assign LUT_2[44184] = 32'b11111111111111101101111011110100;
assign LUT_2[44185] = 32'b11111111111111101010110100001101;
assign LUT_2[44186] = 32'b11111111111111110100110100110000;
assign LUT_2[44187] = 32'b11111111111111110001101101001001;
assign LUT_2[44188] = 32'b11111111111111101010011001011100;
assign LUT_2[44189] = 32'b11111111111111100111010001110101;
assign LUT_2[44190] = 32'b11111111111111110001010010011000;
assign LUT_2[44191] = 32'b11111111111111101110001010110001;
assign LUT_2[44192] = 32'b11111111111111111001000001110110;
assign LUT_2[44193] = 32'b11111111111111110101111010001111;
assign LUT_2[44194] = 32'b11111111111111111111111010110010;
assign LUT_2[44195] = 32'b11111111111111111100110011001011;
assign LUT_2[44196] = 32'b11111111111111110101011111011110;
assign LUT_2[44197] = 32'b11111111111111110010010111110111;
assign LUT_2[44198] = 32'b11111111111111111100011000011010;
assign LUT_2[44199] = 32'b11111111111111111001010000110011;
assign LUT_2[44200] = 32'b11111111111111110011110011010011;
assign LUT_2[44201] = 32'b11111111111111110000101011101100;
assign LUT_2[44202] = 32'b11111111111111111010101100001111;
assign LUT_2[44203] = 32'b11111111111111110111100100101000;
assign LUT_2[44204] = 32'b11111111111111110000010000111011;
assign LUT_2[44205] = 32'b11111111111111101101001001010100;
assign LUT_2[44206] = 32'b11111111111111110111001001110111;
assign LUT_2[44207] = 32'b11111111111111110100000010010000;
assign LUT_2[44208] = 32'b11111111111111110011100110000000;
assign LUT_2[44209] = 32'b11111111111111110000011110011001;
assign LUT_2[44210] = 32'b11111111111111111010011110111100;
assign LUT_2[44211] = 32'b11111111111111110111010111010101;
assign LUT_2[44212] = 32'b11111111111111110000000011101000;
assign LUT_2[44213] = 32'b11111111111111101100111100000001;
assign LUT_2[44214] = 32'b11111111111111110110111100100100;
assign LUT_2[44215] = 32'b11111111111111110011110100111101;
assign LUT_2[44216] = 32'b11111111111111101110010111011101;
assign LUT_2[44217] = 32'b11111111111111101011001111110110;
assign LUT_2[44218] = 32'b11111111111111110101010000011001;
assign LUT_2[44219] = 32'b11111111111111110010001000110010;
assign LUT_2[44220] = 32'b11111111111111101010110101000101;
assign LUT_2[44221] = 32'b11111111111111100111101101011110;
assign LUT_2[44222] = 32'b11111111111111110001101110000001;
assign LUT_2[44223] = 32'b11111111111111101110100110011010;
assign LUT_2[44224] = 32'b11111111111111110000101110110000;
assign LUT_2[44225] = 32'b11111111111111101101100111001001;
assign LUT_2[44226] = 32'b11111111111111110111100111101100;
assign LUT_2[44227] = 32'b11111111111111110100100000000101;
assign LUT_2[44228] = 32'b11111111111111101101001100011000;
assign LUT_2[44229] = 32'b11111111111111101010000100110001;
assign LUT_2[44230] = 32'b11111111111111110100000101010100;
assign LUT_2[44231] = 32'b11111111111111110000111101101101;
assign LUT_2[44232] = 32'b11111111111111101011100000001101;
assign LUT_2[44233] = 32'b11111111111111101000011000100110;
assign LUT_2[44234] = 32'b11111111111111110010011001001001;
assign LUT_2[44235] = 32'b11111111111111101111010001100010;
assign LUT_2[44236] = 32'b11111111111111100111111101110101;
assign LUT_2[44237] = 32'b11111111111111100100110110001110;
assign LUT_2[44238] = 32'b11111111111111101110110110110001;
assign LUT_2[44239] = 32'b11111111111111101011101111001010;
assign LUT_2[44240] = 32'b11111111111111101011010010111010;
assign LUT_2[44241] = 32'b11111111111111101000001011010011;
assign LUT_2[44242] = 32'b11111111111111110010001011110110;
assign LUT_2[44243] = 32'b11111111111111101111000100001111;
assign LUT_2[44244] = 32'b11111111111111100111110000100010;
assign LUT_2[44245] = 32'b11111111111111100100101000111011;
assign LUT_2[44246] = 32'b11111111111111101110101001011110;
assign LUT_2[44247] = 32'b11111111111111101011100001110111;
assign LUT_2[44248] = 32'b11111111111111100110000100010111;
assign LUT_2[44249] = 32'b11111111111111100010111100110000;
assign LUT_2[44250] = 32'b11111111111111101100111101010011;
assign LUT_2[44251] = 32'b11111111111111101001110101101100;
assign LUT_2[44252] = 32'b11111111111111100010100001111111;
assign LUT_2[44253] = 32'b11111111111111011111011010011000;
assign LUT_2[44254] = 32'b11111111111111101001011010111011;
assign LUT_2[44255] = 32'b11111111111111100110010011010100;
assign LUT_2[44256] = 32'b11111111111111110001001010011001;
assign LUT_2[44257] = 32'b11111111111111101110000010110010;
assign LUT_2[44258] = 32'b11111111111111111000000011010101;
assign LUT_2[44259] = 32'b11111111111111110100111011101110;
assign LUT_2[44260] = 32'b11111111111111101101101000000001;
assign LUT_2[44261] = 32'b11111111111111101010100000011010;
assign LUT_2[44262] = 32'b11111111111111110100100000111101;
assign LUT_2[44263] = 32'b11111111111111110001011001010110;
assign LUT_2[44264] = 32'b11111111111111101011111011110110;
assign LUT_2[44265] = 32'b11111111111111101000110100001111;
assign LUT_2[44266] = 32'b11111111111111110010110100110010;
assign LUT_2[44267] = 32'b11111111111111101111101101001011;
assign LUT_2[44268] = 32'b11111111111111101000011001011110;
assign LUT_2[44269] = 32'b11111111111111100101010001110111;
assign LUT_2[44270] = 32'b11111111111111101111010010011010;
assign LUT_2[44271] = 32'b11111111111111101100001010110011;
assign LUT_2[44272] = 32'b11111111111111101011101110100011;
assign LUT_2[44273] = 32'b11111111111111101000100110111100;
assign LUT_2[44274] = 32'b11111111111111110010100111011111;
assign LUT_2[44275] = 32'b11111111111111101111011111111000;
assign LUT_2[44276] = 32'b11111111111111101000001100001011;
assign LUT_2[44277] = 32'b11111111111111100101000100100100;
assign LUT_2[44278] = 32'b11111111111111101111000101000111;
assign LUT_2[44279] = 32'b11111111111111101011111101100000;
assign LUT_2[44280] = 32'b11111111111111100110100000000000;
assign LUT_2[44281] = 32'b11111111111111100011011000011001;
assign LUT_2[44282] = 32'b11111111111111101101011000111100;
assign LUT_2[44283] = 32'b11111111111111101010010001010101;
assign LUT_2[44284] = 32'b11111111111111100010111101101000;
assign LUT_2[44285] = 32'b11111111111111011111110110000001;
assign LUT_2[44286] = 32'b11111111111111101001110110100100;
assign LUT_2[44287] = 32'b11111111111111100110101110111101;
assign LUT_2[44288] = 32'b11111111111111111000010000100100;
assign LUT_2[44289] = 32'b11111111111111110101001000111101;
assign LUT_2[44290] = 32'b11111111111111111111001001100000;
assign LUT_2[44291] = 32'b11111111111111111100000001111001;
assign LUT_2[44292] = 32'b11111111111111110100101110001100;
assign LUT_2[44293] = 32'b11111111111111110001100110100101;
assign LUT_2[44294] = 32'b11111111111111111011100111001000;
assign LUT_2[44295] = 32'b11111111111111111000011111100001;
assign LUT_2[44296] = 32'b11111111111111110011000010000001;
assign LUT_2[44297] = 32'b11111111111111101111111010011010;
assign LUT_2[44298] = 32'b11111111111111111001111010111101;
assign LUT_2[44299] = 32'b11111111111111110110110011010110;
assign LUT_2[44300] = 32'b11111111111111101111011111101001;
assign LUT_2[44301] = 32'b11111111111111101100011000000010;
assign LUT_2[44302] = 32'b11111111111111110110011000100101;
assign LUT_2[44303] = 32'b11111111111111110011010000111110;
assign LUT_2[44304] = 32'b11111111111111110010110100101110;
assign LUT_2[44305] = 32'b11111111111111101111101101000111;
assign LUT_2[44306] = 32'b11111111111111111001101101101010;
assign LUT_2[44307] = 32'b11111111111111110110100110000011;
assign LUT_2[44308] = 32'b11111111111111101111010010010110;
assign LUT_2[44309] = 32'b11111111111111101100001010101111;
assign LUT_2[44310] = 32'b11111111111111110110001011010010;
assign LUT_2[44311] = 32'b11111111111111110011000011101011;
assign LUT_2[44312] = 32'b11111111111111101101100110001011;
assign LUT_2[44313] = 32'b11111111111111101010011110100100;
assign LUT_2[44314] = 32'b11111111111111110100011111000111;
assign LUT_2[44315] = 32'b11111111111111110001010111100000;
assign LUT_2[44316] = 32'b11111111111111101010000011110011;
assign LUT_2[44317] = 32'b11111111111111100110111100001100;
assign LUT_2[44318] = 32'b11111111111111110000111100101111;
assign LUT_2[44319] = 32'b11111111111111101101110101001000;
assign LUT_2[44320] = 32'b11111111111111111000101100001101;
assign LUT_2[44321] = 32'b11111111111111110101100100100110;
assign LUT_2[44322] = 32'b11111111111111111111100101001001;
assign LUT_2[44323] = 32'b11111111111111111100011101100010;
assign LUT_2[44324] = 32'b11111111111111110101001001110101;
assign LUT_2[44325] = 32'b11111111111111110010000010001110;
assign LUT_2[44326] = 32'b11111111111111111100000010110001;
assign LUT_2[44327] = 32'b11111111111111111000111011001010;
assign LUT_2[44328] = 32'b11111111111111110011011101101010;
assign LUT_2[44329] = 32'b11111111111111110000010110000011;
assign LUT_2[44330] = 32'b11111111111111111010010110100110;
assign LUT_2[44331] = 32'b11111111111111110111001110111111;
assign LUT_2[44332] = 32'b11111111111111101111111011010010;
assign LUT_2[44333] = 32'b11111111111111101100110011101011;
assign LUT_2[44334] = 32'b11111111111111110110110100001110;
assign LUT_2[44335] = 32'b11111111111111110011101100100111;
assign LUT_2[44336] = 32'b11111111111111110011010000010111;
assign LUT_2[44337] = 32'b11111111111111110000001000110000;
assign LUT_2[44338] = 32'b11111111111111111010001001010011;
assign LUT_2[44339] = 32'b11111111111111110111000001101100;
assign LUT_2[44340] = 32'b11111111111111101111101101111111;
assign LUT_2[44341] = 32'b11111111111111101100100110011000;
assign LUT_2[44342] = 32'b11111111111111110110100110111011;
assign LUT_2[44343] = 32'b11111111111111110011011111010100;
assign LUT_2[44344] = 32'b11111111111111101110000001110100;
assign LUT_2[44345] = 32'b11111111111111101010111010001101;
assign LUT_2[44346] = 32'b11111111111111110100111010110000;
assign LUT_2[44347] = 32'b11111111111111110001110011001001;
assign LUT_2[44348] = 32'b11111111111111101010011111011100;
assign LUT_2[44349] = 32'b11111111111111100111010111110101;
assign LUT_2[44350] = 32'b11111111111111110001011000011000;
assign LUT_2[44351] = 32'b11111111111111101110010000110001;
assign LUT_2[44352] = 32'b11111111111111110000011001000111;
assign LUT_2[44353] = 32'b11111111111111101101010001100000;
assign LUT_2[44354] = 32'b11111111111111110111010010000011;
assign LUT_2[44355] = 32'b11111111111111110100001010011100;
assign LUT_2[44356] = 32'b11111111111111101100110110101111;
assign LUT_2[44357] = 32'b11111111111111101001101111001000;
assign LUT_2[44358] = 32'b11111111111111110011101111101011;
assign LUT_2[44359] = 32'b11111111111111110000101000000100;
assign LUT_2[44360] = 32'b11111111111111101011001010100100;
assign LUT_2[44361] = 32'b11111111111111101000000010111101;
assign LUT_2[44362] = 32'b11111111111111110010000011100000;
assign LUT_2[44363] = 32'b11111111111111101110111011111001;
assign LUT_2[44364] = 32'b11111111111111100111101000001100;
assign LUT_2[44365] = 32'b11111111111111100100100000100101;
assign LUT_2[44366] = 32'b11111111111111101110100001001000;
assign LUT_2[44367] = 32'b11111111111111101011011001100001;
assign LUT_2[44368] = 32'b11111111111111101010111101010001;
assign LUT_2[44369] = 32'b11111111111111100111110101101010;
assign LUT_2[44370] = 32'b11111111111111110001110110001101;
assign LUT_2[44371] = 32'b11111111111111101110101110100110;
assign LUT_2[44372] = 32'b11111111111111100111011010111001;
assign LUT_2[44373] = 32'b11111111111111100100010011010010;
assign LUT_2[44374] = 32'b11111111111111101110010011110101;
assign LUT_2[44375] = 32'b11111111111111101011001100001110;
assign LUT_2[44376] = 32'b11111111111111100101101110101110;
assign LUT_2[44377] = 32'b11111111111111100010100111000111;
assign LUT_2[44378] = 32'b11111111111111101100100111101010;
assign LUT_2[44379] = 32'b11111111111111101001100000000011;
assign LUT_2[44380] = 32'b11111111111111100010001100010110;
assign LUT_2[44381] = 32'b11111111111111011111000100101111;
assign LUT_2[44382] = 32'b11111111111111101001000101010010;
assign LUT_2[44383] = 32'b11111111111111100101111101101011;
assign LUT_2[44384] = 32'b11111111111111110000110100110000;
assign LUT_2[44385] = 32'b11111111111111101101101101001001;
assign LUT_2[44386] = 32'b11111111111111110111101101101100;
assign LUT_2[44387] = 32'b11111111111111110100100110000101;
assign LUT_2[44388] = 32'b11111111111111101101010010011000;
assign LUT_2[44389] = 32'b11111111111111101010001010110001;
assign LUT_2[44390] = 32'b11111111111111110100001011010100;
assign LUT_2[44391] = 32'b11111111111111110001000011101101;
assign LUT_2[44392] = 32'b11111111111111101011100110001101;
assign LUT_2[44393] = 32'b11111111111111101000011110100110;
assign LUT_2[44394] = 32'b11111111111111110010011111001001;
assign LUT_2[44395] = 32'b11111111111111101111010111100010;
assign LUT_2[44396] = 32'b11111111111111101000000011110101;
assign LUT_2[44397] = 32'b11111111111111100100111100001110;
assign LUT_2[44398] = 32'b11111111111111101110111100110001;
assign LUT_2[44399] = 32'b11111111111111101011110101001010;
assign LUT_2[44400] = 32'b11111111111111101011011000111010;
assign LUT_2[44401] = 32'b11111111111111101000010001010011;
assign LUT_2[44402] = 32'b11111111111111110010010001110110;
assign LUT_2[44403] = 32'b11111111111111101111001010001111;
assign LUT_2[44404] = 32'b11111111111111100111110110100010;
assign LUT_2[44405] = 32'b11111111111111100100101110111011;
assign LUT_2[44406] = 32'b11111111111111101110101111011110;
assign LUT_2[44407] = 32'b11111111111111101011100111110111;
assign LUT_2[44408] = 32'b11111111111111100110001010010111;
assign LUT_2[44409] = 32'b11111111111111100011000010110000;
assign LUT_2[44410] = 32'b11111111111111101101000011010011;
assign LUT_2[44411] = 32'b11111111111111101001111011101100;
assign LUT_2[44412] = 32'b11111111111111100010100111111111;
assign LUT_2[44413] = 32'b11111111111111011111100000011000;
assign LUT_2[44414] = 32'b11111111111111101001100000111011;
assign LUT_2[44415] = 32'b11111111111111100110011001010100;
assign LUT_2[44416] = 32'b11111111111111111100100100110011;
assign LUT_2[44417] = 32'b11111111111111111001011101001100;
assign LUT_2[44418] = 32'b00000000000000000011011101101111;
assign LUT_2[44419] = 32'b00000000000000000000010110001000;
assign LUT_2[44420] = 32'b11111111111111111001000010011011;
assign LUT_2[44421] = 32'b11111111111111110101111010110100;
assign LUT_2[44422] = 32'b11111111111111111111111011010111;
assign LUT_2[44423] = 32'b11111111111111111100110011110000;
assign LUT_2[44424] = 32'b11111111111111110111010110010000;
assign LUT_2[44425] = 32'b11111111111111110100001110101001;
assign LUT_2[44426] = 32'b11111111111111111110001111001100;
assign LUT_2[44427] = 32'b11111111111111111011000111100101;
assign LUT_2[44428] = 32'b11111111111111110011110011111000;
assign LUT_2[44429] = 32'b11111111111111110000101100010001;
assign LUT_2[44430] = 32'b11111111111111111010101100110100;
assign LUT_2[44431] = 32'b11111111111111110111100101001101;
assign LUT_2[44432] = 32'b11111111111111110111001000111101;
assign LUT_2[44433] = 32'b11111111111111110100000001010110;
assign LUT_2[44434] = 32'b11111111111111111110000001111001;
assign LUT_2[44435] = 32'b11111111111111111010111010010010;
assign LUT_2[44436] = 32'b11111111111111110011100110100101;
assign LUT_2[44437] = 32'b11111111111111110000011110111110;
assign LUT_2[44438] = 32'b11111111111111111010011111100001;
assign LUT_2[44439] = 32'b11111111111111110111010111111010;
assign LUT_2[44440] = 32'b11111111111111110001111010011010;
assign LUT_2[44441] = 32'b11111111111111101110110010110011;
assign LUT_2[44442] = 32'b11111111111111111000110011010110;
assign LUT_2[44443] = 32'b11111111111111110101101011101111;
assign LUT_2[44444] = 32'b11111111111111101110011000000010;
assign LUT_2[44445] = 32'b11111111111111101011010000011011;
assign LUT_2[44446] = 32'b11111111111111110101010000111110;
assign LUT_2[44447] = 32'b11111111111111110010001001010111;
assign LUT_2[44448] = 32'b11111111111111111101000000011100;
assign LUT_2[44449] = 32'b11111111111111111001111000110101;
assign LUT_2[44450] = 32'b00000000000000000011111001011000;
assign LUT_2[44451] = 32'b00000000000000000000110001110001;
assign LUT_2[44452] = 32'b11111111111111111001011110000100;
assign LUT_2[44453] = 32'b11111111111111110110010110011101;
assign LUT_2[44454] = 32'b00000000000000000000010111000000;
assign LUT_2[44455] = 32'b11111111111111111101001111011001;
assign LUT_2[44456] = 32'b11111111111111110111110001111001;
assign LUT_2[44457] = 32'b11111111111111110100101010010010;
assign LUT_2[44458] = 32'b11111111111111111110101010110101;
assign LUT_2[44459] = 32'b11111111111111111011100011001110;
assign LUT_2[44460] = 32'b11111111111111110100001111100001;
assign LUT_2[44461] = 32'b11111111111111110001000111111010;
assign LUT_2[44462] = 32'b11111111111111111011001000011101;
assign LUT_2[44463] = 32'b11111111111111111000000000110110;
assign LUT_2[44464] = 32'b11111111111111110111100100100110;
assign LUT_2[44465] = 32'b11111111111111110100011100111111;
assign LUT_2[44466] = 32'b11111111111111111110011101100010;
assign LUT_2[44467] = 32'b11111111111111111011010101111011;
assign LUT_2[44468] = 32'b11111111111111110100000010001110;
assign LUT_2[44469] = 32'b11111111111111110000111010100111;
assign LUT_2[44470] = 32'b11111111111111111010111011001010;
assign LUT_2[44471] = 32'b11111111111111110111110011100011;
assign LUT_2[44472] = 32'b11111111111111110010010110000011;
assign LUT_2[44473] = 32'b11111111111111101111001110011100;
assign LUT_2[44474] = 32'b11111111111111111001001110111111;
assign LUT_2[44475] = 32'b11111111111111110110000111011000;
assign LUT_2[44476] = 32'b11111111111111101110110011101011;
assign LUT_2[44477] = 32'b11111111111111101011101100000100;
assign LUT_2[44478] = 32'b11111111111111110101101100100111;
assign LUT_2[44479] = 32'b11111111111111110010100101000000;
assign LUT_2[44480] = 32'b11111111111111110100101101010110;
assign LUT_2[44481] = 32'b11111111111111110001100101101111;
assign LUT_2[44482] = 32'b11111111111111111011100110010010;
assign LUT_2[44483] = 32'b11111111111111111000011110101011;
assign LUT_2[44484] = 32'b11111111111111110001001010111110;
assign LUT_2[44485] = 32'b11111111111111101110000011010111;
assign LUT_2[44486] = 32'b11111111111111111000000011111010;
assign LUT_2[44487] = 32'b11111111111111110100111100010011;
assign LUT_2[44488] = 32'b11111111111111101111011110110011;
assign LUT_2[44489] = 32'b11111111111111101100010111001100;
assign LUT_2[44490] = 32'b11111111111111110110010111101111;
assign LUT_2[44491] = 32'b11111111111111110011010000001000;
assign LUT_2[44492] = 32'b11111111111111101011111100011011;
assign LUT_2[44493] = 32'b11111111111111101000110100110100;
assign LUT_2[44494] = 32'b11111111111111110010110101010111;
assign LUT_2[44495] = 32'b11111111111111101111101101110000;
assign LUT_2[44496] = 32'b11111111111111101111010001100000;
assign LUT_2[44497] = 32'b11111111111111101100001001111001;
assign LUT_2[44498] = 32'b11111111111111110110001010011100;
assign LUT_2[44499] = 32'b11111111111111110011000010110101;
assign LUT_2[44500] = 32'b11111111111111101011101111001000;
assign LUT_2[44501] = 32'b11111111111111101000100111100001;
assign LUT_2[44502] = 32'b11111111111111110010101000000100;
assign LUT_2[44503] = 32'b11111111111111101111100000011101;
assign LUT_2[44504] = 32'b11111111111111101010000010111101;
assign LUT_2[44505] = 32'b11111111111111100110111011010110;
assign LUT_2[44506] = 32'b11111111111111110000111011111001;
assign LUT_2[44507] = 32'b11111111111111101101110100010010;
assign LUT_2[44508] = 32'b11111111111111100110100000100101;
assign LUT_2[44509] = 32'b11111111111111100011011000111110;
assign LUT_2[44510] = 32'b11111111111111101101011001100001;
assign LUT_2[44511] = 32'b11111111111111101010010001111010;
assign LUT_2[44512] = 32'b11111111111111110101001000111111;
assign LUT_2[44513] = 32'b11111111111111110010000001011000;
assign LUT_2[44514] = 32'b11111111111111111100000001111011;
assign LUT_2[44515] = 32'b11111111111111111000111010010100;
assign LUT_2[44516] = 32'b11111111111111110001100110100111;
assign LUT_2[44517] = 32'b11111111111111101110011111000000;
assign LUT_2[44518] = 32'b11111111111111111000011111100011;
assign LUT_2[44519] = 32'b11111111111111110101010111111100;
assign LUT_2[44520] = 32'b11111111111111101111111010011100;
assign LUT_2[44521] = 32'b11111111111111101100110010110101;
assign LUT_2[44522] = 32'b11111111111111110110110011011000;
assign LUT_2[44523] = 32'b11111111111111110011101011110001;
assign LUT_2[44524] = 32'b11111111111111101100011000000100;
assign LUT_2[44525] = 32'b11111111111111101001010000011101;
assign LUT_2[44526] = 32'b11111111111111110011010001000000;
assign LUT_2[44527] = 32'b11111111111111110000001001011001;
assign LUT_2[44528] = 32'b11111111111111101111101101001001;
assign LUT_2[44529] = 32'b11111111111111101100100101100010;
assign LUT_2[44530] = 32'b11111111111111110110100110000101;
assign LUT_2[44531] = 32'b11111111111111110011011110011110;
assign LUT_2[44532] = 32'b11111111111111101100001010110001;
assign LUT_2[44533] = 32'b11111111111111101001000011001010;
assign LUT_2[44534] = 32'b11111111111111110011000011101101;
assign LUT_2[44535] = 32'b11111111111111101111111100000110;
assign LUT_2[44536] = 32'b11111111111111101010011110100110;
assign LUT_2[44537] = 32'b11111111111111100111010110111111;
assign LUT_2[44538] = 32'b11111111111111110001010111100010;
assign LUT_2[44539] = 32'b11111111111111101110001111111011;
assign LUT_2[44540] = 32'b11111111111111100110111100001110;
assign LUT_2[44541] = 32'b11111111111111100011110100100111;
assign LUT_2[44542] = 32'b11111111111111101101110101001010;
assign LUT_2[44543] = 32'b11111111111111101010101101100011;
assign LUT_2[44544] = 32'b11111111111111111001000011110000;
assign LUT_2[44545] = 32'b11111111111111110101111100001001;
assign LUT_2[44546] = 32'b11111111111111111111111100101100;
assign LUT_2[44547] = 32'b11111111111111111100110101000101;
assign LUT_2[44548] = 32'b11111111111111110101100001011000;
assign LUT_2[44549] = 32'b11111111111111110010011001110001;
assign LUT_2[44550] = 32'b11111111111111111100011010010100;
assign LUT_2[44551] = 32'b11111111111111111001010010101101;
assign LUT_2[44552] = 32'b11111111111111110011110101001101;
assign LUT_2[44553] = 32'b11111111111111110000101101100110;
assign LUT_2[44554] = 32'b11111111111111111010101110001001;
assign LUT_2[44555] = 32'b11111111111111110111100110100010;
assign LUT_2[44556] = 32'b11111111111111110000010010110101;
assign LUT_2[44557] = 32'b11111111111111101101001011001110;
assign LUT_2[44558] = 32'b11111111111111110111001011110001;
assign LUT_2[44559] = 32'b11111111111111110100000100001010;
assign LUT_2[44560] = 32'b11111111111111110011100111111010;
assign LUT_2[44561] = 32'b11111111111111110000100000010011;
assign LUT_2[44562] = 32'b11111111111111111010100000110110;
assign LUT_2[44563] = 32'b11111111111111110111011001001111;
assign LUT_2[44564] = 32'b11111111111111110000000101100010;
assign LUT_2[44565] = 32'b11111111111111101100111101111011;
assign LUT_2[44566] = 32'b11111111111111110110111110011110;
assign LUT_2[44567] = 32'b11111111111111110011110110110111;
assign LUT_2[44568] = 32'b11111111111111101110011001010111;
assign LUT_2[44569] = 32'b11111111111111101011010001110000;
assign LUT_2[44570] = 32'b11111111111111110101010010010011;
assign LUT_2[44571] = 32'b11111111111111110010001010101100;
assign LUT_2[44572] = 32'b11111111111111101010110110111111;
assign LUT_2[44573] = 32'b11111111111111100111101111011000;
assign LUT_2[44574] = 32'b11111111111111110001101111111011;
assign LUT_2[44575] = 32'b11111111111111101110101000010100;
assign LUT_2[44576] = 32'b11111111111111111001011111011001;
assign LUT_2[44577] = 32'b11111111111111110110010111110010;
assign LUT_2[44578] = 32'b00000000000000000000011000010101;
assign LUT_2[44579] = 32'b11111111111111111101010000101110;
assign LUT_2[44580] = 32'b11111111111111110101111101000001;
assign LUT_2[44581] = 32'b11111111111111110010110101011010;
assign LUT_2[44582] = 32'b11111111111111111100110101111101;
assign LUT_2[44583] = 32'b11111111111111111001101110010110;
assign LUT_2[44584] = 32'b11111111111111110100010000110110;
assign LUT_2[44585] = 32'b11111111111111110001001001001111;
assign LUT_2[44586] = 32'b11111111111111111011001001110010;
assign LUT_2[44587] = 32'b11111111111111111000000010001011;
assign LUT_2[44588] = 32'b11111111111111110000101110011110;
assign LUT_2[44589] = 32'b11111111111111101101100110110111;
assign LUT_2[44590] = 32'b11111111111111110111100111011010;
assign LUT_2[44591] = 32'b11111111111111110100011111110011;
assign LUT_2[44592] = 32'b11111111111111110100000011100011;
assign LUT_2[44593] = 32'b11111111111111110000111011111100;
assign LUT_2[44594] = 32'b11111111111111111010111100011111;
assign LUT_2[44595] = 32'b11111111111111110111110100111000;
assign LUT_2[44596] = 32'b11111111111111110000100001001011;
assign LUT_2[44597] = 32'b11111111111111101101011001100100;
assign LUT_2[44598] = 32'b11111111111111110111011010000111;
assign LUT_2[44599] = 32'b11111111111111110100010010100000;
assign LUT_2[44600] = 32'b11111111111111101110110101000000;
assign LUT_2[44601] = 32'b11111111111111101011101101011001;
assign LUT_2[44602] = 32'b11111111111111110101101101111100;
assign LUT_2[44603] = 32'b11111111111111110010100110010101;
assign LUT_2[44604] = 32'b11111111111111101011010010101000;
assign LUT_2[44605] = 32'b11111111111111101000001011000001;
assign LUT_2[44606] = 32'b11111111111111110010001011100100;
assign LUT_2[44607] = 32'b11111111111111101111000011111101;
assign LUT_2[44608] = 32'b11111111111111110001001100010011;
assign LUT_2[44609] = 32'b11111111111111101110000100101100;
assign LUT_2[44610] = 32'b11111111111111111000000101001111;
assign LUT_2[44611] = 32'b11111111111111110100111101101000;
assign LUT_2[44612] = 32'b11111111111111101101101001111011;
assign LUT_2[44613] = 32'b11111111111111101010100010010100;
assign LUT_2[44614] = 32'b11111111111111110100100010110111;
assign LUT_2[44615] = 32'b11111111111111110001011011010000;
assign LUT_2[44616] = 32'b11111111111111101011111101110000;
assign LUT_2[44617] = 32'b11111111111111101000110110001001;
assign LUT_2[44618] = 32'b11111111111111110010110110101100;
assign LUT_2[44619] = 32'b11111111111111101111101111000101;
assign LUT_2[44620] = 32'b11111111111111101000011011011000;
assign LUT_2[44621] = 32'b11111111111111100101010011110001;
assign LUT_2[44622] = 32'b11111111111111101111010100010100;
assign LUT_2[44623] = 32'b11111111111111101100001100101101;
assign LUT_2[44624] = 32'b11111111111111101011110000011101;
assign LUT_2[44625] = 32'b11111111111111101000101000110110;
assign LUT_2[44626] = 32'b11111111111111110010101001011001;
assign LUT_2[44627] = 32'b11111111111111101111100001110010;
assign LUT_2[44628] = 32'b11111111111111101000001110000101;
assign LUT_2[44629] = 32'b11111111111111100101000110011110;
assign LUT_2[44630] = 32'b11111111111111101111000111000001;
assign LUT_2[44631] = 32'b11111111111111101011111111011010;
assign LUT_2[44632] = 32'b11111111111111100110100001111010;
assign LUT_2[44633] = 32'b11111111111111100011011010010011;
assign LUT_2[44634] = 32'b11111111111111101101011010110110;
assign LUT_2[44635] = 32'b11111111111111101010010011001111;
assign LUT_2[44636] = 32'b11111111111111100010111111100010;
assign LUT_2[44637] = 32'b11111111111111011111110111111011;
assign LUT_2[44638] = 32'b11111111111111101001111000011110;
assign LUT_2[44639] = 32'b11111111111111100110110000110111;
assign LUT_2[44640] = 32'b11111111111111110001100111111100;
assign LUT_2[44641] = 32'b11111111111111101110100000010101;
assign LUT_2[44642] = 32'b11111111111111111000100000111000;
assign LUT_2[44643] = 32'b11111111111111110101011001010001;
assign LUT_2[44644] = 32'b11111111111111101110000101100100;
assign LUT_2[44645] = 32'b11111111111111101010111101111101;
assign LUT_2[44646] = 32'b11111111111111110100111110100000;
assign LUT_2[44647] = 32'b11111111111111110001110110111001;
assign LUT_2[44648] = 32'b11111111111111101100011001011001;
assign LUT_2[44649] = 32'b11111111111111101001010001110010;
assign LUT_2[44650] = 32'b11111111111111110011010010010101;
assign LUT_2[44651] = 32'b11111111111111110000001010101110;
assign LUT_2[44652] = 32'b11111111111111101000110111000001;
assign LUT_2[44653] = 32'b11111111111111100101101111011010;
assign LUT_2[44654] = 32'b11111111111111101111101111111101;
assign LUT_2[44655] = 32'b11111111111111101100101000010110;
assign LUT_2[44656] = 32'b11111111111111101100001100000110;
assign LUT_2[44657] = 32'b11111111111111101001000100011111;
assign LUT_2[44658] = 32'b11111111111111110011000101000010;
assign LUT_2[44659] = 32'b11111111111111101111111101011011;
assign LUT_2[44660] = 32'b11111111111111101000101001101110;
assign LUT_2[44661] = 32'b11111111111111100101100010000111;
assign LUT_2[44662] = 32'b11111111111111101111100010101010;
assign LUT_2[44663] = 32'b11111111111111101100011011000011;
assign LUT_2[44664] = 32'b11111111111111100110111101100011;
assign LUT_2[44665] = 32'b11111111111111100011110101111100;
assign LUT_2[44666] = 32'b11111111111111101101110110011111;
assign LUT_2[44667] = 32'b11111111111111101010101110111000;
assign LUT_2[44668] = 32'b11111111111111100011011011001011;
assign LUT_2[44669] = 32'b11111111111111100000010011100100;
assign LUT_2[44670] = 32'b11111111111111101010010100000111;
assign LUT_2[44671] = 32'b11111111111111100111001100100000;
assign LUT_2[44672] = 32'b11111111111111111101010111111111;
assign LUT_2[44673] = 32'b11111111111111111010010000011000;
assign LUT_2[44674] = 32'b00000000000000000100010000111011;
assign LUT_2[44675] = 32'b00000000000000000001001001010100;
assign LUT_2[44676] = 32'b11111111111111111001110101100111;
assign LUT_2[44677] = 32'b11111111111111110110101110000000;
assign LUT_2[44678] = 32'b00000000000000000000101110100011;
assign LUT_2[44679] = 32'b11111111111111111101100110111100;
assign LUT_2[44680] = 32'b11111111111111111000001001011100;
assign LUT_2[44681] = 32'b11111111111111110101000001110101;
assign LUT_2[44682] = 32'b11111111111111111111000010011000;
assign LUT_2[44683] = 32'b11111111111111111011111010110001;
assign LUT_2[44684] = 32'b11111111111111110100100111000100;
assign LUT_2[44685] = 32'b11111111111111110001011111011101;
assign LUT_2[44686] = 32'b11111111111111111011100000000000;
assign LUT_2[44687] = 32'b11111111111111111000011000011001;
assign LUT_2[44688] = 32'b11111111111111110111111100001001;
assign LUT_2[44689] = 32'b11111111111111110100110100100010;
assign LUT_2[44690] = 32'b11111111111111111110110101000101;
assign LUT_2[44691] = 32'b11111111111111111011101101011110;
assign LUT_2[44692] = 32'b11111111111111110100011001110001;
assign LUT_2[44693] = 32'b11111111111111110001010010001010;
assign LUT_2[44694] = 32'b11111111111111111011010010101101;
assign LUT_2[44695] = 32'b11111111111111111000001011000110;
assign LUT_2[44696] = 32'b11111111111111110010101101100110;
assign LUT_2[44697] = 32'b11111111111111101111100101111111;
assign LUT_2[44698] = 32'b11111111111111111001100110100010;
assign LUT_2[44699] = 32'b11111111111111110110011110111011;
assign LUT_2[44700] = 32'b11111111111111101111001011001110;
assign LUT_2[44701] = 32'b11111111111111101100000011100111;
assign LUT_2[44702] = 32'b11111111111111110110000100001010;
assign LUT_2[44703] = 32'b11111111111111110010111100100011;
assign LUT_2[44704] = 32'b11111111111111111101110011101000;
assign LUT_2[44705] = 32'b11111111111111111010101100000001;
assign LUT_2[44706] = 32'b00000000000000000100101100100100;
assign LUT_2[44707] = 32'b00000000000000000001100100111101;
assign LUT_2[44708] = 32'b11111111111111111010010001010000;
assign LUT_2[44709] = 32'b11111111111111110111001001101001;
assign LUT_2[44710] = 32'b00000000000000000001001010001100;
assign LUT_2[44711] = 32'b11111111111111111110000010100101;
assign LUT_2[44712] = 32'b11111111111111111000100101000101;
assign LUT_2[44713] = 32'b11111111111111110101011101011110;
assign LUT_2[44714] = 32'b11111111111111111111011110000001;
assign LUT_2[44715] = 32'b11111111111111111100010110011010;
assign LUT_2[44716] = 32'b11111111111111110101000010101101;
assign LUT_2[44717] = 32'b11111111111111110001111011000110;
assign LUT_2[44718] = 32'b11111111111111111011111011101001;
assign LUT_2[44719] = 32'b11111111111111111000110100000010;
assign LUT_2[44720] = 32'b11111111111111111000010111110010;
assign LUT_2[44721] = 32'b11111111111111110101010000001011;
assign LUT_2[44722] = 32'b11111111111111111111010000101110;
assign LUT_2[44723] = 32'b11111111111111111100001001000111;
assign LUT_2[44724] = 32'b11111111111111110100110101011010;
assign LUT_2[44725] = 32'b11111111111111110001101101110011;
assign LUT_2[44726] = 32'b11111111111111111011101110010110;
assign LUT_2[44727] = 32'b11111111111111111000100110101111;
assign LUT_2[44728] = 32'b11111111111111110011001001001111;
assign LUT_2[44729] = 32'b11111111111111110000000001101000;
assign LUT_2[44730] = 32'b11111111111111111010000010001011;
assign LUT_2[44731] = 32'b11111111111111110110111010100100;
assign LUT_2[44732] = 32'b11111111111111101111100110110111;
assign LUT_2[44733] = 32'b11111111111111101100011111010000;
assign LUT_2[44734] = 32'b11111111111111110110011111110011;
assign LUT_2[44735] = 32'b11111111111111110011011000001100;
assign LUT_2[44736] = 32'b11111111111111110101100000100010;
assign LUT_2[44737] = 32'b11111111111111110010011000111011;
assign LUT_2[44738] = 32'b11111111111111111100011001011110;
assign LUT_2[44739] = 32'b11111111111111111001010001110111;
assign LUT_2[44740] = 32'b11111111111111110001111110001010;
assign LUT_2[44741] = 32'b11111111111111101110110110100011;
assign LUT_2[44742] = 32'b11111111111111111000110111000110;
assign LUT_2[44743] = 32'b11111111111111110101101111011111;
assign LUT_2[44744] = 32'b11111111111111110000010001111111;
assign LUT_2[44745] = 32'b11111111111111101101001010011000;
assign LUT_2[44746] = 32'b11111111111111110111001010111011;
assign LUT_2[44747] = 32'b11111111111111110100000011010100;
assign LUT_2[44748] = 32'b11111111111111101100101111100111;
assign LUT_2[44749] = 32'b11111111111111101001101000000000;
assign LUT_2[44750] = 32'b11111111111111110011101000100011;
assign LUT_2[44751] = 32'b11111111111111110000100000111100;
assign LUT_2[44752] = 32'b11111111111111110000000100101100;
assign LUT_2[44753] = 32'b11111111111111101100111101000101;
assign LUT_2[44754] = 32'b11111111111111110110111101101000;
assign LUT_2[44755] = 32'b11111111111111110011110110000001;
assign LUT_2[44756] = 32'b11111111111111101100100010010100;
assign LUT_2[44757] = 32'b11111111111111101001011010101101;
assign LUT_2[44758] = 32'b11111111111111110011011011010000;
assign LUT_2[44759] = 32'b11111111111111110000010011101001;
assign LUT_2[44760] = 32'b11111111111111101010110110001001;
assign LUT_2[44761] = 32'b11111111111111100111101110100010;
assign LUT_2[44762] = 32'b11111111111111110001101111000101;
assign LUT_2[44763] = 32'b11111111111111101110100111011110;
assign LUT_2[44764] = 32'b11111111111111100111010011110001;
assign LUT_2[44765] = 32'b11111111111111100100001100001010;
assign LUT_2[44766] = 32'b11111111111111101110001100101101;
assign LUT_2[44767] = 32'b11111111111111101011000101000110;
assign LUT_2[44768] = 32'b11111111111111110101111100001011;
assign LUT_2[44769] = 32'b11111111111111110010110100100100;
assign LUT_2[44770] = 32'b11111111111111111100110101000111;
assign LUT_2[44771] = 32'b11111111111111111001101101100000;
assign LUT_2[44772] = 32'b11111111111111110010011001110011;
assign LUT_2[44773] = 32'b11111111111111101111010010001100;
assign LUT_2[44774] = 32'b11111111111111111001010010101111;
assign LUT_2[44775] = 32'b11111111111111110110001011001000;
assign LUT_2[44776] = 32'b11111111111111110000101101101000;
assign LUT_2[44777] = 32'b11111111111111101101100110000001;
assign LUT_2[44778] = 32'b11111111111111110111100110100100;
assign LUT_2[44779] = 32'b11111111111111110100011110111101;
assign LUT_2[44780] = 32'b11111111111111101101001011010000;
assign LUT_2[44781] = 32'b11111111111111101010000011101001;
assign LUT_2[44782] = 32'b11111111111111110100000100001100;
assign LUT_2[44783] = 32'b11111111111111110000111100100101;
assign LUT_2[44784] = 32'b11111111111111110000100000010101;
assign LUT_2[44785] = 32'b11111111111111101101011000101110;
assign LUT_2[44786] = 32'b11111111111111110111011001010001;
assign LUT_2[44787] = 32'b11111111111111110100010001101010;
assign LUT_2[44788] = 32'b11111111111111101100111101111101;
assign LUT_2[44789] = 32'b11111111111111101001110110010110;
assign LUT_2[44790] = 32'b11111111111111110011110110111001;
assign LUT_2[44791] = 32'b11111111111111110000101111010010;
assign LUT_2[44792] = 32'b11111111111111101011010001110010;
assign LUT_2[44793] = 32'b11111111111111101000001010001011;
assign LUT_2[44794] = 32'b11111111111111110010001010101110;
assign LUT_2[44795] = 32'b11111111111111101111000011000111;
assign LUT_2[44796] = 32'b11111111111111100111101111011010;
assign LUT_2[44797] = 32'b11111111111111100100100111110011;
assign LUT_2[44798] = 32'b11111111111111101110101000010110;
assign LUT_2[44799] = 32'b11111111111111101011100000101111;
assign LUT_2[44800] = 32'b11111111111111111101000010010110;
assign LUT_2[44801] = 32'b11111111111111111001111010101111;
assign LUT_2[44802] = 32'b00000000000000000011111011010010;
assign LUT_2[44803] = 32'b00000000000000000000110011101011;
assign LUT_2[44804] = 32'b11111111111111111001011111111110;
assign LUT_2[44805] = 32'b11111111111111110110011000010111;
assign LUT_2[44806] = 32'b00000000000000000000011000111010;
assign LUT_2[44807] = 32'b11111111111111111101010001010011;
assign LUT_2[44808] = 32'b11111111111111110111110011110011;
assign LUT_2[44809] = 32'b11111111111111110100101100001100;
assign LUT_2[44810] = 32'b11111111111111111110101100101111;
assign LUT_2[44811] = 32'b11111111111111111011100101001000;
assign LUT_2[44812] = 32'b11111111111111110100010001011011;
assign LUT_2[44813] = 32'b11111111111111110001001001110100;
assign LUT_2[44814] = 32'b11111111111111111011001010010111;
assign LUT_2[44815] = 32'b11111111111111111000000010110000;
assign LUT_2[44816] = 32'b11111111111111110111100110100000;
assign LUT_2[44817] = 32'b11111111111111110100011110111001;
assign LUT_2[44818] = 32'b11111111111111111110011111011100;
assign LUT_2[44819] = 32'b11111111111111111011010111110101;
assign LUT_2[44820] = 32'b11111111111111110100000100001000;
assign LUT_2[44821] = 32'b11111111111111110000111100100001;
assign LUT_2[44822] = 32'b11111111111111111010111101000100;
assign LUT_2[44823] = 32'b11111111111111110111110101011101;
assign LUT_2[44824] = 32'b11111111111111110010010111111101;
assign LUT_2[44825] = 32'b11111111111111101111010000010110;
assign LUT_2[44826] = 32'b11111111111111111001010000111001;
assign LUT_2[44827] = 32'b11111111111111110110001001010010;
assign LUT_2[44828] = 32'b11111111111111101110110101100101;
assign LUT_2[44829] = 32'b11111111111111101011101101111110;
assign LUT_2[44830] = 32'b11111111111111110101101110100001;
assign LUT_2[44831] = 32'b11111111111111110010100110111010;
assign LUT_2[44832] = 32'b11111111111111111101011101111111;
assign LUT_2[44833] = 32'b11111111111111111010010110011000;
assign LUT_2[44834] = 32'b00000000000000000100010110111011;
assign LUT_2[44835] = 32'b00000000000000000001001111010100;
assign LUT_2[44836] = 32'b11111111111111111001111011100111;
assign LUT_2[44837] = 32'b11111111111111110110110100000000;
assign LUT_2[44838] = 32'b00000000000000000000110100100011;
assign LUT_2[44839] = 32'b11111111111111111101101100111100;
assign LUT_2[44840] = 32'b11111111111111111000001111011100;
assign LUT_2[44841] = 32'b11111111111111110101000111110101;
assign LUT_2[44842] = 32'b11111111111111111111001000011000;
assign LUT_2[44843] = 32'b11111111111111111100000000110001;
assign LUT_2[44844] = 32'b11111111111111110100101101000100;
assign LUT_2[44845] = 32'b11111111111111110001100101011101;
assign LUT_2[44846] = 32'b11111111111111111011100110000000;
assign LUT_2[44847] = 32'b11111111111111111000011110011001;
assign LUT_2[44848] = 32'b11111111111111111000000010001001;
assign LUT_2[44849] = 32'b11111111111111110100111010100010;
assign LUT_2[44850] = 32'b11111111111111111110111011000101;
assign LUT_2[44851] = 32'b11111111111111111011110011011110;
assign LUT_2[44852] = 32'b11111111111111110100011111110001;
assign LUT_2[44853] = 32'b11111111111111110001011000001010;
assign LUT_2[44854] = 32'b11111111111111111011011000101101;
assign LUT_2[44855] = 32'b11111111111111111000010001000110;
assign LUT_2[44856] = 32'b11111111111111110010110011100110;
assign LUT_2[44857] = 32'b11111111111111101111101011111111;
assign LUT_2[44858] = 32'b11111111111111111001101100100010;
assign LUT_2[44859] = 32'b11111111111111110110100100111011;
assign LUT_2[44860] = 32'b11111111111111101111010001001110;
assign LUT_2[44861] = 32'b11111111111111101100001001100111;
assign LUT_2[44862] = 32'b11111111111111110110001010001010;
assign LUT_2[44863] = 32'b11111111111111110011000010100011;
assign LUT_2[44864] = 32'b11111111111111110101001010111001;
assign LUT_2[44865] = 32'b11111111111111110010000011010010;
assign LUT_2[44866] = 32'b11111111111111111100000011110101;
assign LUT_2[44867] = 32'b11111111111111111000111100001110;
assign LUT_2[44868] = 32'b11111111111111110001101000100001;
assign LUT_2[44869] = 32'b11111111111111101110100000111010;
assign LUT_2[44870] = 32'b11111111111111111000100001011101;
assign LUT_2[44871] = 32'b11111111111111110101011001110110;
assign LUT_2[44872] = 32'b11111111111111101111111100010110;
assign LUT_2[44873] = 32'b11111111111111101100110100101111;
assign LUT_2[44874] = 32'b11111111111111110110110101010010;
assign LUT_2[44875] = 32'b11111111111111110011101101101011;
assign LUT_2[44876] = 32'b11111111111111101100011001111110;
assign LUT_2[44877] = 32'b11111111111111101001010010010111;
assign LUT_2[44878] = 32'b11111111111111110011010010111010;
assign LUT_2[44879] = 32'b11111111111111110000001011010011;
assign LUT_2[44880] = 32'b11111111111111101111101111000011;
assign LUT_2[44881] = 32'b11111111111111101100100111011100;
assign LUT_2[44882] = 32'b11111111111111110110100111111111;
assign LUT_2[44883] = 32'b11111111111111110011100000011000;
assign LUT_2[44884] = 32'b11111111111111101100001100101011;
assign LUT_2[44885] = 32'b11111111111111101001000101000100;
assign LUT_2[44886] = 32'b11111111111111110011000101100111;
assign LUT_2[44887] = 32'b11111111111111101111111110000000;
assign LUT_2[44888] = 32'b11111111111111101010100000100000;
assign LUT_2[44889] = 32'b11111111111111100111011000111001;
assign LUT_2[44890] = 32'b11111111111111110001011001011100;
assign LUT_2[44891] = 32'b11111111111111101110010001110101;
assign LUT_2[44892] = 32'b11111111111111100110111110001000;
assign LUT_2[44893] = 32'b11111111111111100011110110100001;
assign LUT_2[44894] = 32'b11111111111111101101110111000100;
assign LUT_2[44895] = 32'b11111111111111101010101111011101;
assign LUT_2[44896] = 32'b11111111111111110101100110100010;
assign LUT_2[44897] = 32'b11111111111111110010011110111011;
assign LUT_2[44898] = 32'b11111111111111111100011111011110;
assign LUT_2[44899] = 32'b11111111111111111001010111110111;
assign LUT_2[44900] = 32'b11111111111111110010000100001010;
assign LUT_2[44901] = 32'b11111111111111101110111100100011;
assign LUT_2[44902] = 32'b11111111111111111000111101000110;
assign LUT_2[44903] = 32'b11111111111111110101110101011111;
assign LUT_2[44904] = 32'b11111111111111110000010111111111;
assign LUT_2[44905] = 32'b11111111111111101101010000011000;
assign LUT_2[44906] = 32'b11111111111111110111010000111011;
assign LUT_2[44907] = 32'b11111111111111110100001001010100;
assign LUT_2[44908] = 32'b11111111111111101100110101100111;
assign LUT_2[44909] = 32'b11111111111111101001101110000000;
assign LUT_2[44910] = 32'b11111111111111110011101110100011;
assign LUT_2[44911] = 32'b11111111111111110000100110111100;
assign LUT_2[44912] = 32'b11111111111111110000001010101100;
assign LUT_2[44913] = 32'b11111111111111101101000011000101;
assign LUT_2[44914] = 32'b11111111111111110111000011101000;
assign LUT_2[44915] = 32'b11111111111111110011111100000001;
assign LUT_2[44916] = 32'b11111111111111101100101000010100;
assign LUT_2[44917] = 32'b11111111111111101001100000101101;
assign LUT_2[44918] = 32'b11111111111111110011100001010000;
assign LUT_2[44919] = 32'b11111111111111110000011001101001;
assign LUT_2[44920] = 32'b11111111111111101010111100001001;
assign LUT_2[44921] = 32'b11111111111111100111110100100010;
assign LUT_2[44922] = 32'b11111111111111110001110101000101;
assign LUT_2[44923] = 32'b11111111111111101110101101011110;
assign LUT_2[44924] = 32'b11111111111111100111011001110001;
assign LUT_2[44925] = 32'b11111111111111100100010010001010;
assign LUT_2[44926] = 32'b11111111111111101110010010101101;
assign LUT_2[44927] = 32'b11111111111111101011001011000110;
assign LUT_2[44928] = 32'b00000000000000000001010110100101;
assign LUT_2[44929] = 32'b11111111111111111110001110111110;
assign LUT_2[44930] = 32'b00000000000000001000001111100001;
assign LUT_2[44931] = 32'b00000000000000000101000111111010;
assign LUT_2[44932] = 32'b11111111111111111101110100001101;
assign LUT_2[44933] = 32'b11111111111111111010101100100110;
assign LUT_2[44934] = 32'b00000000000000000100101101001001;
assign LUT_2[44935] = 32'b00000000000000000001100101100010;
assign LUT_2[44936] = 32'b11111111111111111100001000000010;
assign LUT_2[44937] = 32'b11111111111111111001000000011011;
assign LUT_2[44938] = 32'b00000000000000000011000000111110;
assign LUT_2[44939] = 32'b11111111111111111111111001010111;
assign LUT_2[44940] = 32'b11111111111111111000100101101010;
assign LUT_2[44941] = 32'b11111111111111110101011110000011;
assign LUT_2[44942] = 32'b11111111111111111111011110100110;
assign LUT_2[44943] = 32'b11111111111111111100010110111111;
assign LUT_2[44944] = 32'b11111111111111111011111010101111;
assign LUT_2[44945] = 32'b11111111111111111000110011001000;
assign LUT_2[44946] = 32'b00000000000000000010110011101011;
assign LUT_2[44947] = 32'b11111111111111111111101100000100;
assign LUT_2[44948] = 32'b11111111111111111000011000010111;
assign LUT_2[44949] = 32'b11111111111111110101010000110000;
assign LUT_2[44950] = 32'b11111111111111111111010001010011;
assign LUT_2[44951] = 32'b11111111111111111100001001101100;
assign LUT_2[44952] = 32'b11111111111111110110101100001100;
assign LUT_2[44953] = 32'b11111111111111110011100100100101;
assign LUT_2[44954] = 32'b11111111111111111101100101001000;
assign LUT_2[44955] = 32'b11111111111111111010011101100001;
assign LUT_2[44956] = 32'b11111111111111110011001001110100;
assign LUT_2[44957] = 32'b11111111111111110000000010001101;
assign LUT_2[44958] = 32'b11111111111111111010000010110000;
assign LUT_2[44959] = 32'b11111111111111110110111011001001;
assign LUT_2[44960] = 32'b00000000000000000001110010001110;
assign LUT_2[44961] = 32'b11111111111111111110101010100111;
assign LUT_2[44962] = 32'b00000000000000001000101011001010;
assign LUT_2[44963] = 32'b00000000000000000101100011100011;
assign LUT_2[44964] = 32'b11111111111111111110001111110110;
assign LUT_2[44965] = 32'b11111111111111111011001000001111;
assign LUT_2[44966] = 32'b00000000000000000101001000110010;
assign LUT_2[44967] = 32'b00000000000000000010000001001011;
assign LUT_2[44968] = 32'b11111111111111111100100011101011;
assign LUT_2[44969] = 32'b11111111111111111001011100000100;
assign LUT_2[44970] = 32'b00000000000000000011011100100111;
assign LUT_2[44971] = 32'b00000000000000000000010101000000;
assign LUT_2[44972] = 32'b11111111111111111001000001010011;
assign LUT_2[44973] = 32'b11111111111111110101111001101100;
assign LUT_2[44974] = 32'b11111111111111111111111010001111;
assign LUT_2[44975] = 32'b11111111111111111100110010101000;
assign LUT_2[44976] = 32'b11111111111111111100010110011000;
assign LUT_2[44977] = 32'b11111111111111111001001110110001;
assign LUT_2[44978] = 32'b00000000000000000011001111010100;
assign LUT_2[44979] = 32'b00000000000000000000000111101101;
assign LUT_2[44980] = 32'b11111111111111111000110100000000;
assign LUT_2[44981] = 32'b11111111111111110101101100011001;
assign LUT_2[44982] = 32'b11111111111111111111101100111100;
assign LUT_2[44983] = 32'b11111111111111111100100101010101;
assign LUT_2[44984] = 32'b11111111111111110111000111110101;
assign LUT_2[44985] = 32'b11111111111111110100000000001110;
assign LUT_2[44986] = 32'b11111111111111111110000000110001;
assign LUT_2[44987] = 32'b11111111111111111010111001001010;
assign LUT_2[44988] = 32'b11111111111111110011100101011101;
assign LUT_2[44989] = 32'b11111111111111110000011101110110;
assign LUT_2[44990] = 32'b11111111111111111010011110011001;
assign LUT_2[44991] = 32'b11111111111111110111010110110010;
assign LUT_2[44992] = 32'b11111111111111111001011111001000;
assign LUT_2[44993] = 32'b11111111111111110110010111100001;
assign LUT_2[44994] = 32'b00000000000000000000011000000100;
assign LUT_2[44995] = 32'b11111111111111111101010000011101;
assign LUT_2[44996] = 32'b11111111111111110101111100110000;
assign LUT_2[44997] = 32'b11111111111111110010110101001001;
assign LUT_2[44998] = 32'b11111111111111111100110101101100;
assign LUT_2[44999] = 32'b11111111111111111001101110000101;
assign LUT_2[45000] = 32'b11111111111111110100010000100101;
assign LUT_2[45001] = 32'b11111111111111110001001000111110;
assign LUT_2[45002] = 32'b11111111111111111011001001100001;
assign LUT_2[45003] = 32'b11111111111111111000000001111010;
assign LUT_2[45004] = 32'b11111111111111110000101110001101;
assign LUT_2[45005] = 32'b11111111111111101101100110100110;
assign LUT_2[45006] = 32'b11111111111111110111100111001001;
assign LUT_2[45007] = 32'b11111111111111110100011111100010;
assign LUT_2[45008] = 32'b11111111111111110100000011010010;
assign LUT_2[45009] = 32'b11111111111111110000111011101011;
assign LUT_2[45010] = 32'b11111111111111111010111100001110;
assign LUT_2[45011] = 32'b11111111111111110111110100100111;
assign LUT_2[45012] = 32'b11111111111111110000100000111010;
assign LUT_2[45013] = 32'b11111111111111101101011001010011;
assign LUT_2[45014] = 32'b11111111111111110111011001110110;
assign LUT_2[45015] = 32'b11111111111111110100010010001111;
assign LUT_2[45016] = 32'b11111111111111101110110100101111;
assign LUT_2[45017] = 32'b11111111111111101011101101001000;
assign LUT_2[45018] = 32'b11111111111111110101101101101011;
assign LUT_2[45019] = 32'b11111111111111110010100110000100;
assign LUT_2[45020] = 32'b11111111111111101011010010010111;
assign LUT_2[45021] = 32'b11111111111111101000001010110000;
assign LUT_2[45022] = 32'b11111111111111110010001011010011;
assign LUT_2[45023] = 32'b11111111111111101111000011101100;
assign LUT_2[45024] = 32'b11111111111111111001111010110001;
assign LUT_2[45025] = 32'b11111111111111110110110011001010;
assign LUT_2[45026] = 32'b00000000000000000000110011101101;
assign LUT_2[45027] = 32'b11111111111111111101101100000110;
assign LUT_2[45028] = 32'b11111111111111110110011000011001;
assign LUT_2[45029] = 32'b11111111111111110011010000110010;
assign LUT_2[45030] = 32'b11111111111111111101010001010101;
assign LUT_2[45031] = 32'b11111111111111111010001001101110;
assign LUT_2[45032] = 32'b11111111111111110100101100001110;
assign LUT_2[45033] = 32'b11111111111111110001100100100111;
assign LUT_2[45034] = 32'b11111111111111111011100101001010;
assign LUT_2[45035] = 32'b11111111111111111000011101100011;
assign LUT_2[45036] = 32'b11111111111111110001001001110110;
assign LUT_2[45037] = 32'b11111111111111101110000010001111;
assign LUT_2[45038] = 32'b11111111111111111000000010110010;
assign LUT_2[45039] = 32'b11111111111111110100111011001011;
assign LUT_2[45040] = 32'b11111111111111110100011110111011;
assign LUT_2[45041] = 32'b11111111111111110001010111010100;
assign LUT_2[45042] = 32'b11111111111111111011010111110111;
assign LUT_2[45043] = 32'b11111111111111111000010000010000;
assign LUT_2[45044] = 32'b11111111111111110000111100100011;
assign LUT_2[45045] = 32'b11111111111111101101110100111100;
assign LUT_2[45046] = 32'b11111111111111110111110101011111;
assign LUT_2[45047] = 32'b11111111111111110100101101111000;
assign LUT_2[45048] = 32'b11111111111111101111010000011000;
assign LUT_2[45049] = 32'b11111111111111101100001000110001;
assign LUT_2[45050] = 32'b11111111111111110110001001010100;
assign LUT_2[45051] = 32'b11111111111111110011000001101101;
assign LUT_2[45052] = 32'b11111111111111101011101110000000;
assign LUT_2[45053] = 32'b11111111111111101000100110011001;
assign LUT_2[45054] = 32'b11111111111111110010100110111100;
assign LUT_2[45055] = 32'b11111111111111101111011111010101;
assign LUT_2[45056] = 32'b11111111111111110000110100001000;
assign LUT_2[45057] = 32'b11111111111111101101101100100001;
assign LUT_2[45058] = 32'b11111111111111110111101101000100;
assign LUT_2[45059] = 32'b11111111111111110100100101011101;
assign LUT_2[45060] = 32'b11111111111111101101010001110000;
assign LUT_2[45061] = 32'b11111111111111101010001010001001;
assign LUT_2[45062] = 32'b11111111111111110100001010101100;
assign LUT_2[45063] = 32'b11111111111111110001000011000101;
assign LUT_2[45064] = 32'b11111111111111101011100101100101;
assign LUT_2[45065] = 32'b11111111111111101000011101111110;
assign LUT_2[45066] = 32'b11111111111111110010011110100001;
assign LUT_2[45067] = 32'b11111111111111101111010110111010;
assign LUT_2[45068] = 32'b11111111111111101000000011001101;
assign LUT_2[45069] = 32'b11111111111111100100111011100110;
assign LUT_2[45070] = 32'b11111111111111101110111100001001;
assign LUT_2[45071] = 32'b11111111111111101011110100100010;
assign LUT_2[45072] = 32'b11111111111111101011011000010010;
assign LUT_2[45073] = 32'b11111111111111101000010000101011;
assign LUT_2[45074] = 32'b11111111111111110010010001001110;
assign LUT_2[45075] = 32'b11111111111111101111001001100111;
assign LUT_2[45076] = 32'b11111111111111100111110101111010;
assign LUT_2[45077] = 32'b11111111111111100100101110010011;
assign LUT_2[45078] = 32'b11111111111111101110101110110110;
assign LUT_2[45079] = 32'b11111111111111101011100111001111;
assign LUT_2[45080] = 32'b11111111111111100110001001101111;
assign LUT_2[45081] = 32'b11111111111111100011000010001000;
assign LUT_2[45082] = 32'b11111111111111101101000010101011;
assign LUT_2[45083] = 32'b11111111111111101001111011000100;
assign LUT_2[45084] = 32'b11111111111111100010100111010111;
assign LUT_2[45085] = 32'b11111111111111011111011111110000;
assign LUT_2[45086] = 32'b11111111111111101001100000010011;
assign LUT_2[45087] = 32'b11111111111111100110011000101100;
assign LUT_2[45088] = 32'b11111111111111110001001111110001;
assign LUT_2[45089] = 32'b11111111111111101110001000001010;
assign LUT_2[45090] = 32'b11111111111111111000001000101101;
assign LUT_2[45091] = 32'b11111111111111110101000001000110;
assign LUT_2[45092] = 32'b11111111111111101101101101011001;
assign LUT_2[45093] = 32'b11111111111111101010100101110010;
assign LUT_2[45094] = 32'b11111111111111110100100110010101;
assign LUT_2[45095] = 32'b11111111111111110001011110101110;
assign LUT_2[45096] = 32'b11111111111111101100000001001110;
assign LUT_2[45097] = 32'b11111111111111101000111001100111;
assign LUT_2[45098] = 32'b11111111111111110010111010001010;
assign LUT_2[45099] = 32'b11111111111111101111110010100011;
assign LUT_2[45100] = 32'b11111111111111101000011110110110;
assign LUT_2[45101] = 32'b11111111111111100101010111001111;
assign LUT_2[45102] = 32'b11111111111111101111010111110010;
assign LUT_2[45103] = 32'b11111111111111101100010000001011;
assign LUT_2[45104] = 32'b11111111111111101011110011111011;
assign LUT_2[45105] = 32'b11111111111111101000101100010100;
assign LUT_2[45106] = 32'b11111111111111110010101100110111;
assign LUT_2[45107] = 32'b11111111111111101111100101010000;
assign LUT_2[45108] = 32'b11111111111111101000010001100011;
assign LUT_2[45109] = 32'b11111111111111100101001001111100;
assign LUT_2[45110] = 32'b11111111111111101111001010011111;
assign LUT_2[45111] = 32'b11111111111111101100000010111000;
assign LUT_2[45112] = 32'b11111111111111100110100101011000;
assign LUT_2[45113] = 32'b11111111111111100011011101110001;
assign LUT_2[45114] = 32'b11111111111111101101011110010100;
assign LUT_2[45115] = 32'b11111111111111101010010110101101;
assign LUT_2[45116] = 32'b11111111111111100011000011000000;
assign LUT_2[45117] = 32'b11111111111111011111111011011001;
assign LUT_2[45118] = 32'b11111111111111101001111011111100;
assign LUT_2[45119] = 32'b11111111111111100110110100010101;
assign LUT_2[45120] = 32'b11111111111111101000111100101011;
assign LUT_2[45121] = 32'b11111111111111100101110101000100;
assign LUT_2[45122] = 32'b11111111111111101111110101100111;
assign LUT_2[45123] = 32'b11111111111111101100101110000000;
assign LUT_2[45124] = 32'b11111111111111100101011010010011;
assign LUT_2[45125] = 32'b11111111111111100010010010101100;
assign LUT_2[45126] = 32'b11111111111111101100010011001111;
assign LUT_2[45127] = 32'b11111111111111101001001011101000;
assign LUT_2[45128] = 32'b11111111111111100011101110001000;
assign LUT_2[45129] = 32'b11111111111111100000100110100001;
assign LUT_2[45130] = 32'b11111111111111101010100111000100;
assign LUT_2[45131] = 32'b11111111111111100111011111011101;
assign LUT_2[45132] = 32'b11111111111111100000001011110000;
assign LUT_2[45133] = 32'b11111111111111011101000100001001;
assign LUT_2[45134] = 32'b11111111111111100111000100101100;
assign LUT_2[45135] = 32'b11111111111111100011111101000101;
assign LUT_2[45136] = 32'b11111111111111100011100000110101;
assign LUT_2[45137] = 32'b11111111111111100000011001001110;
assign LUT_2[45138] = 32'b11111111111111101010011001110001;
assign LUT_2[45139] = 32'b11111111111111100111010010001010;
assign LUT_2[45140] = 32'b11111111111111011111111110011101;
assign LUT_2[45141] = 32'b11111111111111011100110110110110;
assign LUT_2[45142] = 32'b11111111111111100110110111011001;
assign LUT_2[45143] = 32'b11111111111111100011101111110010;
assign LUT_2[45144] = 32'b11111111111111011110010010010010;
assign LUT_2[45145] = 32'b11111111111111011011001010101011;
assign LUT_2[45146] = 32'b11111111111111100101001011001110;
assign LUT_2[45147] = 32'b11111111111111100010000011100111;
assign LUT_2[45148] = 32'b11111111111111011010101111111010;
assign LUT_2[45149] = 32'b11111111111111010111101000010011;
assign LUT_2[45150] = 32'b11111111111111100001101000110110;
assign LUT_2[45151] = 32'b11111111111111011110100001001111;
assign LUT_2[45152] = 32'b11111111111111101001011000010100;
assign LUT_2[45153] = 32'b11111111111111100110010000101101;
assign LUT_2[45154] = 32'b11111111111111110000010001010000;
assign LUT_2[45155] = 32'b11111111111111101101001001101001;
assign LUT_2[45156] = 32'b11111111111111100101110101111100;
assign LUT_2[45157] = 32'b11111111111111100010101110010101;
assign LUT_2[45158] = 32'b11111111111111101100101110111000;
assign LUT_2[45159] = 32'b11111111111111101001100111010001;
assign LUT_2[45160] = 32'b11111111111111100100001001110001;
assign LUT_2[45161] = 32'b11111111111111100001000010001010;
assign LUT_2[45162] = 32'b11111111111111101011000010101101;
assign LUT_2[45163] = 32'b11111111111111100111111011000110;
assign LUT_2[45164] = 32'b11111111111111100000100111011001;
assign LUT_2[45165] = 32'b11111111111111011101011111110010;
assign LUT_2[45166] = 32'b11111111111111100111100000010101;
assign LUT_2[45167] = 32'b11111111111111100100011000101110;
assign LUT_2[45168] = 32'b11111111111111100011111100011110;
assign LUT_2[45169] = 32'b11111111111111100000110100110111;
assign LUT_2[45170] = 32'b11111111111111101010110101011010;
assign LUT_2[45171] = 32'b11111111111111100111101101110011;
assign LUT_2[45172] = 32'b11111111111111100000011010000110;
assign LUT_2[45173] = 32'b11111111111111011101010010011111;
assign LUT_2[45174] = 32'b11111111111111100111010011000010;
assign LUT_2[45175] = 32'b11111111111111100100001011011011;
assign LUT_2[45176] = 32'b11111111111111011110101101111011;
assign LUT_2[45177] = 32'b11111111111111011011100110010100;
assign LUT_2[45178] = 32'b11111111111111100101100110110111;
assign LUT_2[45179] = 32'b11111111111111100010011111010000;
assign LUT_2[45180] = 32'b11111111111111011011001011100011;
assign LUT_2[45181] = 32'b11111111111111011000000011111100;
assign LUT_2[45182] = 32'b11111111111111100010000100011111;
assign LUT_2[45183] = 32'b11111111111111011110111100111000;
assign LUT_2[45184] = 32'b11111111111111110101001000010111;
assign LUT_2[45185] = 32'b11111111111111110010000000110000;
assign LUT_2[45186] = 32'b11111111111111111100000001010011;
assign LUT_2[45187] = 32'b11111111111111111000111001101100;
assign LUT_2[45188] = 32'b11111111111111110001100101111111;
assign LUT_2[45189] = 32'b11111111111111101110011110011000;
assign LUT_2[45190] = 32'b11111111111111111000011110111011;
assign LUT_2[45191] = 32'b11111111111111110101010111010100;
assign LUT_2[45192] = 32'b11111111111111101111111001110100;
assign LUT_2[45193] = 32'b11111111111111101100110010001101;
assign LUT_2[45194] = 32'b11111111111111110110110010110000;
assign LUT_2[45195] = 32'b11111111111111110011101011001001;
assign LUT_2[45196] = 32'b11111111111111101100010111011100;
assign LUT_2[45197] = 32'b11111111111111101001001111110101;
assign LUT_2[45198] = 32'b11111111111111110011010000011000;
assign LUT_2[45199] = 32'b11111111111111110000001000110001;
assign LUT_2[45200] = 32'b11111111111111101111101100100001;
assign LUT_2[45201] = 32'b11111111111111101100100100111010;
assign LUT_2[45202] = 32'b11111111111111110110100101011101;
assign LUT_2[45203] = 32'b11111111111111110011011101110110;
assign LUT_2[45204] = 32'b11111111111111101100001010001001;
assign LUT_2[45205] = 32'b11111111111111101001000010100010;
assign LUT_2[45206] = 32'b11111111111111110011000011000101;
assign LUT_2[45207] = 32'b11111111111111101111111011011110;
assign LUT_2[45208] = 32'b11111111111111101010011101111110;
assign LUT_2[45209] = 32'b11111111111111100111010110010111;
assign LUT_2[45210] = 32'b11111111111111110001010110111010;
assign LUT_2[45211] = 32'b11111111111111101110001111010011;
assign LUT_2[45212] = 32'b11111111111111100110111011100110;
assign LUT_2[45213] = 32'b11111111111111100011110011111111;
assign LUT_2[45214] = 32'b11111111111111101101110100100010;
assign LUT_2[45215] = 32'b11111111111111101010101100111011;
assign LUT_2[45216] = 32'b11111111111111110101100100000000;
assign LUT_2[45217] = 32'b11111111111111110010011100011001;
assign LUT_2[45218] = 32'b11111111111111111100011100111100;
assign LUT_2[45219] = 32'b11111111111111111001010101010101;
assign LUT_2[45220] = 32'b11111111111111110010000001101000;
assign LUT_2[45221] = 32'b11111111111111101110111010000001;
assign LUT_2[45222] = 32'b11111111111111111000111010100100;
assign LUT_2[45223] = 32'b11111111111111110101110010111101;
assign LUT_2[45224] = 32'b11111111111111110000010101011101;
assign LUT_2[45225] = 32'b11111111111111101101001101110110;
assign LUT_2[45226] = 32'b11111111111111110111001110011001;
assign LUT_2[45227] = 32'b11111111111111110100000110110010;
assign LUT_2[45228] = 32'b11111111111111101100110011000101;
assign LUT_2[45229] = 32'b11111111111111101001101011011110;
assign LUT_2[45230] = 32'b11111111111111110011101100000001;
assign LUT_2[45231] = 32'b11111111111111110000100100011010;
assign LUT_2[45232] = 32'b11111111111111110000001000001010;
assign LUT_2[45233] = 32'b11111111111111101101000000100011;
assign LUT_2[45234] = 32'b11111111111111110111000001000110;
assign LUT_2[45235] = 32'b11111111111111110011111001011111;
assign LUT_2[45236] = 32'b11111111111111101100100101110010;
assign LUT_2[45237] = 32'b11111111111111101001011110001011;
assign LUT_2[45238] = 32'b11111111111111110011011110101110;
assign LUT_2[45239] = 32'b11111111111111110000010111000111;
assign LUT_2[45240] = 32'b11111111111111101010111001100111;
assign LUT_2[45241] = 32'b11111111111111100111110010000000;
assign LUT_2[45242] = 32'b11111111111111110001110010100011;
assign LUT_2[45243] = 32'b11111111111111101110101010111100;
assign LUT_2[45244] = 32'b11111111111111100111010111001111;
assign LUT_2[45245] = 32'b11111111111111100100001111101000;
assign LUT_2[45246] = 32'b11111111111111101110010000001011;
assign LUT_2[45247] = 32'b11111111111111101011001000100100;
assign LUT_2[45248] = 32'b11111111111111101101010000111010;
assign LUT_2[45249] = 32'b11111111111111101010001001010011;
assign LUT_2[45250] = 32'b11111111111111110100001001110110;
assign LUT_2[45251] = 32'b11111111111111110001000010001111;
assign LUT_2[45252] = 32'b11111111111111101001101110100010;
assign LUT_2[45253] = 32'b11111111111111100110100110111011;
assign LUT_2[45254] = 32'b11111111111111110000100111011110;
assign LUT_2[45255] = 32'b11111111111111101101011111110111;
assign LUT_2[45256] = 32'b11111111111111101000000010010111;
assign LUT_2[45257] = 32'b11111111111111100100111010110000;
assign LUT_2[45258] = 32'b11111111111111101110111011010011;
assign LUT_2[45259] = 32'b11111111111111101011110011101100;
assign LUT_2[45260] = 32'b11111111111111100100011111111111;
assign LUT_2[45261] = 32'b11111111111111100001011000011000;
assign LUT_2[45262] = 32'b11111111111111101011011000111011;
assign LUT_2[45263] = 32'b11111111111111101000010001010100;
assign LUT_2[45264] = 32'b11111111111111100111110101000100;
assign LUT_2[45265] = 32'b11111111111111100100101101011101;
assign LUT_2[45266] = 32'b11111111111111101110101110000000;
assign LUT_2[45267] = 32'b11111111111111101011100110011001;
assign LUT_2[45268] = 32'b11111111111111100100010010101100;
assign LUT_2[45269] = 32'b11111111111111100001001011000101;
assign LUT_2[45270] = 32'b11111111111111101011001011101000;
assign LUT_2[45271] = 32'b11111111111111101000000100000001;
assign LUT_2[45272] = 32'b11111111111111100010100110100001;
assign LUT_2[45273] = 32'b11111111111111011111011110111010;
assign LUT_2[45274] = 32'b11111111111111101001011111011101;
assign LUT_2[45275] = 32'b11111111111111100110010111110110;
assign LUT_2[45276] = 32'b11111111111111011111000100001001;
assign LUT_2[45277] = 32'b11111111111111011011111100100010;
assign LUT_2[45278] = 32'b11111111111111100101111101000101;
assign LUT_2[45279] = 32'b11111111111111100010110101011110;
assign LUT_2[45280] = 32'b11111111111111101101101100100011;
assign LUT_2[45281] = 32'b11111111111111101010100100111100;
assign LUT_2[45282] = 32'b11111111111111110100100101011111;
assign LUT_2[45283] = 32'b11111111111111110001011101111000;
assign LUT_2[45284] = 32'b11111111111111101010001010001011;
assign LUT_2[45285] = 32'b11111111111111100111000010100100;
assign LUT_2[45286] = 32'b11111111111111110001000011000111;
assign LUT_2[45287] = 32'b11111111111111101101111011100000;
assign LUT_2[45288] = 32'b11111111111111101000011110000000;
assign LUT_2[45289] = 32'b11111111111111100101010110011001;
assign LUT_2[45290] = 32'b11111111111111101111010110111100;
assign LUT_2[45291] = 32'b11111111111111101100001111010101;
assign LUT_2[45292] = 32'b11111111111111100100111011101000;
assign LUT_2[45293] = 32'b11111111111111100001110100000001;
assign LUT_2[45294] = 32'b11111111111111101011110100100100;
assign LUT_2[45295] = 32'b11111111111111101000101100111101;
assign LUT_2[45296] = 32'b11111111111111101000010000101101;
assign LUT_2[45297] = 32'b11111111111111100101001001000110;
assign LUT_2[45298] = 32'b11111111111111101111001001101001;
assign LUT_2[45299] = 32'b11111111111111101100000010000010;
assign LUT_2[45300] = 32'b11111111111111100100101110010101;
assign LUT_2[45301] = 32'b11111111111111100001100110101110;
assign LUT_2[45302] = 32'b11111111111111101011100111010001;
assign LUT_2[45303] = 32'b11111111111111101000011111101010;
assign LUT_2[45304] = 32'b11111111111111100011000010001010;
assign LUT_2[45305] = 32'b11111111111111011111111010100011;
assign LUT_2[45306] = 32'b11111111111111101001111011000110;
assign LUT_2[45307] = 32'b11111111111111100110110011011111;
assign LUT_2[45308] = 32'b11111111111111011111011111110010;
assign LUT_2[45309] = 32'b11111111111111011100011000001011;
assign LUT_2[45310] = 32'b11111111111111100110011000101110;
assign LUT_2[45311] = 32'b11111111111111100011010001000111;
assign LUT_2[45312] = 32'b11111111111111110100110010101110;
assign LUT_2[45313] = 32'b11111111111111110001101011000111;
assign LUT_2[45314] = 32'b11111111111111111011101011101010;
assign LUT_2[45315] = 32'b11111111111111111000100100000011;
assign LUT_2[45316] = 32'b11111111111111110001010000010110;
assign LUT_2[45317] = 32'b11111111111111101110001000101111;
assign LUT_2[45318] = 32'b11111111111111111000001001010010;
assign LUT_2[45319] = 32'b11111111111111110101000001101011;
assign LUT_2[45320] = 32'b11111111111111101111100100001011;
assign LUT_2[45321] = 32'b11111111111111101100011100100100;
assign LUT_2[45322] = 32'b11111111111111110110011101000111;
assign LUT_2[45323] = 32'b11111111111111110011010101100000;
assign LUT_2[45324] = 32'b11111111111111101100000001110011;
assign LUT_2[45325] = 32'b11111111111111101000111010001100;
assign LUT_2[45326] = 32'b11111111111111110010111010101111;
assign LUT_2[45327] = 32'b11111111111111101111110011001000;
assign LUT_2[45328] = 32'b11111111111111101111010110111000;
assign LUT_2[45329] = 32'b11111111111111101100001111010001;
assign LUT_2[45330] = 32'b11111111111111110110001111110100;
assign LUT_2[45331] = 32'b11111111111111110011001000001101;
assign LUT_2[45332] = 32'b11111111111111101011110100100000;
assign LUT_2[45333] = 32'b11111111111111101000101100111001;
assign LUT_2[45334] = 32'b11111111111111110010101101011100;
assign LUT_2[45335] = 32'b11111111111111101111100101110101;
assign LUT_2[45336] = 32'b11111111111111101010001000010101;
assign LUT_2[45337] = 32'b11111111111111100111000000101110;
assign LUT_2[45338] = 32'b11111111111111110001000001010001;
assign LUT_2[45339] = 32'b11111111111111101101111001101010;
assign LUT_2[45340] = 32'b11111111111111100110100101111101;
assign LUT_2[45341] = 32'b11111111111111100011011110010110;
assign LUT_2[45342] = 32'b11111111111111101101011110111001;
assign LUT_2[45343] = 32'b11111111111111101010010111010010;
assign LUT_2[45344] = 32'b11111111111111110101001110010111;
assign LUT_2[45345] = 32'b11111111111111110010000110110000;
assign LUT_2[45346] = 32'b11111111111111111100000111010011;
assign LUT_2[45347] = 32'b11111111111111111000111111101100;
assign LUT_2[45348] = 32'b11111111111111110001101011111111;
assign LUT_2[45349] = 32'b11111111111111101110100100011000;
assign LUT_2[45350] = 32'b11111111111111111000100100111011;
assign LUT_2[45351] = 32'b11111111111111110101011101010100;
assign LUT_2[45352] = 32'b11111111111111101111111111110100;
assign LUT_2[45353] = 32'b11111111111111101100111000001101;
assign LUT_2[45354] = 32'b11111111111111110110111000110000;
assign LUT_2[45355] = 32'b11111111111111110011110001001001;
assign LUT_2[45356] = 32'b11111111111111101100011101011100;
assign LUT_2[45357] = 32'b11111111111111101001010101110101;
assign LUT_2[45358] = 32'b11111111111111110011010110011000;
assign LUT_2[45359] = 32'b11111111111111110000001110110001;
assign LUT_2[45360] = 32'b11111111111111101111110010100001;
assign LUT_2[45361] = 32'b11111111111111101100101010111010;
assign LUT_2[45362] = 32'b11111111111111110110101011011101;
assign LUT_2[45363] = 32'b11111111111111110011100011110110;
assign LUT_2[45364] = 32'b11111111111111101100010000001001;
assign LUT_2[45365] = 32'b11111111111111101001001000100010;
assign LUT_2[45366] = 32'b11111111111111110011001001000101;
assign LUT_2[45367] = 32'b11111111111111110000000001011110;
assign LUT_2[45368] = 32'b11111111111111101010100011111110;
assign LUT_2[45369] = 32'b11111111111111100111011100010111;
assign LUT_2[45370] = 32'b11111111111111110001011100111010;
assign LUT_2[45371] = 32'b11111111111111101110010101010011;
assign LUT_2[45372] = 32'b11111111111111100111000001100110;
assign LUT_2[45373] = 32'b11111111111111100011111001111111;
assign LUT_2[45374] = 32'b11111111111111101101111010100010;
assign LUT_2[45375] = 32'b11111111111111101010110010111011;
assign LUT_2[45376] = 32'b11111111111111101100111011010001;
assign LUT_2[45377] = 32'b11111111111111101001110011101010;
assign LUT_2[45378] = 32'b11111111111111110011110100001101;
assign LUT_2[45379] = 32'b11111111111111110000101100100110;
assign LUT_2[45380] = 32'b11111111111111101001011000111001;
assign LUT_2[45381] = 32'b11111111111111100110010001010010;
assign LUT_2[45382] = 32'b11111111111111110000010001110101;
assign LUT_2[45383] = 32'b11111111111111101101001010001110;
assign LUT_2[45384] = 32'b11111111111111100111101100101110;
assign LUT_2[45385] = 32'b11111111111111100100100101000111;
assign LUT_2[45386] = 32'b11111111111111101110100101101010;
assign LUT_2[45387] = 32'b11111111111111101011011110000011;
assign LUT_2[45388] = 32'b11111111111111100100001010010110;
assign LUT_2[45389] = 32'b11111111111111100001000010101111;
assign LUT_2[45390] = 32'b11111111111111101011000011010010;
assign LUT_2[45391] = 32'b11111111111111100111111011101011;
assign LUT_2[45392] = 32'b11111111111111100111011111011011;
assign LUT_2[45393] = 32'b11111111111111100100010111110100;
assign LUT_2[45394] = 32'b11111111111111101110011000010111;
assign LUT_2[45395] = 32'b11111111111111101011010000110000;
assign LUT_2[45396] = 32'b11111111111111100011111101000011;
assign LUT_2[45397] = 32'b11111111111111100000110101011100;
assign LUT_2[45398] = 32'b11111111111111101010110101111111;
assign LUT_2[45399] = 32'b11111111111111100111101110011000;
assign LUT_2[45400] = 32'b11111111111111100010010000111000;
assign LUT_2[45401] = 32'b11111111111111011111001001010001;
assign LUT_2[45402] = 32'b11111111111111101001001001110100;
assign LUT_2[45403] = 32'b11111111111111100110000010001101;
assign LUT_2[45404] = 32'b11111111111111011110101110100000;
assign LUT_2[45405] = 32'b11111111111111011011100110111001;
assign LUT_2[45406] = 32'b11111111111111100101100111011100;
assign LUT_2[45407] = 32'b11111111111111100010011111110101;
assign LUT_2[45408] = 32'b11111111111111101101010110111010;
assign LUT_2[45409] = 32'b11111111111111101010001111010011;
assign LUT_2[45410] = 32'b11111111111111110100001111110110;
assign LUT_2[45411] = 32'b11111111111111110001001000001111;
assign LUT_2[45412] = 32'b11111111111111101001110100100010;
assign LUT_2[45413] = 32'b11111111111111100110101100111011;
assign LUT_2[45414] = 32'b11111111111111110000101101011110;
assign LUT_2[45415] = 32'b11111111111111101101100101110111;
assign LUT_2[45416] = 32'b11111111111111101000001000010111;
assign LUT_2[45417] = 32'b11111111111111100101000000110000;
assign LUT_2[45418] = 32'b11111111111111101111000001010011;
assign LUT_2[45419] = 32'b11111111111111101011111001101100;
assign LUT_2[45420] = 32'b11111111111111100100100101111111;
assign LUT_2[45421] = 32'b11111111111111100001011110011000;
assign LUT_2[45422] = 32'b11111111111111101011011110111011;
assign LUT_2[45423] = 32'b11111111111111101000010111010100;
assign LUT_2[45424] = 32'b11111111111111100111111011000100;
assign LUT_2[45425] = 32'b11111111111111100100110011011101;
assign LUT_2[45426] = 32'b11111111111111101110110100000000;
assign LUT_2[45427] = 32'b11111111111111101011101100011001;
assign LUT_2[45428] = 32'b11111111111111100100011000101100;
assign LUT_2[45429] = 32'b11111111111111100001010001000101;
assign LUT_2[45430] = 32'b11111111111111101011010001101000;
assign LUT_2[45431] = 32'b11111111111111101000001010000001;
assign LUT_2[45432] = 32'b11111111111111100010101100100001;
assign LUT_2[45433] = 32'b11111111111111011111100100111010;
assign LUT_2[45434] = 32'b11111111111111101001100101011101;
assign LUT_2[45435] = 32'b11111111111111100110011101110110;
assign LUT_2[45436] = 32'b11111111111111011111001010001001;
assign LUT_2[45437] = 32'b11111111111111011100000010100010;
assign LUT_2[45438] = 32'b11111111111111100110000011000101;
assign LUT_2[45439] = 32'b11111111111111100010111011011110;
assign LUT_2[45440] = 32'b11111111111111111001000110111101;
assign LUT_2[45441] = 32'b11111111111111110101111111010110;
assign LUT_2[45442] = 32'b11111111111111111111111111111001;
assign LUT_2[45443] = 32'b11111111111111111100111000010010;
assign LUT_2[45444] = 32'b11111111111111110101100100100101;
assign LUT_2[45445] = 32'b11111111111111110010011100111110;
assign LUT_2[45446] = 32'b11111111111111111100011101100001;
assign LUT_2[45447] = 32'b11111111111111111001010101111010;
assign LUT_2[45448] = 32'b11111111111111110011111000011010;
assign LUT_2[45449] = 32'b11111111111111110000110000110011;
assign LUT_2[45450] = 32'b11111111111111111010110001010110;
assign LUT_2[45451] = 32'b11111111111111110111101001101111;
assign LUT_2[45452] = 32'b11111111111111110000010110000010;
assign LUT_2[45453] = 32'b11111111111111101101001110011011;
assign LUT_2[45454] = 32'b11111111111111110111001110111110;
assign LUT_2[45455] = 32'b11111111111111110100000111010111;
assign LUT_2[45456] = 32'b11111111111111110011101011000111;
assign LUT_2[45457] = 32'b11111111111111110000100011100000;
assign LUT_2[45458] = 32'b11111111111111111010100100000011;
assign LUT_2[45459] = 32'b11111111111111110111011100011100;
assign LUT_2[45460] = 32'b11111111111111110000001000101111;
assign LUT_2[45461] = 32'b11111111111111101101000001001000;
assign LUT_2[45462] = 32'b11111111111111110111000001101011;
assign LUT_2[45463] = 32'b11111111111111110011111010000100;
assign LUT_2[45464] = 32'b11111111111111101110011100100100;
assign LUT_2[45465] = 32'b11111111111111101011010100111101;
assign LUT_2[45466] = 32'b11111111111111110101010101100000;
assign LUT_2[45467] = 32'b11111111111111110010001101111001;
assign LUT_2[45468] = 32'b11111111111111101010111010001100;
assign LUT_2[45469] = 32'b11111111111111100111110010100101;
assign LUT_2[45470] = 32'b11111111111111110001110011001000;
assign LUT_2[45471] = 32'b11111111111111101110101011100001;
assign LUT_2[45472] = 32'b11111111111111111001100010100110;
assign LUT_2[45473] = 32'b11111111111111110110011010111111;
assign LUT_2[45474] = 32'b00000000000000000000011011100010;
assign LUT_2[45475] = 32'b11111111111111111101010011111011;
assign LUT_2[45476] = 32'b11111111111111110110000000001110;
assign LUT_2[45477] = 32'b11111111111111110010111000100111;
assign LUT_2[45478] = 32'b11111111111111111100111001001010;
assign LUT_2[45479] = 32'b11111111111111111001110001100011;
assign LUT_2[45480] = 32'b11111111111111110100010100000011;
assign LUT_2[45481] = 32'b11111111111111110001001100011100;
assign LUT_2[45482] = 32'b11111111111111111011001100111111;
assign LUT_2[45483] = 32'b11111111111111111000000101011000;
assign LUT_2[45484] = 32'b11111111111111110000110001101011;
assign LUT_2[45485] = 32'b11111111111111101101101010000100;
assign LUT_2[45486] = 32'b11111111111111110111101010100111;
assign LUT_2[45487] = 32'b11111111111111110100100011000000;
assign LUT_2[45488] = 32'b11111111111111110100000110110000;
assign LUT_2[45489] = 32'b11111111111111110000111111001001;
assign LUT_2[45490] = 32'b11111111111111111010111111101100;
assign LUT_2[45491] = 32'b11111111111111110111111000000101;
assign LUT_2[45492] = 32'b11111111111111110000100100011000;
assign LUT_2[45493] = 32'b11111111111111101101011100110001;
assign LUT_2[45494] = 32'b11111111111111110111011101010100;
assign LUT_2[45495] = 32'b11111111111111110100010101101101;
assign LUT_2[45496] = 32'b11111111111111101110111000001101;
assign LUT_2[45497] = 32'b11111111111111101011110000100110;
assign LUT_2[45498] = 32'b11111111111111110101110001001001;
assign LUT_2[45499] = 32'b11111111111111110010101001100010;
assign LUT_2[45500] = 32'b11111111111111101011010101110101;
assign LUT_2[45501] = 32'b11111111111111101000001110001110;
assign LUT_2[45502] = 32'b11111111111111110010001110110001;
assign LUT_2[45503] = 32'b11111111111111101111000111001010;
assign LUT_2[45504] = 32'b11111111111111110001001111100000;
assign LUT_2[45505] = 32'b11111111111111101110000111111001;
assign LUT_2[45506] = 32'b11111111111111111000001000011100;
assign LUT_2[45507] = 32'b11111111111111110101000000110101;
assign LUT_2[45508] = 32'b11111111111111101101101101001000;
assign LUT_2[45509] = 32'b11111111111111101010100101100001;
assign LUT_2[45510] = 32'b11111111111111110100100110000100;
assign LUT_2[45511] = 32'b11111111111111110001011110011101;
assign LUT_2[45512] = 32'b11111111111111101100000000111101;
assign LUT_2[45513] = 32'b11111111111111101000111001010110;
assign LUT_2[45514] = 32'b11111111111111110010111001111001;
assign LUT_2[45515] = 32'b11111111111111101111110010010010;
assign LUT_2[45516] = 32'b11111111111111101000011110100101;
assign LUT_2[45517] = 32'b11111111111111100101010110111110;
assign LUT_2[45518] = 32'b11111111111111101111010111100001;
assign LUT_2[45519] = 32'b11111111111111101100001111111010;
assign LUT_2[45520] = 32'b11111111111111101011110011101010;
assign LUT_2[45521] = 32'b11111111111111101000101100000011;
assign LUT_2[45522] = 32'b11111111111111110010101100100110;
assign LUT_2[45523] = 32'b11111111111111101111100100111111;
assign LUT_2[45524] = 32'b11111111111111101000010001010010;
assign LUT_2[45525] = 32'b11111111111111100101001001101011;
assign LUT_2[45526] = 32'b11111111111111101111001010001110;
assign LUT_2[45527] = 32'b11111111111111101100000010100111;
assign LUT_2[45528] = 32'b11111111111111100110100101000111;
assign LUT_2[45529] = 32'b11111111111111100011011101100000;
assign LUT_2[45530] = 32'b11111111111111101101011110000011;
assign LUT_2[45531] = 32'b11111111111111101010010110011100;
assign LUT_2[45532] = 32'b11111111111111100011000010101111;
assign LUT_2[45533] = 32'b11111111111111011111111011001000;
assign LUT_2[45534] = 32'b11111111111111101001111011101011;
assign LUT_2[45535] = 32'b11111111111111100110110100000100;
assign LUT_2[45536] = 32'b11111111111111110001101011001001;
assign LUT_2[45537] = 32'b11111111111111101110100011100010;
assign LUT_2[45538] = 32'b11111111111111111000100100000101;
assign LUT_2[45539] = 32'b11111111111111110101011100011110;
assign LUT_2[45540] = 32'b11111111111111101110001000110001;
assign LUT_2[45541] = 32'b11111111111111101011000001001010;
assign LUT_2[45542] = 32'b11111111111111110101000001101101;
assign LUT_2[45543] = 32'b11111111111111110001111010000110;
assign LUT_2[45544] = 32'b11111111111111101100011100100110;
assign LUT_2[45545] = 32'b11111111111111101001010100111111;
assign LUT_2[45546] = 32'b11111111111111110011010101100010;
assign LUT_2[45547] = 32'b11111111111111110000001101111011;
assign LUT_2[45548] = 32'b11111111111111101000111010001110;
assign LUT_2[45549] = 32'b11111111111111100101110010100111;
assign LUT_2[45550] = 32'b11111111111111101111110011001010;
assign LUT_2[45551] = 32'b11111111111111101100101011100011;
assign LUT_2[45552] = 32'b11111111111111101100001111010011;
assign LUT_2[45553] = 32'b11111111111111101001000111101100;
assign LUT_2[45554] = 32'b11111111111111110011001000001111;
assign LUT_2[45555] = 32'b11111111111111110000000000101000;
assign LUT_2[45556] = 32'b11111111111111101000101100111011;
assign LUT_2[45557] = 32'b11111111111111100101100101010100;
assign LUT_2[45558] = 32'b11111111111111101111100101110111;
assign LUT_2[45559] = 32'b11111111111111101100011110010000;
assign LUT_2[45560] = 32'b11111111111111100111000000110000;
assign LUT_2[45561] = 32'b11111111111111100011111001001001;
assign LUT_2[45562] = 32'b11111111111111101101111001101100;
assign LUT_2[45563] = 32'b11111111111111101010110010000101;
assign LUT_2[45564] = 32'b11111111111111100011011110011000;
assign LUT_2[45565] = 32'b11111111111111100000010110110001;
assign LUT_2[45566] = 32'b11111111111111101010010111010100;
assign LUT_2[45567] = 32'b11111111111111100111001111101101;
assign LUT_2[45568] = 32'b11111111111111110101100101111010;
assign LUT_2[45569] = 32'b11111111111111110010011110010011;
assign LUT_2[45570] = 32'b11111111111111111100011110110110;
assign LUT_2[45571] = 32'b11111111111111111001010111001111;
assign LUT_2[45572] = 32'b11111111111111110010000011100010;
assign LUT_2[45573] = 32'b11111111111111101110111011111011;
assign LUT_2[45574] = 32'b11111111111111111000111100011110;
assign LUT_2[45575] = 32'b11111111111111110101110100110111;
assign LUT_2[45576] = 32'b11111111111111110000010111010111;
assign LUT_2[45577] = 32'b11111111111111101101001111110000;
assign LUT_2[45578] = 32'b11111111111111110111010000010011;
assign LUT_2[45579] = 32'b11111111111111110100001000101100;
assign LUT_2[45580] = 32'b11111111111111101100110100111111;
assign LUT_2[45581] = 32'b11111111111111101001101101011000;
assign LUT_2[45582] = 32'b11111111111111110011101101111011;
assign LUT_2[45583] = 32'b11111111111111110000100110010100;
assign LUT_2[45584] = 32'b11111111111111110000001010000100;
assign LUT_2[45585] = 32'b11111111111111101101000010011101;
assign LUT_2[45586] = 32'b11111111111111110111000011000000;
assign LUT_2[45587] = 32'b11111111111111110011111011011001;
assign LUT_2[45588] = 32'b11111111111111101100100111101100;
assign LUT_2[45589] = 32'b11111111111111101001100000000101;
assign LUT_2[45590] = 32'b11111111111111110011100000101000;
assign LUT_2[45591] = 32'b11111111111111110000011001000001;
assign LUT_2[45592] = 32'b11111111111111101010111011100001;
assign LUT_2[45593] = 32'b11111111111111100111110011111010;
assign LUT_2[45594] = 32'b11111111111111110001110100011101;
assign LUT_2[45595] = 32'b11111111111111101110101100110110;
assign LUT_2[45596] = 32'b11111111111111100111011001001001;
assign LUT_2[45597] = 32'b11111111111111100100010001100010;
assign LUT_2[45598] = 32'b11111111111111101110010010000101;
assign LUT_2[45599] = 32'b11111111111111101011001010011110;
assign LUT_2[45600] = 32'b11111111111111110110000001100011;
assign LUT_2[45601] = 32'b11111111111111110010111001111100;
assign LUT_2[45602] = 32'b11111111111111111100111010011111;
assign LUT_2[45603] = 32'b11111111111111111001110010111000;
assign LUT_2[45604] = 32'b11111111111111110010011111001011;
assign LUT_2[45605] = 32'b11111111111111101111010111100100;
assign LUT_2[45606] = 32'b11111111111111111001011000000111;
assign LUT_2[45607] = 32'b11111111111111110110010000100000;
assign LUT_2[45608] = 32'b11111111111111110000110011000000;
assign LUT_2[45609] = 32'b11111111111111101101101011011001;
assign LUT_2[45610] = 32'b11111111111111110111101011111100;
assign LUT_2[45611] = 32'b11111111111111110100100100010101;
assign LUT_2[45612] = 32'b11111111111111101101010000101000;
assign LUT_2[45613] = 32'b11111111111111101010001001000001;
assign LUT_2[45614] = 32'b11111111111111110100001001100100;
assign LUT_2[45615] = 32'b11111111111111110001000001111101;
assign LUT_2[45616] = 32'b11111111111111110000100101101101;
assign LUT_2[45617] = 32'b11111111111111101101011110000110;
assign LUT_2[45618] = 32'b11111111111111110111011110101001;
assign LUT_2[45619] = 32'b11111111111111110100010111000010;
assign LUT_2[45620] = 32'b11111111111111101101000011010101;
assign LUT_2[45621] = 32'b11111111111111101001111011101110;
assign LUT_2[45622] = 32'b11111111111111110011111100010001;
assign LUT_2[45623] = 32'b11111111111111110000110100101010;
assign LUT_2[45624] = 32'b11111111111111101011010111001010;
assign LUT_2[45625] = 32'b11111111111111101000001111100011;
assign LUT_2[45626] = 32'b11111111111111110010010000000110;
assign LUT_2[45627] = 32'b11111111111111101111001000011111;
assign LUT_2[45628] = 32'b11111111111111100111110100110010;
assign LUT_2[45629] = 32'b11111111111111100100101101001011;
assign LUT_2[45630] = 32'b11111111111111101110101101101110;
assign LUT_2[45631] = 32'b11111111111111101011100110000111;
assign LUT_2[45632] = 32'b11111111111111101101101110011101;
assign LUT_2[45633] = 32'b11111111111111101010100110110110;
assign LUT_2[45634] = 32'b11111111111111110100100111011001;
assign LUT_2[45635] = 32'b11111111111111110001011111110010;
assign LUT_2[45636] = 32'b11111111111111101010001100000101;
assign LUT_2[45637] = 32'b11111111111111100111000100011110;
assign LUT_2[45638] = 32'b11111111111111110001000101000001;
assign LUT_2[45639] = 32'b11111111111111101101111101011010;
assign LUT_2[45640] = 32'b11111111111111101000011111111010;
assign LUT_2[45641] = 32'b11111111111111100101011000010011;
assign LUT_2[45642] = 32'b11111111111111101111011000110110;
assign LUT_2[45643] = 32'b11111111111111101100010001001111;
assign LUT_2[45644] = 32'b11111111111111100100111101100010;
assign LUT_2[45645] = 32'b11111111111111100001110101111011;
assign LUT_2[45646] = 32'b11111111111111101011110110011110;
assign LUT_2[45647] = 32'b11111111111111101000101110110111;
assign LUT_2[45648] = 32'b11111111111111101000010010100111;
assign LUT_2[45649] = 32'b11111111111111100101001011000000;
assign LUT_2[45650] = 32'b11111111111111101111001011100011;
assign LUT_2[45651] = 32'b11111111111111101100000011111100;
assign LUT_2[45652] = 32'b11111111111111100100110000001111;
assign LUT_2[45653] = 32'b11111111111111100001101000101000;
assign LUT_2[45654] = 32'b11111111111111101011101001001011;
assign LUT_2[45655] = 32'b11111111111111101000100001100100;
assign LUT_2[45656] = 32'b11111111111111100011000100000100;
assign LUT_2[45657] = 32'b11111111111111011111111100011101;
assign LUT_2[45658] = 32'b11111111111111101001111101000000;
assign LUT_2[45659] = 32'b11111111111111100110110101011001;
assign LUT_2[45660] = 32'b11111111111111011111100001101100;
assign LUT_2[45661] = 32'b11111111111111011100011010000101;
assign LUT_2[45662] = 32'b11111111111111100110011010101000;
assign LUT_2[45663] = 32'b11111111111111100011010011000001;
assign LUT_2[45664] = 32'b11111111111111101110001010000110;
assign LUT_2[45665] = 32'b11111111111111101011000010011111;
assign LUT_2[45666] = 32'b11111111111111110101000011000010;
assign LUT_2[45667] = 32'b11111111111111110001111011011011;
assign LUT_2[45668] = 32'b11111111111111101010100111101110;
assign LUT_2[45669] = 32'b11111111111111100111100000000111;
assign LUT_2[45670] = 32'b11111111111111110001100000101010;
assign LUT_2[45671] = 32'b11111111111111101110011001000011;
assign LUT_2[45672] = 32'b11111111111111101000111011100011;
assign LUT_2[45673] = 32'b11111111111111100101110011111100;
assign LUT_2[45674] = 32'b11111111111111101111110100011111;
assign LUT_2[45675] = 32'b11111111111111101100101100111000;
assign LUT_2[45676] = 32'b11111111111111100101011001001011;
assign LUT_2[45677] = 32'b11111111111111100010010001100100;
assign LUT_2[45678] = 32'b11111111111111101100010010000111;
assign LUT_2[45679] = 32'b11111111111111101001001010100000;
assign LUT_2[45680] = 32'b11111111111111101000101110010000;
assign LUT_2[45681] = 32'b11111111111111100101100110101001;
assign LUT_2[45682] = 32'b11111111111111101111100111001100;
assign LUT_2[45683] = 32'b11111111111111101100011111100101;
assign LUT_2[45684] = 32'b11111111111111100101001011111000;
assign LUT_2[45685] = 32'b11111111111111100010000100010001;
assign LUT_2[45686] = 32'b11111111111111101100000100110100;
assign LUT_2[45687] = 32'b11111111111111101000111101001101;
assign LUT_2[45688] = 32'b11111111111111100011011111101101;
assign LUT_2[45689] = 32'b11111111111111100000011000000110;
assign LUT_2[45690] = 32'b11111111111111101010011000101001;
assign LUT_2[45691] = 32'b11111111111111100111010001000010;
assign LUT_2[45692] = 32'b11111111111111011111111101010101;
assign LUT_2[45693] = 32'b11111111111111011100110101101110;
assign LUT_2[45694] = 32'b11111111111111100110110110010001;
assign LUT_2[45695] = 32'b11111111111111100011101110101010;
assign LUT_2[45696] = 32'b11111111111111111001111010001001;
assign LUT_2[45697] = 32'b11111111111111110110110010100010;
assign LUT_2[45698] = 32'b00000000000000000000110011000101;
assign LUT_2[45699] = 32'b11111111111111111101101011011110;
assign LUT_2[45700] = 32'b11111111111111110110010111110001;
assign LUT_2[45701] = 32'b11111111111111110011010000001010;
assign LUT_2[45702] = 32'b11111111111111111101010000101101;
assign LUT_2[45703] = 32'b11111111111111111010001001000110;
assign LUT_2[45704] = 32'b11111111111111110100101011100110;
assign LUT_2[45705] = 32'b11111111111111110001100011111111;
assign LUT_2[45706] = 32'b11111111111111111011100100100010;
assign LUT_2[45707] = 32'b11111111111111111000011100111011;
assign LUT_2[45708] = 32'b11111111111111110001001001001110;
assign LUT_2[45709] = 32'b11111111111111101110000001100111;
assign LUT_2[45710] = 32'b11111111111111111000000010001010;
assign LUT_2[45711] = 32'b11111111111111110100111010100011;
assign LUT_2[45712] = 32'b11111111111111110100011110010011;
assign LUT_2[45713] = 32'b11111111111111110001010110101100;
assign LUT_2[45714] = 32'b11111111111111111011010111001111;
assign LUT_2[45715] = 32'b11111111111111111000001111101000;
assign LUT_2[45716] = 32'b11111111111111110000111011111011;
assign LUT_2[45717] = 32'b11111111111111101101110100010100;
assign LUT_2[45718] = 32'b11111111111111110111110100110111;
assign LUT_2[45719] = 32'b11111111111111110100101101010000;
assign LUT_2[45720] = 32'b11111111111111101111001111110000;
assign LUT_2[45721] = 32'b11111111111111101100001000001001;
assign LUT_2[45722] = 32'b11111111111111110110001000101100;
assign LUT_2[45723] = 32'b11111111111111110011000001000101;
assign LUT_2[45724] = 32'b11111111111111101011101101011000;
assign LUT_2[45725] = 32'b11111111111111101000100101110001;
assign LUT_2[45726] = 32'b11111111111111110010100110010100;
assign LUT_2[45727] = 32'b11111111111111101111011110101101;
assign LUT_2[45728] = 32'b11111111111111111010010101110010;
assign LUT_2[45729] = 32'b11111111111111110111001110001011;
assign LUT_2[45730] = 32'b00000000000000000001001110101110;
assign LUT_2[45731] = 32'b11111111111111111110000111000111;
assign LUT_2[45732] = 32'b11111111111111110110110011011010;
assign LUT_2[45733] = 32'b11111111111111110011101011110011;
assign LUT_2[45734] = 32'b11111111111111111101101100010110;
assign LUT_2[45735] = 32'b11111111111111111010100100101111;
assign LUT_2[45736] = 32'b11111111111111110101000111001111;
assign LUT_2[45737] = 32'b11111111111111110001111111101000;
assign LUT_2[45738] = 32'b11111111111111111100000000001011;
assign LUT_2[45739] = 32'b11111111111111111000111000100100;
assign LUT_2[45740] = 32'b11111111111111110001100100110111;
assign LUT_2[45741] = 32'b11111111111111101110011101010000;
assign LUT_2[45742] = 32'b11111111111111111000011101110011;
assign LUT_2[45743] = 32'b11111111111111110101010110001100;
assign LUT_2[45744] = 32'b11111111111111110100111001111100;
assign LUT_2[45745] = 32'b11111111111111110001110010010101;
assign LUT_2[45746] = 32'b11111111111111111011110010111000;
assign LUT_2[45747] = 32'b11111111111111111000101011010001;
assign LUT_2[45748] = 32'b11111111111111110001010111100100;
assign LUT_2[45749] = 32'b11111111111111101110001111111101;
assign LUT_2[45750] = 32'b11111111111111111000010000100000;
assign LUT_2[45751] = 32'b11111111111111110101001000111001;
assign LUT_2[45752] = 32'b11111111111111101111101011011001;
assign LUT_2[45753] = 32'b11111111111111101100100011110010;
assign LUT_2[45754] = 32'b11111111111111110110100100010101;
assign LUT_2[45755] = 32'b11111111111111110011011100101110;
assign LUT_2[45756] = 32'b11111111111111101100001001000001;
assign LUT_2[45757] = 32'b11111111111111101001000001011010;
assign LUT_2[45758] = 32'b11111111111111110011000001111101;
assign LUT_2[45759] = 32'b11111111111111101111111010010110;
assign LUT_2[45760] = 32'b11111111111111110010000010101100;
assign LUT_2[45761] = 32'b11111111111111101110111011000101;
assign LUT_2[45762] = 32'b11111111111111111000111011101000;
assign LUT_2[45763] = 32'b11111111111111110101110100000001;
assign LUT_2[45764] = 32'b11111111111111101110100000010100;
assign LUT_2[45765] = 32'b11111111111111101011011000101101;
assign LUT_2[45766] = 32'b11111111111111110101011001010000;
assign LUT_2[45767] = 32'b11111111111111110010010001101001;
assign LUT_2[45768] = 32'b11111111111111101100110100001001;
assign LUT_2[45769] = 32'b11111111111111101001101100100010;
assign LUT_2[45770] = 32'b11111111111111110011101101000101;
assign LUT_2[45771] = 32'b11111111111111110000100101011110;
assign LUT_2[45772] = 32'b11111111111111101001010001110001;
assign LUT_2[45773] = 32'b11111111111111100110001010001010;
assign LUT_2[45774] = 32'b11111111111111110000001010101101;
assign LUT_2[45775] = 32'b11111111111111101101000011000110;
assign LUT_2[45776] = 32'b11111111111111101100100110110110;
assign LUT_2[45777] = 32'b11111111111111101001011111001111;
assign LUT_2[45778] = 32'b11111111111111110011011111110010;
assign LUT_2[45779] = 32'b11111111111111110000011000001011;
assign LUT_2[45780] = 32'b11111111111111101001000100011110;
assign LUT_2[45781] = 32'b11111111111111100101111100110111;
assign LUT_2[45782] = 32'b11111111111111101111111101011010;
assign LUT_2[45783] = 32'b11111111111111101100110101110011;
assign LUT_2[45784] = 32'b11111111111111100111011000010011;
assign LUT_2[45785] = 32'b11111111111111100100010000101100;
assign LUT_2[45786] = 32'b11111111111111101110010001001111;
assign LUT_2[45787] = 32'b11111111111111101011001001101000;
assign LUT_2[45788] = 32'b11111111111111100011110101111011;
assign LUT_2[45789] = 32'b11111111111111100000101110010100;
assign LUT_2[45790] = 32'b11111111111111101010101110110111;
assign LUT_2[45791] = 32'b11111111111111100111100111010000;
assign LUT_2[45792] = 32'b11111111111111110010011110010101;
assign LUT_2[45793] = 32'b11111111111111101111010110101110;
assign LUT_2[45794] = 32'b11111111111111111001010111010001;
assign LUT_2[45795] = 32'b11111111111111110110001111101010;
assign LUT_2[45796] = 32'b11111111111111101110111011111101;
assign LUT_2[45797] = 32'b11111111111111101011110100010110;
assign LUT_2[45798] = 32'b11111111111111110101110100111001;
assign LUT_2[45799] = 32'b11111111111111110010101101010010;
assign LUT_2[45800] = 32'b11111111111111101101001111110010;
assign LUT_2[45801] = 32'b11111111111111101010001000001011;
assign LUT_2[45802] = 32'b11111111111111110100001000101110;
assign LUT_2[45803] = 32'b11111111111111110001000001000111;
assign LUT_2[45804] = 32'b11111111111111101001101101011010;
assign LUT_2[45805] = 32'b11111111111111100110100101110011;
assign LUT_2[45806] = 32'b11111111111111110000100110010110;
assign LUT_2[45807] = 32'b11111111111111101101011110101111;
assign LUT_2[45808] = 32'b11111111111111101101000010011111;
assign LUT_2[45809] = 32'b11111111111111101001111010111000;
assign LUT_2[45810] = 32'b11111111111111110011111011011011;
assign LUT_2[45811] = 32'b11111111111111110000110011110100;
assign LUT_2[45812] = 32'b11111111111111101001100000000111;
assign LUT_2[45813] = 32'b11111111111111100110011000100000;
assign LUT_2[45814] = 32'b11111111111111110000011001000011;
assign LUT_2[45815] = 32'b11111111111111101101010001011100;
assign LUT_2[45816] = 32'b11111111111111100111110011111100;
assign LUT_2[45817] = 32'b11111111111111100100101100010101;
assign LUT_2[45818] = 32'b11111111111111101110101100111000;
assign LUT_2[45819] = 32'b11111111111111101011100101010001;
assign LUT_2[45820] = 32'b11111111111111100100010001100100;
assign LUT_2[45821] = 32'b11111111111111100001001001111101;
assign LUT_2[45822] = 32'b11111111111111101011001010100000;
assign LUT_2[45823] = 32'b11111111111111101000000010111001;
assign LUT_2[45824] = 32'b11111111111111111001100100100000;
assign LUT_2[45825] = 32'b11111111111111110110011100111001;
assign LUT_2[45826] = 32'b00000000000000000000011101011100;
assign LUT_2[45827] = 32'b11111111111111111101010101110101;
assign LUT_2[45828] = 32'b11111111111111110110000010001000;
assign LUT_2[45829] = 32'b11111111111111110010111010100001;
assign LUT_2[45830] = 32'b11111111111111111100111011000100;
assign LUT_2[45831] = 32'b11111111111111111001110011011101;
assign LUT_2[45832] = 32'b11111111111111110100010101111101;
assign LUT_2[45833] = 32'b11111111111111110001001110010110;
assign LUT_2[45834] = 32'b11111111111111111011001110111001;
assign LUT_2[45835] = 32'b11111111111111111000000111010010;
assign LUT_2[45836] = 32'b11111111111111110000110011100101;
assign LUT_2[45837] = 32'b11111111111111101101101011111110;
assign LUT_2[45838] = 32'b11111111111111110111101100100001;
assign LUT_2[45839] = 32'b11111111111111110100100100111010;
assign LUT_2[45840] = 32'b11111111111111110100001000101010;
assign LUT_2[45841] = 32'b11111111111111110001000001000011;
assign LUT_2[45842] = 32'b11111111111111111011000001100110;
assign LUT_2[45843] = 32'b11111111111111110111111001111111;
assign LUT_2[45844] = 32'b11111111111111110000100110010010;
assign LUT_2[45845] = 32'b11111111111111101101011110101011;
assign LUT_2[45846] = 32'b11111111111111110111011111001110;
assign LUT_2[45847] = 32'b11111111111111110100010111100111;
assign LUT_2[45848] = 32'b11111111111111101110111010000111;
assign LUT_2[45849] = 32'b11111111111111101011110010100000;
assign LUT_2[45850] = 32'b11111111111111110101110011000011;
assign LUT_2[45851] = 32'b11111111111111110010101011011100;
assign LUT_2[45852] = 32'b11111111111111101011010111101111;
assign LUT_2[45853] = 32'b11111111111111101000010000001000;
assign LUT_2[45854] = 32'b11111111111111110010010000101011;
assign LUT_2[45855] = 32'b11111111111111101111001001000100;
assign LUT_2[45856] = 32'b11111111111111111010000000001001;
assign LUT_2[45857] = 32'b11111111111111110110111000100010;
assign LUT_2[45858] = 32'b00000000000000000000111001000101;
assign LUT_2[45859] = 32'b11111111111111111101110001011110;
assign LUT_2[45860] = 32'b11111111111111110110011101110001;
assign LUT_2[45861] = 32'b11111111111111110011010110001010;
assign LUT_2[45862] = 32'b11111111111111111101010110101101;
assign LUT_2[45863] = 32'b11111111111111111010001111000110;
assign LUT_2[45864] = 32'b11111111111111110100110001100110;
assign LUT_2[45865] = 32'b11111111111111110001101001111111;
assign LUT_2[45866] = 32'b11111111111111111011101010100010;
assign LUT_2[45867] = 32'b11111111111111111000100010111011;
assign LUT_2[45868] = 32'b11111111111111110001001111001110;
assign LUT_2[45869] = 32'b11111111111111101110000111100111;
assign LUT_2[45870] = 32'b11111111111111111000001000001010;
assign LUT_2[45871] = 32'b11111111111111110101000000100011;
assign LUT_2[45872] = 32'b11111111111111110100100100010011;
assign LUT_2[45873] = 32'b11111111111111110001011100101100;
assign LUT_2[45874] = 32'b11111111111111111011011101001111;
assign LUT_2[45875] = 32'b11111111111111111000010101101000;
assign LUT_2[45876] = 32'b11111111111111110001000001111011;
assign LUT_2[45877] = 32'b11111111111111101101111010010100;
assign LUT_2[45878] = 32'b11111111111111110111111010110111;
assign LUT_2[45879] = 32'b11111111111111110100110011010000;
assign LUT_2[45880] = 32'b11111111111111101111010101110000;
assign LUT_2[45881] = 32'b11111111111111101100001110001001;
assign LUT_2[45882] = 32'b11111111111111110110001110101100;
assign LUT_2[45883] = 32'b11111111111111110011000111000101;
assign LUT_2[45884] = 32'b11111111111111101011110011011000;
assign LUT_2[45885] = 32'b11111111111111101000101011110001;
assign LUT_2[45886] = 32'b11111111111111110010101100010100;
assign LUT_2[45887] = 32'b11111111111111101111100100101101;
assign LUT_2[45888] = 32'b11111111111111110001101101000011;
assign LUT_2[45889] = 32'b11111111111111101110100101011100;
assign LUT_2[45890] = 32'b11111111111111111000100101111111;
assign LUT_2[45891] = 32'b11111111111111110101011110011000;
assign LUT_2[45892] = 32'b11111111111111101110001010101011;
assign LUT_2[45893] = 32'b11111111111111101011000011000100;
assign LUT_2[45894] = 32'b11111111111111110101000011100111;
assign LUT_2[45895] = 32'b11111111111111110001111100000000;
assign LUT_2[45896] = 32'b11111111111111101100011110100000;
assign LUT_2[45897] = 32'b11111111111111101001010110111001;
assign LUT_2[45898] = 32'b11111111111111110011010111011100;
assign LUT_2[45899] = 32'b11111111111111110000001111110101;
assign LUT_2[45900] = 32'b11111111111111101000111100001000;
assign LUT_2[45901] = 32'b11111111111111100101110100100001;
assign LUT_2[45902] = 32'b11111111111111101111110101000100;
assign LUT_2[45903] = 32'b11111111111111101100101101011101;
assign LUT_2[45904] = 32'b11111111111111101100010001001101;
assign LUT_2[45905] = 32'b11111111111111101001001001100110;
assign LUT_2[45906] = 32'b11111111111111110011001010001001;
assign LUT_2[45907] = 32'b11111111111111110000000010100010;
assign LUT_2[45908] = 32'b11111111111111101000101110110101;
assign LUT_2[45909] = 32'b11111111111111100101100111001110;
assign LUT_2[45910] = 32'b11111111111111101111100111110001;
assign LUT_2[45911] = 32'b11111111111111101100100000001010;
assign LUT_2[45912] = 32'b11111111111111100111000010101010;
assign LUT_2[45913] = 32'b11111111111111100011111011000011;
assign LUT_2[45914] = 32'b11111111111111101101111011100110;
assign LUT_2[45915] = 32'b11111111111111101010110011111111;
assign LUT_2[45916] = 32'b11111111111111100011100000010010;
assign LUT_2[45917] = 32'b11111111111111100000011000101011;
assign LUT_2[45918] = 32'b11111111111111101010011001001110;
assign LUT_2[45919] = 32'b11111111111111100111010001100111;
assign LUT_2[45920] = 32'b11111111111111110010001000101100;
assign LUT_2[45921] = 32'b11111111111111101111000001000101;
assign LUT_2[45922] = 32'b11111111111111111001000001101000;
assign LUT_2[45923] = 32'b11111111111111110101111010000001;
assign LUT_2[45924] = 32'b11111111111111101110100110010100;
assign LUT_2[45925] = 32'b11111111111111101011011110101101;
assign LUT_2[45926] = 32'b11111111111111110101011111010000;
assign LUT_2[45927] = 32'b11111111111111110010010111101001;
assign LUT_2[45928] = 32'b11111111111111101100111010001001;
assign LUT_2[45929] = 32'b11111111111111101001110010100010;
assign LUT_2[45930] = 32'b11111111111111110011110011000101;
assign LUT_2[45931] = 32'b11111111111111110000101011011110;
assign LUT_2[45932] = 32'b11111111111111101001010111110001;
assign LUT_2[45933] = 32'b11111111111111100110010000001010;
assign LUT_2[45934] = 32'b11111111111111110000010000101101;
assign LUT_2[45935] = 32'b11111111111111101101001001000110;
assign LUT_2[45936] = 32'b11111111111111101100101100110110;
assign LUT_2[45937] = 32'b11111111111111101001100101001111;
assign LUT_2[45938] = 32'b11111111111111110011100101110010;
assign LUT_2[45939] = 32'b11111111111111110000011110001011;
assign LUT_2[45940] = 32'b11111111111111101001001010011110;
assign LUT_2[45941] = 32'b11111111111111100110000010110111;
assign LUT_2[45942] = 32'b11111111111111110000000011011010;
assign LUT_2[45943] = 32'b11111111111111101100111011110011;
assign LUT_2[45944] = 32'b11111111111111100111011110010011;
assign LUT_2[45945] = 32'b11111111111111100100010110101100;
assign LUT_2[45946] = 32'b11111111111111101110010111001111;
assign LUT_2[45947] = 32'b11111111111111101011001111101000;
assign LUT_2[45948] = 32'b11111111111111100011111011111011;
assign LUT_2[45949] = 32'b11111111111111100000110100010100;
assign LUT_2[45950] = 32'b11111111111111101010110100110111;
assign LUT_2[45951] = 32'b11111111111111100111101101010000;
assign LUT_2[45952] = 32'b11111111111111111101111000101111;
assign LUT_2[45953] = 32'b11111111111111111010110001001000;
assign LUT_2[45954] = 32'b00000000000000000100110001101011;
assign LUT_2[45955] = 32'b00000000000000000001101010000100;
assign LUT_2[45956] = 32'b11111111111111111010010110010111;
assign LUT_2[45957] = 32'b11111111111111110111001110110000;
assign LUT_2[45958] = 32'b00000000000000000001001111010011;
assign LUT_2[45959] = 32'b11111111111111111110000111101100;
assign LUT_2[45960] = 32'b11111111111111111000101010001100;
assign LUT_2[45961] = 32'b11111111111111110101100010100101;
assign LUT_2[45962] = 32'b11111111111111111111100011001000;
assign LUT_2[45963] = 32'b11111111111111111100011011100001;
assign LUT_2[45964] = 32'b11111111111111110101000111110100;
assign LUT_2[45965] = 32'b11111111111111110010000000001101;
assign LUT_2[45966] = 32'b11111111111111111100000000110000;
assign LUT_2[45967] = 32'b11111111111111111000111001001001;
assign LUT_2[45968] = 32'b11111111111111111000011100111001;
assign LUT_2[45969] = 32'b11111111111111110101010101010010;
assign LUT_2[45970] = 32'b11111111111111111111010101110101;
assign LUT_2[45971] = 32'b11111111111111111100001110001110;
assign LUT_2[45972] = 32'b11111111111111110100111010100001;
assign LUT_2[45973] = 32'b11111111111111110001110010111010;
assign LUT_2[45974] = 32'b11111111111111111011110011011101;
assign LUT_2[45975] = 32'b11111111111111111000101011110110;
assign LUT_2[45976] = 32'b11111111111111110011001110010110;
assign LUT_2[45977] = 32'b11111111111111110000000110101111;
assign LUT_2[45978] = 32'b11111111111111111010000111010010;
assign LUT_2[45979] = 32'b11111111111111110110111111101011;
assign LUT_2[45980] = 32'b11111111111111101111101011111110;
assign LUT_2[45981] = 32'b11111111111111101100100100010111;
assign LUT_2[45982] = 32'b11111111111111110110100100111010;
assign LUT_2[45983] = 32'b11111111111111110011011101010011;
assign LUT_2[45984] = 32'b11111111111111111110010100011000;
assign LUT_2[45985] = 32'b11111111111111111011001100110001;
assign LUT_2[45986] = 32'b00000000000000000101001101010100;
assign LUT_2[45987] = 32'b00000000000000000010000101101101;
assign LUT_2[45988] = 32'b11111111111111111010110010000000;
assign LUT_2[45989] = 32'b11111111111111110111101010011001;
assign LUT_2[45990] = 32'b00000000000000000001101010111100;
assign LUT_2[45991] = 32'b11111111111111111110100011010101;
assign LUT_2[45992] = 32'b11111111111111111001000101110101;
assign LUT_2[45993] = 32'b11111111111111110101111110001110;
assign LUT_2[45994] = 32'b11111111111111111111111110110001;
assign LUT_2[45995] = 32'b11111111111111111100110111001010;
assign LUT_2[45996] = 32'b11111111111111110101100011011101;
assign LUT_2[45997] = 32'b11111111111111110010011011110110;
assign LUT_2[45998] = 32'b11111111111111111100011100011001;
assign LUT_2[45999] = 32'b11111111111111111001010100110010;
assign LUT_2[46000] = 32'b11111111111111111000111000100010;
assign LUT_2[46001] = 32'b11111111111111110101110000111011;
assign LUT_2[46002] = 32'b11111111111111111111110001011110;
assign LUT_2[46003] = 32'b11111111111111111100101001110111;
assign LUT_2[46004] = 32'b11111111111111110101010110001010;
assign LUT_2[46005] = 32'b11111111111111110010001110100011;
assign LUT_2[46006] = 32'b11111111111111111100001111000110;
assign LUT_2[46007] = 32'b11111111111111111001000111011111;
assign LUT_2[46008] = 32'b11111111111111110011101001111111;
assign LUT_2[46009] = 32'b11111111111111110000100010011000;
assign LUT_2[46010] = 32'b11111111111111111010100010111011;
assign LUT_2[46011] = 32'b11111111111111110111011011010100;
assign LUT_2[46012] = 32'b11111111111111110000000111100111;
assign LUT_2[46013] = 32'b11111111111111101101000000000000;
assign LUT_2[46014] = 32'b11111111111111110111000000100011;
assign LUT_2[46015] = 32'b11111111111111110011111000111100;
assign LUT_2[46016] = 32'b11111111111111110110000001010010;
assign LUT_2[46017] = 32'b11111111111111110010111001101011;
assign LUT_2[46018] = 32'b11111111111111111100111010001110;
assign LUT_2[46019] = 32'b11111111111111111001110010100111;
assign LUT_2[46020] = 32'b11111111111111110010011110111010;
assign LUT_2[46021] = 32'b11111111111111101111010111010011;
assign LUT_2[46022] = 32'b11111111111111111001010111110110;
assign LUT_2[46023] = 32'b11111111111111110110010000001111;
assign LUT_2[46024] = 32'b11111111111111110000110010101111;
assign LUT_2[46025] = 32'b11111111111111101101101011001000;
assign LUT_2[46026] = 32'b11111111111111110111101011101011;
assign LUT_2[46027] = 32'b11111111111111110100100100000100;
assign LUT_2[46028] = 32'b11111111111111101101010000010111;
assign LUT_2[46029] = 32'b11111111111111101010001000110000;
assign LUT_2[46030] = 32'b11111111111111110100001001010011;
assign LUT_2[46031] = 32'b11111111111111110001000001101100;
assign LUT_2[46032] = 32'b11111111111111110000100101011100;
assign LUT_2[46033] = 32'b11111111111111101101011101110101;
assign LUT_2[46034] = 32'b11111111111111110111011110011000;
assign LUT_2[46035] = 32'b11111111111111110100010110110001;
assign LUT_2[46036] = 32'b11111111111111101101000011000100;
assign LUT_2[46037] = 32'b11111111111111101001111011011101;
assign LUT_2[46038] = 32'b11111111111111110011111100000000;
assign LUT_2[46039] = 32'b11111111111111110000110100011001;
assign LUT_2[46040] = 32'b11111111111111101011010110111001;
assign LUT_2[46041] = 32'b11111111111111101000001111010010;
assign LUT_2[46042] = 32'b11111111111111110010001111110101;
assign LUT_2[46043] = 32'b11111111111111101111001000001110;
assign LUT_2[46044] = 32'b11111111111111100111110100100001;
assign LUT_2[46045] = 32'b11111111111111100100101100111010;
assign LUT_2[46046] = 32'b11111111111111101110101101011101;
assign LUT_2[46047] = 32'b11111111111111101011100101110110;
assign LUT_2[46048] = 32'b11111111111111110110011100111011;
assign LUT_2[46049] = 32'b11111111111111110011010101010100;
assign LUT_2[46050] = 32'b11111111111111111101010101110111;
assign LUT_2[46051] = 32'b11111111111111111010001110010000;
assign LUT_2[46052] = 32'b11111111111111110010111010100011;
assign LUT_2[46053] = 32'b11111111111111101111110010111100;
assign LUT_2[46054] = 32'b11111111111111111001110011011111;
assign LUT_2[46055] = 32'b11111111111111110110101011111000;
assign LUT_2[46056] = 32'b11111111111111110001001110011000;
assign LUT_2[46057] = 32'b11111111111111101110000110110001;
assign LUT_2[46058] = 32'b11111111111111111000000111010100;
assign LUT_2[46059] = 32'b11111111111111110100111111101101;
assign LUT_2[46060] = 32'b11111111111111101101101100000000;
assign LUT_2[46061] = 32'b11111111111111101010100100011001;
assign LUT_2[46062] = 32'b11111111111111110100100100111100;
assign LUT_2[46063] = 32'b11111111111111110001011101010101;
assign LUT_2[46064] = 32'b11111111111111110001000001000101;
assign LUT_2[46065] = 32'b11111111111111101101111001011110;
assign LUT_2[46066] = 32'b11111111111111110111111010000001;
assign LUT_2[46067] = 32'b11111111111111110100110010011010;
assign LUT_2[46068] = 32'b11111111111111101101011110101101;
assign LUT_2[46069] = 32'b11111111111111101010010111000110;
assign LUT_2[46070] = 32'b11111111111111110100010111101001;
assign LUT_2[46071] = 32'b11111111111111110001010000000010;
assign LUT_2[46072] = 32'b11111111111111101011110010100010;
assign LUT_2[46073] = 32'b11111111111111101000101010111011;
assign LUT_2[46074] = 32'b11111111111111110010101011011110;
assign LUT_2[46075] = 32'b11111111111111101111100011110111;
assign LUT_2[46076] = 32'b11111111111111101000010000001010;
assign LUT_2[46077] = 32'b11111111111111100101001000100011;
assign LUT_2[46078] = 32'b11111111111111101111001001000110;
assign LUT_2[46079] = 32'b11111111111111101100000001011111;
assign LUT_2[46080] = 32'b11111111111111110111100000001101;
assign LUT_2[46081] = 32'b11111111111111110100011000100110;
assign LUT_2[46082] = 32'b11111111111111111110011001001001;
assign LUT_2[46083] = 32'b11111111111111111011010001100010;
assign LUT_2[46084] = 32'b11111111111111110011111101110101;
assign LUT_2[46085] = 32'b11111111111111110000110110001110;
assign LUT_2[46086] = 32'b11111111111111111010110110110001;
assign LUT_2[46087] = 32'b11111111111111110111101111001010;
assign LUT_2[46088] = 32'b11111111111111110010010001101010;
assign LUT_2[46089] = 32'b11111111111111101111001010000011;
assign LUT_2[46090] = 32'b11111111111111111001001010100110;
assign LUT_2[46091] = 32'b11111111111111110110000010111111;
assign LUT_2[46092] = 32'b11111111111111101110101111010010;
assign LUT_2[46093] = 32'b11111111111111101011100111101011;
assign LUT_2[46094] = 32'b11111111111111110101101000001110;
assign LUT_2[46095] = 32'b11111111111111110010100000100111;
assign LUT_2[46096] = 32'b11111111111111110010000100010111;
assign LUT_2[46097] = 32'b11111111111111101110111100110000;
assign LUT_2[46098] = 32'b11111111111111111000111101010011;
assign LUT_2[46099] = 32'b11111111111111110101110101101100;
assign LUT_2[46100] = 32'b11111111111111101110100001111111;
assign LUT_2[46101] = 32'b11111111111111101011011010011000;
assign LUT_2[46102] = 32'b11111111111111110101011010111011;
assign LUT_2[46103] = 32'b11111111111111110010010011010100;
assign LUT_2[46104] = 32'b11111111111111101100110101110100;
assign LUT_2[46105] = 32'b11111111111111101001101110001101;
assign LUT_2[46106] = 32'b11111111111111110011101110110000;
assign LUT_2[46107] = 32'b11111111111111110000100111001001;
assign LUT_2[46108] = 32'b11111111111111101001010011011100;
assign LUT_2[46109] = 32'b11111111111111100110001011110101;
assign LUT_2[46110] = 32'b11111111111111110000001100011000;
assign LUT_2[46111] = 32'b11111111111111101101000100110001;
assign LUT_2[46112] = 32'b11111111111111110111111011110110;
assign LUT_2[46113] = 32'b11111111111111110100110100001111;
assign LUT_2[46114] = 32'b11111111111111111110110100110010;
assign LUT_2[46115] = 32'b11111111111111111011101101001011;
assign LUT_2[46116] = 32'b11111111111111110100011001011110;
assign LUT_2[46117] = 32'b11111111111111110001010001110111;
assign LUT_2[46118] = 32'b11111111111111111011010010011010;
assign LUT_2[46119] = 32'b11111111111111111000001010110011;
assign LUT_2[46120] = 32'b11111111111111110010101101010011;
assign LUT_2[46121] = 32'b11111111111111101111100101101100;
assign LUT_2[46122] = 32'b11111111111111111001100110001111;
assign LUT_2[46123] = 32'b11111111111111110110011110101000;
assign LUT_2[46124] = 32'b11111111111111101111001010111011;
assign LUT_2[46125] = 32'b11111111111111101100000011010100;
assign LUT_2[46126] = 32'b11111111111111110110000011110111;
assign LUT_2[46127] = 32'b11111111111111110010111100010000;
assign LUT_2[46128] = 32'b11111111111111110010100000000000;
assign LUT_2[46129] = 32'b11111111111111101111011000011001;
assign LUT_2[46130] = 32'b11111111111111111001011000111100;
assign LUT_2[46131] = 32'b11111111111111110110010001010101;
assign LUT_2[46132] = 32'b11111111111111101110111101101000;
assign LUT_2[46133] = 32'b11111111111111101011110110000001;
assign LUT_2[46134] = 32'b11111111111111110101110110100100;
assign LUT_2[46135] = 32'b11111111111111110010101110111101;
assign LUT_2[46136] = 32'b11111111111111101101010001011101;
assign LUT_2[46137] = 32'b11111111111111101010001001110110;
assign LUT_2[46138] = 32'b11111111111111110100001010011001;
assign LUT_2[46139] = 32'b11111111111111110001000010110010;
assign LUT_2[46140] = 32'b11111111111111101001101111000101;
assign LUT_2[46141] = 32'b11111111111111100110100111011110;
assign LUT_2[46142] = 32'b11111111111111110000101000000001;
assign LUT_2[46143] = 32'b11111111111111101101100000011010;
assign LUT_2[46144] = 32'b11111111111111101111101000110000;
assign LUT_2[46145] = 32'b11111111111111101100100001001001;
assign LUT_2[46146] = 32'b11111111111111110110100001101100;
assign LUT_2[46147] = 32'b11111111111111110011011010000101;
assign LUT_2[46148] = 32'b11111111111111101100000110011000;
assign LUT_2[46149] = 32'b11111111111111101000111110110001;
assign LUT_2[46150] = 32'b11111111111111110010111111010100;
assign LUT_2[46151] = 32'b11111111111111101111110111101101;
assign LUT_2[46152] = 32'b11111111111111101010011010001101;
assign LUT_2[46153] = 32'b11111111111111100111010010100110;
assign LUT_2[46154] = 32'b11111111111111110001010011001001;
assign LUT_2[46155] = 32'b11111111111111101110001011100010;
assign LUT_2[46156] = 32'b11111111111111100110110111110101;
assign LUT_2[46157] = 32'b11111111111111100011110000001110;
assign LUT_2[46158] = 32'b11111111111111101101110000110001;
assign LUT_2[46159] = 32'b11111111111111101010101001001010;
assign LUT_2[46160] = 32'b11111111111111101010001100111010;
assign LUT_2[46161] = 32'b11111111111111100111000101010011;
assign LUT_2[46162] = 32'b11111111111111110001000101110110;
assign LUT_2[46163] = 32'b11111111111111101101111110001111;
assign LUT_2[46164] = 32'b11111111111111100110101010100010;
assign LUT_2[46165] = 32'b11111111111111100011100010111011;
assign LUT_2[46166] = 32'b11111111111111101101100011011110;
assign LUT_2[46167] = 32'b11111111111111101010011011110111;
assign LUT_2[46168] = 32'b11111111111111100100111110010111;
assign LUT_2[46169] = 32'b11111111111111100001110110110000;
assign LUT_2[46170] = 32'b11111111111111101011110111010011;
assign LUT_2[46171] = 32'b11111111111111101000101111101100;
assign LUT_2[46172] = 32'b11111111111111100001011011111111;
assign LUT_2[46173] = 32'b11111111111111011110010100011000;
assign LUT_2[46174] = 32'b11111111111111101000010100111011;
assign LUT_2[46175] = 32'b11111111111111100101001101010100;
assign LUT_2[46176] = 32'b11111111111111110000000100011001;
assign LUT_2[46177] = 32'b11111111111111101100111100110010;
assign LUT_2[46178] = 32'b11111111111111110110111101010101;
assign LUT_2[46179] = 32'b11111111111111110011110101101110;
assign LUT_2[46180] = 32'b11111111111111101100100010000001;
assign LUT_2[46181] = 32'b11111111111111101001011010011010;
assign LUT_2[46182] = 32'b11111111111111110011011010111101;
assign LUT_2[46183] = 32'b11111111111111110000010011010110;
assign LUT_2[46184] = 32'b11111111111111101010110101110110;
assign LUT_2[46185] = 32'b11111111111111100111101110001111;
assign LUT_2[46186] = 32'b11111111111111110001101110110010;
assign LUT_2[46187] = 32'b11111111111111101110100111001011;
assign LUT_2[46188] = 32'b11111111111111100111010011011110;
assign LUT_2[46189] = 32'b11111111111111100100001011110111;
assign LUT_2[46190] = 32'b11111111111111101110001100011010;
assign LUT_2[46191] = 32'b11111111111111101011000100110011;
assign LUT_2[46192] = 32'b11111111111111101010101000100011;
assign LUT_2[46193] = 32'b11111111111111100111100000111100;
assign LUT_2[46194] = 32'b11111111111111110001100001011111;
assign LUT_2[46195] = 32'b11111111111111101110011001111000;
assign LUT_2[46196] = 32'b11111111111111100111000110001011;
assign LUT_2[46197] = 32'b11111111111111100011111110100100;
assign LUT_2[46198] = 32'b11111111111111101101111111000111;
assign LUT_2[46199] = 32'b11111111111111101010110111100000;
assign LUT_2[46200] = 32'b11111111111111100101011010000000;
assign LUT_2[46201] = 32'b11111111111111100010010010011001;
assign LUT_2[46202] = 32'b11111111111111101100010010111100;
assign LUT_2[46203] = 32'b11111111111111101001001011010101;
assign LUT_2[46204] = 32'b11111111111111100001110111101000;
assign LUT_2[46205] = 32'b11111111111111011110110000000001;
assign LUT_2[46206] = 32'b11111111111111101000110000100100;
assign LUT_2[46207] = 32'b11111111111111100101101000111101;
assign LUT_2[46208] = 32'b11111111111111111011110100011100;
assign LUT_2[46209] = 32'b11111111111111111000101100110101;
assign LUT_2[46210] = 32'b00000000000000000010101101011000;
assign LUT_2[46211] = 32'b11111111111111111111100101110001;
assign LUT_2[46212] = 32'b11111111111111111000010010000100;
assign LUT_2[46213] = 32'b11111111111111110101001010011101;
assign LUT_2[46214] = 32'b11111111111111111111001011000000;
assign LUT_2[46215] = 32'b11111111111111111100000011011001;
assign LUT_2[46216] = 32'b11111111111111110110100101111001;
assign LUT_2[46217] = 32'b11111111111111110011011110010010;
assign LUT_2[46218] = 32'b11111111111111111101011110110101;
assign LUT_2[46219] = 32'b11111111111111111010010111001110;
assign LUT_2[46220] = 32'b11111111111111110011000011100001;
assign LUT_2[46221] = 32'b11111111111111101111111011111010;
assign LUT_2[46222] = 32'b11111111111111111001111100011101;
assign LUT_2[46223] = 32'b11111111111111110110110100110110;
assign LUT_2[46224] = 32'b11111111111111110110011000100110;
assign LUT_2[46225] = 32'b11111111111111110011010000111111;
assign LUT_2[46226] = 32'b11111111111111111101010001100010;
assign LUT_2[46227] = 32'b11111111111111111010001001111011;
assign LUT_2[46228] = 32'b11111111111111110010110110001110;
assign LUT_2[46229] = 32'b11111111111111101111101110100111;
assign LUT_2[46230] = 32'b11111111111111111001101111001010;
assign LUT_2[46231] = 32'b11111111111111110110100111100011;
assign LUT_2[46232] = 32'b11111111111111110001001010000011;
assign LUT_2[46233] = 32'b11111111111111101110000010011100;
assign LUT_2[46234] = 32'b11111111111111111000000010111111;
assign LUT_2[46235] = 32'b11111111111111110100111011011000;
assign LUT_2[46236] = 32'b11111111111111101101100111101011;
assign LUT_2[46237] = 32'b11111111111111101010100000000100;
assign LUT_2[46238] = 32'b11111111111111110100100000100111;
assign LUT_2[46239] = 32'b11111111111111110001011001000000;
assign LUT_2[46240] = 32'b11111111111111111100010000000101;
assign LUT_2[46241] = 32'b11111111111111111001001000011110;
assign LUT_2[46242] = 32'b00000000000000000011001001000001;
assign LUT_2[46243] = 32'b00000000000000000000000001011010;
assign LUT_2[46244] = 32'b11111111111111111000101101101101;
assign LUT_2[46245] = 32'b11111111111111110101100110000110;
assign LUT_2[46246] = 32'b11111111111111111111100110101001;
assign LUT_2[46247] = 32'b11111111111111111100011111000010;
assign LUT_2[46248] = 32'b11111111111111110111000001100010;
assign LUT_2[46249] = 32'b11111111111111110011111001111011;
assign LUT_2[46250] = 32'b11111111111111111101111010011110;
assign LUT_2[46251] = 32'b11111111111111111010110010110111;
assign LUT_2[46252] = 32'b11111111111111110011011111001010;
assign LUT_2[46253] = 32'b11111111111111110000010111100011;
assign LUT_2[46254] = 32'b11111111111111111010011000000110;
assign LUT_2[46255] = 32'b11111111111111110111010000011111;
assign LUT_2[46256] = 32'b11111111111111110110110100001111;
assign LUT_2[46257] = 32'b11111111111111110011101100101000;
assign LUT_2[46258] = 32'b11111111111111111101101101001011;
assign LUT_2[46259] = 32'b11111111111111111010100101100100;
assign LUT_2[46260] = 32'b11111111111111110011010001110111;
assign LUT_2[46261] = 32'b11111111111111110000001010010000;
assign LUT_2[46262] = 32'b11111111111111111010001010110011;
assign LUT_2[46263] = 32'b11111111111111110111000011001100;
assign LUT_2[46264] = 32'b11111111111111110001100101101100;
assign LUT_2[46265] = 32'b11111111111111101110011110000101;
assign LUT_2[46266] = 32'b11111111111111111000011110101000;
assign LUT_2[46267] = 32'b11111111111111110101010111000001;
assign LUT_2[46268] = 32'b11111111111111101110000011010100;
assign LUT_2[46269] = 32'b11111111111111101010111011101101;
assign LUT_2[46270] = 32'b11111111111111110100111100010000;
assign LUT_2[46271] = 32'b11111111111111110001110100101001;
assign LUT_2[46272] = 32'b11111111111111110011111100111111;
assign LUT_2[46273] = 32'b11111111111111110000110101011000;
assign LUT_2[46274] = 32'b11111111111111111010110101111011;
assign LUT_2[46275] = 32'b11111111111111110111101110010100;
assign LUT_2[46276] = 32'b11111111111111110000011010100111;
assign LUT_2[46277] = 32'b11111111111111101101010011000000;
assign LUT_2[46278] = 32'b11111111111111110111010011100011;
assign LUT_2[46279] = 32'b11111111111111110100001011111100;
assign LUT_2[46280] = 32'b11111111111111101110101110011100;
assign LUT_2[46281] = 32'b11111111111111101011100110110101;
assign LUT_2[46282] = 32'b11111111111111110101100111011000;
assign LUT_2[46283] = 32'b11111111111111110010011111110001;
assign LUT_2[46284] = 32'b11111111111111101011001100000100;
assign LUT_2[46285] = 32'b11111111111111101000000100011101;
assign LUT_2[46286] = 32'b11111111111111110010000101000000;
assign LUT_2[46287] = 32'b11111111111111101110111101011001;
assign LUT_2[46288] = 32'b11111111111111101110100001001001;
assign LUT_2[46289] = 32'b11111111111111101011011001100010;
assign LUT_2[46290] = 32'b11111111111111110101011010000101;
assign LUT_2[46291] = 32'b11111111111111110010010010011110;
assign LUT_2[46292] = 32'b11111111111111101010111110110001;
assign LUT_2[46293] = 32'b11111111111111100111110111001010;
assign LUT_2[46294] = 32'b11111111111111110001110111101101;
assign LUT_2[46295] = 32'b11111111111111101110110000000110;
assign LUT_2[46296] = 32'b11111111111111101001010010100110;
assign LUT_2[46297] = 32'b11111111111111100110001010111111;
assign LUT_2[46298] = 32'b11111111111111110000001011100010;
assign LUT_2[46299] = 32'b11111111111111101101000011111011;
assign LUT_2[46300] = 32'b11111111111111100101110000001110;
assign LUT_2[46301] = 32'b11111111111111100010101000100111;
assign LUT_2[46302] = 32'b11111111111111101100101001001010;
assign LUT_2[46303] = 32'b11111111111111101001100001100011;
assign LUT_2[46304] = 32'b11111111111111110100011000101000;
assign LUT_2[46305] = 32'b11111111111111110001010001000001;
assign LUT_2[46306] = 32'b11111111111111111011010001100100;
assign LUT_2[46307] = 32'b11111111111111111000001001111101;
assign LUT_2[46308] = 32'b11111111111111110000110110010000;
assign LUT_2[46309] = 32'b11111111111111101101101110101001;
assign LUT_2[46310] = 32'b11111111111111110111101111001100;
assign LUT_2[46311] = 32'b11111111111111110100100111100101;
assign LUT_2[46312] = 32'b11111111111111101111001010000101;
assign LUT_2[46313] = 32'b11111111111111101100000010011110;
assign LUT_2[46314] = 32'b11111111111111110110000011000001;
assign LUT_2[46315] = 32'b11111111111111110010111011011010;
assign LUT_2[46316] = 32'b11111111111111101011100111101101;
assign LUT_2[46317] = 32'b11111111111111101000100000000110;
assign LUT_2[46318] = 32'b11111111111111110010100000101001;
assign LUT_2[46319] = 32'b11111111111111101111011001000010;
assign LUT_2[46320] = 32'b11111111111111101110111100110010;
assign LUT_2[46321] = 32'b11111111111111101011110101001011;
assign LUT_2[46322] = 32'b11111111111111110101110101101110;
assign LUT_2[46323] = 32'b11111111111111110010101110000111;
assign LUT_2[46324] = 32'b11111111111111101011011010011010;
assign LUT_2[46325] = 32'b11111111111111101000010010110011;
assign LUT_2[46326] = 32'b11111111111111110010010011010110;
assign LUT_2[46327] = 32'b11111111111111101111001011101111;
assign LUT_2[46328] = 32'b11111111111111101001101110001111;
assign LUT_2[46329] = 32'b11111111111111100110100110101000;
assign LUT_2[46330] = 32'b11111111111111110000100111001011;
assign LUT_2[46331] = 32'b11111111111111101101011111100100;
assign LUT_2[46332] = 32'b11111111111111100110001011110111;
assign LUT_2[46333] = 32'b11111111111111100011000100010000;
assign LUT_2[46334] = 32'b11111111111111101101000100110011;
assign LUT_2[46335] = 32'b11111111111111101001111101001100;
assign LUT_2[46336] = 32'b11111111111111111011011110110011;
assign LUT_2[46337] = 32'b11111111111111111000010111001100;
assign LUT_2[46338] = 32'b00000000000000000010010111101111;
assign LUT_2[46339] = 32'b11111111111111111111010000001000;
assign LUT_2[46340] = 32'b11111111111111110111111100011011;
assign LUT_2[46341] = 32'b11111111111111110100110100110100;
assign LUT_2[46342] = 32'b11111111111111111110110101010111;
assign LUT_2[46343] = 32'b11111111111111111011101101110000;
assign LUT_2[46344] = 32'b11111111111111110110010000010000;
assign LUT_2[46345] = 32'b11111111111111110011001000101001;
assign LUT_2[46346] = 32'b11111111111111111101001001001100;
assign LUT_2[46347] = 32'b11111111111111111010000001100101;
assign LUT_2[46348] = 32'b11111111111111110010101101111000;
assign LUT_2[46349] = 32'b11111111111111101111100110010001;
assign LUT_2[46350] = 32'b11111111111111111001100110110100;
assign LUT_2[46351] = 32'b11111111111111110110011111001101;
assign LUT_2[46352] = 32'b11111111111111110110000010111101;
assign LUT_2[46353] = 32'b11111111111111110010111011010110;
assign LUT_2[46354] = 32'b11111111111111111100111011111001;
assign LUT_2[46355] = 32'b11111111111111111001110100010010;
assign LUT_2[46356] = 32'b11111111111111110010100000100101;
assign LUT_2[46357] = 32'b11111111111111101111011000111110;
assign LUT_2[46358] = 32'b11111111111111111001011001100001;
assign LUT_2[46359] = 32'b11111111111111110110010001111010;
assign LUT_2[46360] = 32'b11111111111111110000110100011010;
assign LUT_2[46361] = 32'b11111111111111101101101100110011;
assign LUT_2[46362] = 32'b11111111111111110111101101010110;
assign LUT_2[46363] = 32'b11111111111111110100100101101111;
assign LUT_2[46364] = 32'b11111111111111101101010010000010;
assign LUT_2[46365] = 32'b11111111111111101010001010011011;
assign LUT_2[46366] = 32'b11111111111111110100001010111110;
assign LUT_2[46367] = 32'b11111111111111110001000011010111;
assign LUT_2[46368] = 32'b11111111111111111011111010011100;
assign LUT_2[46369] = 32'b11111111111111111000110010110101;
assign LUT_2[46370] = 32'b00000000000000000010110011011000;
assign LUT_2[46371] = 32'b11111111111111111111101011110001;
assign LUT_2[46372] = 32'b11111111111111111000011000000100;
assign LUT_2[46373] = 32'b11111111111111110101010000011101;
assign LUT_2[46374] = 32'b11111111111111111111010001000000;
assign LUT_2[46375] = 32'b11111111111111111100001001011001;
assign LUT_2[46376] = 32'b11111111111111110110101011111001;
assign LUT_2[46377] = 32'b11111111111111110011100100010010;
assign LUT_2[46378] = 32'b11111111111111111101100100110101;
assign LUT_2[46379] = 32'b11111111111111111010011101001110;
assign LUT_2[46380] = 32'b11111111111111110011001001100001;
assign LUT_2[46381] = 32'b11111111111111110000000001111010;
assign LUT_2[46382] = 32'b11111111111111111010000010011101;
assign LUT_2[46383] = 32'b11111111111111110110111010110110;
assign LUT_2[46384] = 32'b11111111111111110110011110100110;
assign LUT_2[46385] = 32'b11111111111111110011010110111111;
assign LUT_2[46386] = 32'b11111111111111111101010111100010;
assign LUT_2[46387] = 32'b11111111111111111010001111111011;
assign LUT_2[46388] = 32'b11111111111111110010111100001110;
assign LUT_2[46389] = 32'b11111111111111101111110100100111;
assign LUT_2[46390] = 32'b11111111111111111001110101001010;
assign LUT_2[46391] = 32'b11111111111111110110101101100011;
assign LUT_2[46392] = 32'b11111111111111110001010000000011;
assign LUT_2[46393] = 32'b11111111111111101110001000011100;
assign LUT_2[46394] = 32'b11111111111111111000001000111111;
assign LUT_2[46395] = 32'b11111111111111110101000001011000;
assign LUT_2[46396] = 32'b11111111111111101101101101101011;
assign LUT_2[46397] = 32'b11111111111111101010100110000100;
assign LUT_2[46398] = 32'b11111111111111110100100110100111;
assign LUT_2[46399] = 32'b11111111111111110001011111000000;
assign LUT_2[46400] = 32'b11111111111111110011100111010110;
assign LUT_2[46401] = 32'b11111111111111110000011111101111;
assign LUT_2[46402] = 32'b11111111111111111010100000010010;
assign LUT_2[46403] = 32'b11111111111111110111011000101011;
assign LUT_2[46404] = 32'b11111111111111110000000100111110;
assign LUT_2[46405] = 32'b11111111111111101100111101010111;
assign LUT_2[46406] = 32'b11111111111111110110111101111010;
assign LUT_2[46407] = 32'b11111111111111110011110110010011;
assign LUT_2[46408] = 32'b11111111111111101110011000110011;
assign LUT_2[46409] = 32'b11111111111111101011010001001100;
assign LUT_2[46410] = 32'b11111111111111110101010001101111;
assign LUT_2[46411] = 32'b11111111111111110010001010001000;
assign LUT_2[46412] = 32'b11111111111111101010110110011011;
assign LUT_2[46413] = 32'b11111111111111100111101110110100;
assign LUT_2[46414] = 32'b11111111111111110001101111010111;
assign LUT_2[46415] = 32'b11111111111111101110100111110000;
assign LUT_2[46416] = 32'b11111111111111101110001011100000;
assign LUT_2[46417] = 32'b11111111111111101011000011111001;
assign LUT_2[46418] = 32'b11111111111111110101000100011100;
assign LUT_2[46419] = 32'b11111111111111110001111100110101;
assign LUT_2[46420] = 32'b11111111111111101010101001001000;
assign LUT_2[46421] = 32'b11111111111111100111100001100001;
assign LUT_2[46422] = 32'b11111111111111110001100010000100;
assign LUT_2[46423] = 32'b11111111111111101110011010011101;
assign LUT_2[46424] = 32'b11111111111111101000111100111101;
assign LUT_2[46425] = 32'b11111111111111100101110101010110;
assign LUT_2[46426] = 32'b11111111111111101111110101111001;
assign LUT_2[46427] = 32'b11111111111111101100101110010010;
assign LUT_2[46428] = 32'b11111111111111100101011010100101;
assign LUT_2[46429] = 32'b11111111111111100010010010111110;
assign LUT_2[46430] = 32'b11111111111111101100010011100001;
assign LUT_2[46431] = 32'b11111111111111101001001011111010;
assign LUT_2[46432] = 32'b11111111111111110100000010111111;
assign LUT_2[46433] = 32'b11111111111111110000111011011000;
assign LUT_2[46434] = 32'b11111111111111111010111011111011;
assign LUT_2[46435] = 32'b11111111111111110111110100010100;
assign LUT_2[46436] = 32'b11111111111111110000100000100111;
assign LUT_2[46437] = 32'b11111111111111101101011001000000;
assign LUT_2[46438] = 32'b11111111111111110111011001100011;
assign LUT_2[46439] = 32'b11111111111111110100010001111100;
assign LUT_2[46440] = 32'b11111111111111101110110100011100;
assign LUT_2[46441] = 32'b11111111111111101011101100110101;
assign LUT_2[46442] = 32'b11111111111111110101101101011000;
assign LUT_2[46443] = 32'b11111111111111110010100101110001;
assign LUT_2[46444] = 32'b11111111111111101011010010000100;
assign LUT_2[46445] = 32'b11111111111111101000001010011101;
assign LUT_2[46446] = 32'b11111111111111110010001011000000;
assign LUT_2[46447] = 32'b11111111111111101111000011011001;
assign LUT_2[46448] = 32'b11111111111111101110100111001001;
assign LUT_2[46449] = 32'b11111111111111101011011111100010;
assign LUT_2[46450] = 32'b11111111111111110101100000000101;
assign LUT_2[46451] = 32'b11111111111111110010011000011110;
assign LUT_2[46452] = 32'b11111111111111101011000100110001;
assign LUT_2[46453] = 32'b11111111111111100111111101001010;
assign LUT_2[46454] = 32'b11111111111111110001111101101101;
assign LUT_2[46455] = 32'b11111111111111101110110110000110;
assign LUT_2[46456] = 32'b11111111111111101001011000100110;
assign LUT_2[46457] = 32'b11111111111111100110010000111111;
assign LUT_2[46458] = 32'b11111111111111110000010001100010;
assign LUT_2[46459] = 32'b11111111111111101101001001111011;
assign LUT_2[46460] = 32'b11111111111111100101110110001110;
assign LUT_2[46461] = 32'b11111111111111100010101110100111;
assign LUT_2[46462] = 32'b11111111111111101100101111001010;
assign LUT_2[46463] = 32'b11111111111111101001100111100011;
assign LUT_2[46464] = 32'b11111111111111111111110011000010;
assign LUT_2[46465] = 32'b11111111111111111100101011011011;
assign LUT_2[46466] = 32'b00000000000000000110101011111110;
assign LUT_2[46467] = 32'b00000000000000000011100100010111;
assign LUT_2[46468] = 32'b11111111111111111100010000101010;
assign LUT_2[46469] = 32'b11111111111111111001001001000011;
assign LUT_2[46470] = 32'b00000000000000000011001001100110;
assign LUT_2[46471] = 32'b00000000000000000000000001111111;
assign LUT_2[46472] = 32'b11111111111111111010100100011111;
assign LUT_2[46473] = 32'b11111111111111110111011100111000;
assign LUT_2[46474] = 32'b00000000000000000001011101011011;
assign LUT_2[46475] = 32'b11111111111111111110010101110100;
assign LUT_2[46476] = 32'b11111111111111110111000010000111;
assign LUT_2[46477] = 32'b11111111111111110011111010100000;
assign LUT_2[46478] = 32'b11111111111111111101111011000011;
assign LUT_2[46479] = 32'b11111111111111111010110011011100;
assign LUT_2[46480] = 32'b11111111111111111010010111001100;
assign LUT_2[46481] = 32'b11111111111111110111001111100101;
assign LUT_2[46482] = 32'b00000000000000000001010000001000;
assign LUT_2[46483] = 32'b11111111111111111110001000100001;
assign LUT_2[46484] = 32'b11111111111111110110110100110100;
assign LUT_2[46485] = 32'b11111111111111110011101101001101;
assign LUT_2[46486] = 32'b11111111111111111101101101110000;
assign LUT_2[46487] = 32'b11111111111111111010100110001001;
assign LUT_2[46488] = 32'b11111111111111110101001000101001;
assign LUT_2[46489] = 32'b11111111111111110010000001000010;
assign LUT_2[46490] = 32'b11111111111111111100000001100101;
assign LUT_2[46491] = 32'b11111111111111111000111001111110;
assign LUT_2[46492] = 32'b11111111111111110001100110010001;
assign LUT_2[46493] = 32'b11111111111111101110011110101010;
assign LUT_2[46494] = 32'b11111111111111111000011111001101;
assign LUT_2[46495] = 32'b11111111111111110101010111100110;
assign LUT_2[46496] = 32'b00000000000000000000001110101011;
assign LUT_2[46497] = 32'b11111111111111111101000111000100;
assign LUT_2[46498] = 32'b00000000000000000111000111100111;
assign LUT_2[46499] = 32'b00000000000000000100000000000000;
assign LUT_2[46500] = 32'b11111111111111111100101100010011;
assign LUT_2[46501] = 32'b11111111111111111001100100101100;
assign LUT_2[46502] = 32'b00000000000000000011100101001111;
assign LUT_2[46503] = 32'b00000000000000000000011101101000;
assign LUT_2[46504] = 32'b11111111111111111011000000001000;
assign LUT_2[46505] = 32'b11111111111111110111111000100001;
assign LUT_2[46506] = 32'b00000000000000000001111001000100;
assign LUT_2[46507] = 32'b11111111111111111110110001011101;
assign LUT_2[46508] = 32'b11111111111111110111011101110000;
assign LUT_2[46509] = 32'b11111111111111110100010110001001;
assign LUT_2[46510] = 32'b11111111111111111110010110101100;
assign LUT_2[46511] = 32'b11111111111111111011001111000101;
assign LUT_2[46512] = 32'b11111111111111111010110010110101;
assign LUT_2[46513] = 32'b11111111111111110111101011001110;
assign LUT_2[46514] = 32'b00000000000000000001101011110001;
assign LUT_2[46515] = 32'b11111111111111111110100100001010;
assign LUT_2[46516] = 32'b11111111111111110111010000011101;
assign LUT_2[46517] = 32'b11111111111111110100001000110110;
assign LUT_2[46518] = 32'b11111111111111111110001001011001;
assign LUT_2[46519] = 32'b11111111111111111011000001110010;
assign LUT_2[46520] = 32'b11111111111111110101100100010010;
assign LUT_2[46521] = 32'b11111111111111110010011100101011;
assign LUT_2[46522] = 32'b11111111111111111100011101001110;
assign LUT_2[46523] = 32'b11111111111111111001010101100111;
assign LUT_2[46524] = 32'b11111111111111110010000001111010;
assign LUT_2[46525] = 32'b11111111111111101110111010010011;
assign LUT_2[46526] = 32'b11111111111111111000111010110110;
assign LUT_2[46527] = 32'b11111111111111110101110011001111;
assign LUT_2[46528] = 32'b11111111111111110111111011100101;
assign LUT_2[46529] = 32'b11111111111111110100110011111110;
assign LUT_2[46530] = 32'b11111111111111111110110100100001;
assign LUT_2[46531] = 32'b11111111111111111011101100111010;
assign LUT_2[46532] = 32'b11111111111111110100011001001101;
assign LUT_2[46533] = 32'b11111111111111110001010001100110;
assign LUT_2[46534] = 32'b11111111111111111011010010001001;
assign LUT_2[46535] = 32'b11111111111111111000001010100010;
assign LUT_2[46536] = 32'b11111111111111110010101101000010;
assign LUT_2[46537] = 32'b11111111111111101111100101011011;
assign LUT_2[46538] = 32'b11111111111111111001100101111110;
assign LUT_2[46539] = 32'b11111111111111110110011110010111;
assign LUT_2[46540] = 32'b11111111111111101111001010101010;
assign LUT_2[46541] = 32'b11111111111111101100000011000011;
assign LUT_2[46542] = 32'b11111111111111110110000011100110;
assign LUT_2[46543] = 32'b11111111111111110010111011111111;
assign LUT_2[46544] = 32'b11111111111111110010011111101111;
assign LUT_2[46545] = 32'b11111111111111101111011000001000;
assign LUT_2[46546] = 32'b11111111111111111001011000101011;
assign LUT_2[46547] = 32'b11111111111111110110010001000100;
assign LUT_2[46548] = 32'b11111111111111101110111101010111;
assign LUT_2[46549] = 32'b11111111111111101011110101110000;
assign LUT_2[46550] = 32'b11111111111111110101110110010011;
assign LUT_2[46551] = 32'b11111111111111110010101110101100;
assign LUT_2[46552] = 32'b11111111111111101101010001001100;
assign LUT_2[46553] = 32'b11111111111111101010001001100101;
assign LUT_2[46554] = 32'b11111111111111110100001010001000;
assign LUT_2[46555] = 32'b11111111111111110001000010100001;
assign LUT_2[46556] = 32'b11111111111111101001101110110100;
assign LUT_2[46557] = 32'b11111111111111100110100111001101;
assign LUT_2[46558] = 32'b11111111111111110000100111110000;
assign LUT_2[46559] = 32'b11111111111111101101100000001001;
assign LUT_2[46560] = 32'b11111111111111111000010111001110;
assign LUT_2[46561] = 32'b11111111111111110101001111100111;
assign LUT_2[46562] = 32'b11111111111111111111010000001010;
assign LUT_2[46563] = 32'b11111111111111111100001000100011;
assign LUT_2[46564] = 32'b11111111111111110100110100110110;
assign LUT_2[46565] = 32'b11111111111111110001101101001111;
assign LUT_2[46566] = 32'b11111111111111111011101101110010;
assign LUT_2[46567] = 32'b11111111111111111000100110001011;
assign LUT_2[46568] = 32'b11111111111111110011001000101011;
assign LUT_2[46569] = 32'b11111111111111110000000001000100;
assign LUT_2[46570] = 32'b11111111111111111010000001100111;
assign LUT_2[46571] = 32'b11111111111111110110111010000000;
assign LUT_2[46572] = 32'b11111111111111101111100110010011;
assign LUT_2[46573] = 32'b11111111111111101100011110101100;
assign LUT_2[46574] = 32'b11111111111111110110011111001111;
assign LUT_2[46575] = 32'b11111111111111110011010111101000;
assign LUT_2[46576] = 32'b11111111111111110010111011011000;
assign LUT_2[46577] = 32'b11111111111111101111110011110001;
assign LUT_2[46578] = 32'b11111111111111111001110100010100;
assign LUT_2[46579] = 32'b11111111111111110110101100101101;
assign LUT_2[46580] = 32'b11111111111111101111011001000000;
assign LUT_2[46581] = 32'b11111111111111101100010001011001;
assign LUT_2[46582] = 32'b11111111111111110110010001111100;
assign LUT_2[46583] = 32'b11111111111111110011001010010101;
assign LUT_2[46584] = 32'b11111111111111101101101100110101;
assign LUT_2[46585] = 32'b11111111111111101010100101001110;
assign LUT_2[46586] = 32'b11111111111111110100100101110001;
assign LUT_2[46587] = 32'b11111111111111110001011110001010;
assign LUT_2[46588] = 32'b11111111111111101010001010011101;
assign LUT_2[46589] = 32'b11111111111111100111000010110110;
assign LUT_2[46590] = 32'b11111111111111110001000011011001;
assign LUT_2[46591] = 32'b11111111111111101101111011110010;
assign LUT_2[46592] = 32'b11111111111111111100010001111111;
assign LUT_2[46593] = 32'b11111111111111111001001010011000;
assign LUT_2[46594] = 32'b00000000000000000011001010111011;
assign LUT_2[46595] = 32'b00000000000000000000000011010100;
assign LUT_2[46596] = 32'b11111111111111111000101111100111;
assign LUT_2[46597] = 32'b11111111111111110101101000000000;
assign LUT_2[46598] = 32'b11111111111111111111101000100011;
assign LUT_2[46599] = 32'b11111111111111111100100000111100;
assign LUT_2[46600] = 32'b11111111111111110111000011011100;
assign LUT_2[46601] = 32'b11111111111111110011111011110101;
assign LUT_2[46602] = 32'b11111111111111111101111100011000;
assign LUT_2[46603] = 32'b11111111111111111010110100110001;
assign LUT_2[46604] = 32'b11111111111111110011100001000100;
assign LUT_2[46605] = 32'b11111111111111110000011001011101;
assign LUT_2[46606] = 32'b11111111111111111010011010000000;
assign LUT_2[46607] = 32'b11111111111111110111010010011001;
assign LUT_2[46608] = 32'b11111111111111110110110110001001;
assign LUT_2[46609] = 32'b11111111111111110011101110100010;
assign LUT_2[46610] = 32'b11111111111111111101101111000101;
assign LUT_2[46611] = 32'b11111111111111111010100111011110;
assign LUT_2[46612] = 32'b11111111111111110011010011110001;
assign LUT_2[46613] = 32'b11111111111111110000001100001010;
assign LUT_2[46614] = 32'b11111111111111111010001100101101;
assign LUT_2[46615] = 32'b11111111111111110111000101000110;
assign LUT_2[46616] = 32'b11111111111111110001100111100110;
assign LUT_2[46617] = 32'b11111111111111101110011111111111;
assign LUT_2[46618] = 32'b11111111111111111000100000100010;
assign LUT_2[46619] = 32'b11111111111111110101011000111011;
assign LUT_2[46620] = 32'b11111111111111101110000101001110;
assign LUT_2[46621] = 32'b11111111111111101010111101100111;
assign LUT_2[46622] = 32'b11111111111111110100111110001010;
assign LUT_2[46623] = 32'b11111111111111110001110110100011;
assign LUT_2[46624] = 32'b11111111111111111100101101101000;
assign LUT_2[46625] = 32'b11111111111111111001100110000001;
assign LUT_2[46626] = 32'b00000000000000000011100110100100;
assign LUT_2[46627] = 32'b00000000000000000000011110111101;
assign LUT_2[46628] = 32'b11111111111111111001001011010000;
assign LUT_2[46629] = 32'b11111111111111110110000011101001;
assign LUT_2[46630] = 32'b00000000000000000000000100001100;
assign LUT_2[46631] = 32'b11111111111111111100111100100101;
assign LUT_2[46632] = 32'b11111111111111110111011111000101;
assign LUT_2[46633] = 32'b11111111111111110100010111011110;
assign LUT_2[46634] = 32'b11111111111111111110011000000001;
assign LUT_2[46635] = 32'b11111111111111111011010000011010;
assign LUT_2[46636] = 32'b11111111111111110011111100101101;
assign LUT_2[46637] = 32'b11111111111111110000110101000110;
assign LUT_2[46638] = 32'b11111111111111111010110101101001;
assign LUT_2[46639] = 32'b11111111111111110111101110000010;
assign LUT_2[46640] = 32'b11111111111111110111010001110010;
assign LUT_2[46641] = 32'b11111111111111110100001010001011;
assign LUT_2[46642] = 32'b11111111111111111110001010101110;
assign LUT_2[46643] = 32'b11111111111111111011000011000111;
assign LUT_2[46644] = 32'b11111111111111110011101111011010;
assign LUT_2[46645] = 32'b11111111111111110000100111110011;
assign LUT_2[46646] = 32'b11111111111111111010101000010110;
assign LUT_2[46647] = 32'b11111111111111110111100000101111;
assign LUT_2[46648] = 32'b11111111111111110010000011001111;
assign LUT_2[46649] = 32'b11111111111111101110111011101000;
assign LUT_2[46650] = 32'b11111111111111111000111100001011;
assign LUT_2[46651] = 32'b11111111111111110101110100100100;
assign LUT_2[46652] = 32'b11111111111111101110100000110111;
assign LUT_2[46653] = 32'b11111111111111101011011001010000;
assign LUT_2[46654] = 32'b11111111111111110101011001110011;
assign LUT_2[46655] = 32'b11111111111111110010010010001100;
assign LUT_2[46656] = 32'b11111111111111110100011010100010;
assign LUT_2[46657] = 32'b11111111111111110001010010111011;
assign LUT_2[46658] = 32'b11111111111111111011010011011110;
assign LUT_2[46659] = 32'b11111111111111111000001011110111;
assign LUT_2[46660] = 32'b11111111111111110000111000001010;
assign LUT_2[46661] = 32'b11111111111111101101110000100011;
assign LUT_2[46662] = 32'b11111111111111110111110001000110;
assign LUT_2[46663] = 32'b11111111111111110100101001011111;
assign LUT_2[46664] = 32'b11111111111111101111001011111111;
assign LUT_2[46665] = 32'b11111111111111101100000100011000;
assign LUT_2[46666] = 32'b11111111111111110110000100111011;
assign LUT_2[46667] = 32'b11111111111111110010111101010100;
assign LUT_2[46668] = 32'b11111111111111101011101001100111;
assign LUT_2[46669] = 32'b11111111111111101000100010000000;
assign LUT_2[46670] = 32'b11111111111111110010100010100011;
assign LUT_2[46671] = 32'b11111111111111101111011010111100;
assign LUT_2[46672] = 32'b11111111111111101110111110101100;
assign LUT_2[46673] = 32'b11111111111111101011110111000101;
assign LUT_2[46674] = 32'b11111111111111110101110111101000;
assign LUT_2[46675] = 32'b11111111111111110010110000000001;
assign LUT_2[46676] = 32'b11111111111111101011011100010100;
assign LUT_2[46677] = 32'b11111111111111101000010100101101;
assign LUT_2[46678] = 32'b11111111111111110010010101010000;
assign LUT_2[46679] = 32'b11111111111111101111001101101001;
assign LUT_2[46680] = 32'b11111111111111101001110000001001;
assign LUT_2[46681] = 32'b11111111111111100110101000100010;
assign LUT_2[46682] = 32'b11111111111111110000101001000101;
assign LUT_2[46683] = 32'b11111111111111101101100001011110;
assign LUT_2[46684] = 32'b11111111111111100110001101110001;
assign LUT_2[46685] = 32'b11111111111111100011000110001010;
assign LUT_2[46686] = 32'b11111111111111101101000110101101;
assign LUT_2[46687] = 32'b11111111111111101001111111000110;
assign LUT_2[46688] = 32'b11111111111111110100110110001011;
assign LUT_2[46689] = 32'b11111111111111110001101110100100;
assign LUT_2[46690] = 32'b11111111111111111011101111000111;
assign LUT_2[46691] = 32'b11111111111111111000100111100000;
assign LUT_2[46692] = 32'b11111111111111110001010011110011;
assign LUT_2[46693] = 32'b11111111111111101110001100001100;
assign LUT_2[46694] = 32'b11111111111111111000001100101111;
assign LUT_2[46695] = 32'b11111111111111110101000101001000;
assign LUT_2[46696] = 32'b11111111111111101111100111101000;
assign LUT_2[46697] = 32'b11111111111111101100100000000001;
assign LUT_2[46698] = 32'b11111111111111110110100000100100;
assign LUT_2[46699] = 32'b11111111111111110011011000111101;
assign LUT_2[46700] = 32'b11111111111111101100000101010000;
assign LUT_2[46701] = 32'b11111111111111101000111101101001;
assign LUT_2[46702] = 32'b11111111111111110010111110001100;
assign LUT_2[46703] = 32'b11111111111111101111110110100101;
assign LUT_2[46704] = 32'b11111111111111101111011010010101;
assign LUT_2[46705] = 32'b11111111111111101100010010101110;
assign LUT_2[46706] = 32'b11111111111111110110010011010001;
assign LUT_2[46707] = 32'b11111111111111110011001011101010;
assign LUT_2[46708] = 32'b11111111111111101011110111111101;
assign LUT_2[46709] = 32'b11111111111111101000110000010110;
assign LUT_2[46710] = 32'b11111111111111110010110000111001;
assign LUT_2[46711] = 32'b11111111111111101111101001010010;
assign LUT_2[46712] = 32'b11111111111111101010001011110010;
assign LUT_2[46713] = 32'b11111111111111100111000100001011;
assign LUT_2[46714] = 32'b11111111111111110001000100101110;
assign LUT_2[46715] = 32'b11111111111111101101111101000111;
assign LUT_2[46716] = 32'b11111111111111100110101001011010;
assign LUT_2[46717] = 32'b11111111111111100011100001110011;
assign LUT_2[46718] = 32'b11111111111111101101100010010110;
assign LUT_2[46719] = 32'b11111111111111101010011010101111;
assign LUT_2[46720] = 32'b00000000000000000000100110001110;
assign LUT_2[46721] = 32'b11111111111111111101011110100111;
assign LUT_2[46722] = 32'b00000000000000000111011111001010;
assign LUT_2[46723] = 32'b00000000000000000100010111100011;
assign LUT_2[46724] = 32'b11111111111111111101000011110110;
assign LUT_2[46725] = 32'b11111111111111111001111100001111;
assign LUT_2[46726] = 32'b00000000000000000011111100110010;
assign LUT_2[46727] = 32'b00000000000000000000110101001011;
assign LUT_2[46728] = 32'b11111111111111111011010111101011;
assign LUT_2[46729] = 32'b11111111111111111000010000000100;
assign LUT_2[46730] = 32'b00000000000000000010010000100111;
assign LUT_2[46731] = 32'b11111111111111111111001001000000;
assign LUT_2[46732] = 32'b11111111111111110111110101010011;
assign LUT_2[46733] = 32'b11111111111111110100101101101100;
assign LUT_2[46734] = 32'b11111111111111111110101110001111;
assign LUT_2[46735] = 32'b11111111111111111011100110101000;
assign LUT_2[46736] = 32'b11111111111111111011001010011000;
assign LUT_2[46737] = 32'b11111111111111111000000010110001;
assign LUT_2[46738] = 32'b00000000000000000010000011010100;
assign LUT_2[46739] = 32'b11111111111111111110111011101101;
assign LUT_2[46740] = 32'b11111111111111110111101000000000;
assign LUT_2[46741] = 32'b11111111111111110100100000011001;
assign LUT_2[46742] = 32'b11111111111111111110100000111100;
assign LUT_2[46743] = 32'b11111111111111111011011001010101;
assign LUT_2[46744] = 32'b11111111111111110101111011110101;
assign LUT_2[46745] = 32'b11111111111111110010110100001110;
assign LUT_2[46746] = 32'b11111111111111111100110100110001;
assign LUT_2[46747] = 32'b11111111111111111001101101001010;
assign LUT_2[46748] = 32'b11111111111111110010011001011101;
assign LUT_2[46749] = 32'b11111111111111101111010001110110;
assign LUT_2[46750] = 32'b11111111111111111001010010011001;
assign LUT_2[46751] = 32'b11111111111111110110001010110010;
assign LUT_2[46752] = 32'b00000000000000000001000001110111;
assign LUT_2[46753] = 32'b11111111111111111101111010010000;
assign LUT_2[46754] = 32'b00000000000000000111111010110011;
assign LUT_2[46755] = 32'b00000000000000000100110011001100;
assign LUT_2[46756] = 32'b11111111111111111101011111011111;
assign LUT_2[46757] = 32'b11111111111111111010010111111000;
assign LUT_2[46758] = 32'b00000000000000000100011000011011;
assign LUT_2[46759] = 32'b00000000000000000001010000110100;
assign LUT_2[46760] = 32'b11111111111111111011110011010100;
assign LUT_2[46761] = 32'b11111111111111111000101011101101;
assign LUT_2[46762] = 32'b00000000000000000010101100010000;
assign LUT_2[46763] = 32'b11111111111111111111100100101001;
assign LUT_2[46764] = 32'b11111111111111111000010000111100;
assign LUT_2[46765] = 32'b11111111111111110101001001010101;
assign LUT_2[46766] = 32'b11111111111111111111001001111000;
assign LUT_2[46767] = 32'b11111111111111111100000010010001;
assign LUT_2[46768] = 32'b11111111111111111011100110000001;
assign LUT_2[46769] = 32'b11111111111111111000011110011010;
assign LUT_2[46770] = 32'b00000000000000000010011110111101;
assign LUT_2[46771] = 32'b11111111111111111111010111010110;
assign LUT_2[46772] = 32'b11111111111111111000000011101001;
assign LUT_2[46773] = 32'b11111111111111110100111100000010;
assign LUT_2[46774] = 32'b11111111111111111110111100100101;
assign LUT_2[46775] = 32'b11111111111111111011110100111110;
assign LUT_2[46776] = 32'b11111111111111110110010111011110;
assign LUT_2[46777] = 32'b11111111111111110011001111110111;
assign LUT_2[46778] = 32'b11111111111111111101010000011010;
assign LUT_2[46779] = 32'b11111111111111111010001000110011;
assign LUT_2[46780] = 32'b11111111111111110010110101000110;
assign LUT_2[46781] = 32'b11111111111111101111101101011111;
assign LUT_2[46782] = 32'b11111111111111111001101110000010;
assign LUT_2[46783] = 32'b11111111111111110110100110011011;
assign LUT_2[46784] = 32'b11111111111111111000101110110001;
assign LUT_2[46785] = 32'b11111111111111110101100111001010;
assign LUT_2[46786] = 32'b11111111111111111111100111101101;
assign LUT_2[46787] = 32'b11111111111111111100100000000110;
assign LUT_2[46788] = 32'b11111111111111110101001100011001;
assign LUT_2[46789] = 32'b11111111111111110010000100110010;
assign LUT_2[46790] = 32'b11111111111111111100000101010101;
assign LUT_2[46791] = 32'b11111111111111111000111101101110;
assign LUT_2[46792] = 32'b11111111111111110011100000001110;
assign LUT_2[46793] = 32'b11111111111111110000011000100111;
assign LUT_2[46794] = 32'b11111111111111111010011001001010;
assign LUT_2[46795] = 32'b11111111111111110111010001100011;
assign LUT_2[46796] = 32'b11111111111111101111111101110110;
assign LUT_2[46797] = 32'b11111111111111101100110110001111;
assign LUT_2[46798] = 32'b11111111111111110110110110110010;
assign LUT_2[46799] = 32'b11111111111111110011101111001011;
assign LUT_2[46800] = 32'b11111111111111110011010010111011;
assign LUT_2[46801] = 32'b11111111111111110000001011010100;
assign LUT_2[46802] = 32'b11111111111111111010001011110111;
assign LUT_2[46803] = 32'b11111111111111110111000100010000;
assign LUT_2[46804] = 32'b11111111111111101111110000100011;
assign LUT_2[46805] = 32'b11111111111111101100101000111100;
assign LUT_2[46806] = 32'b11111111111111110110101001011111;
assign LUT_2[46807] = 32'b11111111111111110011100001111000;
assign LUT_2[46808] = 32'b11111111111111101110000100011000;
assign LUT_2[46809] = 32'b11111111111111101010111100110001;
assign LUT_2[46810] = 32'b11111111111111110100111101010100;
assign LUT_2[46811] = 32'b11111111111111110001110101101101;
assign LUT_2[46812] = 32'b11111111111111101010100010000000;
assign LUT_2[46813] = 32'b11111111111111100111011010011001;
assign LUT_2[46814] = 32'b11111111111111110001011010111100;
assign LUT_2[46815] = 32'b11111111111111101110010011010101;
assign LUT_2[46816] = 32'b11111111111111111001001010011010;
assign LUT_2[46817] = 32'b11111111111111110110000010110011;
assign LUT_2[46818] = 32'b00000000000000000000000011010110;
assign LUT_2[46819] = 32'b11111111111111111100111011101111;
assign LUT_2[46820] = 32'b11111111111111110101101000000010;
assign LUT_2[46821] = 32'b11111111111111110010100000011011;
assign LUT_2[46822] = 32'b11111111111111111100100000111110;
assign LUT_2[46823] = 32'b11111111111111111001011001010111;
assign LUT_2[46824] = 32'b11111111111111110011111011110111;
assign LUT_2[46825] = 32'b11111111111111110000110100010000;
assign LUT_2[46826] = 32'b11111111111111111010110100110011;
assign LUT_2[46827] = 32'b11111111111111110111101101001100;
assign LUT_2[46828] = 32'b11111111111111110000011001011111;
assign LUT_2[46829] = 32'b11111111111111101101010001111000;
assign LUT_2[46830] = 32'b11111111111111110111010010011011;
assign LUT_2[46831] = 32'b11111111111111110100001010110100;
assign LUT_2[46832] = 32'b11111111111111110011101110100100;
assign LUT_2[46833] = 32'b11111111111111110000100110111101;
assign LUT_2[46834] = 32'b11111111111111111010100111100000;
assign LUT_2[46835] = 32'b11111111111111110111011111111001;
assign LUT_2[46836] = 32'b11111111111111110000001100001100;
assign LUT_2[46837] = 32'b11111111111111101101000100100101;
assign LUT_2[46838] = 32'b11111111111111110111000101001000;
assign LUT_2[46839] = 32'b11111111111111110011111101100001;
assign LUT_2[46840] = 32'b11111111111111101110100000000001;
assign LUT_2[46841] = 32'b11111111111111101011011000011010;
assign LUT_2[46842] = 32'b11111111111111110101011000111101;
assign LUT_2[46843] = 32'b11111111111111110010010001010110;
assign LUT_2[46844] = 32'b11111111111111101010111101101001;
assign LUT_2[46845] = 32'b11111111111111100111110110000010;
assign LUT_2[46846] = 32'b11111111111111110001110110100101;
assign LUT_2[46847] = 32'b11111111111111101110101110111110;
assign LUT_2[46848] = 32'b00000000000000000000010000100101;
assign LUT_2[46849] = 32'b11111111111111111101001000111110;
assign LUT_2[46850] = 32'b00000000000000000111001001100001;
assign LUT_2[46851] = 32'b00000000000000000100000001111010;
assign LUT_2[46852] = 32'b11111111111111111100101110001101;
assign LUT_2[46853] = 32'b11111111111111111001100110100110;
assign LUT_2[46854] = 32'b00000000000000000011100111001001;
assign LUT_2[46855] = 32'b00000000000000000000011111100010;
assign LUT_2[46856] = 32'b11111111111111111011000010000010;
assign LUT_2[46857] = 32'b11111111111111110111111010011011;
assign LUT_2[46858] = 32'b00000000000000000001111010111110;
assign LUT_2[46859] = 32'b11111111111111111110110011010111;
assign LUT_2[46860] = 32'b11111111111111110111011111101010;
assign LUT_2[46861] = 32'b11111111111111110100011000000011;
assign LUT_2[46862] = 32'b11111111111111111110011000100110;
assign LUT_2[46863] = 32'b11111111111111111011010000111111;
assign LUT_2[46864] = 32'b11111111111111111010110100101111;
assign LUT_2[46865] = 32'b11111111111111110111101101001000;
assign LUT_2[46866] = 32'b00000000000000000001101101101011;
assign LUT_2[46867] = 32'b11111111111111111110100110000100;
assign LUT_2[46868] = 32'b11111111111111110111010010010111;
assign LUT_2[46869] = 32'b11111111111111110100001010110000;
assign LUT_2[46870] = 32'b11111111111111111110001011010011;
assign LUT_2[46871] = 32'b11111111111111111011000011101100;
assign LUT_2[46872] = 32'b11111111111111110101100110001100;
assign LUT_2[46873] = 32'b11111111111111110010011110100101;
assign LUT_2[46874] = 32'b11111111111111111100011111001000;
assign LUT_2[46875] = 32'b11111111111111111001010111100001;
assign LUT_2[46876] = 32'b11111111111111110010000011110100;
assign LUT_2[46877] = 32'b11111111111111101110111100001101;
assign LUT_2[46878] = 32'b11111111111111111000111100110000;
assign LUT_2[46879] = 32'b11111111111111110101110101001001;
assign LUT_2[46880] = 32'b00000000000000000000101100001110;
assign LUT_2[46881] = 32'b11111111111111111101100100100111;
assign LUT_2[46882] = 32'b00000000000000000111100101001010;
assign LUT_2[46883] = 32'b00000000000000000100011101100011;
assign LUT_2[46884] = 32'b11111111111111111101001001110110;
assign LUT_2[46885] = 32'b11111111111111111010000010001111;
assign LUT_2[46886] = 32'b00000000000000000100000010110010;
assign LUT_2[46887] = 32'b00000000000000000000111011001011;
assign LUT_2[46888] = 32'b11111111111111111011011101101011;
assign LUT_2[46889] = 32'b11111111111111111000010110000100;
assign LUT_2[46890] = 32'b00000000000000000010010110100111;
assign LUT_2[46891] = 32'b11111111111111111111001111000000;
assign LUT_2[46892] = 32'b11111111111111110111111011010011;
assign LUT_2[46893] = 32'b11111111111111110100110011101100;
assign LUT_2[46894] = 32'b11111111111111111110110100001111;
assign LUT_2[46895] = 32'b11111111111111111011101100101000;
assign LUT_2[46896] = 32'b11111111111111111011010000011000;
assign LUT_2[46897] = 32'b11111111111111111000001000110001;
assign LUT_2[46898] = 32'b00000000000000000010001001010100;
assign LUT_2[46899] = 32'b11111111111111111111000001101101;
assign LUT_2[46900] = 32'b11111111111111110111101110000000;
assign LUT_2[46901] = 32'b11111111111111110100100110011001;
assign LUT_2[46902] = 32'b11111111111111111110100110111100;
assign LUT_2[46903] = 32'b11111111111111111011011111010101;
assign LUT_2[46904] = 32'b11111111111111110110000001110101;
assign LUT_2[46905] = 32'b11111111111111110010111010001110;
assign LUT_2[46906] = 32'b11111111111111111100111010110001;
assign LUT_2[46907] = 32'b11111111111111111001110011001010;
assign LUT_2[46908] = 32'b11111111111111110010011111011101;
assign LUT_2[46909] = 32'b11111111111111101111010111110110;
assign LUT_2[46910] = 32'b11111111111111111001011000011001;
assign LUT_2[46911] = 32'b11111111111111110110010000110010;
assign LUT_2[46912] = 32'b11111111111111111000011001001000;
assign LUT_2[46913] = 32'b11111111111111110101010001100001;
assign LUT_2[46914] = 32'b11111111111111111111010010000100;
assign LUT_2[46915] = 32'b11111111111111111100001010011101;
assign LUT_2[46916] = 32'b11111111111111110100110110110000;
assign LUT_2[46917] = 32'b11111111111111110001101111001001;
assign LUT_2[46918] = 32'b11111111111111111011101111101100;
assign LUT_2[46919] = 32'b11111111111111111000101000000101;
assign LUT_2[46920] = 32'b11111111111111110011001010100101;
assign LUT_2[46921] = 32'b11111111111111110000000010111110;
assign LUT_2[46922] = 32'b11111111111111111010000011100001;
assign LUT_2[46923] = 32'b11111111111111110110111011111010;
assign LUT_2[46924] = 32'b11111111111111101111101000001101;
assign LUT_2[46925] = 32'b11111111111111101100100000100110;
assign LUT_2[46926] = 32'b11111111111111110110100001001001;
assign LUT_2[46927] = 32'b11111111111111110011011001100010;
assign LUT_2[46928] = 32'b11111111111111110010111101010010;
assign LUT_2[46929] = 32'b11111111111111101111110101101011;
assign LUT_2[46930] = 32'b11111111111111111001110110001110;
assign LUT_2[46931] = 32'b11111111111111110110101110100111;
assign LUT_2[46932] = 32'b11111111111111101111011010111010;
assign LUT_2[46933] = 32'b11111111111111101100010011010011;
assign LUT_2[46934] = 32'b11111111111111110110010011110110;
assign LUT_2[46935] = 32'b11111111111111110011001100001111;
assign LUT_2[46936] = 32'b11111111111111101101101110101111;
assign LUT_2[46937] = 32'b11111111111111101010100111001000;
assign LUT_2[46938] = 32'b11111111111111110100100111101011;
assign LUT_2[46939] = 32'b11111111111111110001100000000100;
assign LUT_2[46940] = 32'b11111111111111101010001100010111;
assign LUT_2[46941] = 32'b11111111111111100111000100110000;
assign LUT_2[46942] = 32'b11111111111111110001000101010011;
assign LUT_2[46943] = 32'b11111111111111101101111101101100;
assign LUT_2[46944] = 32'b11111111111111111000110100110001;
assign LUT_2[46945] = 32'b11111111111111110101101101001010;
assign LUT_2[46946] = 32'b11111111111111111111101101101101;
assign LUT_2[46947] = 32'b11111111111111111100100110000110;
assign LUT_2[46948] = 32'b11111111111111110101010010011001;
assign LUT_2[46949] = 32'b11111111111111110010001010110010;
assign LUT_2[46950] = 32'b11111111111111111100001011010101;
assign LUT_2[46951] = 32'b11111111111111111001000011101110;
assign LUT_2[46952] = 32'b11111111111111110011100110001110;
assign LUT_2[46953] = 32'b11111111111111110000011110100111;
assign LUT_2[46954] = 32'b11111111111111111010011111001010;
assign LUT_2[46955] = 32'b11111111111111110111010111100011;
assign LUT_2[46956] = 32'b11111111111111110000000011110110;
assign LUT_2[46957] = 32'b11111111111111101100111100001111;
assign LUT_2[46958] = 32'b11111111111111110110111100110010;
assign LUT_2[46959] = 32'b11111111111111110011110101001011;
assign LUT_2[46960] = 32'b11111111111111110011011000111011;
assign LUT_2[46961] = 32'b11111111111111110000010001010100;
assign LUT_2[46962] = 32'b11111111111111111010010001110111;
assign LUT_2[46963] = 32'b11111111111111110111001010010000;
assign LUT_2[46964] = 32'b11111111111111101111110110100011;
assign LUT_2[46965] = 32'b11111111111111101100101110111100;
assign LUT_2[46966] = 32'b11111111111111110110101111011111;
assign LUT_2[46967] = 32'b11111111111111110011100111111000;
assign LUT_2[46968] = 32'b11111111111111101110001010011000;
assign LUT_2[46969] = 32'b11111111111111101011000010110001;
assign LUT_2[46970] = 32'b11111111111111110101000011010100;
assign LUT_2[46971] = 32'b11111111111111110001111011101101;
assign LUT_2[46972] = 32'b11111111111111101010101000000000;
assign LUT_2[46973] = 32'b11111111111111100111100000011001;
assign LUT_2[46974] = 32'b11111111111111110001100000111100;
assign LUT_2[46975] = 32'b11111111111111101110011001010101;
assign LUT_2[46976] = 32'b00000000000000000100100100110100;
assign LUT_2[46977] = 32'b00000000000000000001011101001101;
assign LUT_2[46978] = 32'b00000000000000001011011101110000;
assign LUT_2[46979] = 32'b00000000000000001000010110001001;
assign LUT_2[46980] = 32'b00000000000000000001000010011100;
assign LUT_2[46981] = 32'b11111111111111111101111010110101;
assign LUT_2[46982] = 32'b00000000000000000111111011011000;
assign LUT_2[46983] = 32'b00000000000000000100110011110001;
assign LUT_2[46984] = 32'b11111111111111111111010110010001;
assign LUT_2[46985] = 32'b11111111111111111100001110101010;
assign LUT_2[46986] = 32'b00000000000000000110001111001101;
assign LUT_2[46987] = 32'b00000000000000000011000111100110;
assign LUT_2[46988] = 32'b11111111111111111011110011111001;
assign LUT_2[46989] = 32'b11111111111111111000101100010010;
assign LUT_2[46990] = 32'b00000000000000000010101100110101;
assign LUT_2[46991] = 32'b11111111111111111111100101001110;
assign LUT_2[46992] = 32'b11111111111111111111001000111110;
assign LUT_2[46993] = 32'b11111111111111111100000001010111;
assign LUT_2[46994] = 32'b00000000000000000110000001111010;
assign LUT_2[46995] = 32'b00000000000000000010111010010011;
assign LUT_2[46996] = 32'b11111111111111111011100110100110;
assign LUT_2[46997] = 32'b11111111111111111000011110111111;
assign LUT_2[46998] = 32'b00000000000000000010011111100010;
assign LUT_2[46999] = 32'b11111111111111111111010111111011;
assign LUT_2[47000] = 32'b11111111111111111001111010011011;
assign LUT_2[47001] = 32'b11111111111111110110110010110100;
assign LUT_2[47002] = 32'b00000000000000000000110011010111;
assign LUT_2[47003] = 32'b11111111111111111101101011110000;
assign LUT_2[47004] = 32'b11111111111111110110011000000011;
assign LUT_2[47005] = 32'b11111111111111110011010000011100;
assign LUT_2[47006] = 32'b11111111111111111101010000111111;
assign LUT_2[47007] = 32'b11111111111111111010001001011000;
assign LUT_2[47008] = 32'b00000000000000000101000000011101;
assign LUT_2[47009] = 32'b00000000000000000001111000110110;
assign LUT_2[47010] = 32'b00000000000000001011111001011001;
assign LUT_2[47011] = 32'b00000000000000001000110001110010;
assign LUT_2[47012] = 32'b00000000000000000001011110000101;
assign LUT_2[47013] = 32'b11111111111111111110010110011110;
assign LUT_2[47014] = 32'b00000000000000001000010111000001;
assign LUT_2[47015] = 32'b00000000000000000101001111011010;
assign LUT_2[47016] = 32'b11111111111111111111110001111010;
assign LUT_2[47017] = 32'b11111111111111111100101010010011;
assign LUT_2[47018] = 32'b00000000000000000110101010110110;
assign LUT_2[47019] = 32'b00000000000000000011100011001111;
assign LUT_2[47020] = 32'b11111111111111111100001111100010;
assign LUT_2[47021] = 32'b11111111111111111001000111111011;
assign LUT_2[47022] = 32'b00000000000000000011001000011110;
assign LUT_2[47023] = 32'b00000000000000000000000000110111;
assign LUT_2[47024] = 32'b11111111111111111111100100100111;
assign LUT_2[47025] = 32'b11111111111111111100011101000000;
assign LUT_2[47026] = 32'b00000000000000000110011101100011;
assign LUT_2[47027] = 32'b00000000000000000011010101111100;
assign LUT_2[47028] = 32'b11111111111111111100000010001111;
assign LUT_2[47029] = 32'b11111111111111111000111010101000;
assign LUT_2[47030] = 32'b00000000000000000010111011001011;
assign LUT_2[47031] = 32'b11111111111111111111110011100100;
assign LUT_2[47032] = 32'b11111111111111111010010110000100;
assign LUT_2[47033] = 32'b11111111111111110111001110011101;
assign LUT_2[47034] = 32'b00000000000000000001001111000000;
assign LUT_2[47035] = 32'b11111111111111111110000111011001;
assign LUT_2[47036] = 32'b11111111111111110110110011101100;
assign LUT_2[47037] = 32'b11111111111111110011101100000101;
assign LUT_2[47038] = 32'b11111111111111111101101100101000;
assign LUT_2[47039] = 32'b11111111111111111010100101000001;
assign LUT_2[47040] = 32'b11111111111111111100101101010111;
assign LUT_2[47041] = 32'b11111111111111111001100101110000;
assign LUT_2[47042] = 32'b00000000000000000011100110010011;
assign LUT_2[47043] = 32'b00000000000000000000011110101100;
assign LUT_2[47044] = 32'b11111111111111111001001010111111;
assign LUT_2[47045] = 32'b11111111111111110110000011011000;
assign LUT_2[47046] = 32'b00000000000000000000000011111011;
assign LUT_2[47047] = 32'b11111111111111111100111100010100;
assign LUT_2[47048] = 32'b11111111111111110111011110110100;
assign LUT_2[47049] = 32'b11111111111111110100010111001101;
assign LUT_2[47050] = 32'b11111111111111111110010111110000;
assign LUT_2[47051] = 32'b11111111111111111011010000001001;
assign LUT_2[47052] = 32'b11111111111111110011111100011100;
assign LUT_2[47053] = 32'b11111111111111110000110100110101;
assign LUT_2[47054] = 32'b11111111111111111010110101011000;
assign LUT_2[47055] = 32'b11111111111111110111101101110001;
assign LUT_2[47056] = 32'b11111111111111110111010001100001;
assign LUT_2[47057] = 32'b11111111111111110100001001111010;
assign LUT_2[47058] = 32'b11111111111111111110001010011101;
assign LUT_2[47059] = 32'b11111111111111111011000010110110;
assign LUT_2[47060] = 32'b11111111111111110011101111001001;
assign LUT_2[47061] = 32'b11111111111111110000100111100010;
assign LUT_2[47062] = 32'b11111111111111111010101000000101;
assign LUT_2[47063] = 32'b11111111111111110111100000011110;
assign LUT_2[47064] = 32'b11111111111111110010000010111110;
assign LUT_2[47065] = 32'b11111111111111101110111011010111;
assign LUT_2[47066] = 32'b11111111111111111000111011111010;
assign LUT_2[47067] = 32'b11111111111111110101110100010011;
assign LUT_2[47068] = 32'b11111111111111101110100000100110;
assign LUT_2[47069] = 32'b11111111111111101011011000111111;
assign LUT_2[47070] = 32'b11111111111111110101011001100010;
assign LUT_2[47071] = 32'b11111111111111110010010001111011;
assign LUT_2[47072] = 32'b11111111111111111101001001000000;
assign LUT_2[47073] = 32'b11111111111111111010000001011001;
assign LUT_2[47074] = 32'b00000000000000000100000001111100;
assign LUT_2[47075] = 32'b00000000000000000000111010010101;
assign LUT_2[47076] = 32'b11111111111111111001100110101000;
assign LUT_2[47077] = 32'b11111111111111110110011111000001;
assign LUT_2[47078] = 32'b00000000000000000000011111100100;
assign LUT_2[47079] = 32'b11111111111111111101010111111101;
assign LUT_2[47080] = 32'b11111111111111110111111010011101;
assign LUT_2[47081] = 32'b11111111111111110100110010110110;
assign LUT_2[47082] = 32'b11111111111111111110110011011001;
assign LUT_2[47083] = 32'b11111111111111111011101011110010;
assign LUT_2[47084] = 32'b11111111111111110100011000000101;
assign LUT_2[47085] = 32'b11111111111111110001010000011110;
assign LUT_2[47086] = 32'b11111111111111111011010001000001;
assign LUT_2[47087] = 32'b11111111111111111000001001011010;
assign LUT_2[47088] = 32'b11111111111111110111101101001010;
assign LUT_2[47089] = 32'b11111111111111110100100101100011;
assign LUT_2[47090] = 32'b11111111111111111110100110000110;
assign LUT_2[47091] = 32'b11111111111111111011011110011111;
assign LUT_2[47092] = 32'b11111111111111110100001010110010;
assign LUT_2[47093] = 32'b11111111111111110001000011001011;
assign LUT_2[47094] = 32'b11111111111111111011000011101110;
assign LUT_2[47095] = 32'b11111111111111110111111100000111;
assign LUT_2[47096] = 32'b11111111111111110010011110100111;
assign LUT_2[47097] = 32'b11111111111111101111010111000000;
assign LUT_2[47098] = 32'b11111111111111111001010111100011;
assign LUT_2[47099] = 32'b11111111111111110110001111111100;
assign LUT_2[47100] = 32'b11111111111111101110111100001111;
assign LUT_2[47101] = 32'b11111111111111101011110100101000;
assign LUT_2[47102] = 32'b11111111111111110101110101001011;
assign LUT_2[47103] = 32'b11111111111111110010101101100100;
assign LUT_2[47104] = 32'b11111111111111101100101010000100;
assign LUT_2[47105] = 32'b11111111111111101001100010011101;
assign LUT_2[47106] = 32'b11111111111111110011100011000000;
assign LUT_2[47107] = 32'b11111111111111110000011011011001;
assign LUT_2[47108] = 32'b11111111111111101001000111101100;
assign LUT_2[47109] = 32'b11111111111111100110000000000101;
assign LUT_2[47110] = 32'b11111111111111110000000000101000;
assign LUT_2[47111] = 32'b11111111111111101100111001000001;
assign LUT_2[47112] = 32'b11111111111111100111011011100001;
assign LUT_2[47113] = 32'b11111111111111100100010011111010;
assign LUT_2[47114] = 32'b11111111111111101110010100011101;
assign LUT_2[47115] = 32'b11111111111111101011001100110110;
assign LUT_2[47116] = 32'b11111111111111100011111001001001;
assign LUT_2[47117] = 32'b11111111111111100000110001100010;
assign LUT_2[47118] = 32'b11111111111111101010110010000101;
assign LUT_2[47119] = 32'b11111111111111100111101010011110;
assign LUT_2[47120] = 32'b11111111111111100111001110001110;
assign LUT_2[47121] = 32'b11111111111111100100000110100111;
assign LUT_2[47122] = 32'b11111111111111101110000111001010;
assign LUT_2[47123] = 32'b11111111111111101010111111100011;
assign LUT_2[47124] = 32'b11111111111111100011101011110110;
assign LUT_2[47125] = 32'b11111111111111100000100100001111;
assign LUT_2[47126] = 32'b11111111111111101010100100110010;
assign LUT_2[47127] = 32'b11111111111111100111011101001011;
assign LUT_2[47128] = 32'b11111111111111100001111111101011;
assign LUT_2[47129] = 32'b11111111111111011110111000000100;
assign LUT_2[47130] = 32'b11111111111111101000111000100111;
assign LUT_2[47131] = 32'b11111111111111100101110001000000;
assign LUT_2[47132] = 32'b11111111111111011110011101010011;
assign LUT_2[47133] = 32'b11111111111111011011010101101100;
assign LUT_2[47134] = 32'b11111111111111100101010110001111;
assign LUT_2[47135] = 32'b11111111111111100010001110101000;
assign LUT_2[47136] = 32'b11111111111111101101000101101101;
assign LUT_2[47137] = 32'b11111111111111101001111110000110;
assign LUT_2[47138] = 32'b11111111111111110011111110101001;
assign LUT_2[47139] = 32'b11111111111111110000110111000010;
assign LUT_2[47140] = 32'b11111111111111101001100011010101;
assign LUT_2[47141] = 32'b11111111111111100110011011101110;
assign LUT_2[47142] = 32'b11111111111111110000011100010001;
assign LUT_2[47143] = 32'b11111111111111101101010100101010;
assign LUT_2[47144] = 32'b11111111111111100111110111001010;
assign LUT_2[47145] = 32'b11111111111111100100101111100011;
assign LUT_2[47146] = 32'b11111111111111101110110000000110;
assign LUT_2[47147] = 32'b11111111111111101011101000011111;
assign LUT_2[47148] = 32'b11111111111111100100010100110010;
assign LUT_2[47149] = 32'b11111111111111100001001101001011;
assign LUT_2[47150] = 32'b11111111111111101011001101101110;
assign LUT_2[47151] = 32'b11111111111111101000000110000111;
assign LUT_2[47152] = 32'b11111111111111100111101001110111;
assign LUT_2[47153] = 32'b11111111111111100100100010010000;
assign LUT_2[47154] = 32'b11111111111111101110100010110011;
assign LUT_2[47155] = 32'b11111111111111101011011011001100;
assign LUT_2[47156] = 32'b11111111111111100100000111011111;
assign LUT_2[47157] = 32'b11111111111111100000111111111000;
assign LUT_2[47158] = 32'b11111111111111101011000000011011;
assign LUT_2[47159] = 32'b11111111111111100111111000110100;
assign LUT_2[47160] = 32'b11111111111111100010011011010100;
assign LUT_2[47161] = 32'b11111111111111011111010011101101;
assign LUT_2[47162] = 32'b11111111111111101001010100010000;
assign LUT_2[47163] = 32'b11111111111111100110001100101001;
assign LUT_2[47164] = 32'b11111111111111011110111000111100;
assign LUT_2[47165] = 32'b11111111111111011011110001010101;
assign LUT_2[47166] = 32'b11111111111111100101110001111000;
assign LUT_2[47167] = 32'b11111111111111100010101010010001;
assign LUT_2[47168] = 32'b11111111111111100100110010100111;
assign LUT_2[47169] = 32'b11111111111111100001101011000000;
assign LUT_2[47170] = 32'b11111111111111101011101011100011;
assign LUT_2[47171] = 32'b11111111111111101000100011111100;
assign LUT_2[47172] = 32'b11111111111111100001010000001111;
assign LUT_2[47173] = 32'b11111111111111011110001000101000;
assign LUT_2[47174] = 32'b11111111111111101000001001001011;
assign LUT_2[47175] = 32'b11111111111111100101000001100100;
assign LUT_2[47176] = 32'b11111111111111011111100100000100;
assign LUT_2[47177] = 32'b11111111111111011100011100011101;
assign LUT_2[47178] = 32'b11111111111111100110011101000000;
assign LUT_2[47179] = 32'b11111111111111100011010101011001;
assign LUT_2[47180] = 32'b11111111111111011100000001101100;
assign LUT_2[47181] = 32'b11111111111111011000111010000101;
assign LUT_2[47182] = 32'b11111111111111100010111010101000;
assign LUT_2[47183] = 32'b11111111111111011111110011000001;
assign LUT_2[47184] = 32'b11111111111111011111010110110001;
assign LUT_2[47185] = 32'b11111111111111011100001111001010;
assign LUT_2[47186] = 32'b11111111111111100110001111101101;
assign LUT_2[47187] = 32'b11111111111111100011001000000110;
assign LUT_2[47188] = 32'b11111111111111011011110100011001;
assign LUT_2[47189] = 32'b11111111111111011000101100110010;
assign LUT_2[47190] = 32'b11111111111111100010101101010101;
assign LUT_2[47191] = 32'b11111111111111011111100101101110;
assign LUT_2[47192] = 32'b11111111111111011010001000001110;
assign LUT_2[47193] = 32'b11111111111111010111000000100111;
assign LUT_2[47194] = 32'b11111111111111100001000001001010;
assign LUT_2[47195] = 32'b11111111111111011101111001100011;
assign LUT_2[47196] = 32'b11111111111111010110100101110110;
assign LUT_2[47197] = 32'b11111111111111010011011110001111;
assign LUT_2[47198] = 32'b11111111111111011101011110110010;
assign LUT_2[47199] = 32'b11111111111111011010010111001011;
assign LUT_2[47200] = 32'b11111111111111100101001110010000;
assign LUT_2[47201] = 32'b11111111111111100010000110101001;
assign LUT_2[47202] = 32'b11111111111111101100000111001100;
assign LUT_2[47203] = 32'b11111111111111101000111111100101;
assign LUT_2[47204] = 32'b11111111111111100001101011111000;
assign LUT_2[47205] = 32'b11111111111111011110100100010001;
assign LUT_2[47206] = 32'b11111111111111101000100100110100;
assign LUT_2[47207] = 32'b11111111111111100101011101001101;
assign LUT_2[47208] = 32'b11111111111111011111111111101101;
assign LUT_2[47209] = 32'b11111111111111011100111000000110;
assign LUT_2[47210] = 32'b11111111111111100110111000101001;
assign LUT_2[47211] = 32'b11111111111111100011110001000010;
assign LUT_2[47212] = 32'b11111111111111011100011101010101;
assign LUT_2[47213] = 32'b11111111111111011001010101101110;
assign LUT_2[47214] = 32'b11111111111111100011010110010001;
assign LUT_2[47215] = 32'b11111111111111100000001110101010;
assign LUT_2[47216] = 32'b11111111111111011111110010011010;
assign LUT_2[47217] = 32'b11111111111111011100101010110011;
assign LUT_2[47218] = 32'b11111111111111100110101011010110;
assign LUT_2[47219] = 32'b11111111111111100011100011101111;
assign LUT_2[47220] = 32'b11111111111111011100010000000010;
assign LUT_2[47221] = 32'b11111111111111011001001000011011;
assign LUT_2[47222] = 32'b11111111111111100011001000111110;
assign LUT_2[47223] = 32'b11111111111111100000000001010111;
assign LUT_2[47224] = 32'b11111111111111011010100011110111;
assign LUT_2[47225] = 32'b11111111111111010111011100010000;
assign LUT_2[47226] = 32'b11111111111111100001011100110011;
assign LUT_2[47227] = 32'b11111111111111011110010101001100;
assign LUT_2[47228] = 32'b11111111111111010111000001011111;
assign LUT_2[47229] = 32'b11111111111111010011111001111000;
assign LUT_2[47230] = 32'b11111111111111011101111010011011;
assign LUT_2[47231] = 32'b11111111111111011010110010110100;
assign LUT_2[47232] = 32'b11111111111111110000111110010011;
assign LUT_2[47233] = 32'b11111111111111101101110110101100;
assign LUT_2[47234] = 32'b11111111111111110111110111001111;
assign LUT_2[47235] = 32'b11111111111111110100101111101000;
assign LUT_2[47236] = 32'b11111111111111101101011011111011;
assign LUT_2[47237] = 32'b11111111111111101010010100010100;
assign LUT_2[47238] = 32'b11111111111111110100010100110111;
assign LUT_2[47239] = 32'b11111111111111110001001101010000;
assign LUT_2[47240] = 32'b11111111111111101011101111110000;
assign LUT_2[47241] = 32'b11111111111111101000101000001001;
assign LUT_2[47242] = 32'b11111111111111110010101000101100;
assign LUT_2[47243] = 32'b11111111111111101111100001000101;
assign LUT_2[47244] = 32'b11111111111111101000001101011000;
assign LUT_2[47245] = 32'b11111111111111100101000101110001;
assign LUT_2[47246] = 32'b11111111111111101111000110010100;
assign LUT_2[47247] = 32'b11111111111111101011111110101101;
assign LUT_2[47248] = 32'b11111111111111101011100010011101;
assign LUT_2[47249] = 32'b11111111111111101000011010110110;
assign LUT_2[47250] = 32'b11111111111111110010011011011001;
assign LUT_2[47251] = 32'b11111111111111101111010011110010;
assign LUT_2[47252] = 32'b11111111111111101000000000000101;
assign LUT_2[47253] = 32'b11111111111111100100111000011110;
assign LUT_2[47254] = 32'b11111111111111101110111001000001;
assign LUT_2[47255] = 32'b11111111111111101011110001011010;
assign LUT_2[47256] = 32'b11111111111111100110010011111010;
assign LUT_2[47257] = 32'b11111111111111100011001100010011;
assign LUT_2[47258] = 32'b11111111111111101101001100110110;
assign LUT_2[47259] = 32'b11111111111111101010000101001111;
assign LUT_2[47260] = 32'b11111111111111100010110001100010;
assign LUT_2[47261] = 32'b11111111111111011111101001111011;
assign LUT_2[47262] = 32'b11111111111111101001101010011110;
assign LUT_2[47263] = 32'b11111111111111100110100010110111;
assign LUT_2[47264] = 32'b11111111111111110001011001111100;
assign LUT_2[47265] = 32'b11111111111111101110010010010101;
assign LUT_2[47266] = 32'b11111111111111111000010010111000;
assign LUT_2[47267] = 32'b11111111111111110101001011010001;
assign LUT_2[47268] = 32'b11111111111111101101110111100100;
assign LUT_2[47269] = 32'b11111111111111101010101111111101;
assign LUT_2[47270] = 32'b11111111111111110100110000100000;
assign LUT_2[47271] = 32'b11111111111111110001101000111001;
assign LUT_2[47272] = 32'b11111111111111101100001011011001;
assign LUT_2[47273] = 32'b11111111111111101001000011110010;
assign LUT_2[47274] = 32'b11111111111111110011000100010101;
assign LUT_2[47275] = 32'b11111111111111101111111100101110;
assign LUT_2[47276] = 32'b11111111111111101000101001000001;
assign LUT_2[47277] = 32'b11111111111111100101100001011010;
assign LUT_2[47278] = 32'b11111111111111101111100001111101;
assign LUT_2[47279] = 32'b11111111111111101100011010010110;
assign LUT_2[47280] = 32'b11111111111111101011111110000110;
assign LUT_2[47281] = 32'b11111111111111101000110110011111;
assign LUT_2[47282] = 32'b11111111111111110010110111000010;
assign LUT_2[47283] = 32'b11111111111111101111101111011011;
assign LUT_2[47284] = 32'b11111111111111101000011011101110;
assign LUT_2[47285] = 32'b11111111111111100101010100000111;
assign LUT_2[47286] = 32'b11111111111111101111010100101010;
assign LUT_2[47287] = 32'b11111111111111101100001101000011;
assign LUT_2[47288] = 32'b11111111111111100110101111100011;
assign LUT_2[47289] = 32'b11111111111111100011100111111100;
assign LUT_2[47290] = 32'b11111111111111101101101000011111;
assign LUT_2[47291] = 32'b11111111111111101010100000111000;
assign LUT_2[47292] = 32'b11111111111111100011001101001011;
assign LUT_2[47293] = 32'b11111111111111100000000101100100;
assign LUT_2[47294] = 32'b11111111111111101010000110000111;
assign LUT_2[47295] = 32'b11111111111111100110111110100000;
assign LUT_2[47296] = 32'b11111111111111101001000110110110;
assign LUT_2[47297] = 32'b11111111111111100101111111001111;
assign LUT_2[47298] = 32'b11111111111111101111111111110010;
assign LUT_2[47299] = 32'b11111111111111101100111000001011;
assign LUT_2[47300] = 32'b11111111111111100101100100011110;
assign LUT_2[47301] = 32'b11111111111111100010011100110111;
assign LUT_2[47302] = 32'b11111111111111101100011101011010;
assign LUT_2[47303] = 32'b11111111111111101001010101110011;
assign LUT_2[47304] = 32'b11111111111111100011111000010011;
assign LUT_2[47305] = 32'b11111111111111100000110000101100;
assign LUT_2[47306] = 32'b11111111111111101010110001001111;
assign LUT_2[47307] = 32'b11111111111111100111101001101000;
assign LUT_2[47308] = 32'b11111111111111100000010101111011;
assign LUT_2[47309] = 32'b11111111111111011101001110010100;
assign LUT_2[47310] = 32'b11111111111111100111001110110111;
assign LUT_2[47311] = 32'b11111111111111100100000111010000;
assign LUT_2[47312] = 32'b11111111111111100011101011000000;
assign LUT_2[47313] = 32'b11111111111111100000100011011001;
assign LUT_2[47314] = 32'b11111111111111101010100011111100;
assign LUT_2[47315] = 32'b11111111111111100111011100010101;
assign LUT_2[47316] = 32'b11111111111111100000001000101000;
assign LUT_2[47317] = 32'b11111111111111011101000001000001;
assign LUT_2[47318] = 32'b11111111111111100111000001100100;
assign LUT_2[47319] = 32'b11111111111111100011111001111101;
assign LUT_2[47320] = 32'b11111111111111011110011100011101;
assign LUT_2[47321] = 32'b11111111111111011011010100110110;
assign LUT_2[47322] = 32'b11111111111111100101010101011001;
assign LUT_2[47323] = 32'b11111111111111100010001101110010;
assign LUT_2[47324] = 32'b11111111111111011010111010000101;
assign LUT_2[47325] = 32'b11111111111111010111110010011110;
assign LUT_2[47326] = 32'b11111111111111100001110011000001;
assign LUT_2[47327] = 32'b11111111111111011110101011011010;
assign LUT_2[47328] = 32'b11111111111111101001100010011111;
assign LUT_2[47329] = 32'b11111111111111100110011010111000;
assign LUT_2[47330] = 32'b11111111111111110000011011011011;
assign LUT_2[47331] = 32'b11111111111111101101010011110100;
assign LUT_2[47332] = 32'b11111111111111100110000000000111;
assign LUT_2[47333] = 32'b11111111111111100010111000100000;
assign LUT_2[47334] = 32'b11111111111111101100111001000011;
assign LUT_2[47335] = 32'b11111111111111101001110001011100;
assign LUT_2[47336] = 32'b11111111111111100100010011111100;
assign LUT_2[47337] = 32'b11111111111111100001001100010101;
assign LUT_2[47338] = 32'b11111111111111101011001100111000;
assign LUT_2[47339] = 32'b11111111111111101000000101010001;
assign LUT_2[47340] = 32'b11111111111111100000110001100100;
assign LUT_2[47341] = 32'b11111111111111011101101001111101;
assign LUT_2[47342] = 32'b11111111111111100111101010100000;
assign LUT_2[47343] = 32'b11111111111111100100100010111001;
assign LUT_2[47344] = 32'b11111111111111100100000110101001;
assign LUT_2[47345] = 32'b11111111111111100000111111000010;
assign LUT_2[47346] = 32'b11111111111111101010111111100101;
assign LUT_2[47347] = 32'b11111111111111100111110111111110;
assign LUT_2[47348] = 32'b11111111111111100000100100010001;
assign LUT_2[47349] = 32'b11111111111111011101011100101010;
assign LUT_2[47350] = 32'b11111111111111100111011101001101;
assign LUT_2[47351] = 32'b11111111111111100100010101100110;
assign LUT_2[47352] = 32'b11111111111111011110111000000110;
assign LUT_2[47353] = 32'b11111111111111011011110000011111;
assign LUT_2[47354] = 32'b11111111111111100101110001000010;
assign LUT_2[47355] = 32'b11111111111111100010101001011011;
assign LUT_2[47356] = 32'b11111111111111011011010101101110;
assign LUT_2[47357] = 32'b11111111111111011000001110000111;
assign LUT_2[47358] = 32'b11111111111111100010001110101010;
assign LUT_2[47359] = 32'b11111111111111011111000111000011;
assign LUT_2[47360] = 32'b11111111111111110000101000101010;
assign LUT_2[47361] = 32'b11111111111111101101100001000011;
assign LUT_2[47362] = 32'b11111111111111110111100001100110;
assign LUT_2[47363] = 32'b11111111111111110100011001111111;
assign LUT_2[47364] = 32'b11111111111111101101000110010010;
assign LUT_2[47365] = 32'b11111111111111101001111110101011;
assign LUT_2[47366] = 32'b11111111111111110011111111001110;
assign LUT_2[47367] = 32'b11111111111111110000110111100111;
assign LUT_2[47368] = 32'b11111111111111101011011010000111;
assign LUT_2[47369] = 32'b11111111111111101000010010100000;
assign LUT_2[47370] = 32'b11111111111111110010010011000011;
assign LUT_2[47371] = 32'b11111111111111101111001011011100;
assign LUT_2[47372] = 32'b11111111111111100111110111101111;
assign LUT_2[47373] = 32'b11111111111111100100110000001000;
assign LUT_2[47374] = 32'b11111111111111101110110000101011;
assign LUT_2[47375] = 32'b11111111111111101011101001000100;
assign LUT_2[47376] = 32'b11111111111111101011001100110100;
assign LUT_2[47377] = 32'b11111111111111101000000101001101;
assign LUT_2[47378] = 32'b11111111111111110010000101110000;
assign LUT_2[47379] = 32'b11111111111111101110111110001001;
assign LUT_2[47380] = 32'b11111111111111100111101010011100;
assign LUT_2[47381] = 32'b11111111111111100100100010110101;
assign LUT_2[47382] = 32'b11111111111111101110100011011000;
assign LUT_2[47383] = 32'b11111111111111101011011011110001;
assign LUT_2[47384] = 32'b11111111111111100101111110010001;
assign LUT_2[47385] = 32'b11111111111111100010110110101010;
assign LUT_2[47386] = 32'b11111111111111101100110111001101;
assign LUT_2[47387] = 32'b11111111111111101001101111100110;
assign LUT_2[47388] = 32'b11111111111111100010011011111001;
assign LUT_2[47389] = 32'b11111111111111011111010100010010;
assign LUT_2[47390] = 32'b11111111111111101001010100110101;
assign LUT_2[47391] = 32'b11111111111111100110001101001110;
assign LUT_2[47392] = 32'b11111111111111110001000100010011;
assign LUT_2[47393] = 32'b11111111111111101101111100101100;
assign LUT_2[47394] = 32'b11111111111111110111111101001111;
assign LUT_2[47395] = 32'b11111111111111110100110101101000;
assign LUT_2[47396] = 32'b11111111111111101101100001111011;
assign LUT_2[47397] = 32'b11111111111111101010011010010100;
assign LUT_2[47398] = 32'b11111111111111110100011010110111;
assign LUT_2[47399] = 32'b11111111111111110001010011010000;
assign LUT_2[47400] = 32'b11111111111111101011110101110000;
assign LUT_2[47401] = 32'b11111111111111101000101110001001;
assign LUT_2[47402] = 32'b11111111111111110010101110101100;
assign LUT_2[47403] = 32'b11111111111111101111100111000101;
assign LUT_2[47404] = 32'b11111111111111101000010011011000;
assign LUT_2[47405] = 32'b11111111111111100101001011110001;
assign LUT_2[47406] = 32'b11111111111111101111001100010100;
assign LUT_2[47407] = 32'b11111111111111101100000100101101;
assign LUT_2[47408] = 32'b11111111111111101011101000011101;
assign LUT_2[47409] = 32'b11111111111111101000100000110110;
assign LUT_2[47410] = 32'b11111111111111110010100001011001;
assign LUT_2[47411] = 32'b11111111111111101111011001110010;
assign LUT_2[47412] = 32'b11111111111111101000000110000101;
assign LUT_2[47413] = 32'b11111111111111100100111110011110;
assign LUT_2[47414] = 32'b11111111111111101110111111000001;
assign LUT_2[47415] = 32'b11111111111111101011110111011010;
assign LUT_2[47416] = 32'b11111111111111100110011001111010;
assign LUT_2[47417] = 32'b11111111111111100011010010010011;
assign LUT_2[47418] = 32'b11111111111111101101010010110110;
assign LUT_2[47419] = 32'b11111111111111101010001011001111;
assign LUT_2[47420] = 32'b11111111111111100010110111100010;
assign LUT_2[47421] = 32'b11111111111111011111101111111011;
assign LUT_2[47422] = 32'b11111111111111101001110000011110;
assign LUT_2[47423] = 32'b11111111111111100110101000110111;
assign LUT_2[47424] = 32'b11111111111111101000110001001101;
assign LUT_2[47425] = 32'b11111111111111100101101001100110;
assign LUT_2[47426] = 32'b11111111111111101111101010001001;
assign LUT_2[47427] = 32'b11111111111111101100100010100010;
assign LUT_2[47428] = 32'b11111111111111100101001110110101;
assign LUT_2[47429] = 32'b11111111111111100010000111001110;
assign LUT_2[47430] = 32'b11111111111111101100000111110001;
assign LUT_2[47431] = 32'b11111111111111101001000000001010;
assign LUT_2[47432] = 32'b11111111111111100011100010101010;
assign LUT_2[47433] = 32'b11111111111111100000011011000011;
assign LUT_2[47434] = 32'b11111111111111101010011011100110;
assign LUT_2[47435] = 32'b11111111111111100111010011111111;
assign LUT_2[47436] = 32'b11111111111111100000000000010010;
assign LUT_2[47437] = 32'b11111111111111011100111000101011;
assign LUT_2[47438] = 32'b11111111111111100110111001001110;
assign LUT_2[47439] = 32'b11111111111111100011110001100111;
assign LUT_2[47440] = 32'b11111111111111100011010101010111;
assign LUT_2[47441] = 32'b11111111111111100000001101110000;
assign LUT_2[47442] = 32'b11111111111111101010001110010011;
assign LUT_2[47443] = 32'b11111111111111100111000110101100;
assign LUT_2[47444] = 32'b11111111111111011111110010111111;
assign LUT_2[47445] = 32'b11111111111111011100101011011000;
assign LUT_2[47446] = 32'b11111111111111100110101011111011;
assign LUT_2[47447] = 32'b11111111111111100011100100010100;
assign LUT_2[47448] = 32'b11111111111111011110000110110100;
assign LUT_2[47449] = 32'b11111111111111011010111111001101;
assign LUT_2[47450] = 32'b11111111111111100100111111110000;
assign LUT_2[47451] = 32'b11111111111111100001111000001001;
assign LUT_2[47452] = 32'b11111111111111011010100100011100;
assign LUT_2[47453] = 32'b11111111111111010111011100110101;
assign LUT_2[47454] = 32'b11111111111111100001011101011000;
assign LUT_2[47455] = 32'b11111111111111011110010101110001;
assign LUT_2[47456] = 32'b11111111111111101001001100110110;
assign LUT_2[47457] = 32'b11111111111111100110000101001111;
assign LUT_2[47458] = 32'b11111111111111110000000101110010;
assign LUT_2[47459] = 32'b11111111111111101100111110001011;
assign LUT_2[47460] = 32'b11111111111111100101101010011110;
assign LUT_2[47461] = 32'b11111111111111100010100010110111;
assign LUT_2[47462] = 32'b11111111111111101100100011011010;
assign LUT_2[47463] = 32'b11111111111111101001011011110011;
assign LUT_2[47464] = 32'b11111111111111100011111110010011;
assign LUT_2[47465] = 32'b11111111111111100000110110101100;
assign LUT_2[47466] = 32'b11111111111111101010110111001111;
assign LUT_2[47467] = 32'b11111111111111100111101111101000;
assign LUT_2[47468] = 32'b11111111111111100000011011111011;
assign LUT_2[47469] = 32'b11111111111111011101010100010100;
assign LUT_2[47470] = 32'b11111111111111100111010100110111;
assign LUT_2[47471] = 32'b11111111111111100100001101010000;
assign LUT_2[47472] = 32'b11111111111111100011110001000000;
assign LUT_2[47473] = 32'b11111111111111100000101001011001;
assign LUT_2[47474] = 32'b11111111111111101010101001111100;
assign LUT_2[47475] = 32'b11111111111111100111100010010101;
assign LUT_2[47476] = 32'b11111111111111100000001110101000;
assign LUT_2[47477] = 32'b11111111111111011101000111000001;
assign LUT_2[47478] = 32'b11111111111111100111000111100100;
assign LUT_2[47479] = 32'b11111111111111100011111111111101;
assign LUT_2[47480] = 32'b11111111111111011110100010011101;
assign LUT_2[47481] = 32'b11111111111111011011011010110110;
assign LUT_2[47482] = 32'b11111111111111100101011011011001;
assign LUT_2[47483] = 32'b11111111111111100010010011110010;
assign LUT_2[47484] = 32'b11111111111111011011000000000101;
assign LUT_2[47485] = 32'b11111111111111010111111000011110;
assign LUT_2[47486] = 32'b11111111111111100001111001000001;
assign LUT_2[47487] = 32'b11111111111111011110110001011010;
assign LUT_2[47488] = 32'b11111111111111110100111100111001;
assign LUT_2[47489] = 32'b11111111111111110001110101010010;
assign LUT_2[47490] = 32'b11111111111111111011110101110101;
assign LUT_2[47491] = 32'b11111111111111111000101110001110;
assign LUT_2[47492] = 32'b11111111111111110001011010100001;
assign LUT_2[47493] = 32'b11111111111111101110010010111010;
assign LUT_2[47494] = 32'b11111111111111111000010011011101;
assign LUT_2[47495] = 32'b11111111111111110101001011110110;
assign LUT_2[47496] = 32'b11111111111111101111101110010110;
assign LUT_2[47497] = 32'b11111111111111101100100110101111;
assign LUT_2[47498] = 32'b11111111111111110110100111010010;
assign LUT_2[47499] = 32'b11111111111111110011011111101011;
assign LUT_2[47500] = 32'b11111111111111101100001011111110;
assign LUT_2[47501] = 32'b11111111111111101001000100010111;
assign LUT_2[47502] = 32'b11111111111111110011000100111010;
assign LUT_2[47503] = 32'b11111111111111101111111101010011;
assign LUT_2[47504] = 32'b11111111111111101111100001000011;
assign LUT_2[47505] = 32'b11111111111111101100011001011100;
assign LUT_2[47506] = 32'b11111111111111110110011001111111;
assign LUT_2[47507] = 32'b11111111111111110011010010011000;
assign LUT_2[47508] = 32'b11111111111111101011111110101011;
assign LUT_2[47509] = 32'b11111111111111101000110111000100;
assign LUT_2[47510] = 32'b11111111111111110010110111100111;
assign LUT_2[47511] = 32'b11111111111111101111110000000000;
assign LUT_2[47512] = 32'b11111111111111101010010010100000;
assign LUT_2[47513] = 32'b11111111111111100111001010111001;
assign LUT_2[47514] = 32'b11111111111111110001001011011100;
assign LUT_2[47515] = 32'b11111111111111101110000011110101;
assign LUT_2[47516] = 32'b11111111111111100110110000001000;
assign LUT_2[47517] = 32'b11111111111111100011101000100001;
assign LUT_2[47518] = 32'b11111111111111101101101001000100;
assign LUT_2[47519] = 32'b11111111111111101010100001011101;
assign LUT_2[47520] = 32'b11111111111111110101011000100010;
assign LUT_2[47521] = 32'b11111111111111110010010000111011;
assign LUT_2[47522] = 32'b11111111111111111100010001011110;
assign LUT_2[47523] = 32'b11111111111111111001001001110111;
assign LUT_2[47524] = 32'b11111111111111110001110110001010;
assign LUT_2[47525] = 32'b11111111111111101110101110100011;
assign LUT_2[47526] = 32'b11111111111111111000101111000110;
assign LUT_2[47527] = 32'b11111111111111110101100111011111;
assign LUT_2[47528] = 32'b11111111111111110000001001111111;
assign LUT_2[47529] = 32'b11111111111111101101000010011000;
assign LUT_2[47530] = 32'b11111111111111110111000010111011;
assign LUT_2[47531] = 32'b11111111111111110011111011010100;
assign LUT_2[47532] = 32'b11111111111111101100100111100111;
assign LUT_2[47533] = 32'b11111111111111101001100000000000;
assign LUT_2[47534] = 32'b11111111111111110011100000100011;
assign LUT_2[47535] = 32'b11111111111111110000011000111100;
assign LUT_2[47536] = 32'b11111111111111101111111100101100;
assign LUT_2[47537] = 32'b11111111111111101100110101000101;
assign LUT_2[47538] = 32'b11111111111111110110110101101000;
assign LUT_2[47539] = 32'b11111111111111110011101110000001;
assign LUT_2[47540] = 32'b11111111111111101100011010010100;
assign LUT_2[47541] = 32'b11111111111111101001010010101101;
assign LUT_2[47542] = 32'b11111111111111110011010011010000;
assign LUT_2[47543] = 32'b11111111111111110000001011101001;
assign LUT_2[47544] = 32'b11111111111111101010101110001001;
assign LUT_2[47545] = 32'b11111111111111100111100110100010;
assign LUT_2[47546] = 32'b11111111111111110001100111000101;
assign LUT_2[47547] = 32'b11111111111111101110011111011110;
assign LUT_2[47548] = 32'b11111111111111100111001011110001;
assign LUT_2[47549] = 32'b11111111111111100100000100001010;
assign LUT_2[47550] = 32'b11111111111111101110000100101101;
assign LUT_2[47551] = 32'b11111111111111101010111101000110;
assign LUT_2[47552] = 32'b11111111111111101101000101011100;
assign LUT_2[47553] = 32'b11111111111111101001111101110101;
assign LUT_2[47554] = 32'b11111111111111110011111110011000;
assign LUT_2[47555] = 32'b11111111111111110000110110110001;
assign LUT_2[47556] = 32'b11111111111111101001100011000100;
assign LUT_2[47557] = 32'b11111111111111100110011011011101;
assign LUT_2[47558] = 32'b11111111111111110000011100000000;
assign LUT_2[47559] = 32'b11111111111111101101010100011001;
assign LUT_2[47560] = 32'b11111111111111100111110110111001;
assign LUT_2[47561] = 32'b11111111111111100100101111010010;
assign LUT_2[47562] = 32'b11111111111111101110101111110101;
assign LUT_2[47563] = 32'b11111111111111101011101000001110;
assign LUT_2[47564] = 32'b11111111111111100100010100100001;
assign LUT_2[47565] = 32'b11111111111111100001001100111010;
assign LUT_2[47566] = 32'b11111111111111101011001101011101;
assign LUT_2[47567] = 32'b11111111111111101000000101110110;
assign LUT_2[47568] = 32'b11111111111111100111101001100110;
assign LUT_2[47569] = 32'b11111111111111100100100001111111;
assign LUT_2[47570] = 32'b11111111111111101110100010100010;
assign LUT_2[47571] = 32'b11111111111111101011011010111011;
assign LUT_2[47572] = 32'b11111111111111100100000111001110;
assign LUT_2[47573] = 32'b11111111111111100000111111100111;
assign LUT_2[47574] = 32'b11111111111111101011000000001010;
assign LUT_2[47575] = 32'b11111111111111100111111000100011;
assign LUT_2[47576] = 32'b11111111111111100010011011000011;
assign LUT_2[47577] = 32'b11111111111111011111010011011100;
assign LUT_2[47578] = 32'b11111111111111101001010011111111;
assign LUT_2[47579] = 32'b11111111111111100110001100011000;
assign LUT_2[47580] = 32'b11111111111111011110111000101011;
assign LUT_2[47581] = 32'b11111111111111011011110001000100;
assign LUT_2[47582] = 32'b11111111111111100101110001100111;
assign LUT_2[47583] = 32'b11111111111111100010101010000000;
assign LUT_2[47584] = 32'b11111111111111101101100001000101;
assign LUT_2[47585] = 32'b11111111111111101010011001011110;
assign LUT_2[47586] = 32'b11111111111111110100011010000001;
assign LUT_2[47587] = 32'b11111111111111110001010010011010;
assign LUT_2[47588] = 32'b11111111111111101001111110101101;
assign LUT_2[47589] = 32'b11111111111111100110110111000110;
assign LUT_2[47590] = 32'b11111111111111110000110111101001;
assign LUT_2[47591] = 32'b11111111111111101101110000000010;
assign LUT_2[47592] = 32'b11111111111111101000010010100010;
assign LUT_2[47593] = 32'b11111111111111100101001010111011;
assign LUT_2[47594] = 32'b11111111111111101111001011011110;
assign LUT_2[47595] = 32'b11111111111111101100000011110111;
assign LUT_2[47596] = 32'b11111111111111100100110000001010;
assign LUT_2[47597] = 32'b11111111111111100001101000100011;
assign LUT_2[47598] = 32'b11111111111111101011101001000110;
assign LUT_2[47599] = 32'b11111111111111101000100001011111;
assign LUT_2[47600] = 32'b11111111111111101000000101001111;
assign LUT_2[47601] = 32'b11111111111111100100111101101000;
assign LUT_2[47602] = 32'b11111111111111101110111110001011;
assign LUT_2[47603] = 32'b11111111111111101011110110100100;
assign LUT_2[47604] = 32'b11111111111111100100100010110111;
assign LUT_2[47605] = 32'b11111111111111100001011011010000;
assign LUT_2[47606] = 32'b11111111111111101011011011110011;
assign LUT_2[47607] = 32'b11111111111111101000010100001100;
assign LUT_2[47608] = 32'b11111111111111100010110110101100;
assign LUT_2[47609] = 32'b11111111111111011111101111000101;
assign LUT_2[47610] = 32'b11111111111111101001101111101000;
assign LUT_2[47611] = 32'b11111111111111100110101000000001;
assign LUT_2[47612] = 32'b11111111111111011111010100010100;
assign LUT_2[47613] = 32'b11111111111111011100001100101101;
assign LUT_2[47614] = 32'b11111111111111100110001101010000;
assign LUT_2[47615] = 32'b11111111111111100011000101101001;
assign LUT_2[47616] = 32'b11111111111111110001011011110110;
assign LUT_2[47617] = 32'b11111111111111101110010100001111;
assign LUT_2[47618] = 32'b11111111111111111000010100110010;
assign LUT_2[47619] = 32'b11111111111111110101001101001011;
assign LUT_2[47620] = 32'b11111111111111101101111001011110;
assign LUT_2[47621] = 32'b11111111111111101010110001110111;
assign LUT_2[47622] = 32'b11111111111111110100110010011010;
assign LUT_2[47623] = 32'b11111111111111110001101010110011;
assign LUT_2[47624] = 32'b11111111111111101100001101010011;
assign LUT_2[47625] = 32'b11111111111111101001000101101100;
assign LUT_2[47626] = 32'b11111111111111110011000110001111;
assign LUT_2[47627] = 32'b11111111111111101111111110101000;
assign LUT_2[47628] = 32'b11111111111111101000101010111011;
assign LUT_2[47629] = 32'b11111111111111100101100011010100;
assign LUT_2[47630] = 32'b11111111111111101111100011110111;
assign LUT_2[47631] = 32'b11111111111111101100011100010000;
assign LUT_2[47632] = 32'b11111111111111101100000000000000;
assign LUT_2[47633] = 32'b11111111111111101000111000011001;
assign LUT_2[47634] = 32'b11111111111111110010111000111100;
assign LUT_2[47635] = 32'b11111111111111101111110001010101;
assign LUT_2[47636] = 32'b11111111111111101000011101101000;
assign LUT_2[47637] = 32'b11111111111111100101010110000001;
assign LUT_2[47638] = 32'b11111111111111101111010110100100;
assign LUT_2[47639] = 32'b11111111111111101100001110111101;
assign LUT_2[47640] = 32'b11111111111111100110110001011101;
assign LUT_2[47641] = 32'b11111111111111100011101001110110;
assign LUT_2[47642] = 32'b11111111111111101101101010011001;
assign LUT_2[47643] = 32'b11111111111111101010100010110010;
assign LUT_2[47644] = 32'b11111111111111100011001111000101;
assign LUT_2[47645] = 32'b11111111111111100000000111011110;
assign LUT_2[47646] = 32'b11111111111111101010001000000001;
assign LUT_2[47647] = 32'b11111111111111100111000000011010;
assign LUT_2[47648] = 32'b11111111111111110001110111011111;
assign LUT_2[47649] = 32'b11111111111111101110101111111000;
assign LUT_2[47650] = 32'b11111111111111111000110000011011;
assign LUT_2[47651] = 32'b11111111111111110101101000110100;
assign LUT_2[47652] = 32'b11111111111111101110010101000111;
assign LUT_2[47653] = 32'b11111111111111101011001101100000;
assign LUT_2[47654] = 32'b11111111111111110101001110000011;
assign LUT_2[47655] = 32'b11111111111111110010000110011100;
assign LUT_2[47656] = 32'b11111111111111101100101000111100;
assign LUT_2[47657] = 32'b11111111111111101001100001010101;
assign LUT_2[47658] = 32'b11111111111111110011100001111000;
assign LUT_2[47659] = 32'b11111111111111110000011010010001;
assign LUT_2[47660] = 32'b11111111111111101001000110100100;
assign LUT_2[47661] = 32'b11111111111111100101111110111101;
assign LUT_2[47662] = 32'b11111111111111101111111111100000;
assign LUT_2[47663] = 32'b11111111111111101100110111111001;
assign LUT_2[47664] = 32'b11111111111111101100011011101001;
assign LUT_2[47665] = 32'b11111111111111101001010100000010;
assign LUT_2[47666] = 32'b11111111111111110011010100100101;
assign LUT_2[47667] = 32'b11111111111111110000001100111110;
assign LUT_2[47668] = 32'b11111111111111101000111001010001;
assign LUT_2[47669] = 32'b11111111111111100101110001101010;
assign LUT_2[47670] = 32'b11111111111111101111110010001101;
assign LUT_2[47671] = 32'b11111111111111101100101010100110;
assign LUT_2[47672] = 32'b11111111111111100111001101000110;
assign LUT_2[47673] = 32'b11111111111111100100000101011111;
assign LUT_2[47674] = 32'b11111111111111101110000110000010;
assign LUT_2[47675] = 32'b11111111111111101010111110011011;
assign LUT_2[47676] = 32'b11111111111111100011101010101110;
assign LUT_2[47677] = 32'b11111111111111100000100011000111;
assign LUT_2[47678] = 32'b11111111111111101010100011101010;
assign LUT_2[47679] = 32'b11111111111111100111011100000011;
assign LUT_2[47680] = 32'b11111111111111101001100100011001;
assign LUT_2[47681] = 32'b11111111111111100110011100110010;
assign LUT_2[47682] = 32'b11111111111111110000011101010101;
assign LUT_2[47683] = 32'b11111111111111101101010101101110;
assign LUT_2[47684] = 32'b11111111111111100110000010000001;
assign LUT_2[47685] = 32'b11111111111111100010111010011010;
assign LUT_2[47686] = 32'b11111111111111101100111010111101;
assign LUT_2[47687] = 32'b11111111111111101001110011010110;
assign LUT_2[47688] = 32'b11111111111111100100010101110110;
assign LUT_2[47689] = 32'b11111111111111100001001110001111;
assign LUT_2[47690] = 32'b11111111111111101011001110110010;
assign LUT_2[47691] = 32'b11111111111111101000000111001011;
assign LUT_2[47692] = 32'b11111111111111100000110011011110;
assign LUT_2[47693] = 32'b11111111111111011101101011110111;
assign LUT_2[47694] = 32'b11111111111111100111101100011010;
assign LUT_2[47695] = 32'b11111111111111100100100100110011;
assign LUT_2[47696] = 32'b11111111111111100100001000100011;
assign LUT_2[47697] = 32'b11111111111111100001000000111100;
assign LUT_2[47698] = 32'b11111111111111101011000001011111;
assign LUT_2[47699] = 32'b11111111111111100111111001111000;
assign LUT_2[47700] = 32'b11111111111111100000100110001011;
assign LUT_2[47701] = 32'b11111111111111011101011110100100;
assign LUT_2[47702] = 32'b11111111111111100111011111000111;
assign LUT_2[47703] = 32'b11111111111111100100010111100000;
assign LUT_2[47704] = 32'b11111111111111011110111010000000;
assign LUT_2[47705] = 32'b11111111111111011011110010011001;
assign LUT_2[47706] = 32'b11111111111111100101110010111100;
assign LUT_2[47707] = 32'b11111111111111100010101011010101;
assign LUT_2[47708] = 32'b11111111111111011011010111101000;
assign LUT_2[47709] = 32'b11111111111111011000010000000001;
assign LUT_2[47710] = 32'b11111111111111100010010000100100;
assign LUT_2[47711] = 32'b11111111111111011111001000111101;
assign LUT_2[47712] = 32'b11111111111111101010000000000010;
assign LUT_2[47713] = 32'b11111111111111100110111000011011;
assign LUT_2[47714] = 32'b11111111111111110000111000111110;
assign LUT_2[47715] = 32'b11111111111111101101110001010111;
assign LUT_2[47716] = 32'b11111111111111100110011101101010;
assign LUT_2[47717] = 32'b11111111111111100011010110000011;
assign LUT_2[47718] = 32'b11111111111111101101010110100110;
assign LUT_2[47719] = 32'b11111111111111101010001110111111;
assign LUT_2[47720] = 32'b11111111111111100100110001011111;
assign LUT_2[47721] = 32'b11111111111111100001101001111000;
assign LUT_2[47722] = 32'b11111111111111101011101010011011;
assign LUT_2[47723] = 32'b11111111111111101000100010110100;
assign LUT_2[47724] = 32'b11111111111111100001001111000111;
assign LUT_2[47725] = 32'b11111111111111011110000111100000;
assign LUT_2[47726] = 32'b11111111111111101000001000000011;
assign LUT_2[47727] = 32'b11111111111111100101000000011100;
assign LUT_2[47728] = 32'b11111111111111100100100100001100;
assign LUT_2[47729] = 32'b11111111111111100001011100100101;
assign LUT_2[47730] = 32'b11111111111111101011011101001000;
assign LUT_2[47731] = 32'b11111111111111101000010101100001;
assign LUT_2[47732] = 32'b11111111111111100001000001110100;
assign LUT_2[47733] = 32'b11111111111111011101111010001101;
assign LUT_2[47734] = 32'b11111111111111100111111010110000;
assign LUT_2[47735] = 32'b11111111111111100100110011001001;
assign LUT_2[47736] = 32'b11111111111111011111010101101001;
assign LUT_2[47737] = 32'b11111111111111011100001110000010;
assign LUT_2[47738] = 32'b11111111111111100110001110100101;
assign LUT_2[47739] = 32'b11111111111111100011000110111110;
assign LUT_2[47740] = 32'b11111111111111011011110011010001;
assign LUT_2[47741] = 32'b11111111111111011000101011101010;
assign LUT_2[47742] = 32'b11111111111111100010101100001101;
assign LUT_2[47743] = 32'b11111111111111011111100100100110;
assign LUT_2[47744] = 32'b11111111111111110101110000000101;
assign LUT_2[47745] = 32'b11111111111111110010101000011110;
assign LUT_2[47746] = 32'b11111111111111111100101001000001;
assign LUT_2[47747] = 32'b11111111111111111001100001011010;
assign LUT_2[47748] = 32'b11111111111111110010001101101101;
assign LUT_2[47749] = 32'b11111111111111101111000110000110;
assign LUT_2[47750] = 32'b11111111111111111001000110101001;
assign LUT_2[47751] = 32'b11111111111111110101111111000010;
assign LUT_2[47752] = 32'b11111111111111110000100001100010;
assign LUT_2[47753] = 32'b11111111111111101101011001111011;
assign LUT_2[47754] = 32'b11111111111111110111011010011110;
assign LUT_2[47755] = 32'b11111111111111110100010010110111;
assign LUT_2[47756] = 32'b11111111111111101100111111001010;
assign LUT_2[47757] = 32'b11111111111111101001110111100011;
assign LUT_2[47758] = 32'b11111111111111110011111000000110;
assign LUT_2[47759] = 32'b11111111111111110000110000011111;
assign LUT_2[47760] = 32'b11111111111111110000010100001111;
assign LUT_2[47761] = 32'b11111111111111101101001100101000;
assign LUT_2[47762] = 32'b11111111111111110111001101001011;
assign LUT_2[47763] = 32'b11111111111111110100000101100100;
assign LUT_2[47764] = 32'b11111111111111101100110001110111;
assign LUT_2[47765] = 32'b11111111111111101001101010010000;
assign LUT_2[47766] = 32'b11111111111111110011101010110011;
assign LUT_2[47767] = 32'b11111111111111110000100011001100;
assign LUT_2[47768] = 32'b11111111111111101011000101101100;
assign LUT_2[47769] = 32'b11111111111111100111111110000101;
assign LUT_2[47770] = 32'b11111111111111110001111110101000;
assign LUT_2[47771] = 32'b11111111111111101110110111000001;
assign LUT_2[47772] = 32'b11111111111111100111100011010100;
assign LUT_2[47773] = 32'b11111111111111100100011011101101;
assign LUT_2[47774] = 32'b11111111111111101110011100010000;
assign LUT_2[47775] = 32'b11111111111111101011010100101001;
assign LUT_2[47776] = 32'b11111111111111110110001011101110;
assign LUT_2[47777] = 32'b11111111111111110011000100000111;
assign LUT_2[47778] = 32'b11111111111111111101000100101010;
assign LUT_2[47779] = 32'b11111111111111111001111101000011;
assign LUT_2[47780] = 32'b11111111111111110010101001010110;
assign LUT_2[47781] = 32'b11111111111111101111100001101111;
assign LUT_2[47782] = 32'b11111111111111111001100010010010;
assign LUT_2[47783] = 32'b11111111111111110110011010101011;
assign LUT_2[47784] = 32'b11111111111111110000111101001011;
assign LUT_2[47785] = 32'b11111111111111101101110101100100;
assign LUT_2[47786] = 32'b11111111111111110111110110000111;
assign LUT_2[47787] = 32'b11111111111111110100101110100000;
assign LUT_2[47788] = 32'b11111111111111101101011010110011;
assign LUT_2[47789] = 32'b11111111111111101010010011001100;
assign LUT_2[47790] = 32'b11111111111111110100010011101111;
assign LUT_2[47791] = 32'b11111111111111110001001100001000;
assign LUT_2[47792] = 32'b11111111111111110000101111111000;
assign LUT_2[47793] = 32'b11111111111111101101101000010001;
assign LUT_2[47794] = 32'b11111111111111110111101000110100;
assign LUT_2[47795] = 32'b11111111111111110100100001001101;
assign LUT_2[47796] = 32'b11111111111111101101001101100000;
assign LUT_2[47797] = 32'b11111111111111101010000101111001;
assign LUT_2[47798] = 32'b11111111111111110100000110011100;
assign LUT_2[47799] = 32'b11111111111111110000111110110101;
assign LUT_2[47800] = 32'b11111111111111101011100001010101;
assign LUT_2[47801] = 32'b11111111111111101000011001101110;
assign LUT_2[47802] = 32'b11111111111111110010011010010001;
assign LUT_2[47803] = 32'b11111111111111101111010010101010;
assign LUT_2[47804] = 32'b11111111111111100111111110111101;
assign LUT_2[47805] = 32'b11111111111111100100110111010110;
assign LUT_2[47806] = 32'b11111111111111101110110111111001;
assign LUT_2[47807] = 32'b11111111111111101011110000010010;
assign LUT_2[47808] = 32'b11111111111111101101111000101000;
assign LUT_2[47809] = 32'b11111111111111101010110001000001;
assign LUT_2[47810] = 32'b11111111111111110100110001100100;
assign LUT_2[47811] = 32'b11111111111111110001101001111101;
assign LUT_2[47812] = 32'b11111111111111101010010110010000;
assign LUT_2[47813] = 32'b11111111111111100111001110101001;
assign LUT_2[47814] = 32'b11111111111111110001001111001100;
assign LUT_2[47815] = 32'b11111111111111101110000111100101;
assign LUT_2[47816] = 32'b11111111111111101000101010000101;
assign LUT_2[47817] = 32'b11111111111111100101100010011110;
assign LUT_2[47818] = 32'b11111111111111101111100011000001;
assign LUT_2[47819] = 32'b11111111111111101100011011011010;
assign LUT_2[47820] = 32'b11111111111111100101000111101101;
assign LUT_2[47821] = 32'b11111111111111100010000000000110;
assign LUT_2[47822] = 32'b11111111111111101100000000101001;
assign LUT_2[47823] = 32'b11111111111111101000111001000010;
assign LUT_2[47824] = 32'b11111111111111101000011100110010;
assign LUT_2[47825] = 32'b11111111111111100101010101001011;
assign LUT_2[47826] = 32'b11111111111111101111010101101110;
assign LUT_2[47827] = 32'b11111111111111101100001110000111;
assign LUT_2[47828] = 32'b11111111111111100100111010011010;
assign LUT_2[47829] = 32'b11111111111111100001110010110011;
assign LUT_2[47830] = 32'b11111111111111101011110011010110;
assign LUT_2[47831] = 32'b11111111111111101000101011101111;
assign LUT_2[47832] = 32'b11111111111111100011001110001111;
assign LUT_2[47833] = 32'b11111111111111100000000110101000;
assign LUT_2[47834] = 32'b11111111111111101010000111001011;
assign LUT_2[47835] = 32'b11111111111111100110111111100100;
assign LUT_2[47836] = 32'b11111111111111011111101011110111;
assign LUT_2[47837] = 32'b11111111111111011100100100010000;
assign LUT_2[47838] = 32'b11111111111111100110100100110011;
assign LUT_2[47839] = 32'b11111111111111100011011101001100;
assign LUT_2[47840] = 32'b11111111111111101110010100010001;
assign LUT_2[47841] = 32'b11111111111111101011001100101010;
assign LUT_2[47842] = 32'b11111111111111110101001101001101;
assign LUT_2[47843] = 32'b11111111111111110010000101100110;
assign LUT_2[47844] = 32'b11111111111111101010110001111001;
assign LUT_2[47845] = 32'b11111111111111100111101010010010;
assign LUT_2[47846] = 32'b11111111111111110001101010110101;
assign LUT_2[47847] = 32'b11111111111111101110100011001110;
assign LUT_2[47848] = 32'b11111111111111101001000101101110;
assign LUT_2[47849] = 32'b11111111111111100101111110000111;
assign LUT_2[47850] = 32'b11111111111111101111111110101010;
assign LUT_2[47851] = 32'b11111111111111101100110111000011;
assign LUT_2[47852] = 32'b11111111111111100101100011010110;
assign LUT_2[47853] = 32'b11111111111111100010011011101111;
assign LUT_2[47854] = 32'b11111111111111101100011100010010;
assign LUT_2[47855] = 32'b11111111111111101001010100101011;
assign LUT_2[47856] = 32'b11111111111111101000111000011011;
assign LUT_2[47857] = 32'b11111111111111100101110000110100;
assign LUT_2[47858] = 32'b11111111111111101111110001010111;
assign LUT_2[47859] = 32'b11111111111111101100101001110000;
assign LUT_2[47860] = 32'b11111111111111100101010110000011;
assign LUT_2[47861] = 32'b11111111111111100010001110011100;
assign LUT_2[47862] = 32'b11111111111111101100001110111111;
assign LUT_2[47863] = 32'b11111111111111101001000111011000;
assign LUT_2[47864] = 32'b11111111111111100011101001111000;
assign LUT_2[47865] = 32'b11111111111111100000100010010001;
assign LUT_2[47866] = 32'b11111111111111101010100010110100;
assign LUT_2[47867] = 32'b11111111111111100111011011001101;
assign LUT_2[47868] = 32'b11111111111111100000000111100000;
assign LUT_2[47869] = 32'b11111111111111011100111111111001;
assign LUT_2[47870] = 32'b11111111111111100111000000011100;
assign LUT_2[47871] = 32'b11111111111111100011111000110101;
assign LUT_2[47872] = 32'b11111111111111110101011010011100;
assign LUT_2[47873] = 32'b11111111111111110010010010110101;
assign LUT_2[47874] = 32'b11111111111111111100010011011000;
assign LUT_2[47875] = 32'b11111111111111111001001011110001;
assign LUT_2[47876] = 32'b11111111111111110001111000000100;
assign LUT_2[47877] = 32'b11111111111111101110110000011101;
assign LUT_2[47878] = 32'b11111111111111111000110001000000;
assign LUT_2[47879] = 32'b11111111111111110101101001011001;
assign LUT_2[47880] = 32'b11111111111111110000001011111001;
assign LUT_2[47881] = 32'b11111111111111101101000100010010;
assign LUT_2[47882] = 32'b11111111111111110111000100110101;
assign LUT_2[47883] = 32'b11111111111111110011111101001110;
assign LUT_2[47884] = 32'b11111111111111101100101001100001;
assign LUT_2[47885] = 32'b11111111111111101001100001111010;
assign LUT_2[47886] = 32'b11111111111111110011100010011101;
assign LUT_2[47887] = 32'b11111111111111110000011010110110;
assign LUT_2[47888] = 32'b11111111111111101111111110100110;
assign LUT_2[47889] = 32'b11111111111111101100110110111111;
assign LUT_2[47890] = 32'b11111111111111110110110111100010;
assign LUT_2[47891] = 32'b11111111111111110011101111111011;
assign LUT_2[47892] = 32'b11111111111111101100011100001110;
assign LUT_2[47893] = 32'b11111111111111101001010100100111;
assign LUT_2[47894] = 32'b11111111111111110011010101001010;
assign LUT_2[47895] = 32'b11111111111111110000001101100011;
assign LUT_2[47896] = 32'b11111111111111101010110000000011;
assign LUT_2[47897] = 32'b11111111111111100111101000011100;
assign LUT_2[47898] = 32'b11111111111111110001101000111111;
assign LUT_2[47899] = 32'b11111111111111101110100001011000;
assign LUT_2[47900] = 32'b11111111111111100111001101101011;
assign LUT_2[47901] = 32'b11111111111111100100000110000100;
assign LUT_2[47902] = 32'b11111111111111101110000110100111;
assign LUT_2[47903] = 32'b11111111111111101010111111000000;
assign LUT_2[47904] = 32'b11111111111111110101110110000101;
assign LUT_2[47905] = 32'b11111111111111110010101110011110;
assign LUT_2[47906] = 32'b11111111111111111100101111000001;
assign LUT_2[47907] = 32'b11111111111111111001100111011010;
assign LUT_2[47908] = 32'b11111111111111110010010011101101;
assign LUT_2[47909] = 32'b11111111111111101111001100000110;
assign LUT_2[47910] = 32'b11111111111111111001001100101001;
assign LUT_2[47911] = 32'b11111111111111110110000101000010;
assign LUT_2[47912] = 32'b11111111111111110000100111100010;
assign LUT_2[47913] = 32'b11111111111111101101011111111011;
assign LUT_2[47914] = 32'b11111111111111110111100000011110;
assign LUT_2[47915] = 32'b11111111111111110100011000110111;
assign LUT_2[47916] = 32'b11111111111111101101000101001010;
assign LUT_2[47917] = 32'b11111111111111101001111101100011;
assign LUT_2[47918] = 32'b11111111111111110011111110000110;
assign LUT_2[47919] = 32'b11111111111111110000110110011111;
assign LUT_2[47920] = 32'b11111111111111110000011010001111;
assign LUT_2[47921] = 32'b11111111111111101101010010101000;
assign LUT_2[47922] = 32'b11111111111111110111010011001011;
assign LUT_2[47923] = 32'b11111111111111110100001011100100;
assign LUT_2[47924] = 32'b11111111111111101100110111110111;
assign LUT_2[47925] = 32'b11111111111111101001110000010000;
assign LUT_2[47926] = 32'b11111111111111110011110000110011;
assign LUT_2[47927] = 32'b11111111111111110000101001001100;
assign LUT_2[47928] = 32'b11111111111111101011001011101100;
assign LUT_2[47929] = 32'b11111111111111101000000100000101;
assign LUT_2[47930] = 32'b11111111111111110010000100101000;
assign LUT_2[47931] = 32'b11111111111111101110111101000001;
assign LUT_2[47932] = 32'b11111111111111100111101001010100;
assign LUT_2[47933] = 32'b11111111111111100100100001101101;
assign LUT_2[47934] = 32'b11111111111111101110100010010000;
assign LUT_2[47935] = 32'b11111111111111101011011010101001;
assign LUT_2[47936] = 32'b11111111111111101101100010111111;
assign LUT_2[47937] = 32'b11111111111111101010011011011000;
assign LUT_2[47938] = 32'b11111111111111110100011011111011;
assign LUT_2[47939] = 32'b11111111111111110001010100010100;
assign LUT_2[47940] = 32'b11111111111111101010000000100111;
assign LUT_2[47941] = 32'b11111111111111100110111001000000;
assign LUT_2[47942] = 32'b11111111111111110000111001100011;
assign LUT_2[47943] = 32'b11111111111111101101110001111100;
assign LUT_2[47944] = 32'b11111111111111101000010100011100;
assign LUT_2[47945] = 32'b11111111111111100101001100110101;
assign LUT_2[47946] = 32'b11111111111111101111001101011000;
assign LUT_2[47947] = 32'b11111111111111101100000101110001;
assign LUT_2[47948] = 32'b11111111111111100100110010000100;
assign LUT_2[47949] = 32'b11111111111111100001101010011101;
assign LUT_2[47950] = 32'b11111111111111101011101011000000;
assign LUT_2[47951] = 32'b11111111111111101000100011011001;
assign LUT_2[47952] = 32'b11111111111111101000000111001001;
assign LUT_2[47953] = 32'b11111111111111100100111111100010;
assign LUT_2[47954] = 32'b11111111111111101111000000000101;
assign LUT_2[47955] = 32'b11111111111111101011111000011110;
assign LUT_2[47956] = 32'b11111111111111100100100100110001;
assign LUT_2[47957] = 32'b11111111111111100001011101001010;
assign LUT_2[47958] = 32'b11111111111111101011011101101101;
assign LUT_2[47959] = 32'b11111111111111101000010110000110;
assign LUT_2[47960] = 32'b11111111111111100010111000100110;
assign LUT_2[47961] = 32'b11111111111111011111110000111111;
assign LUT_2[47962] = 32'b11111111111111101001110001100010;
assign LUT_2[47963] = 32'b11111111111111100110101001111011;
assign LUT_2[47964] = 32'b11111111111111011111010110001110;
assign LUT_2[47965] = 32'b11111111111111011100001110100111;
assign LUT_2[47966] = 32'b11111111111111100110001111001010;
assign LUT_2[47967] = 32'b11111111111111100011000111100011;
assign LUT_2[47968] = 32'b11111111111111101101111110101000;
assign LUT_2[47969] = 32'b11111111111111101010110111000001;
assign LUT_2[47970] = 32'b11111111111111110100110111100100;
assign LUT_2[47971] = 32'b11111111111111110001101111111101;
assign LUT_2[47972] = 32'b11111111111111101010011100010000;
assign LUT_2[47973] = 32'b11111111111111100111010100101001;
assign LUT_2[47974] = 32'b11111111111111110001010101001100;
assign LUT_2[47975] = 32'b11111111111111101110001101100101;
assign LUT_2[47976] = 32'b11111111111111101000110000000101;
assign LUT_2[47977] = 32'b11111111111111100101101000011110;
assign LUT_2[47978] = 32'b11111111111111101111101001000001;
assign LUT_2[47979] = 32'b11111111111111101100100001011010;
assign LUT_2[47980] = 32'b11111111111111100101001101101101;
assign LUT_2[47981] = 32'b11111111111111100010000110000110;
assign LUT_2[47982] = 32'b11111111111111101100000110101001;
assign LUT_2[47983] = 32'b11111111111111101000111111000010;
assign LUT_2[47984] = 32'b11111111111111101000100010110010;
assign LUT_2[47985] = 32'b11111111111111100101011011001011;
assign LUT_2[47986] = 32'b11111111111111101111011011101110;
assign LUT_2[47987] = 32'b11111111111111101100010100000111;
assign LUT_2[47988] = 32'b11111111111111100101000000011010;
assign LUT_2[47989] = 32'b11111111111111100001111000110011;
assign LUT_2[47990] = 32'b11111111111111101011111001010110;
assign LUT_2[47991] = 32'b11111111111111101000110001101111;
assign LUT_2[47992] = 32'b11111111111111100011010100001111;
assign LUT_2[47993] = 32'b11111111111111100000001100101000;
assign LUT_2[47994] = 32'b11111111111111101010001101001011;
assign LUT_2[47995] = 32'b11111111111111100111000101100100;
assign LUT_2[47996] = 32'b11111111111111011111110001110111;
assign LUT_2[47997] = 32'b11111111111111011100101010010000;
assign LUT_2[47998] = 32'b11111111111111100110101010110011;
assign LUT_2[47999] = 32'b11111111111111100011100011001100;
assign LUT_2[48000] = 32'b11111111111111111001101110101011;
assign LUT_2[48001] = 32'b11111111111111110110100111000100;
assign LUT_2[48002] = 32'b00000000000000000000100111100111;
assign LUT_2[48003] = 32'b11111111111111111101100000000000;
assign LUT_2[48004] = 32'b11111111111111110110001100010011;
assign LUT_2[48005] = 32'b11111111111111110011000100101100;
assign LUT_2[48006] = 32'b11111111111111111101000101001111;
assign LUT_2[48007] = 32'b11111111111111111001111101101000;
assign LUT_2[48008] = 32'b11111111111111110100100000001000;
assign LUT_2[48009] = 32'b11111111111111110001011000100001;
assign LUT_2[48010] = 32'b11111111111111111011011001000100;
assign LUT_2[48011] = 32'b11111111111111111000010001011101;
assign LUT_2[48012] = 32'b11111111111111110000111101110000;
assign LUT_2[48013] = 32'b11111111111111101101110110001001;
assign LUT_2[48014] = 32'b11111111111111110111110110101100;
assign LUT_2[48015] = 32'b11111111111111110100101111000101;
assign LUT_2[48016] = 32'b11111111111111110100010010110101;
assign LUT_2[48017] = 32'b11111111111111110001001011001110;
assign LUT_2[48018] = 32'b11111111111111111011001011110001;
assign LUT_2[48019] = 32'b11111111111111111000000100001010;
assign LUT_2[48020] = 32'b11111111111111110000110000011101;
assign LUT_2[48021] = 32'b11111111111111101101101000110110;
assign LUT_2[48022] = 32'b11111111111111110111101001011001;
assign LUT_2[48023] = 32'b11111111111111110100100001110010;
assign LUT_2[48024] = 32'b11111111111111101111000100010010;
assign LUT_2[48025] = 32'b11111111111111101011111100101011;
assign LUT_2[48026] = 32'b11111111111111110101111101001110;
assign LUT_2[48027] = 32'b11111111111111110010110101100111;
assign LUT_2[48028] = 32'b11111111111111101011100001111010;
assign LUT_2[48029] = 32'b11111111111111101000011010010011;
assign LUT_2[48030] = 32'b11111111111111110010011010110110;
assign LUT_2[48031] = 32'b11111111111111101111010011001111;
assign LUT_2[48032] = 32'b11111111111111111010001010010100;
assign LUT_2[48033] = 32'b11111111111111110111000010101101;
assign LUT_2[48034] = 32'b00000000000000000001000011010000;
assign LUT_2[48035] = 32'b11111111111111111101111011101001;
assign LUT_2[48036] = 32'b11111111111111110110100111111100;
assign LUT_2[48037] = 32'b11111111111111110011100000010101;
assign LUT_2[48038] = 32'b11111111111111111101100000111000;
assign LUT_2[48039] = 32'b11111111111111111010011001010001;
assign LUT_2[48040] = 32'b11111111111111110100111011110001;
assign LUT_2[48041] = 32'b11111111111111110001110100001010;
assign LUT_2[48042] = 32'b11111111111111111011110100101101;
assign LUT_2[48043] = 32'b11111111111111111000101101000110;
assign LUT_2[48044] = 32'b11111111111111110001011001011001;
assign LUT_2[48045] = 32'b11111111111111101110010001110010;
assign LUT_2[48046] = 32'b11111111111111111000010010010101;
assign LUT_2[48047] = 32'b11111111111111110101001010101110;
assign LUT_2[48048] = 32'b11111111111111110100101110011110;
assign LUT_2[48049] = 32'b11111111111111110001100110110111;
assign LUT_2[48050] = 32'b11111111111111111011100111011010;
assign LUT_2[48051] = 32'b11111111111111111000011111110011;
assign LUT_2[48052] = 32'b11111111111111110001001100000110;
assign LUT_2[48053] = 32'b11111111111111101110000100011111;
assign LUT_2[48054] = 32'b11111111111111111000000101000010;
assign LUT_2[48055] = 32'b11111111111111110100111101011011;
assign LUT_2[48056] = 32'b11111111111111101111011111111011;
assign LUT_2[48057] = 32'b11111111111111101100011000010100;
assign LUT_2[48058] = 32'b11111111111111110110011000110111;
assign LUT_2[48059] = 32'b11111111111111110011010001010000;
assign LUT_2[48060] = 32'b11111111111111101011111101100011;
assign LUT_2[48061] = 32'b11111111111111101000110101111100;
assign LUT_2[48062] = 32'b11111111111111110010110110011111;
assign LUT_2[48063] = 32'b11111111111111101111101110111000;
assign LUT_2[48064] = 32'b11111111111111110001110111001110;
assign LUT_2[48065] = 32'b11111111111111101110101111100111;
assign LUT_2[48066] = 32'b11111111111111111000110000001010;
assign LUT_2[48067] = 32'b11111111111111110101101000100011;
assign LUT_2[48068] = 32'b11111111111111101110010100110110;
assign LUT_2[48069] = 32'b11111111111111101011001101001111;
assign LUT_2[48070] = 32'b11111111111111110101001101110010;
assign LUT_2[48071] = 32'b11111111111111110010000110001011;
assign LUT_2[48072] = 32'b11111111111111101100101000101011;
assign LUT_2[48073] = 32'b11111111111111101001100001000100;
assign LUT_2[48074] = 32'b11111111111111110011100001100111;
assign LUT_2[48075] = 32'b11111111111111110000011010000000;
assign LUT_2[48076] = 32'b11111111111111101001000110010011;
assign LUT_2[48077] = 32'b11111111111111100101111110101100;
assign LUT_2[48078] = 32'b11111111111111101111111111001111;
assign LUT_2[48079] = 32'b11111111111111101100110111101000;
assign LUT_2[48080] = 32'b11111111111111101100011011011000;
assign LUT_2[48081] = 32'b11111111111111101001010011110001;
assign LUT_2[48082] = 32'b11111111111111110011010100010100;
assign LUT_2[48083] = 32'b11111111111111110000001100101101;
assign LUT_2[48084] = 32'b11111111111111101000111001000000;
assign LUT_2[48085] = 32'b11111111111111100101110001011001;
assign LUT_2[48086] = 32'b11111111111111101111110001111100;
assign LUT_2[48087] = 32'b11111111111111101100101010010101;
assign LUT_2[48088] = 32'b11111111111111100111001100110101;
assign LUT_2[48089] = 32'b11111111111111100100000101001110;
assign LUT_2[48090] = 32'b11111111111111101110000101110001;
assign LUT_2[48091] = 32'b11111111111111101010111110001010;
assign LUT_2[48092] = 32'b11111111111111100011101010011101;
assign LUT_2[48093] = 32'b11111111111111100000100010110110;
assign LUT_2[48094] = 32'b11111111111111101010100011011001;
assign LUT_2[48095] = 32'b11111111111111100111011011110010;
assign LUT_2[48096] = 32'b11111111111111110010010010110111;
assign LUT_2[48097] = 32'b11111111111111101111001011010000;
assign LUT_2[48098] = 32'b11111111111111111001001011110011;
assign LUT_2[48099] = 32'b11111111111111110110000100001100;
assign LUT_2[48100] = 32'b11111111111111101110110000011111;
assign LUT_2[48101] = 32'b11111111111111101011101000111000;
assign LUT_2[48102] = 32'b11111111111111110101101001011011;
assign LUT_2[48103] = 32'b11111111111111110010100001110100;
assign LUT_2[48104] = 32'b11111111111111101101000100010100;
assign LUT_2[48105] = 32'b11111111111111101001111100101101;
assign LUT_2[48106] = 32'b11111111111111110011111101010000;
assign LUT_2[48107] = 32'b11111111111111110000110101101001;
assign LUT_2[48108] = 32'b11111111111111101001100001111100;
assign LUT_2[48109] = 32'b11111111111111100110011010010101;
assign LUT_2[48110] = 32'b11111111111111110000011010111000;
assign LUT_2[48111] = 32'b11111111111111101101010011010001;
assign LUT_2[48112] = 32'b11111111111111101100110111000001;
assign LUT_2[48113] = 32'b11111111111111101001101111011010;
assign LUT_2[48114] = 32'b11111111111111110011101111111101;
assign LUT_2[48115] = 32'b11111111111111110000101000010110;
assign LUT_2[48116] = 32'b11111111111111101001010100101001;
assign LUT_2[48117] = 32'b11111111111111100110001101000010;
assign LUT_2[48118] = 32'b11111111111111110000001101100101;
assign LUT_2[48119] = 32'b11111111111111101101000101111110;
assign LUT_2[48120] = 32'b11111111111111100111101000011110;
assign LUT_2[48121] = 32'b11111111111111100100100000110111;
assign LUT_2[48122] = 32'b11111111111111101110100001011010;
assign LUT_2[48123] = 32'b11111111111111101011011001110011;
assign LUT_2[48124] = 32'b11111111111111100100000110000110;
assign LUT_2[48125] = 32'b11111111111111100000111110011111;
assign LUT_2[48126] = 32'b11111111111111101010111111000010;
assign LUT_2[48127] = 32'b11111111111111100111110111011011;
assign LUT_2[48128] = 32'b11111111111111110011010110001001;
assign LUT_2[48129] = 32'b11111111111111110000001110100010;
assign LUT_2[48130] = 32'b11111111111111111010001111000101;
assign LUT_2[48131] = 32'b11111111111111110111000111011110;
assign LUT_2[48132] = 32'b11111111111111101111110011110001;
assign LUT_2[48133] = 32'b11111111111111101100101100001010;
assign LUT_2[48134] = 32'b11111111111111110110101100101101;
assign LUT_2[48135] = 32'b11111111111111110011100101000110;
assign LUT_2[48136] = 32'b11111111111111101110000111100110;
assign LUT_2[48137] = 32'b11111111111111101010111111111111;
assign LUT_2[48138] = 32'b11111111111111110101000000100010;
assign LUT_2[48139] = 32'b11111111111111110001111000111011;
assign LUT_2[48140] = 32'b11111111111111101010100101001110;
assign LUT_2[48141] = 32'b11111111111111100111011101100111;
assign LUT_2[48142] = 32'b11111111111111110001011110001010;
assign LUT_2[48143] = 32'b11111111111111101110010110100011;
assign LUT_2[48144] = 32'b11111111111111101101111010010011;
assign LUT_2[48145] = 32'b11111111111111101010110010101100;
assign LUT_2[48146] = 32'b11111111111111110100110011001111;
assign LUT_2[48147] = 32'b11111111111111110001101011101000;
assign LUT_2[48148] = 32'b11111111111111101010010111111011;
assign LUT_2[48149] = 32'b11111111111111100111010000010100;
assign LUT_2[48150] = 32'b11111111111111110001010000110111;
assign LUT_2[48151] = 32'b11111111111111101110001001010000;
assign LUT_2[48152] = 32'b11111111111111101000101011110000;
assign LUT_2[48153] = 32'b11111111111111100101100100001001;
assign LUT_2[48154] = 32'b11111111111111101111100100101100;
assign LUT_2[48155] = 32'b11111111111111101100011101000101;
assign LUT_2[48156] = 32'b11111111111111100101001001011000;
assign LUT_2[48157] = 32'b11111111111111100010000001110001;
assign LUT_2[48158] = 32'b11111111111111101100000010010100;
assign LUT_2[48159] = 32'b11111111111111101000111010101101;
assign LUT_2[48160] = 32'b11111111111111110011110001110010;
assign LUT_2[48161] = 32'b11111111111111110000101010001011;
assign LUT_2[48162] = 32'b11111111111111111010101010101110;
assign LUT_2[48163] = 32'b11111111111111110111100011000111;
assign LUT_2[48164] = 32'b11111111111111110000001111011010;
assign LUT_2[48165] = 32'b11111111111111101101000111110011;
assign LUT_2[48166] = 32'b11111111111111110111001000010110;
assign LUT_2[48167] = 32'b11111111111111110100000000101111;
assign LUT_2[48168] = 32'b11111111111111101110100011001111;
assign LUT_2[48169] = 32'b11111111111111101011011011101000;
assign LUT_2[48170] = 32'b11111111111111110101011100001011;
assign LUT_2[48171] = 32'b11111111111111110010010100100100;
assign LUT_2[48172] = 32'b11111111111111101011000000110111;
assign LUT_2[48173] = 32'b11111111111111100111111001010000;
assign LUT_2[48174] = 32'b11111111111111110001111001110011;
assign LUT_2[48175] = 32'b11111111111111101110110010001100;
assign LUT_2[48176] = 32'b11111111111111101110010101111100;
assign LUT_2[48177] = 32'b11111111111111101011001110010101;
assign LUT_2[48178] = 32'b11111111111111110101001110111000;
assign LUT_2[48179] = 32'b11111111111111110010000111010001;
assign LUT_2[48180] = 32'b11111111111111101010110011100100;
assign LUT_2[48181] = 32'b11111111111111100111101011111101;
assign LUT_2[48182] = 32'b11111111111111110001101100100000;
assign LUT_2[48183] = 32'b11111111111111101110100100111001;
assign LUT_2[48184] = 32'b11111111111111101001000111011001;
assign LUT_2[48185] = 32'b11111111111111100101111111110010;
assign LUT_2[48186] = 32'b11111111111111110000000000010101;
assign LUT_2[48187] = 32'b11111111111111101100111000101110;
assign LUT_2[48188] = 32'b11111111111111100101100101000001;
assign LUT_2[48189] = 32'b11111111111111100010011101011010;
assign LUT_2[48190] = 32'b11111111111111101100011101111101;
assign LUT_2[48191] = 32'b11111111111111101001010110010110;
assign LUT_2[48192] = 32'b11111111111111101011011110101100;
assign LUT_2[48193] = 32'b11111111111111101000010111000101;
assign LUT_2[48194] = 32'b11111111111111110010010111101000;
assign LUT_2[48195] = 32'b11111111111111101111010000000001;
assign LUT_2[48196] = 32'b11111111111111100111111100010100;
assign LUT_2[48197] = 32'b11111111111111100100110100101101;
assign LUT_2[48198] = 32'b11111111111111101110110101010000;
assign LUT_2[48199] = 32'b11111111111111101011101101101001;
assign LUT_2[48200] = 32'b11111111111111100110010000001001;
assign LUT_2[48201] = 32'b11111111111111100011001000100010;
assign LUT_2[48202] = 32'b11111111111111101101001001000101;
assign LUT_2[48203] = 32'b11111111111111101010000001011110;
assign LUT_2[48204] = 32'b11111111111111100010101101110001;
assign LUT_2[48205] = 32'b11111111111111011111100110001010;
assign LUT_2[48206] = 32'b11111111111111101001100110101101;
assign LUT_2[48207] = 32'b11111111111111100110011111000110;
assign LUT_2[48208] = 32'b11111111111111100110000010110110;
assign LUT_2[48209] = 32'b11111111111111100010111011001111;
assign LUT_2[48210] = 32'b11111111111111101100111011110010;
assign LUT_2[48211] = 32'b11111111111111101001110100001011;
assign LUT_2[48212] = 32'b11111111111111100010100000011110;
assign LUT_2[48213] = 32'b11111111111111011111011000110111;
assign LUT_2[48214] = 32'b11111111111111101001011001011010;
assign LUT_2[48215] = 32'b11111111111111100110010001110011;
assign LUT_2[48216] = 32'b11111111111111100000110100010011;
assign LUT_2[48217] = 32'b11111111111111011101101100101100;
assign LUT_2[48218] = 32'b11111111111111100111101101001111;
assign LUT_2[48219] = 32'b11111111111111100100100101101000;
assign LUT_2[48220] = 32'b11111111111111011101010001111011;
assign LUT_2[48221] = 32'b11111111111111011010001010010100;
assign LUT_2[48222] = 32'b11111111111111100100001010110111;
assign LUT_2[48223] = 32'b11111111111111100001000011010000;
assign LUT_2[48224] = 32'b11111111111111101011111010010101;
assign LUT_2[48225] = 32'b11111111111111101000110010101110;
assign LUT_2[48226] = 32'b11111111111111110010110011010001;
assign LUT_2[48227] = 32'b11111111111111101111101011101010;
assign LUT_2[48228] = 32'b11111111111111101000010111111101;
assign LUT_2[48229] = 32'b11111111111111100101010000010110;
assign LUT_2[48230] = 32'b11111111111111101111010000111001;
assign LUT_2[48231] = 32'b11111111111111101100001001010010;
assign LUT_2[48232] = 32'b11111111111111100110101011110010;
assign LUT_2[48233] = 32'b11111111111111100011100100001011;
assign LUT_2[48234] = 32'b11111111111111101101100100101110;
assign LUT_2[48235] = 32'b11111111111111101010011101000111;
assign LUT_2[48236] = 32'b11111111111111100011001001011010;
assign LUT_2[48237] = 32'b11111111111111100000000001110011;
assign LUT_2[48238] = 32'b11111111111111101010000010010110;
assign LUT_2[48239] = 32'b11111111111111100110111010101111;
assign LUT_2[48240] = 32'b11111111111111100110011110011111;
assign LUT_2[48241] = 32'b11111111111111100011010110111000;
assign LUT_2[48242] = 32'b11111111111111101101010111011011;
assign LUT_2[48243] = 32'b11111111111111101010001111110100;
assign LUT_2[48244] = 32'b11111111111111100010111100000111;
assign LUT_2[48245] = 32'b11111111111111011111110100100000;
assign LUT_2[48246] = 32'b11111111111111101001110101000011;
assign LUT_2[48247] = 32'b11111111111111100110101101011100;
assign LUT_2[48248] = 32'b11111111111111100001001111111100;
assign LUT_2[48249] = 32'b11111111111111011110001000010101;
assign LUT_2[48250] = 32'b11111111111111101000001000111000;
assign LUT_2[48251] = 32'b11111111111111100101000001010001;
assign LUT_2[48252] = 32'b11111111111111011101101101100100;
assign LUT_2[48253] = 32'b11111111111111011010100101111101;
assign LUT_2[48254] = 32'b11111111111111100100100110100000;
assign LUT_2[48255] = 32'b11111111111111100001011110111001;
assign LUT_2[48256] = 32'b11111111111111110111101010011000;
assign LUT_2[48257] = 32'b11111111111111110100100010110001;
assign LUT_2[48258] = 32'b11111111111111111110100011010100;
assign LUT_2[48259] = 32'b11111111111111111011011011101101;
assign LUT_2[48260] = 32'b11111111111111110100001000000000;
assign LUT_2[48261] = 32'b11111111111111110001000000011001;
assign LUT_2[48262] = 32'b11111111111111111011000000111100;
assign LUT_2[48263] = 32'b11111111111111110111111001010101;
assign LUT_2[48264] = 32'b11111111111111110010011011110101;
assign LUT_2[48265] = 32'b11111111111111101111010100001110;
assign LUT_2[48266] = 32'b11111111111111111001010100110001;
assign LUT_2[48267] = 32'b11111111111111110110001101001010;
assign LUT_2[48268] = 32'b11111111111111101110111001011101;
assign LUT_2[48269] = 32'b11111111111111101011110001110110;
assign LUT_2[48270] = 32'b11111111111111110101110010011001;
assign LUT_2[48271] = 32'b11111111111111110010101010110010;
assign LUT_2[48272] = 32'b11111111111111110010001110100010;
assign LUT_2[48273] = 32'b11111111111111101111000110111011;
assign LUT_2[48274] = 32'b11111111111111111001000111011110;
assign LUT_2[48275] = 32'b11111111111111110101111111110111;
assign LUT_2[48276] = 32'b11111111111111101110101100001010;
assign LUT_2[48277] = 32'b11111111111111101011100100100011;
assign LUT_2[48278] = 32'b11111111111111110101100101000110;
assign LUT_2[48279] = 32'b11111111111111110010011101011111;
assign LUT_2[48280] = 32'b11111111111111101100111111111111;
assign LUT_2[48281] = 32'b11111111111111101001111000011000;
assign LUT_2[48282] = 32'b11111111111111110011111000111011;
assign LUT_2[48283] = 32'b11111111111111110000110001010100;
assign LUT_2[48284] = 32'b11111111111111101001011101100111;
assign LUT_2[48285] = 32'b11111111111111100110010110000000;
assign LUT_2[48286] = 32'b11111111111111110000010110100011;
assign LUT_2[48287] = 32'b11111111111111101101001110111100;
assign LUT_2[48288] = 32'b11111111111111111000000110000001;
assign LUT_2[48289] = 32'b11111111111111110100111110011010;
assign LUT_2[48290] = 32'b11111111111111111110111110111101;
assign LUT_2[48291] = 32'b11111111111111111011110111010110;
assign LUT_2[48292] = 32'b11111111111111110100100011101001;
assign LUT_2[48293] = 32'b11111111111111110001011100000010;
assign LUT_2[48294] = 32'b11111111111111111011011100100101;
assign LUT_2[48295] = 32'b11111111111111111000010100111110;
assign LUT_2[48296] = 32'b11111111111111110010110111011110;
assign LUT_2[48297] = 32'b11111111111111101111101111110111;
assign LUT_2[48298] = 32'b11111111111111111001110000011010;
assign LUT_2[48299] = 32'b11111111111111110110101000110011;
assign LUT_2[48300] = 32'b11111111111111101111010101000110;
assign LUT_2[48301] = 32'b11111111111111101100001101011111;
assign LUT_2[48302] = 32'b11111111111111110110001110000010;
assign LUT_2[48303] = 32'b11111111111111110011000110011011;
assign LUT_2[48304] = 32'b11111111111111110010101010001011;
assign LUT_2[48305] = 32'b11111111111111101111100010100100;
assign LUT_2[48306] = 32'b11111111111111111001100011000111;
assign LUT_2[48307] = 32'b11111111111111110110011011100000;
assign LUT_2[48308] = 32'b11111111111111101111000111110011;
assign LUT_2[48309] = 32'b11111111111111101100000000001100;
assign LUT_2[48310] = 32'b11111111111111110110000000101111;
assign LUT_2[48311] = 32'b11111111111111110010111001001000;
assign LUT_2[48312] = 32'b11111111111111101101011011101000;
assign LUT_2[48313] = 32'b11111111111111101010010100000001;
assign LUT_2[48314] = 32'b11111111111111110100010100100100;
assign LUT_2[48315] = 32'b11111111111111110001001100111101;
assign LUT_2[48316] = 32'b11111111111111101001111001010000;
assign LUT_2[48317] = 32'b11111111111111100110110001101001;
assign LUT_2[48318] = 32'b11111111111111110000110010001100;
assign LUT_2[48319] = 32'b11111111111111101101101010100101;
assign LUT_2[48320] = 32'b11111111111111101111110010111011;
assign LUT_2[48321] = 32'b11111111111111101100101011010100;
assign LUT_2[48322] = 32'b11111111111111110110101011110111;
assign LUT_2[48323] = 32'b11111111111111110011100100010000;
assign LUT_2[48324] = 32'b11111111111111101100010000100011;
assign LUT_2[48325] = 32'b11111111111111101001001000111100;
assign LUT_2[48326] = 32'b11111111111111110011001001011111;
assign LUT_2[48327] = 32'b11111111111111110000000001111000;
assign LUT_2[48328] = 32'b11111111111111101010100100011000;
assign LUT_2[48329] = 32'b11111111111111100111011100110001;
assign LUT_2[48330] = 32'b11111111111111110001011101010100;
assign LUT_2[48331] = 32'b11111111111111101110010101101101;
assign LUT_2[48332] = 32'b11111111111111100111000010000000;
assign LUT_2[48333] = 32'b11111111111111100011111010011001;
assign LUT_2[48334] = 32'b11111111111111101101111010111100;
assign LUT_2[48335] = 32'b11111111111111101010110011010101;
assign LUT_2[48336] = 32'b11111111111111101010010111000101;
assign LUT_2[48337] = 32'b11111111111111100111001111011110;
assign LUT_2[48338] = 32'b11111111111111110001010000000001;
assign LUT_2[48339] = 32'b11111111111111101110001000011010;
assign LUT_2[48340] = 32'b11111111111111100110110100101101;
assign LUT_2[48341] = 32'b11111111111111100011101101000110;
assign LUT_2[48342] = 32'b11111111111111101101101101101001;
assign LUT_2[48343] = 32'b11111111111111101010100110000010;
assign LUT_2[48344] = 32'b11111111111111100101001000100010;
assign LUT_2[48345] = 32'b11111111111111100010000000111011;
assign LUT_2[48346] = 32'b11111111111111101100000001011110;
assign LUT_2[48347] = 32'b11111111111111101000111001110111;
assign LUT_2[48348] = 32'b11111111111111100001100110001010;
assign LUT_2[48349] = 32'b11111111111111011110011110100011;
assign LUT_2[48350] = 32'b11111111111111101000011111000110;
assign LUT_2[48351] = 32'b11111111111111100101010111011111;
assign LUT_2[48352] = 32'b11111111111111110000001110100100;
assign LUT_2[48353] = 32'b11111111111111101101000110111101;
assign LUT_2[48354] = 32'b11111111111111110111000111100000;
assign LUT_2[48355] = 32'b11111111111111110011111111111001;
assign LUT_2[48356] = 32'b11111111111111101100101100001100;
assign LUT_2[48357] = 32'b11111111111111101001100100100101;
assign LUT_2[48358] = 32'b11111111111111110011100101001000;
assign LUT_2[48359] = 32'b11111111111111110000011101100001;
assign LUT_2[48360] = 32'b11111111111111101011000000000001;
assign LUT_2[48361] = 32'b11111111111111100111111000011010;
assign LUT_2[48362] = 32'b11111111111111110001111000111101;
assign LUT_2[48363] = 32'b11111111111111101110110001010110;
assign LUT_2[48364] = 32'b11111111111111100111011101101001;
assign LUT_2[48365] = 32'b11111111111111100100010110000010;
assign LUT_2[48366] = 32'b11111111111111101110010110100101;
assign LUT_2[48367] = 32'b11111111111111101011001110111110;
assign LUT_2[48368] = 32'b11111111111111101010110010101110;
assign LUT_2[48369] = 32'b11111111111111100111101011000111;
assign LUT_2[48370] = 32'b11111111111111110001101011101010;
assign LUT_2[48371] = 32'b11111111111111101110100100000011;
assign LUT_2[48372] = 32'b11111111111111100111010000010110;
assign LUT_2[48373] = 32'b11111111111111100100001000101111;
assign LUT_2[48374] = 32'b11111111111111101110001001010010;
assign LUT_2[48375] = 32'b11111111111111101011000001101011;
assign LUT_2[48376] = 32'b11111111111111100101100100001011;
assign LUT_2[48377] = 32'b11111111111111100010011100100100;
assign LUT_2[48378] = 32'b11111111111111101100011101000111;
assign LUT_2[48379] = 32'b11111111111111101001010101100000;
assign LUT_2[48380] = 32'b11111111111111100010000001110011;
assign LUT_2[48381] = 32'b11111111111111011110111010001100;
assign LUT_2[48382] = 32'b11111111111111101000111010101111;
assign LUT_2[48383] = 32'b11111111111111100101110011001000;
assign LUT_2[48384] = 32'b11111111111111110111010100101111;
assign LUT_2[48385] = 32'b11111111111111110100001101001000;
assign LUT_2[48386] = 32'b11111111111111111110001101101011;
assign LUT_2[48387] = 32'b11111111111111111011000110000100;
assign LUT_2[48388] = 32'b11111111111111110011110010010111;
assign LUT_2[48389] = 32'b11111111111111110000101010110000;
assign LUT_2[48390] = 32'b11111111111111111010101011010011;
assign LUT_2[48391] = 32'b11111111111111110111100011101100;
assign LUT_2[48392] = 32'b11111111111111110010000110001100;
assign LUT_2[48393] = 32'b11111111111111101110111110100101;
assign LUT_2[48394] = 32'b11111111111111111000111111001000;
assign LUT_2[48395] = 32'b11111111111111110101110111100001;
assign LUT_2[48396] = 32'b11111111111111101110100011110100;
assign LUT_2[48397] = 32'b11111111111111101011011100001101;
assign LUT_2[48398] = 32'b11111111111111110101011100110000;
assign LUT_2[48399] = 32'b11111111111111110010010101001001;
assign LUT_2[48400] = 32'b11111111111111110001111000111001;
assign LUT_2[48401] = 32'b11111111111111101110110001010010;
assign LUT_2[48402] = 32'b11111111111111111000110001110101;
assign LUT_2[48403] = 32'b11111111111111110101101010001110;
assign LUT_2[48404] = 32'b11111111111111101110010110100001;
assign LUT_2[48405] = 32'b11111111111111101011001110111010;
assign LUT_2[48406] = 32'b11111111111111110101001111011101;
assign LUT_2[48407] = 32'b11111111111111110010000111110110;
assign LUT_2[48408] = 32'b11111111111111101100101010010110;
assign LUT_2[48409] = 32'b11111111111111101001100010101111;
assign LUT_2[48410] = 32'b11111111111111110011100011010010;
assign LUT_2[48411] = 32'b11111111111111110000011011101011;
assign LUT_2[48412] = 32'b11111111111111101001000111111110;
assign LUT_2[48413] = 32'b11111111111111100110000000010111;
assign LUT_2[48414] = 32'b11111111111111110000000000111010;
assign LUT_2[48415] = 32'b11111111111111101100111001010011;
assign LUT_2[48416] = 32'b11111111111111110111110000011000;
assign LUT_2[48417] = 32'b11111111111111110100101000110001;
assign LUT_2[48418] = 32'b11111111111111111110101001010100;
assign LUT_2[48419] = 32'b11111111111111111011100001101101;
assign LUT_2[48420] = 32'b11111111111111110100001110000000;
assign LUT_2[48421] = 32'b11111111111111110001000110011001;
assign LUT_2[48422] = 32'b11111111111111111011000110111100;
assign LUT_2[48423] = 32'b11111111111111110111111111010101;
assign LUT_2[48424] = 32'b11111111111111110010100001110101;
assign LUT_2[48425] = 32'b11111111111111101111011010001110;
assign LUT_2[48426] = 32'b11111111111111111001011010110001;
assign LUT_2[48427] = 32'b11111111111111110110010011001010;
assign LUT_2[48428] = 32'b11111111111111101110111111011101;
assign LUT_2[48429] = 32'b11111111111111101011110111110110;
assign LUT_2[48430] = 32'b11111111111111110101111000011001;
assign LUT_2[48431] = 32'b11111111111111110010110000110010;
assign LUT_2[48432] = 32'b11111111111111110010010100100010;
assign LUT_2[48433] = 32'b11111111111111101111001100111011;
assign LUT_2[48434] = 32'b11111111111111111001001101011110;
assign LUT_2[48435] = 32'b11111111111111110110000101110111;
assign LUT_2[48436] = 32'b11111111111111101110110010001010;
assign LUT_2[48437] = 32'b11111111111111101011101010100011;
assign LUT_2[48438] = 32'b11111111111111110101101011000110;
assign LUT_2[48439] = 32'b11111111111111110010100011011111;
assign LUT_2[48440] = 32'b11111111111111101101000101111111;
assign LUT_2[48441] = 32'b11111111111111101001111110011000;
assign LUT_2[48442] = 32'b11111111111111110011111110111011;
assign LUT_2[48443] = 32'b11111111111111110000110111010100;
assign LUT_2[48444] = 32'b11111111111111101001100011100111;
assign LUT_2[48445] = 32'b11111111111111100110011100000000;
assign LUT_2[48446] = 32'b11111111111111110000011100100011;
assign LUT_2[48447] = 32'b11111111111111101101010100111100;
assign LUT_2[48448] = 32'b11111111111111101111011101010010;
assign LUT_2[48449] = 32'b11111111111111101100010101101011;
assign LUT_2[48450] = 32'b11111111111111110110010110001110;
assign LUT_2[48451] = 32'b11111111111111110011001110100111;
assign LUT_2[48452] = 32'b11111111111111101011111010111010;
assign LUT_2[48453] = 32'b11111111111111101000110011010011;
assign LUT_2[48454] = 32'b11111111111111110010110011110110;
assign LUT_2[48455] = 32'b11111111111111101111101100001111;
assign LUT_2[48456] = 32'b11111111111111101010001110101111;
assign LUT_2[48457] = 32'b11111111111111100111000111001000;
assign LUT_2[48458] = 32'b11111111111111110001000111101011;
assign LUT_2[48459] = 32'b11111111111111101110000000000100;
assign LUT_2[48460] = 32'b11111111111111100110101100010111;
assign LUT_2[48461] = 32'b11111111111111100011100100110000;
assign LUT_2[48462] = 32'b11111111111111101101100101010011;
assign LUT_2[48463] = 32'b11111111111111101010011101101100;
assign LUT_2[48464] = 32'b11111111111111101010000001011100;
assign LUT_2[48465] = 32'b11111111111111100110111001110101;
assign LUT_2[48466] = 32'b11111111111111110000111010011000;
assign LUT_2[48467] = 32'b11111111111111101101110010110001;
assign LUT_2[48468] = 32'b11111111111111100110011111000100;
assign LUT_2[48469] = 32'b11111111111111100011010111011101;
assign LUT_2[48470] = 32'b11111111111111101101011000000000;
assign LUT_2[48471] = 32'b11111111111111101010010000011001;
assign LUT_2[48472] = 32'b11111111111111100100110010111001;
assign LUT_2[48473] = 32'b11111111111111100001101011010010;
assign LUT_2[48474] = 32'b11111111111111101011101011110101;
assign LUT_2[48475] = 32'b11111111111111101000100100001110;
assign LUT_2[48476] = 32'b11111111111111100001010000100001;
assign LUT_2[48477] = 32'b11111111111111011110001000111010;
assign LUT_2[48478] = 32'b11111111111111101000001001011101;
assign LUT_2[48479] = 32'b11111111111111100101000001110110;
assign LUT_2[48480] = 32'b11111111111111101111111000111011;
assign LUT_2[48481] = 32'b11111111111111101100110001010100;
assign LUT_2[48482] = 32'b11111111111111110110110001110111;
assign LUT_2[48483] = 32'b11111111111111110011101010010000;
assign LUT_2[48484] = 32'b11111111111111101100010110100011;
assign LUT_2[48485] = 32'b11111111111111101001001110111100;
assign LUT_2[48486] = 32'b11111111111111110011001111011111;
assign LUT_2[48487] = 32'b11111111111111110000000111111000;
assign LUT_2[48488] = 32'b11111111111111101010101010011000;
assign LUT_2[48489] = 32'b11111111111111100111100010110001;
assign LUT_2[48490] = 32'b11111111111111110001100011010100;
assign LUT_2[48491] = 32'b11111111111111101110011011101101;
assign LUT_2[48492] = 32'b11111111111111100111001000000000;
assign LUT_2[48493] = 32'b11111111111111100100000000011001;
assign LUT_2[48494] = 32'b11111111111111101110000000111100;
assign LUT_2[48495] = 32'b11111111111111101010111001010101;
assign LUT_2[48496] = 32'b11111111111111101010011101000101;
assign LUT_2[48497] = 32'b11111111111111100111010101011110;
assign LUT_2[48498] = 32'b11111111111111110001010110000001;
assign LUT_2[48499] = 32'b11111111111111101110001110011010;
assign LUT_2[48500] = 32'b11111111111111100110111010101101;
assign LUT_2[48501] = 32'b11111111111111100011110011000110;
assign LUT_2[48502] = 32'b11111111111111101101110011101001;
assign LUT_2[48503] = 32'b11111111111111101010101100000010;
assign LUT_2[48504] = 32'b11111111111111100101001110100010;
assign LUT_2[48505] = 32'b11111111111111100010000110111011;
assign LUT_2[48506] = 32'b11111111111111101100000111011110;
assign LUT_2[48507] = 32'b11111111111111101000111111110111;
assign LUT_2[48508] = 32'b11111111111111100001101100001010;
assign LUT_2[48509] = 32'b11111111111111011110100100100011;
assign LUT_2[48510] = 32'b11111111111111101000100101000110;
assign LUT_2[48511] = 32'b11111111111111100101011101011111;
assign LUT_2[48512] = 32'b11111111111111111011101000111110;
assign LUT_2[48513] = 32'b11111111111111111000100001010111;
assign LUT_2[48514] = 32'b00000000000000000010100001111010;
assign LUT_2[48515] = 32'b11111111111111111111011010010011;
assign LUT_2[48516] = 32'b11111111111111111000000110100110;
assign LUT_2[48517] = 32'b11111111111111110100111110111111;
assign LUT_2[48518] = 32'b11111111111111111110111111100010;
assign LUT_2[48519] = 32'b11111111111111111011110111111011;
assign LUT_2[48520] = 32'b11111111111111110110011010011011;
assign LUT_2[48521] = 32'b11111111111111110011010010110100;
assign LUT_2[48522] = 32'b11111111111111111101010011010111;
assign LUT_2[48523] = 32'b11111111111111111010001011110000;
assign LUT_2[48524] = 32'b11111111111111110010111000000011;
assign LUT_2[48525] = 32'b11111111111111101111110000011100;
assign LUT_2[48526] = 32'b11111111111111111001110000111111;
assign LUT_2[48527] = 32'b11111111111111110110101001011000;
assign LUT_2[48528] = 32'b11111111111111110110001101001000;
assign LUT_2[48529] = 32'b11111111111111110011000101100001;
assign LUT_2[48530] = 32'b11111111111111111101000110000100;
assign LUT_2[48531] = 32'b11111111111111111001111110011101;
assign LUT_2[48532] = 32'b11111111111111110010101010110000;
assign LUT_2[48533] = 32'b11111111111111101111100011001001;
assign LUT_2[48534] = 32'b11111111111111111001100011101100;
assign LUT_2[48535] = 32'b11111111111111110110011100000101;
assign LUT_2[48536] = 32'b11111111111111110000111110100101;
assign LUT_2[48537] = 32'b11111111111111101101110110111110;
assign LUT_2[48538] = 32'b11111111111111110111110111100001;
assign LUT_2[48539] = 32'b11111111111111110100101111111010;
assign LUT_2[48540] = 32'b11111111111111101101011100001101;
assign LUT_2[48541] = 32'b11111111111111101010010100100110;
assign LUT_2[48542] = 32'b11111111111111110100010101001001;
assign LUT_2[48543] = 32'b11111111111111110001001101100010;
assign LUT_2[48544] = 32'b11111111111111111100000100100111;
assign LUT_2[48545] = 32'b11111111111111111000111101000000;
assign LUT_2[48546] = 32'b00000000000000000010111101100011;
assign LUT_2[48547] = 32'b11111111111111111111110101111100;
assign LUT_2[48548] = 32'b11111111111111111000100010001111;
assign LUT_2[48549] = 32'b11111111111111110101011010101000;
assign LUT_2[48550] = 32'b11111111111111111111011011001011;
assign LUT_2[48551] = 32'b11111111111111111100010011100100;
assign LUT_2[48552] = 32'b11111111111111110110110110000100;
assign LUT_2[48553] = 32'b11111111111111110011101110011101;
assign LUT_2[48554] = 32'b11111111111111111101101111000000;
assign LUT_2[48555] = 32'b11111111111111111010100111011001;
assign LUT_2[48556] = 32'b11111111111111110011010011101100;
assign LUT_2[48557] = 32'b11111111111111110000001100000101;
assign LUT_2[48558] = 32'b11111111111111111010001100101000;
assign LUT_2[48559] = 32'b11111111111111110111000101000001;
assign LUT_2[48560] = 32'b11111111111111110110101000110001;
assign LUT_2[48561] = 32'b11111111111111110011100001001010;
assign LUT_2[48562] = 32'b11111111111111111101100001101101;
assign LUT_2[48563] = 32'b11111111111111111010011010000110;
assign LUT_2[48564] = 32'b11111111111111110011000110011001;
assign LUT_2[48565] = 32'b11111111111111101111111110110010;
assign LUT_2[48566] = 32'b11111111111111111001111111010101;
assign LUT_2[48567] = 32'b11111111111111110110110111101110;
assign LUT_2[48568] = 32'b11111111111111110001011010001110;
assign LUT_2[48569] = 32'b11111111111111101110010010100111;
assign LUT_2[48570] = 32'b11111111111111111000010011001010;
assign LUT_2[48571] = 32'b11111111111111110101001011100011;
assign LUT_2[48572] = 32'b11111111111111101101110111110110;
assign LUT_2[48573] = 32'b11111111111111101010110000001111;
assign LUT_2[48574] = 32'b11111111111111110100110000110010;
assign LUT_2[48575] = 32'b11111111111111110001101001001011;
assign LUT_2[48576] = 32'b11111111111111110011110001100001;
assign LUT_2[48577] = 32'b11111111111111110000101001111010;
assign LUT_2[48578] = 32'b11111111111111111010101010011101;
assign LUT_2[48579] = 32'b11111111111111110111100010110110;
assign LUT_2[48580] = 32'b11111111111111110000001111001001;
assign LUT_2[48581] = 32'b11111111111111101101000111100010;
assign LUT_2[48582] = 32'b11111111111111110111001000000101;
assign LUT_2[48583] = 32'b11111111111111110100000000011110;
assign LUT_2[48584] = 32'b11111111111111101110100010111110;
assign LUT_2[48585] = 32'b11111111111111101011011011010111;
assign LUT_2[48586] = 32'b11111111111111110101011011111010;
assign LUT_2[48587] = 32'b11111111111111110010010100010011;
assign LUT_2[48588] = 32'b11111111111111101011000000100110;
assign LUT_2[48589] = 32'b11111111111111100111111000111111;
assign LUT_2[48590] = 32'b11111111111111110001111001100010;
assign LUT_2[48591] = 32'b11111111111111101110110001111011;
assign LUT_2[48592] = 32'b11111111111111101110010101101011;
assign LUT_2[48593] = 32'b11111111111111101011001110000100;
assign LUT_2[48594] = 32'b11111111111111110101001110100111;
assign LUT_2[48595] = 32'b11111111111111110010000111000000;
assign LUT_2[48596] = 32'b11111111111111101010110011010011;
assign LUT_2[48597] = 32'b11111111111111100111101011101100;
assign LUT_2[48598] = 32'b11111111111111110001101100001111;
assign LUT_2[48599] = 32'b11111111111111101110100100101000;
assign LUT_2[48600] = 32'b11111111111111101001000111001000;
assign LUT_2[48601] = 32'b11111111111111100101111111100001;
assign LUT_2[48602] = 32'b11111111111111110000000000000100;
assign LUT_2[48603] = 32'b11111111111111101100111000011101;
assign LUT_2[48604] = 32'b11111111111111100101100100110000;
assign LUT_2[48605] = 32'b11111111111111100010011101001001;
assign LUT_2[48606] = 32'b11111111111111101100011101101100;
assign LUT_2[48607] = 32'b11111111111111101001010110000101;
assign LUT_2[48608] = 32'b11111111111111110100001101001010;
assign LUT_2[48609] = 32'b11111111111111110001000101100011;
assign LUT_2[48610] = 32'b11111111111111111011000110000110;
assign LUT_2[48611] = 32'b11111111111111110111111110011111;
assign LUT_2[48612] = 32'b11111111111111110000101010110010;
assign LUT_2[48613] = 32'b11111111111111101101100011001011;
assign LUT_2[48614] = 32'b11111111111111110111100011101110;
assign LUT_2[48615] = 32'b11111111111111110100011100000111;
assign LUT_2[48616] = 32'b11111111111111101110111110100111;
assign LUT_2[48617] = 32'b11111111111111101011110111000000;
assign LUT_2[48618] = 32'b11111111111111110101110111100011;
assign LUT_2[48619] = 32'b11111111111111110010101111111100;
assign LUT_2[48620] = 32'b11111111111111101011011100001111;
assign LUT_2[48621] = 32'b11111111111111101000010100101000;
assign LUT_2[48622] = 32'b11111111111111110010010101001011;
assign LUT_2[48623] = 32'b11111111111111101111001101100100;
assign LUT_2[48624] = 32'b11111111111111101110110001010100;
assign LUT_2[48625] = 32'b11111111111111101011101001101101;
assign LUT_2[48626] = 32'b11111111111111110101101010010000;
assign LUT_2[48627] = 32'b11111111111111110010100010101001;
assign LUT_2[48628] = 32'b11111111111111101011001110111100;
assign LUT_2[48629] = 32'b11111111111111101000000111010101;
assign LUT_2[48630] = 32'b11111111111111110010000111111000;
assign LUT_2[48631] = 32'b11111111111111101111000000010001;
assign LUT_2[48632] = 32'b11111111111111101001100010110001;
assign LUT_2[48633] = 32'b11111111111111100110011011001010;
assign LUT_2[48634] = 32'b11111111111111110000011011101101;
assign LUT_2[48635] = 32'b11111111111111101101010100000110;
assign LUT_2[48636] = 32'b11111111111111100110000000011001;
assign LUT_2[48637] = 32'b11111111111111100010111000110010;
assign LUT_2[48638] = 32'b11111111111111101100111001010101;
assign LUT_2[48639] = 32'b11111111111111101001110001101110;
assign LUT_2[48640] = 32'b11111111111111111000000111111011;
assign LUT_2[48641] = 32'b11111111111111110101000000010100;
assign LUT_2[48642] = 32'b11111111111111111111000000110111;
assign LUT_2[48643] = 32'b11111111111111111011111001010000;
assign LUT_2[48644] = 32'b11111111111111110100100101100011;
assign LUT_2[48645] = 32'b11111111111111110001011101111100;
assign LUT_2[48646] = 32'b11111111111111111011011110011111;
assign LUT_2[48647] = 32'b11111111111111111000010110111000;
assign LUT_2[48648] = 32'b11111111111111110010111001011000;
assign LUT_2[48649] = 32'b11111111111111101111110001110001;
assign LUT_2[48650] = 32'b11111111111111111001110010010100;
assign LUT_2[48651] = 32'b11111111111111110110101010101101;
assign LUT_2[48652] = 32'b11111111111111101111010111000000;
assign LUT_2[48653] = 32'b11111111111111101100001111011001;
assign LUT_2[48654] = 32'b11111111111111110110001111111100;
assign LUT_2[48655] = 32'b11111111111111110011001000010101;
assign LUT_2[48656] = 32'b11111111111111110010101100000101;
assign LUT_2[48657] = 32'b11111111111111101111100100011110;
assign LUT_2[48658] = 32'b11111111111111111001100101000001;
assign LUT_2[48659] = 32'b11111111111111110110011101011010;
assign LUT_2[48660] = 32'b11111111111111101111001001101101;
assign LUT_2[48661] = 32'b11111111111111101100000010000110;
assign LUT_2[48662] = 32'b11111111111111110110000010101001;
assign LUT_2[48663] = 32'b11111111111111110010111011000010;
assign LUT_2[48664] = 32'b11111111111111101101011101100010;
assign LUT_2[48665] = 32'b11111111111111101010010101111011;
assign LUT_2[48666] = 32'b11111111111111110100010110011110;
assign LUT_2[48667] = 32'b11111111111111110001001110110111;
assign LUT_2[48668] = 32'b11111111111111101001111011001010;
assign LUT_2[48669] = 32'b11111111111111100110110011100011;
assign LUT_2[48670] = 32'b11111111111111110000110100000110;
assign LUT_2[48671] = 32'b11111111111111101101101100011111;
assign LUT_2[48672] = 32'b11111111111111111000100011100100;
assign LUT_2[48673] = 32'b11111111111111110101011011111101;
assign LUT_2[48674] = 32'b11111111111111111111011100100000;
assign LUT_2[48675] = 32'b11111111111111111100010100111001;
assign LUT_2[48676] = 32'b11111111111111110101000001001100;
assign LUT_2[48677] = 32'b11111111111111110001111001100101;
assign LUT_2[48678] = 32'b11111111111111111011111010001000;
assign LUT_2[48679] = 32'b11111111111111111000110010100001;
assign LUT_2[48680] = 32'b11111111111111110011010101000001;
assign LUT_2[48681] = 32'b11111111111111110000001101011010;
assign LUT_2[48682] = 32'b11111111111111111010001101111101;
assign LUT_2[48683] = 32'b11111111111111110111000110010110;
assign LUT_2[48684] = 32'b11111111111111101111110010101001;
assign LUT_2[48685] = 32'b11111111111111101100101011000010;
assign LUT_2[48686] = 32'b11111111111111110110101011100101;
assign LUT_2[48687] = 32'b11111111111111110011100011111110;
assign LUT_2[48688] = 32'b11111111111111110011000111101110;
assign LUT_2[48689] = 32'b11111111111111110000000000000111;
assign LUT_2[48690] = 32'b11111111111111111010000000101010;
assign LUT_2[48691] = 32'b11111111111111110110111001000011;
assign LUT_2[48692] = 32'b11111111111111101111100101010110;
assign LUT_2[48693] = 32'b11111111111111101100011101101111;
assign LUT_2[48694] = 32'b11111111111111110110011110010010;
assign LUT_2[48695] = 32'b11111111111111110011010110101011;
assign LUT_2[48696] = 32'b11111111111111101101111001001011;
assign LUT_2[48697] = 32'b11111111111111101010110001100100;
assign LUT_2[48698] = 32'b11111111111111110100110010000111;
assign LUT_2[48699] = 32'b11111111111111110001101010100000;
assign LUT_2[48700] = 32'b11111111111111101010010110110011;
assign LUT_2[48701] = 32'b11111111111111100111001111001100;
assign LUT_2[48702] = 32'b11111111111111110001001111101111;
assign LUT_2[48703] = 32'b11111111111111101110001000001000;
assign LUT_2[48704] = 32'b11111111111111110000010000011110;
assign LUT_2[48705] = 32'b11111111111111101101001000110111;
assign LUT_2[48706] = 32'b11111111111111110111001001011010;
assign LUT_2[48707] = 32'b11111111111111110100000001110011;
assign LUT_2[48708] = 32'b11111111111111101100101110000110;
assign LUT_2[48709] = 32'b11111111111111101001100110011111;
assign LUT_2[48710] = 32'b11111111111111110011100111000010;
assign LUT_2[48711] = 32'b11111111111111110000011111011011;
assign LUT_2[48712] = 32'b11111111111111101011000001111011;
assign LUT_2[48713] = 32'b11111111111111100111111010010100;
assign LUT_2[48714] = 32'b11111111111111110001111010110111;
assign LUT_2[48715] = 32'b11111111111111101110110011010000;
assign LUT_2[48716] = 32'b11111111111111100111011111100011;
assign LUT_2[48717] = 32'b11111111111111100100010111111100;
assign LUT_2[48718] = 32'b11111111111111101110011000011111;
assign LUT_2[48719] = 32'b11111111111111101011010000111000;
assign LUT_2[48720] = 32'b11111111111111101010110100101000;
assign LUT_2[48721] = 32'b11111111111111100111101101000001;
assign LUT_2[48722] = 32'b11111111111111110001101101100100;
assign LUT_2[48723] = 32'b11111111111111101110100101111101;
assign LUT_2[48724] = 32'b11111111111111100111010010010000;
assign LUT_2[48725] = 32'b11111111111111100100001010101001;
assign LUT_2[48726] = 32'b11111111111111101110001011001100;
assign LUT_2[48727] = 32'b11111111111111101011000011100101;
assign LUT_2[48728] = 32'b11111111111111100101100110000101;
assign LUT_2[48729] = 32'b11111111111111100010011110011110;
assign LUT_2[48730] = 32'b11111111111111101100011111000001;
assign LUT_2[48731] = 32'b11111111111111101001010111011010;
assign LUT_2[48732] = 32'b11111111111111100010000011101101;
assign LUT_2[48733] = 32'b11111111111111011110111100000110;
assign LUT_2[48734] = 32'b11111111111111101000111100101001;
assign LUT_2[48735] = 32'b11111111111111100101110101000010;
assign LUT_2[48736] = 32'b11111111111111110000101100000111;
assign LUT_2[48737] = 32'b11111111111111101101100100100000;
assign LUT_2[48738] = 32'b11111111111111110111100101000011;
assign LUT_2[48739] = 32'b11111111111111110100011101011100;
assign LUT_2[48740] = 32'b11111111111111101101001001101111;
assign LUT_2[48741] = 32'b11111111111111101010000010001000;
assign LUT_2[48742] = 32'b11111111111111110100000010101011;
assign LUT_2[48743] = 32'b11111111111111110000111011000100;
assign LUT_2[48744] = 32'b11111111111111101011011101100100;
assign LUT_2[48745] = 32'b11111111111111101000010101111101;
assign LUT_2[48746] = 32'b11111111111111110010010110100000;
assign LUT_2[48747] = 32'b11111111111111101111001110111001;
assign LUT_2[48748] = 32'b11111111111111100111111011001100;
assign LUT_2[48749] = 32'b11111111111111100100110011100101;
assign LUT_2[48750] = 32'b11111111111111101110110100001000;
assign LUT_2[48751] = 32'b11111111111111101011101100100001;
assign LUT_2[48752] = 32'b11111111111111101011010000010001;
assign LUT_2[48753] = 32'b11111111111111101000001000101010;
assign LUT_2[48754] = 32'b11111111111111110010001001001101;
assign LUT_2[48755] = 32'b11111111111111101111000001100110;
assign LUT_2[48756] = 32'b11111111111111100111101101111001;
assign LUT_2[48757] = 32'b11111111111111100100100110010010;
assign LUT_2[48758] = 32'b11111111111111101110100110110101;
assign LUT_2[48759] = 32'b11111111111111101011011111001110;
assign LUT_2[48760] = 32'b11111111111111100110000001101110;
assign LUT_2[48761] = 32'b11111111111111100010111010000111;
assign LUT_2[48762] = 32'b11111111111111101100111010101010;
assign LUT_2[48763] = 32'b11111111111111101001110011000011;
assign LUT_2[48764] = 32'b11111111111111100010011111010110;
assign LUT_2[48765] = 32'b11111111111111011111010111101111;
assign LUT_2[48766] = 32'b11111111111111101001011000010010;
assign LUT_2[48767] = 32'b11111111111111100110010000101011;
assign LUT_2[48768] = 32'b11111111111111111100011100001010;
assign LUT_2[48769] = 32'b11111111111111111001010100100011;
assign LUT_2[48770] = 32'b00000000000000000011010101000110;
assign LUT_2[48771] = 32'b00000000000000000000001101011111;
assign LUT_2[48772] = 32'b11111111111111111000111001110010;
assign LUT_2[48773] = 32'b11111111111111110101110010001011;
assign LUT_2[48774] = 32'b11111111111111111111110010101110;
assign LUT_2[48775] = 32'b11111111111111111100101011000111;
assign LUT_2[48776] = 32'b11111111111111110111001101100111;
assign LUT_2[48777] = 32'b11111111111111110100000110000000;
assign LUT_2[48778] = 32'b11111111111111111110000110100011;
assign LUT_2[48779] = 32'b11111111111111111010111110111100;
assign LUT_2[48780] = 32'b11111111111111110011101011001111;
assign LUT_2[48781] = 32'b11111111111111110000100011101000;
assign LUT_2[48782] = 32'b11111111111111111010100100001011;
assign LUT_2[48783] = 32'b11111111111111110111011100100100;
assign LUT_2[48784] = 32'b11111111111111110111000000010100;
assign LUT_2[48785] = 32'b11111111111111110011111000101101;
assign LUT_2[48786] = 32'b11111111111111111101111001010000;
assign LUT_2[48787] = 32'b11111111111111111010110001101001;
assign LUT_2[48788] = 32'b11111111111111110011011101111100;
assign LUT_2[48789] = 32'b11111111111111110000010110010101;
assign LUT_2[48790] = 32'b11111111111111111010010110111000;
assign LUT_2[48791] = 32'b11111111111111110111001111010001;
assign LUT_2[48792] = 32'b11111111111111110001110001110001;
assign LUT_2[48793] = 32'b11111111111111101110101010001010;
assign LUT_2[48794] = 32'b11111111111111111000101010101101;
assign LUT_2[48795] = 32'b11111111111111110101100011000110;
assign LUT_2[48796] = 32'b11111111111111101110001111011001;
assign LUT_2[48797] = 32'b11111111111111101011000111110010;
assign LUT_2[48798] = 32'b11111111111111110101001000010101;
assign LUT_2[48799] = 32'b11111111111111110010000000101110;
assign LUT_2[48800] = 32'b11111111111111111100110111110011;
assign LUT_2[48801] = 32'b11111111111111111001110000001100;
assign LUT_2[48802] = 32'b00000000000000000011110000101111;
assign LUT_2[48803] = 32'b00000000000000000000101001001000;
assign LUT_2[48804] = 32'b11111111111111111001010101011011;
assign LUT_2[48805] = 32'b11111111111111110110001101110100;
assign LUT_2[48806] = 32'b00000000000000000000001110010111;
assign LUT_2[48807] = 32'b11111111111111111101000110110000;
assign LUT_2[48808] = 32'b11111111111111110111101001010000;
assign LUT_2[48809] = 32'b11111111111111110100100001101001;
assign LUT_2[48810] = 32'b11111111111111111110100010001100;
assign LUT_2[48811] = 32'b11111111111111111011011010100101;
assign LUT_2[48812] = 32'b11111111111111110100000110111000;
assign LUT_2[48813] = 32'b11111111111111110000111111010001;
assign LUT_2[48814] = 32'b11111111111111111010111111110100;
assign LUT_2[48815] = 32'b11111111111111110111111000001101;
assign LUT_2[48816] = 32'b11111111111111110111011011111101;
assign LUT_2[48817] = 32'b11111111111111110100010100010110;
assign LUT_2[48818] = 32'b11111111111111111110010100111001;
assign LUT_2[48819] = 32'b11111111111111111011001101010010;
assign LUT_2[48820] = 32'b11111111111111110011111001100101;
assign LUT_2[48821] = 32'b11111111111111110000110001111110;
assign LUT_2[48822] = 32'b11111111111111111010110010100001;
assign LUT_2[48823] = 32'b11111111111111110111101010111010;
assign LUT_2[48824] = 32'b11111111111111110010001101011010;
assign LUT_2[48825] = 32'b11111111111111101111000101110011;
assign LUT_2[48826] = 32'b11111111111111111001000110010110;
assign LUT_2[48827] = 32'b11111111111111110101111110101111;
assign LUT_2[48828] = 32'b11111111111111101110101011000010;
assign LUT_2[48829] = 32'b11111111111111101011100011011011;
assign LUT_2[48830] = 32'b11111111111111110101100011111110;
assign LUT_2[48831] = 32'b11111111111111110010011100010111;
assign LUT_2[48832] = 32'b11111111111111110100100100101101;
assign LUT_2[48833] = 32'b11111111111111110001011101000110;
assign LUT_2[48834] = 32'b11111111111111111011011101101001;
assign LUT_2[48835] = 32'b11111111111111111000010110000010;
assign LUT_2[48836] = 32'b11111111111111110001000010010101;
assign LUT_2[48837] = 32'b11111111111111101101111010101110;
assign LUT_2[48838] = 32'b11111111111111110111111011010001;
assign LUT_2[48839] = 32'b11111111111111110100110011101010;
assign LUT_2[48840] = 32'b11111111111111101111010110001010;
assign LUT_2[48841] = 32'b11111111111111101100001110100011;
assign LUT_2[48842] = 32'b11111111111111110110001111000110;
assign LUT_2[48843] = 32'b11111111111111110011000111011111;
assign LUT_2[48844] = 32'b11111111111111101011110011110010;
assign LUT_2[48845] = 32'b11111111111111101000101100001011;
assign LUT_2[48846] = 32'b11111111111111110010101100101110;
assign LUT_2[48847] = 32'b11111111111111101111100101000111;
assign LUT_2[48848] = 32'b11111111111111101111001000110111;
assign LUT_2[48849] = 32'b11111111111111101100000001010000;
assign LUT_2[48850] = 32'b11111111111111110110000001110011;
assign LUT_2[48851] = 32'b11111111111111110010111010001100;
assign LUT_2[48852] = 32'b11111111111111101011100110011111;
assign LUT_2[48853] = 32'b11111111111111101000011110111000;
assign LUT_2[48854] = 32'b11111111111111110010011111011011;
assign LUT_2[48855] = 32'b11111111111111101111010111110100;
assign LUT_2[48856] = 32'b11111111111111101001111010010100;
assign LUT_2[48857] = 32'b11111111111111100110110010101101;
assign LUT_2[48858] = 32'b11111111111111110000110011010000;
assign LUT_2[48859] = 32'b11111111111111101101101011101001;
assign LUT_2[48860] = 32'b11111111111111100110010111111100;
assign LUT_2[48861] = 32'b11111111111111100011010000010101;
assign LUT_2[48862] = 32'b11111111111111101101010000111000;
assign LUT_2[48863] = 32'b11111111111111101010001001010001;
assign LUT_2[48864] = 32'b11111111111111110101000000010110;
assign LUT_2[48865] = 32'b11111111111111110001111000101111;
assign LUT_2[48866] = 32'b11111111111111111011111001010010;
assign LUT_2[48867] = 32'b11111111111111111000110001101011;
assign LUT_2[48868] = 32'b11111111111111110001011101111110;
assign LUT_2[48869] = 32'b11111111111111101110010110010111;
assign LUT_2[48870] = 32'b11111111111111111000010110111010;
assign LUT_2[48871] = 32'b11111111111111110101001111010011;
assign LUT_2[48872] = 32'b11111111111111101111110001110011;
assign LUT_2[48873] = 32'b11111111111111101100101010001100;
assign LUT_2[48874] = 32'b11111111111111110110101010101111;
assign LUT_2[48875] = 32'b11111111111111110011100011001000;
assign LUT_2[48876] = 32'b11111111111111101100001111011011;
assign LUT_2[48877] = 32'b11111111111111101001000111110100;
assign LUT_2[48878] = 32'b11111111111111110011001000010111;
assign LUT_2[48879] = 32'b11111111111111110000000000110000;
assign LUT_2[48880] = 32'b11111111111111101111100100100000;
assign LUT_2[48881] = 32'b11111111111111101100011100111001;
assign LUT_2[48882] = 32'b11111111111111110110011101011100;
assign LUT_2[48883] = 32'b11111111111111110011010101110101;
assign LUT_2[48884] = 32'b11111111111111101100000010001000;
assign LUT_2[48885] = 32'b11111111111111101000111010100001;
assign LUT_2[48886] = 32'b11111111111111110010111011000100;
assign LUT_2[48887] = 32'b11111111111111101111110011011101;
assign LUT_2[48888] = 32'b11111111111111101010010101111101;
assign LUT_2[48889] = 32'b11111111111111100111001110010110;
assign LUT_2[48890] = 32'b11111111111111110001001110111001;
assign LUT_2[48891] = 32'b11111111111111101110000111010010;
assign LUT_2[48892] = 32'b11111111111111100110110011100101;
assign LUT_2[48893] = 32'b11111111111111100011101011111110;
assign LUT_2[48894] = 32'b11111111111111101101101100100001;
assign LUT_2[48895] = 32'b11111111111111101010100100111010;
assign LUT_2[48896] = 32'b11111111111111111100000110100001;
assign LUT_2[48897] = 32'b11111111111111111000111110111010;
assign LUT_2[48898] = 32'b00000000000000000010111111011101;
assign LUT_2[48899] = 32'b11111111111111111111110111110110;
assign LUT_2[48900] = 32'b11111111111111111000100100001001;
assign LUT_2[48901] = 32'b11111111111111110101011100100010;
assign LUT_2[48902] = 32'b11111111111111111111011101000101;
assign LUT_2[48903] = 32'b11111111111111111100010101011110;
assign LUT_2[48904] = 32'b11111111111111110110110111111110;
assign LUT_2[48905] = 32'b11111111111111110011110000010111;
assign LUT_2[48906] = 32'b11111111111111111101110000111010;
assign LUT_2[48907] = 32'b11111111111111111010101001010011;
assign LUT_2[48908] = 32'b11111111111111110011010101100110;
assign LUT_2[48909] = 32'b11111111111111110000001101111111;
assign LUT_2[48910] = 32'b11111111111111111010001110100010;
assign LUT_2[48911] = 32'b11111111111111110111000110111011;
assign LUT_2[48912] = 32'b11111111111111110110101010101011;
assign LUT_2[48913] = 32'b11111111111111110011100011000100;
assign LUT_2[48914] = 32'b11111111111111111101100011100111;
assign LUT_2[48915] = 32'b11111111111111111010011100000000;
assign LUT_2[48916] = 32'b11111111111111110011001000010011;
assign LUT_2[48917] = 32'b11111111111111110000000000101100;
assign LUT_2[48918] = 32'b11111111111111111010000001001111;
assign LUT_2[48919] = 32'b11111111111111110110111001101000;
assign LUT_2[48920] = 32'b11111111111111110001011100001000;
assign LUT_2[48921] = 32'b11111111111111101110010100100001;
assign LUT_2[48922] = 32'b11111111111111111000010101000100;
assign LUT_2[48923] = 32'b11111111111111110101001101011101;
assign LUT_2[48924] = 32'b11111111111111101101111001110000;
assign LUT_2[48925] = 32'b11111111111111101010110010001001;
assign LUT_2[48926] = 32'b11111111111111110100110010101100;
assign LUT_2[48927] = 32'b11111111111111110001101011000101;
assign LUT_2[48928] = 32'b11111111111111111100100010001010;
assign LUT_2[48929] = 32'b11111111111111111001011010100011;
assign LUT_2[48930] = 32'b00000000000000000011011011000110;
assign LUT_2[48931] = 32'b00000000000000000000010011011111;
assign LUT_2[48932] = 32'b11111111111111111000111111110010;
assign LUT_2[48933] = 32'b11111111111111110101111000001011;
assign LUT_2[48934] = 32'b11111111111111111111111000101110;
assign LUT_2[48935] = 32'b11111111111111111100110001000111;
assign LUT_2[48936] = 32'b11111111111111110111010011100111;
assign LUT_2[48937] = 32'b11111111111111110100001100000000;
assign LUT_2[48938] = 32'b11111111111111111110001100100011;
assign LUT_2[48939] = 32'b11111111111111111011000100111100;
assign LUT_2[48940] = 32'b11111111111111110011110001001111;
assign LUT_2[48941] = 32'b11111111111111110000101001101000;
assign LUT_2[48942] = 32'b11111111111111111010101010001011;
assign LUT_2[48943] = 32'b11111111111111110111100010100100;
assign LUT_2[48944] = 32'b11111111111111110111000110010100;
assign LUT_2[48945] = 32'b11111111111111110011111110101101;
assign LUT_2[48946] = 32'b11111111111111111101111111010000;
assign LUT_2[48947] = 32'b11111111111111111010110111101001;
assign LUT_2[48948] = 32'b11111111111111110011100011111100;
assign LUT_2[48949] = 32'b11111111111111110000011100010101;
assign LUT_2[48950] = 32'b11111111111111111010011100111000;
assign LUT_2[48951] = 32'b11111111111111110111010101010001;
assign LUT_2[48952] = 32'b11111111111111110001110111110001;
assign LUT_2[48953] = 32'b11111111111111101110110000001010;
assign LUT_2[48954] = 32'b11111111111111111000110000101101;
assign LUT_2[48955] = 32'b11111111111111110101101001000110;
assign LUT_2[48956] = 32'b11111111111111101110010101011001;
assign LUT_2[48957] = 32'b11111111111111101011001101110010;
assign LUT_2[48958] = 32'b11111111111111110101001110010101;
assign LUT_2[48959] = 32'b11111111111111110010000110101110;
assign LUT_2[48960] = 32'b11111111111111110100001111000100;
assign LUT_2[48961] = 32'b11111111111111110001000111011101;
assign LUT_2[48962] = 32'b11111111111111111011001000000000;
assign LUT_2[48963] = 32'b11111111111111111000000000011001;
assign LUT_2[48964] = 32'b11111111111111110000101100101100;
assign LUT_2[48965] = 32'b11111111111111101101100101000101;
assign LUT_2[48966] = 32'b11111111111111110111100101101000;
assign LUT_2[48967] = 32'b11111111111111110100011110000001;
assign LUT_2[48968] = 32'b11111111111111101111000000100001;
assign LUT_2[48969] = 32'b11111111111111101011111000111010;
assign LUT_2[48970] = 32'b11111111111111110101111001011101;
assign LUT_2[48971] = 32'b11111111111111110010110001110110;
assign LUT_2[48972] = 32'b11111111111111101011011110001001;
assign LUT_2[48973] = 32'b11111111111111101000010110100010;
assign LUT_2[48974] = 32'b11111111111111110010010111000101;
assign LUT_2[48975] = 32'b11111111111111101111001111011110;
assign LUT_2[48976] = 32'b11111111111111101110110011001110;
assign LUT_2[48977] = 32'b11111111111111101011101011100111;
assign LUT_2[48978] = 32'b11111111111111110101101100001010;
assign LUT_2[48979] = 32'b11111111111111110010100100100011;
assign LUT_2[48980] = 32'b11111111111111101011010000110110;
assign LUT_2[48981] = 32'b11111111111111101000001001001111;
assign LUT_2[48982] = 32'b11111111111111110010001001110010;
assign LUT_2[48983] = 32'b11111111111111101111000010001011;
assign LUT_2[48984] = 32'b11111111111111101001100100101011;
assign LUT_2[48985] = 32'b11111111111111100110011101000100;
assign LUT_2[48986] = 32'b11111111111111110000011101100111;
assign LUT_2[48987] = 32'b11111111111111101101010110000000;
assign LUT_2[48988] = 32'b11111111111111100110000010010011;
assign LUT_2[48989] = 32'b11111111111111100010111010101100;
assign LUT_2[48990] = 32'b11111111111111101100111011001111;
assign LUT_2[48991] = 32'b11111111111111101001110011101000;
assign LUT_2[48992] = 32'b11111111111111110100101010101101;
assign LUT_2[48993] = 32'b11111111111111110001100011000110;
assign LUT_2[48994] = 32'b11111111111111111011100011101001;
assign LUT_2[48995] = 32'b11111111111111111000011100000010;
assign LUT_2[48996] = 32'b11111111111111110001001000010101;
assign LUT_2[48997] = 32'b11111111111111101110000000101110;
assign LUT_2[48998] = 32'b11111111111111111000000001010001;
assign LUT_2[48999] = 32'b11111111111111110100111001101010;
assign LUT_2[49000] = 32'b11111111111111101111011100001010;
assign LUT_2[49001] = 32'b11111111111111101100010100100011;
assign LUT_2[49002] = 32'b11111111111111110110010101000110;
assign LUT_2[49003] = 32'b11111111111111110011001101011111;
assign LUT_2[49004] = 32'b11111111111111101011111001110010;
assign LUT_2[49005] = 32'b11111111111111101000110010001011;
assign LUT_2[49006] = 32'b11111111111111110010110010101110;
assign LUT_2[49007] = 32'b11111111111111101111101011000111;
assign LUT_2[49008] = 32'b11111111111111101111001110110111;
assign LUT_2[49009] = 32'b11111111111111101100000111010000;
assign LUT_2[49010] = 32'b11111111111111110110000111110011;
assign LUT_2[49011] = 32'b11111111111111110011000000001100;
assign LUT_2[49012] = 32'b11111111111111101011101100011111;
assign LUT_2[49013] = 32'b11111111111111101000100100111000;
assign LUT_2[49014] = 32'b11111111111111110010100101011011;
assign LUT_2[49015] = 32'b11111111111111101111011101110100;
assign LUT_2[49016] = 32'b11111111111111101010000000010100;
assign LUT_2[49017] = 32'b11111111111111100110111000101101;
assign LUT_2[49018] = 32'b11111111111111110000111001010000;
assign LUT_2[49019] = 32'b11111111111111101101110001101001;
assign LUT_2[49020] = 32'b11111111111111100110011101111100;
assign LUT_2[49021] = 32'b11111111111111100011010110010101;
assign LUT_2[49022] = 32'b11111111111111101101010110111000;
assign LUT_2[49023] = 32'b11111111111111101010001111010001;
assign LUT_2[49024] = 32'b00000000000000000000011010110000;
assign LUT_2[49025] = 32'b11111111111111111101010011001001;
assign LUT_2[49026] = 32'b00000000000000000111010011101100;
assign LUT_2[49027] = 32'b00000000000000000100001100000101;
assign LUT_2[49028] = 32'b11111111111111111100111000011000;
assign LUT_2[49029] = 32'b11111111111111111001110000110001;
assign LUT_2[49030] = 32'b00000000000000000011110001010100;
assign LUT_2[49031] = 32'b00000000000000000000101001101101;
assign LUT_2[49032] = 32'b11111111111111111011001100001101;
assign LUT_2[49033] = 32'b11111111111111111000000100100110;
assign LUT_2[49034] = 32'b00000000000000000010000101001001;
assign LUT_2[49035] = 32'b11111111111111111110111101100010;
assign LUT_2[49036] = 32'b11111111111111110111101001110101;
assign LUT_2[49037] = 32'b11111111111111110100100010001110;
assign LUT_2[49038] = 32'b11111111111111111110100010110001;
assign LUT_2[49039] = 32'b11111111111111111011011011001010;
assign LUT_2[49040] = 32'b11111111111111111010111110111010;
assign LUT_2[49041] = 32'b11111111111111110111110111010011;
assign LUT_2[49042] = 32'b00000000000000000001110111110110;
assign LUT_2[49043] = 32'b11111111111111111110110000001111;
assign LUT_2[49044] = 32'b11111111111111110111011100100010;
assign LUT_2[49045] = 32'b11111111111111110100010100111011;
assign LUT_2[49046] = 32'b11111111111111111110010101011110;
assign LUT_2[49047] = 32'b11111111111111111011001101110111;
assign LUT_2[49048] = 32'b11111111111111110101110000010111;
assign LUT_2[49049] = 32'b11111111111111110010101000110000;
assign LUT_2[49050] = 32'b11111111111111111100101001010011;
assign LUT_2[49051] = 32'b11111111111111111001100001101100;
assign LUT_2[49052] = 32'b11111111111111110010001101111111;
assign LUT_2[49053] = 32'b11111111111111101111000110011000;
assign LUT_2[49054] = 32'b11111111111111111001000110111011;
assign LUT_2[49055] = 32'b11111111111111110101111111010100;
assign LUT_2[49056] = 32'b00000000000000000000110110011001;
assign LUT_2[49057] = 32'b11111111111111111101101110110010;
assign LUT_2[49058] = 32'b00000000000000000111101111010101;
assign LUT_2[49059] = 32'b00000000000000000100100111101110;
assign LUT_2[49060] = 32'b11111111111111111101010100000001;
assign LUT_2[49061] = 32'b11111111111111111010001100011010;
assign LUT_2[49062] = 32'b00000000000000000100001100111101;
assign LUT_2[49063] = 32'b00000000000000000001000101010110;
assign LUT_2[49064] = 32'b11111111111111111011100111110110;
assign LUT_2[49065] = 32'b11111111111111111000100000001111;
assign LUT_2[49066] = 32'b00000000000000000010100000110010;
assign LUT_2[49067] = 32'b11111111111111111111011001001011;
assign LUT_2[49068] = 32'b11111111111111111000000101011110;
assign LUT_2[49069] = 32'b11111111111111110100111101110111;
assign LUT_2[49070] = 32'b11111111111111111110111110011010;
assign LUT_2[49071] = 32'b11111111111111111011110110110011;
assign LUT_2[49072] = 32'b11111111111111111011011010100011;
assign LUT_2[49073] = 32'b11111111111111111000010010111100;
assign LUT_2[49074] = 32'b00000000000000000010010011011111;
assign LUT_2[49075] = 32'b11111111111111111111001011111000;
assign LUT_2[49076] = 32'b11111111111111110111111000001011;
assign LUT_2[49077] = 32'b11111111111111110100110000100100;
assign LUT_2[49078] = 32'b11111111111111111110110001000111;
assign LUT_2[49079] = 32'b11111111111111111011101001100000;
assign LUT_2[49080] = 32'b11111111111111110110001100000000;
assign LUT_2[49081] = 32'b11111111111111110011000100011001;
assign LUT_2[49082] = 32'b11111111111111111101000100111100;
assign LUT_2[49083] = 32'b11111111111111111001111101010101;
assign LUT_2[49084] = 32'b11111111111111110010101001101000;
assign LUT_2[49085] = 32'b11111111111111101111100010000001;
assign LUT_2[49086] = 32'b11111111111111111001100010100100;
assign LUT_2[49087] = 32'b11111111111111110110011010111101;
assign LUT_2[49088] = 32'b11111111111111111000100011010011;
assign LUT_2[49089] = 32'b11111111111111110101011011101100;
assign LUT_2[49090] = 32'b11111111111111111111011100001111;
assign LUT_2[49091] = 32'b11111111111111111100010100101000;
assign LUT_2[49092] = 32'b11111111111111110101000000111011;
assign LUT_2[49093] = 32'b11111111111111110001111001010100;
assign LUT_2[49094] = 32'b11111111111111111011111001110111;
assign LUT_2[49095] = 32'b11111111111111111000110010010000;
assign LUT_2[49096] = 32'b11111111111111110011010100110000;
assign LUT_2[49097] = 32'b11111111111111110000001101001001;
assign LUT_2[49098] = 32'b11111111111111111010001101101100;
assign LUT_2[49099] = 32'b11111111111111110111000110000101;
assign LUT_2[49100] = 32'b11111111111111101111110010011000;
assign LUT_2[49101] = 32'b11111111111111101100101010110001;
assign LUT_2[49102] = 32'b11111111111111110110101011010100;
assign LUT_2[49103] = 32'b11111111111111110011100011101101;
assign LUT_2[49104] = 32'b11111111111111110011000111011101;
assign LUT_2[49105] = 32'b11111111111111101111111111110110;
assign LUT_2[49106] = 32'b11111111111111111010000000011001;
assign LUT_2[49107] = 32'b11111111111111110110111000110010;
assign LUT_2[49108] = 32'b11111111111111101111100101000101;
assign LUT_2[49109] = 32'b11111111111111101100011101011110;
assign LUT_2[49110] = 32'b11111111111111110110011110000001;
assign LUT_2[49111] = 32'b11111111111111110011010110011010;
assign LUT_2[49112] = 32'b11111111111111101101111000111010;
assign LUT_2[49113] = 32'b11111111111111101010110001010011;
assign LUT_2[49114] = 32'b11111111111111110100110001110110;
assign LUT_2[49115] = 32'b11111111111111110001101010001111;
assign LUT_2[49116] = 32'b11111111111111101010010110100010;
assign LUT_2[49117] = 32'b11111111111111100111001110111011;
assign LUT_2[49118] = 32'b11111111111111110001001111011110;
assign LUT_2[49119] = 32'b11111111111111101110000111110111;
assign LUT_2[49120] = 32'b11111111111111111000111110111100;
assign LUT_2[49121] = 32'b11111111111111110101110111010101;
assign LUT_2[49122] = 32'b11111111111111111111110111111000;
assign LUT_2[49123] = 32'b11111111111111111100110000010001;
assign LUT_2[49124] = 32'b11111111111111110101011100100100;
assign LUT_2[49125] = 32'b11111111111111110010010100111101;
assign LUT_2[49126] = 32'b11111111111111111100010101100000;
assign LUT_2[49127] = 32'b11111111111111111001001101111001;
assign LUT_2[49128] = 32'b11111111111111110011110000011001;
assign LUT_2[49129] = 32'b11111111111111110000101000110010;
assign LUT_2[49130] = 32'b11111111111111111010101001010101;
assign LUT_2[49131] = 32'b11111111111111110111100001101110;
assign LUT_2[49132] = 32'b11111111111111110000001110000001;
assign LUT_2[49133] = 32'b11111111111111101101000110011010;
assign LUT_2[49134] = 32'b11111111111111110111000110111101;
assign LUT_2[49135] = 32'b11111111111111110011111111010110;
assign LUT_2[49136] = 32'b11111111111111110011100011000110;
assign LUT_2[49137] = 32'b11111111111111110000011011011111;
assign LUT_2[49138] = 32'b11111111111111111010011100000010;
assign LUT_2[49139] = 32'b11111111111111110111010100011011;
assign LUT_2[49140] = 32'b11111111111111110000000000101110;
assign LUT_2[49141] = 32'b11111111111111101100111001000111;
assign LUT_2[49142] = 32'b11111111111111110110111001101010;
assign LUT_2[49143] = 32'b11111111111111110011110010000011;
assign LUT_2[49144] = 32'b11111111111111101110010100100011;
assign LUT_2[49145] = 32'b11111111111111101011001100111100;
assign LUT_2[49146] = 32'b11111111111111110101001101011111;
assign LUT_2[49147] = 32'b11111111111111110010000101111000;
assign LUT_2[49148] = 32'b11111111111111101010110010001011;
assign LUT_2[49149] = 32'b11111111111111100111101010100100;
assign LUT_2[49150] = 32'b11111111111111110001101011000111;
assign LUT_2[49151] = 32'b11111111111111101110100011100000;
assign LUT_2[49152] = 32'b11111111111111110100000011110010;
assign LUT_2[49153] = 32'b11111111111111110000111100001011;
assign LUT_2[49154] = 32'b11111111111111111010111100101110;
assign LUT_2[49155] = 32'b11111111111111110111110101000111;
assign LUT_2[49156] = 32'b11111111111111110000100001011010;
assign LUT_2[49157] = 32'b11111111111111101101011001110011;
assign LUT_2[49158] = 32'b11111111111111110111011010010110;
assign LUT_2[49159] = 32'b11111111111111110100010010101111;
assign LUT_2[49160] = 32'b11111111111111101110110101001111;
assign LUT_2[49161] = 32'b11111111111111101011101101101000;
assign LUT_2[49162] = 32'b11111111111111110101101110001011;
assign LUT_2[49163] = 32'b11111111111111110010100110100100;
assign LUT_2[49164] = 32'b11111111111111101011010010110111;
assign LUT_2[49165] = 32'b11111111111111101000001011010000;
assign LUT_2[49166] = 32'b11111111111111110010001011110011;
assign LUT_2[49167] = 32'b11111111111111101111000100001100;
assign LUT_2[49168] = 32'b11111111111111101110100111111100;
assign LUT_2[49169] = 32'b11111111111111101011100000010101;
assign LUT_2[49170] = 32'b11111111111111110101100000111000;
assign LUT_2[49171] = 32'b11111111111111110010011001010001;
assign LUT_2[49172] = 32'b11111111111111101011000101100100;
assign LUT_2[49173] = 32'b11111111111111100111111101111101;
assign LUT_2[49174] = 32'b11111111111111110001111110100000;
assign LUT_2[49175] = 32'b11111111111111101110110110111001;
assign LUT_2[49176] = 32'b11111111111111101001011001011001;
assign LUT_2[49177] = 32'b11111111111111100110010001110010;
assign LUT_2[49178] = 32'b11111111111111110000010010010101;
assign LUT_2[49179] = 32'b11111111111111101101001010101110;
assign LUT_2[49180] = 32'b11111111111111100101110111000001;
assign LUT_2[49181] = 32'b11111111111111100010101111011010;
assign LUT_2[49182] = 32'b11111111111111101100101111111101;
assign LUT_2[49183] = 32'b11111111111111101001101000010110;
assign LUT_2[49184] = 32'b11111111111111110100011111011011;
assign LUT_2[49185] = 32'b11111111111111110001010111110100;
assign LUT_2[49186] = 32'b11111111111111111011011000010111;
assign LUT_2[49187] = 32'b11111111111111111000010000110000;
assign LUT_2[49188] = 32'b11111111111111110000111101000011;
assign LUT_2[49189] = 32'b11111111111111101101110101011100;
assign LUT_2[49190] = 32'b11111111111111110111110101111111;
assign LUT_2[49191] = 32'b11111111111111110100101110011000;
assign LUT_2[49192] = 32'b11111111111111101111010000111000;
assign LUT_2[49193] = 32'b11111111111111101100001001010001;
assign LUT_2[49194] = 32'b11111111111111110110001001110100;
assign LUT_2[49195] = 32'b11111111111111110011000010001101;
assign LUT_2[49196] = 32'b11111111111111101011101110100000;
assign LUT_2[49197] = 32'b11111111111111101000100110111001;
assign LUT_2[49198] = 32'b11111111111111110010100111011100;
assign LUT_2[49199] = 32'b11111111111111101111011111110101;
assign LUT_2[49200] = 32'b11111111111111101111000011100101;
assign LUT_2[49201] = 32'b11111111111111101011111011111110;
assign LUT_2[49202] = 32'b11111111111111110101111100100001;
assign LUT_2[49203] = 32'b11111111111111110010110100111010;
assign LUT_2[49204] = 32'b11111111111111101011100001001101;
assign LUT_2[49205] = 32'b11111111111111101000011001100110;
assign LUT_2[49206] = 32'b11111111111111110010011010001001;
assign LUT_2[49207] = 32'b11111111111111101111010010100010;
assign LUT_2[49208] = 32'b11111111111111101001110101000010;
assign LUT_2[49209] = 32'b11111111111111100110101101011011;
assign LUT_2[49210] = 32'b11111111111111110000101101111110;
assign LUT_2[49211] = 32'b11111111111111101101100110010111;
assign LUT_2[49212] = 32'b11111111111111100110010010101010;
assign LUT_2[49213] = 32'b11111111111111100011001011000011;
assign LUT_2[49214] = 32'b11111111111111101101001011100110;
assign LUT_2[49215] = 32'b11111111111111101010000011111111;
assign LUT_2[49216] = 32'b11111111111111101100001100010101;
assign LUT_2[49217] = 32'b11111111111111101001000100101110;
assign LUT_2[49218] = 32'b11111111111111110011000101010001;
assign LUT_2[49219] = 32'b11111111111111101111111101101010;
assign LUT_2[49220] = 32'b11111111111111101000101001111101;
assign LUT_2[49221] = 32'b11111111111111100101100010010110;
assign LUT_2[49222] = 32'b11111111111111101111100010111001;
assign LUT_2[49223] = 32'b11111111111111101100011011010010;
assign LUT_2[49224] = 32'b11111111111111100110111101110010;
assign LUT_2[49225] = 32'b11111111111111100011110110001011;
assign LUT_2[49226] = 32'b11111111111111101101110110101110;
assign LUT_2[49227] = 32'b11111111111111101010101111000111;
assign LUT_2[49228] = 32'b11111111111111100011011011011010;
assign LUT_2[49229] = 32'b11111111111111100000010011110011;
assign LUT_2[49230] = 32'b11111111111111101010010100010110;
assign LUT_2[49231] = 32'b11111111111111100111001100101111;
assign LUT_2[49232] = 32'b11111111111111100110110000011111;
assign LUT_2[49233] = 32'b11111111111111100011101000111000;
assign LUT_2[49234] = 32'b11111111111111101101101001011011;
assign LUT_2[49235] = 32'b11111111111111101010100001110100;
assign LUT_2[49236] = 32'b11111111111111100011001110000111;
assign LUT_2[49237] = 32'b11111111111111100000000110100000;
assign LUT_2[49238] = 32'b11111111111111101010000111000011;
assign LUT_2[49239] = 32'b11111111111111100110111111011100;
assign LUT_2[49240] = 32'b11111111111111100001100001111100;
assign LUT_2[49241] = 32'b11111111111111011110011010010101;
assign LUT_2[49242] = 32'b11111111111111101000011010111000;
assign LUT_2[49243] = 32'b11111111111111100101010011010001;
assign LUT_2[49244] = 32'b11111111111111011101111111100100;
assign LUT_2[49245] = 32'b11111111111111011010110111111101;
assign LUT_2[49246] = 32'b11111111111111100100111000100000;
assign LUT_2[49247] = 32'b11111111111111100001110000111001;
assign LUT_2[49248] = 32'b11111111111111101100100111111110;
assign LUT_2[49249] = 32'b11111111111111101001100000010111;
assign LUT_2[49250] = 32'b11111111111111110011100000111010;
assign LUT_2[49251] = 32'b11111111111111110000011001010011;
assign LUT_2[49252] = 32'b11111111111111101001000101100110;
assign LUT_2[49253] = 32'b11111111111111100101111101111111;
assign LUT_2[49254] = 32'b11111111111111101111111110100010;
assign LUT_2[49255] = 32'b11111111111111101100110110111011;
assign LUT_2[49256] = 32'b11111111111111100111011001011011;
assign LUT_2[49257] = 32'b11111111111111100100010001110100;
assign LUT_2[49258] = 32'b11111111111111101110010010010111;
assign LUT_2[49259] = 32'b11111111111111101011001010110000;
assign LUT_2[49260] = 32'b11111111111111100011110111000011;
assign LUT_2[49261] = 32'b11111111111111100000101111011100;
assign LUT_2[49262] = 32'b11111111111111101010101111111111;
assign LUT_2[49263] = 32'b11111111111111100111101000011000;
assign LUT_2[49264] = 32'b11111111111111100111001100001000;
assign LUT_2[49265] = 32'b11111111111111100100000100100001;
assign LUT_2[49266] = 32'b11111111111111101110000101000100;
assign LUT_2[49267] = 32'b11111111111111101010111101011101;
assign LUT_2[49268] = 32'b11111111111111100011101001110000;
assign LUT_2[49269] = 32'b11111111111111100000100010001001;
assign LUT_2[49270] = 32'b11111111111111101010100010101100;
assign LUT_2[49271] = 32'b11111111111111100111011011000101;
assign LUT_2[49272] = 32'b11111111111111100001111101100101;
assign LUT_2[49273] = 32'b11111111111111011110110101111110;
assign LUT_2[49274] = 32'b11111111111111101000110110100001;
assign LUT_2[49275] = 32'b11111111111111100101101110111010;
assign LUT_2[49276] = 32'b11111111111111011110011011001101;
assign LUT_2[49277] = 32'b11111111111111011011010011100110;
assign LUT_2[49278] = 32'b11111111111111100101010100001001;
assign LUT_2[49279] = 32'b11111111111111100010001100100010;
assign LUT_2[49280] = 32'b11111111111111111000011000000001;
assign LUT_2[49281] = 32'b11111111111111110101010000011010;
assign LUT_2[49282] = 32'b11111111111111111111010000111101;
assign LUT_2[49283] = 32'b11111111111111111100001001010110;
assign LUT_2[49284] = 32'b11111111111111110100110101101001;
assign LUT_2[49285] = 32'b11111111111111110001101110000010;
assign LUT_2[49286] = 32'b11111111111111111011101110100101;
assign LUT_2[49287] = 32'b11111111111111111000100110111110;
assign LUT_2[49288] = 32'b11111111111111110011001001011110;
assign LUT_2[49289] = 32'b11111111111111110000000001110111;
assign LUT_2[49290] = 32'b11111111111111111010000010011010;
assign LUT_2[49291] = 32'b11111111111111110110111010110011;
assign LUT_2[49292] = 32'b11111111111111101111100111000110;
assign LUT_2[49293] = 32'b11111111111111101100011111011111;
assign LUT_2[49294] = 32'b11111111111111110110100000000010;
assign LUT_2[49295] = 32'b11111111111111110011011000011011;
assign LUT_2[49296] = 32'b11111111111111110010111100001011;
assign LUT_2[49297] = 32'b11111111111111101111110100100100;
assign LUT_2[49298] = 32'b11111111111111111001110101000111;
assign LUT_2[49299] = 32'b11111111111111110110101101100000;
assign LUT_2[49300] = 32'b11111111111111101111011001110011;
assign LUT_2[49301] = 32'b11111111111111101100010010001100;
assign LUT_2[49302] = 32'b11111111111111110110010010101111;
assign LUT_2[49303] = 32'b11111111111111110011001011001000;
assign LUT_2[49304] = 32'b11111111111111101101101101101000;
assign LUT_2[49305] = 32'b11111111111111101010100110000001;
assign LUT_2[49306] = 32'b11111111111111110100100110100100;
assign LUT_2[49307] = 32'b11111111111111110001011110111101;
assign LUT_2[49308] = 32'b11111111111111101010001011010000;
assign LUT_2[49309] = 32'b11111111111111100111000011101001;
assign LUT_2[49310] = 32'b11111111111111110001000100001100;
assign LUT_2[49311] = 32'b11111111111111101101111100100101;
assign LUT_2[49312] = 32'b11111111111111111000110011101010;
assign LUT_2[49313] = 32'b11111111111111110101101100000011;
assign LUT_2[49314] = 32'b11111111111111111111101100100110;
assign LUT_2[49315] = 32'b11111111111111111100100100111111;
assign LUT_2[49316] = 32'b11111111111111110101010001010010;
assign LUT_2[49317] = 32'b11111111111111110010001001101011;
assign LUT_2[49318] = 32'b11111111111111111100001010001110;
assign LUT_2[49319] = 32'b11111111111111111001000010100111;
assign LUT_2[49320] = 32'b11111111111111110011100101000111;
assign LUT_2[49321] = 32'b11111111111111110000011101100000;
assign LUT_2[49322] = 32'b11111111111111111010011110000011;
assign LUT_2[49323] = 32'b11111111111111110111010110011100;
assign LUT_2[49324] = 32'b11111111111111110000000010101111;
assign LUT_2[49325] = 32'b11111111111111101100111011001000;
assign LUT_2[49326] = 32'b11111111111111110110111011101011;
assign LUT_2[49327] = 32'b11111111111111110011110100000100;
assign LUT_2[49328] = 32'b11111111111111110011010111110100;
assign LUT_2[49329] = 32'b11111111111111110000010000001101;
assign LUT_2[49330] = 32'b11111111111111111010010000110000;
assign LUT_2[49331] = 32'b11111111111111110111001001001001;
assign LUT_2[49332] = 32'b11111111111111101111110101011100;
assign LUT_2[49333] = 32'b11111111111111101100101101110101;
assign LUT_2[49334] = 32'b11111111111111110110101110011000;
assign LUT_2[49335] = 32'b11111111111111110011100110110001;
assign LUT_2[49336] = 32'b11111111111111101110001001010001;
assign LUT_2[49337] = 32'b11111111111111101011000001101010;
assign LUT_2[49338] = 32'b11111111111111110101000010001101;
assign LUT_2[49339] = 32'b11111111111111110001111010100110;
assign LUT_2[49340] = 32'b11111111111111101010100110111001;
assign LUT_2[49341] = 32'b11111111111111100111011111010010;
assign LUT_2[49342] = 32'b11111111111111110001011111110101;
assign LUT_2[49343] = 32'b11111111111111101110011000001110;
assign LUT_2[49344] = 32'b11111111111111110000100000100100;
assign LUT_2[49345] = 32'b11111111111111101101011000111101;
assign LUT_2[49346] = 32'b11111111111111110111011001100000;
assign LUT_2[49347] = 32'b11111111111111110100010001111001;
assign LUT_2[49348] = 32'b11111111111111101100111110001100;
assign LUT_2[49349] = 32'b11111111111111101001110110100101;
assign LUT_2[49350] = 32'b11111111111111110011110111001000;
assign LUT_2[49351] = 32'b11111111111111110000101111100001;
assign LUT_2[49352] = 32'b11111111111111101011010010000001;
assign LUT_2[49353] = 32'b11111111111111101000001010011010;
assign LUT_2[49354] = 32'b11111111111111110010001010111101;
assign LUT_2[49355] = 32'b11111111111111101111000011010110;
assign LUT_2[49356] = 32'b11111111111111100111101111101001;
assign LUT_2[49357] = 32'b11111111111111100100101000000010;
assign LUT_2[49358] = 32'b11111111111111101110101000100101;
assign LUT_2[49359] = 32'b11111111111111101011100000111110;
assign LUT_2[49360] = 32'b11111111111111101011000100101110;
assign LUT_2[49361] = 32'b11111111111111100111111101000111;
assign LUT_2[49362] = 32'b11111111111111110001111101101010;
assign LUT_2[49363] = 32'b11111111111111101110110110000011;
assign LUT_2[49364] = 32'b11111111111111100111100010010110;
assign LUT_2[49365] = 32'b11111111111111100100011010101111;
assign LUT_2[49366] = 32'b11111111111111101110011011010010;
assign LUT_2[49367] = 32'b11111111111111101011010011101011;
assign LUT_2[49368] = 32'b11111111111111100101110110001011;
assign LUT_2[49369] = 32'b11111111111111100010101110100100;
assign LUT_2[49370] = 32'b11111111111111101100101111000111;
assign LUT_2[49371] = 32'b11111111111111101001100111100000;
assign LUT_2[49372] = 32'b11111111111111100010010011110011;
assign LUT_2[49373] = 32'b11111111111111011111001100001100;
assign LUT_2[49374] = 32'b11111111111111101001001100101111;
assign LUT_2[49375] = 32'b11111111111111100110000101001000;
assign LUT_2[49376] = 32'b11111111111111110000111100001101;
assign LUT_2[49377] = 32'b11111111111111101101110100100110;
assign LUT_2[49378] = 32'b11111111111111110111110101001001;
assign LUT_2[49379] = 32'b11111111111111110100101101100010;
assign LUT_2[49380] = 32'b11111111111111101101011001110101;
assign LUT_2[49381] = 32'b11111111111111101010010010001110;
assign LUT_2[49382] = 32'b11111111111111110100010010110001;
assign LUT_2[49383] = 32'b11111111111111110001001011001010;
assign LUT_2[49384] = 32'b11111111111111101011101101101010;
assign LUT_2[49385] = 32'b11111111111111101000100110000011;
assign LUT_2[49386] = 32'b11111111111111110010100110100110;
assign LUT_2[49387] = 32'b11111111111111101111011110111111;
assign LUT_2[49388] = 32'b11111111111111101000001011010010;
assign LUT_2[49389] = 32'b11111111111111100101000011101011;
assign LUT_2[49390] = 32'b11111111111111101111000100001110;
assign LUT_2[49391] = 32'b11111111111111101011111100100111;
assign LUT_2[49392] = 32'b11111111111111101011100000010111;
assign LUT_2[49393] = 32'b11111111111111101000011000110000;
assign LUT_2[49394] = 32'b11111111111111110010011001010011;
assign LUT_2[49395] = 32'b11111111111111101111010001101100;
assign LUT_2[49396] = 32'b11111111111111100111111101111111;
assign LUT_2[49397] = 32'b11111111111111100100110110011000;
assign LUT_2[49398] = 32'b11111111111111101110110110111011;
assign LUT_2[49399] = 32'b11111111111111101011101111010100;
assign LUT_2[49400] = 32'b11111111111111100110010001110100;
assign LUT_2[49401] = 32'b11111111111111100011001010001101;
assign LUT_2[49402] = 32'b11111111111111101101001010110000;
assign LUT_2[49403] = 32'b11111111111111101010000011001001;
assign LUT_2[49404] = 32'b11111111111111100010101111011100;
assign LUT_2[49405] = 32'b11111111111111011111100111110101;
assign LUT_2[49406] = 32'b11111111111111101001101000011000;
assign LUT_2[49407] = 32'b11111111111111100110100000110001;
assign LUT_2[49408] = 32'b11111111111111111000000010011000;
assign LUT_2[49409] = 32'b11111111111111110100111010110001;
assign LUT_2[49410] = 32'b11111111111111111110111011010100;
assign LUT_2[49411] = 32'b11111111111111111011110011101101;
assign LUT_2[49412] = 32'b11111111111111110100100000000000;
assign LUT_2[49413] = 32'b11111111111111110001011000011001;
assign LUT_2[49414] = 32'b11111111111111111011011000111100;
assign LUT_2[49415] = 32'b11111111111111111000010001010101;
assign LUT_2[49416] = 32'b11111111111111110010110011110101;
assign LUT_2[49417] = 32'b11111111111111101111101100001110;
assign LUT_2[49418] = 32'b11111111111111111001101100110001;
assign LUT_2[49419] = 32'b11111111111111110110100101001010;
assign LUT_2[49420] = 32'b11111111111111101111010001011101;
assign LUT_2[49421] = 32'b11111111111111101100001001110110;
assign LUT_2[49422] = 32'b11111111111111110110001010011001;
assign LUT_2[49423] = 32'b11111111111111110011000010110010;
assign LUT_2[49424] = 32'b11111111111111110010100110100010;
assign LUT_2[49425] = 32'b11111111111111101111011110111011;
assign LUT_2[49426] = 32'b11111111111111111001011111011110;
assign LUT_2[49427] = 32'b11111111111111110110010111110111;
assign LUT_2[49428] = 32'b11111111111111101111000100001010;
assign LUT_2[49429] = 32'b11111111111111101011111100100011;
assign LUT_2[49430] = 32'b11111111111111110101111101000110;
assign LUT_2[49431] = 32'b11111111111111110010110101011111;
assign LUT_2[49432] = 32'b11111111111111101101010111111111;
assign LUT_2[49433] = 32'b11111111111111101010010000011000;
assign LUT_2[49434] = 32'b11111111111111110100010000111011;
assign LUT_2[49435] = 32'b11111111111111110001001001010100;
assign LUT_2[49436] = 32'b11111111111111101001110101100111;
assign LUT_2[49437] = 32'b11111111111111100110101110000000;
assign LUT_2[49438] = 32'b11111111111111110000101110100011;
assign LUT_2[49439] = 32'b11111111111111101101100110111100;
assign LUT_2[49440] = 32'b11111111111111111000011110000001;
assign LUT_2[49441] = 32'b11111111111111110101010110011010;
assign LUT_2[49442] = 32'b11111111111111111111010110111101;
assign LUT_2[49443] = 32'b11111111111111111100001111010110;
assign LUT_2[49444] = 32'b11111111111111110100111011101001;
assign LUT_2[49445] = 32'b11111111111111110001110100000010;
assign LUT_2[49446] = 32'b11111111111111111011110100100101;
assign LUT_2[49447] = 32'b11111111111111111000101100111110;
assign LUT_2[49448] = 32'b11111111111111110011001111011110;
assign LUT_2[49449] = 32'b11111111111111110000000111110111;
assign LUT_2[49450] = 32'b11111111111111111010001000011010;
assign LUT_2[49451] = 32'b11111111111111110111000000110011;
assign LUT_2[49452] = 32'b11111111111111101111101101000110;
assign LUT_2[49453] = 32'b11111111111111101100100101011111;
assign LUT_2[49454] = 32'b11111111111111110110100110000010;
assign LUT_2[49455] = 32'b11111111111111110011011110011011;
assign LUT_2[49456] = 32'b11111111111111110011000010001011;
assign LUT_2[49457] = 32'b11111111111111101111111010100100;
assign LUT_2[49458] = 32'b11111111111111111001111011000111;
assign LUT_2[49459] = 32'b11111111111111110110110011100000;
assign LUT_2[49460] = 32'b11111111111111101111011111110011;
assign LUT_2[49461] = 32'b11111111111111101100011000001100;
assign LUT_2[49462] = 32'b11111111111111110110011000101111;
assign LUT_2[49463] = 32'b11111111111111110011010001001000;
assign LUT_2[49464] = 32'b11111111111111101101110011101000;
assign LUT_2[49465] = 32'b11111111111111101010101100000001;
assign LUT_2[49466] = 32'b11111111111111110100101100100100;
assign LUT_2[49467] = 32'b11111111111111110001100100111101;
assign LUT_2[49468] = 32'b11111111111111101010010001010000;
assign LUT_2[49469] = 32'b11111111111111100111001001101001;
assign LUT_2[49470] = 32'b11111111111111110001001010001100;
assign LUT_2[49471] = 32'b11111111111111101110000010100101;
assign LUT_2[49472] = 32'b11111111111111110000001010111011;
assign LUT_2[49473] = 32'b11111111111111101101000011010100;
assign LUT_2[49474] = 32'b11111111111111110111000011110111;
assign LUT_2[49475] = 32'b11111111111111110011111100010000;
assign LUT_2[49476] = 32'b11111111111111101100101000100011;
assign LUT_2[49477] = 32'b11111111111111101001100000111100;
assign LUT_2[49478] = 32'b11111111111111110011100001011111;
assign LUT_2[49479] = 32'b11111111111111110000011001111000;
assign LUT_2[49480] = 32'b11111111111111101010111100011000;
assign LUT_2[49481] = 32'b11111111111111100111110100110001;
assign LUT_2[49482] = 32'b11111111111111110001110101010100;
assign LUT_2[49483] = 32'b11111111111111101110101101101101;
assign LUT_2[49484] = 32'b11111111111111100111011010000000;
assign LUT_2[49485] = 32'b11111111111111100100010010011001;
assign LUT_2[49486] = 32'b11111111111111101110010010111100;
assign LUT_2[49487] = 32'b11111111111111101011001011010101;
assign LUT_2[49488] = 32'b11111111111111101010101111000101;
assign LUT_2[49489] = 32'b11111111111111100111100111011110;
assign LUT_2[49490] = 32'b11111111111111110001101000000001;
assign LUT_2[49491] = 32'b11111111111111101110100000011010;
assign LUT_2[49492] = 32'b11111111111111100111001100101101;
assign LUT_2[49493] = 32'b11111111111111100100000101000110;
assign LUT_2[49494] = 32'b11111111111111101110000101101001;
assign LUT_2[49495] = 32'b11111111111111101010111110000010;
assign LUT_2[49496] = 32'b11111111111111100101100000100010;
assign LUT_2[49497] = 32'b11111111111111100010011000111011;
assign LUT_2[49498] = 32'b11111111111111101100011001011110;
assign LUT_2[49499] = 32'b11111111111111101001010001110111;
assign LUT_2[49500] = 32'b11111111111111100001111110001010;
assign LUT_2[49501] = 32'b11111111111111011110110110100011;
assign LUT_2[49502] = 32'b11111111111111101000110111000110;
assign LUT_2[49503] = 32'b11111111111111100101101111011111;
assign LUT_2[49504] = 32'b11111111111111110000100110100100;
assign LUT_2[49505] = 32'b11111111111111101101011110111101;
assign LUT_2[49506] = 32'b11111111111111110111011111100000;
assign LUT_2[49507] = 32'b11111111111111110100010111111001;
assign LUT_2[49508] = 32'b11111111111111101101000100001100;
assign LUT_2[49509] = 32'b11111111111111101001111100100101;
assign LUT_2[49510] = 32'b11111111111111110011111101001000;
assign LUT_2[49511] = 32'b11111111111111110000110101100001;
assign LUT_2[49512] = 32'b11111111111111101011011000000001;
assign LUT_2[49513] = 32'b11111111111111101000010000011010;
assign LUT_2[49514] = 32'b11111111111111110010010000111101;
assign LUT_2[49515] = 32'b11111111111111101111001001010110;
assign LUT_2[49516] = 32'b11111111111111100111110101101001;
assign LUT_2[49517] = 32'b11111111111111100100101110000010;
assign LUT_2[49518] = 32'b11111111111111101110101110100101;
assign LUT_2[49519] = 32'b11111111111111101011100110111110;
assign LUT_2[49520] = 32'b11111111111111101011001010101110;
assign LUT_2[49521] = 32'b11111111111111101000000011000111;
assign LUT_2[49522] = 32'b11111111111111110010000011101010;
assign LUT_2[49523] = 32'b11111111111111101110111100000011;
assign LUT_2[49524] = 32'b11111111111111100111101000010110;
assign LUT_2[49525] = 32'b11111111111111100100100000101111;
assign LUT_2[49526] = 32'b11111111111111101110100001010010;
assign LUT_2[49527] = 32'b11111111111111101011011001101011;
assign LUT_2[49528] = 32'b11111111111111100101111100001011;
assign LUT_2[49529] = 32'b11111111111111100010110100100100;
assign LUT_2[49530] = 32'b11111111111111101100110101000111;
assign LUT_2[49531] = 32'b11111111111111101001101101100000;
assign LUT_2[49532] = 32'b11111111111111100010011001110011;
assign LUT_2[49533] = 32'b11111111111111011111010010001100;
assign LUT_2[49534] = 32'b11111111111111101001010010101111;
assign LUT_2[49535] = 32'b11111111111111100110001011001000;
assign LUT_2[49536] = 32'b11111111111111111100010110100111;
assign LUT_2[49537] = 32'b11111111111111111001001111000000;
assign LUT_2[49538] = 32'b00000000000000000011001111100011;
assign LUT_2[49539] = 32'b00000000000000000000000111111100;
assign LUT_2[49540] = 32'b11111111111111111000110100001111;
assign LUT_2[49541] = 32'b11111111111111110101101100101000;
assign LUT_2[49542] = 32'b11111111111111111111101101001011;
assign LUT_2[49543] = 32'b11111111111111111100100101100100;
assign LUT_2[49544] = 32'b11111111111111110111001000000100;
assign LUT_2[49545] = 32'b11111111111111110100000000011101;
assign LUT_2[49546] = 32'b11111111111111111110000001000000;
assign LUT_2[49547] = 32'b11111111111111111010111001011001;
assign LUT_2[49548] = 32'b11111111111111110011100101101100;
assign LUT_2[49549] = 32'b11111111111111110000011110000101;
assign LUT_2[49550] = 32'b11111111111111111010011110101000;
assign LUT_2[49551] = 32'b11111111111111110111010111000001;
assign LUT_2[49552] = 32'b11111111111111110110111010110001;
assign LUT_2[49553] = 32'b11111111111111110011110011001010;
assign LUT_2[49554] = 32'b11111111111111111101110011101101;
assign LUT_2[49555] = 32'b11111111111111111010101100000110;
assign LUT_2[49556] = 32'b11111111111111110011011000011001;
assign LUT_2[49557] = 32'b11111111111111110000010000110010;
assign LUT_2[49558] = 32'b11111111111111111010010001010101;
assign LUT_2[49559] = 32'b11111111111111110111001001101110;
assign LUT_2[49560] = 32'b11111111111111110001101100001110;
assign LUT_2[49561] = 32'b11111111111111101110100100100111;
assign LUT_2[49562] = 32'b11111111111111111000100101001010;
assign LUT_2[49563] = 32'b11111111111111110101011101100011;
assign LUT_2[49564] = 32'b11111111111111101110001001110110;
assign LUT_2[49565] = 32'b11111111111111101011000010001111;
assign LUT_2[49566] = 32'b11111111111111110101000010110010;
assign LUT_2[49567] = 32'b11111111111111110001111011001011;
assign LUT_2[49568] = 32'b11111111111111111100110010010000;
assign LUT_2[49569] = 32'b11111111111111111001101010101001;
assign LUT_2[49570] = 32'b00000000000000000011101011001100;
assign LUT_2[49571] = 32'b00000000000000000000100011100101;
assign LUT_2[49572] = 32'b11111111111111111001001111111000;
assign LUT_2[49573] = 32'b11111111111111110110001000010001;
assign LUT_2[49574] = 32'b00000000000000000000001000110100;
assign LUT_2[49575] = 32'b11111111111111111101000001001101;
assign LUT_2[49576] = 32'b11111111111111110111100011101101;
assign LUT_2[49577] = 32'b11111111111111110100011100000110;
assign LUT_2[49578] = 32'b11111111111111111110011100101001;
assign LUT_2[49579] = 32'b11111111111111111011010101000010;
assign LUT_2[49580] = 32'b11111111111111110100000001010101;
assign LUT_2[49581] = 32'b11111111111111110000111001101110;
assign LUT_2[49582] = 32'b11111111111111111010111010010001;
assign LUT_2[49583] = 32'b11111111111111110111110010101010;
assign LUT_2[49584] = 32'b11111111111111110111010110011010;
assign LUT_2[49585] = 32'b11111111111111110100001110110011;
assign LUT_2[49586] = 32'b11111111111111111110001111010110;
assign LUT_2[49587] = 32'b11111111111111111011000111101111;
assign LUT_2[49588] = 32'b11111111111111110011110100000010;
assign LUT_2[49589] = 32'b11111111111111110000101100011011;
assign LUT_2[49590] = 32'b11111111111111111010101100111110;
assign LUT_2[49591] = 32'b11111111111111110111100101010111;
assign LUT_2[49592] = 32'b11111111111111110010000111110111;
assign LUT_2[49593] = 32'b11111111111111101111000000010000;
assign LUT_2[49594] = 32'b11111111111111111001000000110011;
assign LUT_2[49595] = 32'b11111111111111110101111001001100;
assign LUT_2[49596] = 32'b11111111111111101110100101011111;
assign LUT_2[49597] = 32'b11111111111111101011011101111000;
assign LUT_2[49598] = 32'b11111111111111110101011110011011;
assign LUT_2[49599] = 32'b11111111111111110010010110110100;
assign LUT_2[49600] = 32'b11111111111111110100011111001010;
assign LUT_2[49601] = 32'b11111111111111110001010111100011;
assign LUT_2[49602] = 32'b11111111111111111011011000000110;
assign LUT_2[49603] = 32'b11111111111111111000010000011111;
assign LUT_2[49604] = 32'b11111111111111110000111100110010;
assign LUT_2[49605] = 32'b11111111111111101101110101001011;
assign LUT_2[49606] = 32'b11111111111111110111110101101110;
assign LUT_2[49607] = 32'b11111111111111110100101110000111;
assign LUT_2[49608] = 32'b11111111111111101111010000100111;
assign LUT_2[49609] = 32'b11111111111111101100001001000000;
assign LUT_2[49610] = 32'b11111111111111110110001001100011;
assign LUT_2[49611] = 32'b11111111111111110011000001111100;
assign LUT_2[49612] = 32'b11111111111111101011101110001111;
assign LUT_2[49613] = 32'b11111111111111101000100110101000;
assign LUT_2[49614] = 32'b11111111111111110010100111001011;
assign LUT_2[49615] = 32'b11111111111111101111011111100100;
assign LUT_2[49616] = 32'b11111111111111101111000011010100;
assign LUT_2[49617] = 32'b11111111111111101011111011101101;
assign LUT_2[49618] = 32'b11111111111111110101111100010000;
assign LUT_2[49619] = 32'b11111111111111110010110100101001;
assign LUT_2[49620] = 32'b11111111111111101011100000111100;
assign LUT_2[49621] = 32'b11111111111111101000011001010101;
assign LUT_2[49622] = 32'b11111111111111110010011001111000;
assign LUT_2[49623] = 32'b11111111111111101111010010010001;
assign LUT_2[49624] = 32'b11111111111111101001110100110001;
assign LUT_2[49625] = 32'b11111111111111100110101101001010;
assign LUT_2[49626] = 32'b11111111111111110000101101101101;
assign LUT_2[49627] = 32'b11111111111111101101100110000110;
assign LUT_2[49628] = 32'b11111111111111100110010010011001;
assign LUT_2[49629] = 32'b11111111111111100011001010110010;
assign LUT_2[49630] = 32'b11111111111111101101001011010101;
assign LUT_2[49631] = 32'b11111111111111101010000011101110;
assign LUT_2[49632] = 32'b11111111111111110100111010110011;
assign LUT_2[49633] = 32'b11111111111111110001110011001100;
assign LUT_2[49634] = 32'b11111111111111111011110011101111;
assign LUT_2[49635] = 32'b11111111111111111000101100001000;
assign LUT_2[49636] = 32'b11111111111111110001011000011011;
assign LUT_2[49637] = 32'b11111111111111101110010000110100;
assign LUT_2[49638] = 32'b11111111111111111000010001010111;
assign LUT_2[49639] = 32'b11111111111111110101001001110000;
assign LUT_2[49640] = 32'b11111111111111101111101100010000;
assign LUT_2[49641] = 32'b11111111111111101100100100101001;
assign LUT_2[49642] = 32'b11111111111111110110100101001100;
assign LUT_2[49643] = 32'b11111111111111110011011101100101;
assign LUT_2[49644] = 32'b11111111111111101100001001111000;
assign LUT_2[49645] = 32'b11111111111111101001000010010001;
assign LUT_2[49646] = 32'b11111111111111110011000010110100;
assign LUT_2[49647] = 32'b11111111111111101111111011001101;
assign LUT_2[49648] = 32'b11111111111111101111011110111101;
assign LUT_2[49649] = 32'b11111111111111101100010111010110;
assign LUT_2[49650] = 32'b11111111111111110110010111111001;
assign LUT_2[49651] = 32'b11111111111111110011010000010010;
assign LUT_2[49652] = 32'b11111111111111101011111100100101;
assign LUT_2[49653] = 32'b11111111111111101000110100111110;
assign LUT_2[49654] = 32'b11111111111111110010110101100001;
assign LUT_2[49655] = 32'b11111111111111101111101101111010;
assign LUT_2[49656] = 32'b11111111111111101010010000011010;
assign LUT_2[49657] = 32'b11111111111111100111001000110011;
assign LUT_2[49658] = 32'b11111111111111110001001001010110;
assign LUT_2[49659] = 32'b11111111111111101110000001101111;
assign LUT_2[49660] = 32'b11111111111111100110101110000010;
assign LUT_2[49661] = 32'b11111111111111100011100110011011;
assign LUT_2[49662] = 32'b11111111111111101101100110111110;
assign LUT_2[49663] = 32'b11111111111111101010011111010111;
assign LUT_2[49664] = 32'b11111111111111111000110101100100;
assign LUT_2[49665] = 32'b11111111111111110101101101111101;
assign LUT_2[49666] = 32'b11111111111111111111101110100000;
assign LUT_2[49667] = 32'b11111111111111111100100110111001;
assign LUT_2[49668] = 32'b11111111111111110101010011001100;
assign LUT_2[49669] = 32'b11111111111111110010001011100101;
assign LUT_2[49670] = 32'b11111111111111111100001100001000;
assign LUT_2[49671] = 32'b11111111111111111001000100100001;
assign LUT_2[49672] = 32'b11111111111111110011100111000001;
assign LUT_2[49673] = 32'b11111111111111110000011111011010;
assign LUT_2[49674] = 32'b11111111111111111010011111111101;
assign LUT_2[49675] = 32'b11111111111111110111011000010110;
assign LUT_2[49676] = 32'b11111111111111110000000100101001;
assign LUT_2[49677] = 32'b11111111111111101100111101000010;
assign LUT_2[49678] = 32'b11111111111111110110111101100101;
assign LUT_2[49679] = 32'b11111111111111110011110101111110;
assign LUT_2[49680] = 32'b11111111111111110011011001101110;
assign LUT_2[49681] = 32'b11111111111111110000010010000111;
assign LUT_2[49682] = 32'b11111111111111111010010010101010;
assign LUT_2[49683] = 32'b11111111111111110111001011000011;
assign LUT_2[49684] = 32'b11111111111111101111110111010110;
assign LUT_2[49685] = 32'b11111111111111101100101111101111;
assign LUT_2[49686] = 32'b11111111111111110110110000010010;
assign LUT_2[49687] = 32'b11111111111111110011101000101011;
assign LUT_2[49688] = 32'b11111111111111101110001011001011;
assign LUT_2[49689] = 32'b11111111111111101011000011100100;
assign LUT_2[49690] = 32'b11111111111111110101000100000111;
assign LUT_2[49691] = 32'b11111111111111110001111100100000;
assign LUT_2[49692] = 32'b11111111111111101010101000110011;
assign LUT_2[49693] = 32'b11111111111111100111100001001100;
assign LUT_2[49694] = 32'b11111111111111110001100001101111;
assign LUT_2[49695] = 32'b11111111111111101110011010001000;
assign LUT_2[49696] = 32'b11111111111111111001010001001101;
assign LUT_2[49697] = 32'b11111111111111110110001001100110;
assign LUT_2[49698] = 32'b00000000000000000000001010001001;
assign LUT_2[49699] = 32'b11111111111111111101000010100010;
assign LUT_2[49700] = 32'b11111111111111110101101110110101;
assign LUT_2[49701] = 32'b11111111111111110010100111001110;
assign LUT_2[49702] = 32'b11111111111111111100100111110001;
assign LUT_2[49703] = 32'b11111111111111111001100000001010;
assign LUT_2[49704] = 32'b11111111111111110100000010101010;
assign LUT_2[49705] = 32'b11111111111111110000111011000011;
assign LUT_2[49706] = 32'b11111111111111111010111011100110;
assign LUT_2[49707] = 32'b11111111111111110111110011111111;
assign LUT_2[49708] = 32'b11111111111111110000100000010010;
assign LUT_2[49709] = 32'b11111111111111101101011000101011;
assign LUT_2[49710] = 32'b11111111111111110111011001001110;
assign LUT_2[49711] = 32'b11111111111111110100010001100111;
assign LUT_2[49712] = 32'b11111111111111110011110101010111;
assign LUT_2[49713] = 32'b11111111111111110000101101110000;
assign LUT_2[49714] = 32'b11111111111111111010101110010011;
assign LUT_2[49715] = 32'b11111111111111110111100110101100;
assign LUT_2[49716] = 32'b11111111111111110000010010111111;
assign LUT_2[49717] = 32'b11111111111111101101001011011000;
assign LUT_2[49718] = 32'b11111111111111110111001011111011;
assign LUT_2[49719] = 32'b11111111111111110100000100010100;
assign LUT_2[49720] = 32'b11111111111111101110100110110100;
assign LUT_2[49721] = 32'b11111111111111101011011111001101;
assign LUT_2[49722] = 32'b11111111111111110101011111110000;
assign LUT_2[49723] = 32'b11111111111111110010011000001001;
assign LUT_2[49724] = 32'b11111111111111101011000100011100;
assign LUT_2[49725] = 32'b11111111111111100111111100110101;
assign LUT_2[49726] = 32'b11111111111111110001111101011000;
assign LUT_2[49727] = 32'b11111111111111101110110101110001;
assign LUT_2[49728] = 32'b11111111111111110000111110000111;
assign LUT_2[49729] = 32'b11111111111111101101110110100000;
assign LUT_2[49730] = 32'b11111111111111110111110111000011;
assign LUT_2[49731] = 32'b11111111111111110100101111011100;
assign LUT_2[49732] = 32'b11111111111111101101011011101111;
assign LUT_2[49733] = 32'b11111111111111101010010100001000;
assign LUT_2[49734] = 32'b11111111111111110100010100101011;
assign LUT_2[49735] = 32'b11111111111111110001001101000100;
assign LUT_2[49736] = 32'b11111111111111101011101111100100;
assign LUT_2[49737] = 32'b11111111111111101000100111111101;
assign LUT_2[49738] = 32'b11111111111111110010101000100000;
assign LUT_2[49739] = 32'b11111111111111101111100000111001;
assign LUT_2[49740] = 32'b11111111111111101000001101001100;
assign LUT_2[49741] = 32'b11111111111111100101000101100101;
assign LUT_2[49742] = 32'b11111111111111101111000110001000;
assign LUT_2[49743] = 32'b11111111111111101011111110100001;
assign LUT_2[49744] = 32'b11111111111111101011100010010001;
assign LUT_2[49745] = 32'b11111111111111101000011010101010;
assign LUT_2[49746] = 32'b11111111111111110010011011001101;
assign LUT_2[49747] = 32'b11111111111111101111010011100110;
assign LUT_2[49748] = 32'b11111111111111100111111111111001;
assign LUT_2[49749] = 32'b11111111111111100100111000010010;
assign LUT_2[49750] = 32'b11111111111111101110111000110101;
assign LUT_2[49751] = 32'b11111111111111101011110001001110;
assign LUT_2[49752] = 32'b11111111111111100110010011101110;
assign LUT_2[49753] = 32'b11111111111111100011001100000111;
assign LUT_2[49754] = 32'b11111111111111101101001100101010;
assign LUT_2[49755] = 32'b11111111111111101010000101000011;
assign LUT_2[49756] = 32'b11111111111111100010110001010110;
assign LUT_2[49757] = 32'b11111111111111011111101001101111;
assign LUT_2[49758] = 32'b11111111111111101001101010010010;
assign LUT_2[49759] = 32'b11111111111111100110100010101011;
assign LUT_2[49760] = 32'b11111111111111110001011001110000;
assign LUT_2[49761] = 32'b11111111111111101110010010001001;
assign LUT_2[49762] = 32'b11111111111111111000010010101100;
assign LUT_2[49763] = 32'b11111111111111110101001011000101;
assign LUT_2[49764] = 32'b11111111111111101101110111011000;
assign LUT_2[49765] = 32'b11111111111111101010101111110001;
assign LUT_2[49766] = 32'b11111111111111110100110000010100;
assign LUT_2[49767] = 32'b11111111111111110001101000101101;
assign LUT_2[49768] = 32'b11111111111111101100001011001101;
assign LUT_2[49769] = 32'b11111111111111101001000011100110;
assign LUT_2[49770] = 32'b11111111111111110011000100001001;
assign LUT_2[49771] = 32'b11111111111111101111111100100010;
assign LUT_2[49772] = 32'b11111111111111101000101000110101;
assign LUT_2[49773] = 32'b11111111111111100101100001001110;
assign LUT_2[49774] = 32'b11111111111111101111100001110001;
assign LUT_2[49775] = 32'b11111111111111101100011010001010;
assign LUT_2[49776] = 32'b11111111111111101011111101111010;
assign LUT_2[49777] = 32'b11111111111111101000110110010011;
assign LUT_2[49778] = 32'b11111111111111110010110110110110;
assign LUT_2[49779] = 32'b11111111111111101111101111001111;
assign LUT_2[49780] = 32'b11111111111111101000011011100010;
assign LUT_2[49781] = 32'b11111111111111100101010011111011;
assign LUT_2[49782] = 32'b11111111111111101111010100011110;
assign LUT_2[49783] = 32'b11111111111111101100001100110111;
assign LUT_2[49784] = 32'b11111111111111100110101111010111;
assign LUT_2[49785] = 32'b11111111111111100011100111110000;
assign LUT_2[49786] = 32'b11111111111111101101101000010011;
assign LUT_2[49787] = 32'b11111111111111101010100000101100;
assign LUT_2[49788] = 32'b11111111111111100011001100111111;
assign LUT_2[49789] = 32'b11111111111111100000000101011000;
assign LUT_2[49790] = 32'b11111111111111101010000101111011;
assign LUT_2[49791] = 32'b11111111111111100110111110010100;
assign LUT_2[49792] = 32'b11111111111111111101001001110011;
assign LUT_2[49793] = 32'b11111111111111111010000010001100;
assign LUT_2[49794] = 32'b00000000000000000100000010101111;
assign LUT_2[49795] = 32'b00000000000000000000111011001000;
assign LUT_2[49796] = 32'b11111111111111111001100111011011;
assign LUT_2[49797] = 32'b11111111111111110110011111110100;
assign LUT_2[49798] = 32'b00000000000000000000100000010111;
assign LUT_2[49799] = 32'b11111111111111111101011000110000;
assign LUT_2[49800] = 32'b11111111111111110111111011010000;
assign LUT_2[49801] = 32'b11111111111111110100110011101001;
assign LUT_2[49802] = 32'b11111111111111111110110100001100;
assign LUT_2[49803] = 32'b11111111111111111011101100100101;
assign LUT_2[49804] = 32'b11111111111111110100011000111000;
assign LUT_2[49805] = 32'b11111111111111110001010001010001;
assign LUT_2[49806] = 32'b11111111111111111011010001110100;
assign LUT_2[49807] = 32'b11111111111111111000001010001101;
assign LUT_2[49808] = 32'b11111111111111110111101101111101;
assign LUT_2[49809] = 32'b11111111111111110100100110010110;
assign LUT_2[49810] = 32'b11111111111111111110100110111001;
assign LUT_2[49811] = 32'b11111111111111111011011111010010;
assign LUT_2[49812] = 32'b11111111111111110100001011100101;
assign LUT_2[49813] = 32'b11111111111111110001000011111110;
assign LUT_2[49814] = 32'b11111111111111111011000100100001;
assign LUT_2[49815] = 32'b11111111111111110111111100111010;
assign LUT_2[49816] = 32'b11111111111111110010011111011010;
assign LUT_2[49817] = 32'b11111111111111101111010111110011;
assign LUT_2[49818] = 32'b11111111111111111001011000010110;
assign LUT_2[49819] = 32'b11111111111111110110010000101111;
assign LUT_2[49820] = 32'b11111111111111101110111101000010;
assign LUT_2[49821] = 32'b11111111111111101011110101011011;
assign LUT_2[49822] = 32'b11111111111111110101110101111110;
assign LUT_2[49823] = 32'b11111111111111110010101110010111;
assign LUT_2[49824] = 32'b11111111111111111101100101011100;
assign LUT_2[49825] = 32'b11111111111111111010011101110101;
assign LUT_2[49826] = 32'b00000000000000000100011110011000;
assign LUT_2[49827] = 32'b00000000000000000001010110110001;
assign LUT_2[49828] = 32'b11111111111111111010000011000100;
assign LUT_2[49829] = 32'b11111111111111110110111011011101;
assign LUT_2[49830] = 32'b00000000000000000000111100000000;
assign LUT_2[49831] = 32'b11111111111111111101110100011001;
assign LUT_2[49832] = 32'b11111111111111111000010110111001;
assign LUT_2[49833] = 32'b11111111111111110101001111010010;
assign LUT_2[49834] = 32'b11111111111111111111001111110101;
assign LUT_2[49835] = 32'b11111111111111111100001000001110;
assign LUT_2[49836] = 32'b11111111111111110100110100100001;
assign LUT_2[49837] = 32'b11111111111111110001101100111010;
assign LUT_2[49838] = 32'b11111111111111111011101101011101;
assign LUT_2[49839] = 32'b11111111111111111000100101110110;
assign LUT_2[49840] = 32'b11111111111111111000001001100110;
assign LUT_2[49841] = 32'b11111111111111110101000001111111;
assign LUT_2[49842] = 32'b11111111111111111111000010100010;
assign LUT_2[49843] = 32'b11111111111111111011111010111011;
assign LUT_2[49844] = 32'b11111111111111110100100111001110;
assign LUT_2[49845] = 32'b11111111111111110001011111100111;
assign LUT_2[49846] = 32'b11111111111111111011100000001010;
assign LUT_2[49847] = 32'b11111111111111111000011000100011;
assign LUT_2[49848] = 32'b11111111111111110010111011000011;
assign LUT_2[49849] = 32'b11111111111111101111110011011100;
assign LUT_2[49850] = 32'b11111111111111111001110011111111;
assign LUT_2[49851] = 32'b11111111111111110110101100011000;
assign LUT_2[49852] = 32'b11111111111111101111011000101011;
assign LUT_2[49853] = 32'b11111111111111101100010001000100;
assign LUT_2[49854] = 32'b11111111111111110110010001100111;
assign LUT_2[49855] = 32'b11111111111111110011001010000000;
assign LUT_2[49856] = 32'b11111111111111110101010010010110;
assign LUT_2[49857] = 32'b11111111111111110010001010101111;
assign LUT_2[49858] = 32'b11111111111111111100001011010010;
assign LUT_2[49859] = 32'b11111111111111111001000011101011;
assign LUT_2[49860] = 32'b11111111111111110001101111111110;
assign LUT_2[49861] = 32'b11111111111111101110101000010111;
assign LUT_2[49862] = 32'b11111111111111111000101000111010;
assign LUT_2[49863] = 32'b11111111111111110101100001010011;
assign LUT_2[49864] = 32'b11111111111111110000000011110011;
assign LUT_2[49865] = 32'b11111111111111101100111100001100;
assign LUT_2[49866] = 32'b11111111111111110110111100101111;
assign LUT_2[49867] = 32'b11111111111111110011110101001000;
assign LUT_2[49868] = 32'b11111111111111101100100001011011;
assign LUT_2[49869] = 32'b11111111111111101001011001110100;
assign LUT_2[49870] = 32'b11111111111111110011011010010111;
assign LUT_2[49871] = 32'b11111111111111110000010010110000;
assign LUT_2[49872] = 32'b11111111111111101111110110100000;
assign LUT_2[49873] = 32'b11111111111111101100101110111001;
assign LUT_2[49874] = 32'b11111111111111110110101111011100;
assign LUT_2[49875] = 32'b11111111111111110011100111110101;
assign LUT_2[49876] = 32'b11111111111111101100010100001000;
assign LUT_2[49877] = 32'b11111111111111101001001100100001;
assign LUT_2[49878] = 32'b11111111111111110011001101000100;
assign LUT_2[49879] = 32'b11111111111111110000000101011101;
assign LUT_2[49880] = 32'b11111111111111101010100111111101;
assign LUT_2[49881] = 32'b11111111111111100111100000010110;
assign LUT_2[49882] = 32'b11111111111111110001100000111001;
assign LUT_2[49883] = 32'b11111111111111101110011001010010;
assign LUT_2[49884] = 32'b11111111111111100111000101100101;
assign LUT_2[49885] = 32'b11111111111111100011111101111110;
assign LUT_2[49886] = 32'b11111111111111101101111110100001;
assign LUT_2[49887] = 32'b11111111111111101010110110111010;
assign LUT_2[49888] = 32'b11111111111111110101101101111111;
assign LUT_2[49889] = 32'b11111111111111110010100110011000;
assign LUT_2[49890] = 32'b11111111111111111100100110111011;
assign LUT_2[49891] = 32'b11111111111111111001011111010100;
assign LUT_2[49892] = 32'b11111111111111110010001011100111;
assign LUT_2[49893] = 32'b11111111111111101111000100000000;
assign LUT_2[49894] = 32'b11111111111111111001000100100011;
assign LUT_2[49895] = 32'b11111111111111110101111100111100;
assign LUT_2[49896] = 32'b11111111111111110000011111011100;
assign LUT_2[49897] = 32'b11111111111111101101010111110101;
assign LUT_2[49898] = 32'b11111111111111110111011000011000;
assign LUT_2[49899] = 32'b11111111111111110100010000110001;
assign LUT_2[49900] = 32'b11111111111111101100111101000100;
assign LUT_2[49901] = 32'b11111111111111101001110101011101;
assign LUT_2[49902] = 32'b11111111111111110011110110000000;
assign LUT_2[49903] = 32'b11111111111111110000101110011001;
assign LUT_2[49904] = 32'b11111111111111110000010010001001;
assign LUT_2[49905] = 32'b11111111111111101101001010100010;
assign LUT_2[49906] = 32'b11111111111111110111001011000101;
assign LUT_2[49907] = 32'b11111111111111110100000011011110;
assign LUT_2[49908] = 32'b11111111111111101100101111110001;
assign LUT_2[49909] = 32'b11111111111111101001101000001010;
assign LUT_2[49910] = 32'b11111111111111110011101000101101;
assign LUT_2[49911] = 32'b11111111111111110000100001000110;
assign LUT_2[49912] = 32'b11111111111111101011000011100110;
assign LUT_2[49913] = 32'b11111111111111100111111011111111;
assign LUT_2[49914] = 32'b11111111111111110001111100100010;
assign LUT_2[49915] = 32'b11111111111111101110110100111011;
assign LUT_2[49916] = 32'b11111111111111100111100001001110;
assign LUT_2[49917] = 32'b11111111111111100100011001100111;
assign LUT_2[49918] = 32'b11111111111111101110011010001010;
assign LUT_2[49919] = 32'b11111111111111101011010010100011;
assign LUT_2[49920] = 32'b11111111111111111100110100001010;
assign LUT_2[49921] = 32'b11111111111111111001101100100011;
assign LUT_2[49922] = 32'b00000000000000000011101101000110;
assign LUT_2[49923] = 32'b00000000000000000000100101011111;
assign LUT_2[49924] = 32'b11111111111111111001010001110010;
assign LUT_2[49925] = 32'b11111111111111110110001010001011;
assign LUT_2[49926] = 32'b00000000000000000000001010101110;
assign LUT_2[49927] = 32'b11111111111111111101000011000111;
assign LUT_2[49928] = 32'b11111111111111110111100101100111;
assign LUT_2[49929] = 32'b11111111111111110100011110000000;
assign LUT_2[49930] = 32'b11111111111111111110011110100011;
assign LUT_2[49931] = 32'b11111111111111111011010110111100;
assign LUT_2[49932] = 32'b11111111111111110100000011001111;
assign LUT_2[49933] = 32'b11111111111111110000111011101000;
assign LUT_2[49934] = 32'b11111111111111111010111100001011;
assign LUT_2[49935] = 32'b11111111111111110111110100100100;
assign LUT_2[49936] = 32'b11111111111111110111011000010100;
assign LUT_2[49937] = 32'b11111111111111110100010000101101;
assign LUT_2[49938] = 32'b11111111111111111110010001010000;
assign LUT_2[49939] = 32'b11111111111111111011001001101001;
assign LUT_2[49940] = 32'b11111111111111110011110101111100;
assign LUT_2[49941] = 32'b11111111111111110000101110010101;
assign LUT_2[49942] = 32'b11111111111111111010101110111000;
assign LUT_2[49943] = 32'b11111111111111110111100111010001;
assign LUT_2[49944] = 32'b11111111111111110010001001110001;
assign LUT_2[49945] = 32'b11111111111111101111000010001010;
assign LUT_2[49946] = 32'b11111111111111111001000010101101;
assign LUT_2[49947] = 32'b11111111111111110101111011000110;
assign LUT_2[49948] = 32'b11111111111111101110100111011001;
assign LUT_2[49949] = 32'b11111111111111101011011111110010;
assign LUT_2[49950] = 32'b11111111111111110101100000010101;
assign LUT_2[49951] = 32'b11111111111111110010011000101110;
assign LUT_2[49952] = 32'b11111111111111111101001111110011;
assign LUT_2[49953] = 32'b11111111111111111010001000001100;
assign LUT_2[49954] = 32'b00000000000000000100001000101111;
assign LUT_2[49955] = 32'b00000000000000000001000001001000;
assign LUT_2[49956] = 32'b11111111111111111001101101011011;
assign LUT_2[49957] = 32'b11111111111111110110100101110100;
assign LUT_2[49958] = 32'b00000000000000000000100110010111;
assign LUT_2[49959] = 32'b11111111111111111101011110110000;
assign LUT_2[49960] = 32'b11111111111111111000000001010000;
assign LUT_2[49961] = 32'b11111111111111110100111001101001;
assign LUT_2[49962] = 32'b11111111111111111110111010001100;
assign LUT_2[49963] = 32'b11111111111111111011110010100101;
assign LUT_2[49964] = 32'b11111111111111110100011110111000;
assign LUT_2[49965] = 32'b11111111111111110001010111010001;
assign LUT_2[49966] = 32'b11111111111111111011010111110100;
assign LUT_2[49967] = 32'b11111111111111111000010000001101;
assign LUT_2[49968] = 32'b11111111111111110111110011111101;
assign LUT_2[49969] = 32'b11111111111111110100101100010110;
assign LUT_2[49970] = 32'b11111111111111111110101100111001;
assign LUT_2[49971] = 32'b11111111111111111011100101010010;
assign LUT_2[49972] = 32'b11111111111111110100010001100101;
assign LUT_2[49973] = 32'b11111111111111110001001001111110;
assign LUT_2[49974] = 32'b11111111111111111011001010100001;
assign LUT_2[49975] = 32'b11111111111111111000000010111010;
assign LUT_2[49976] = 32'b11111111111111110010100101011010;
assign LUT_2[49977] = 32'b11111111111111101111011101110011;
assign LUT_2[49978] = 32'b11111111111111111001011110010110;
assign LUT_2[49979] = 32'b11111111111111110110010110101111;
assign LUT_2[49980] = 32'b11111111111111101111000011000010;
assign LUT_2[49981] = 32'b11111111111111101011111011011011;
assign LUT_2[49982] = 32'b11111111111111110101111011111110;
assign LUT_2[49983] = 32'b11111111111111110010110100010111;
assign LUT_2[49984] = 32'b11111111111111110100111100101101;
assign LUT_2[49985] = 32'b11111111111111110001110101000110;
assign LUT_2[49986] = 32'b11111111111111111011110101101001;
assign LUT_2[49987] = 32'b11111111111111111000101110000010;
assign LUT_2[49988] = 32'b11111111111111110001011010010101;
assign LUT_2[49989] = 32'b11111111111111101110010010101110;
assign LUT_2[49990] = 32'b11111111111111111000010011010001;
assign LUT_2[49991] = 32'b11111111111111110101001011101010;
assign LUT_2[49992] = 32'b11111111111111101111101110001010;
assign LUT_2[49993] = 32'b11111111111111101100100110100011;
assign LUT_2[49994] = 32'b11111111111111110110100111000110;
assign LUT_2[49995] = 32'b11111111111111110011011111011111;
assign LUT_2[49996] = 32'b11111111111111101100001011110010;
assign LUT_2[49997] = 32'b11111111111111101001000100001011;
assign LUT_2[49998] = 32'b11111111111111110011000100101110;
assign LUT_2[49999] = 32'b11111111111111101111111101000111;
assign LUT_2[50000] = 32'b11111111111111101111100000110111;
assign LUT_2[50001] = 32'b11111111111111101100011001010000;
assign LUT_2[50002] = 32'b11111111111111110110011001110011;
assign LUT_2[50003] = 32'b11111111111111110011010010001100;
assign LUT_2[50004] = 32'b11111111111111101011111110011111;
assign LUT_2[50005] = 32'b11111111111111101000110110111000;
assign LUT_2[50006] = 32'b11111111111111110010110111011011;
assign LUT_2[50007] = 32'b11111111111111101111101111110100;
assign LUT_2[50008] = 32'b11111111111111101010010010010100;
assign LUT_2[50009] = 32'b11111111111111100111001010101101;
assign LUT_2[50010] = 32'b11111111111111110001001011010000;
assign LUT_2[50011] = 32'b11111111111111101110000011101001;
assign LUT_2[50012] = 32'b11111111111111100110101111111100;
assign LUT_2[50013] = 32'b11111111111111100011101000010101;
assign LUT_2[50014] = 32'b11111111111111101101101000111000;
assign LUT_2[50015] = 32'b11111111111111101010100001010001;
assign LUT_2[50016] = 32'b11111111111111110101011000010110;
assign LUT_2[50017] = 32'b11111111111111110010010000101111;
assign LUT_2[50018] = 32'b11111111111111111100010001010010;
assign LUT_2[50019] = 32'b11111111111111111001001001101011;
assign LUT_2[50020] = 32'b11111111111111110001110101111110;
assign LUT_2[50021] = 32'b11111111111111101110101110010111;
assign LUT_2[50022] = 32'b11111111111111111000101110111010;
assign LUT_2[50023] = 32'b11111111111111110101100111010011;
assign LUT_2[50024] = 32'b11111111111111110000001001110011;
assign LUT_2[50025] = 32'b11111111111111101101000010001100;
assign LUT_2[50026] = 32'b11111111111111110111000010101111;
assign LUT_2[50027] = 32'b11111111111111110011111011001000;
assign LUT_2[50028] = 32'b11111111111111101100100111011011;
assign LUT_2[50029] = 32'b11111111111111101001011111110100;
assign LUT_2[50030] = 32'b11111111111111110011100000010111;
assign LUT_2[50031] = 32'b11111111111111110000011000110000;
assign LUT_2[50032] = 32'b11111111111111101111111100100000;
assign LUT_2[50033] = 32'b11111111111111101100110100111001;
assign LUT_2[50034] = 32'b11111111111111110110110101011100;
assign LUT_2[50035] = 32'b11111111111111110011101101110101;
assign LUT_2[50036] = 32'b11111111111111101100011010001000;
assign LUT_2[50037] = 32'b11111111111111101001010010100001;
assign LUT_2[50038] = 32'b11111111111111110011010011000100;
assign LUT_2[50039] = 32'b11111111111111110000001011011101;
assign LUT_2[50040] = 32'b11111111111111101010101101111101;
assign LUT_2[50041] = 32'b11111111111111100111100110010110;
assign LUT_2[50042] = 32'b11111111111111110001100110111001;
assign LUT_2[50043] = 32'b11111111111111101110011111010010;
assign LUT_2[50044] = 32'b11111111111111100111001011100101;
assign LUT_2[50045] = 32'b11111111111111100100000011111110;
assign LUT_2[50046] = 32'b11111111111111101110000100100001;
assign LUT_2[50047] = 32'b11111111111111101010111100111010;
assign LUT_2[50048] = 32'b00000000000000000001001000011001;
assign LUT_2[50049] = 32'b11111111111111111110000000110010;
assign LUT_2[50050] = 32'b00000000000000001000000001010101;
assign LUT_2[50051] = 32'b00000000000000000100111001101110;
assign LUT_2[50052] = 32'b11111111111111111101100110000001;
assign LUT_2[50053] = 32'b11111111111111111010011110011010;
assign LUT_2[50054] = 32'b00000000000000000100011110111101;
assign LUT_2[50055] = 32'b00000000000000000001010111010110;
assign LUT_2[50056] = 32'b11111111111111111011111001110110;
assign LUT_2[50057] = 32'b11111111111111111000110010001111;
assign LUT_2[50058] = 32'b00000000000000000010110010110010;
assign LUT_2[50059] = 32'b11111111111111111111101011001011;
assign LUT_2[50060] = 32'b11111111111111111000010111011110;
assign LUT_2[50061] = 32'b11111111111111110101001111110111;
assign LUT_2[50062] = 32'b11111111111111111111010000011010;
assign LUT_2[50063] = 32'b11111111111111111100001000110011;
assign LUT_2[50064] = 32'b11111111111111111011101100100011;
assign LUT_2[50065] = 32'b11111111111111111000100100111100;
assign LUT_2[50066] = 32'b00000000000000000010100101011111;
assign LUT_2[50067] = 32'b11111111111111111111011101111000;
assign LUT_2[50068] = 32'b11111111111111111000001010001011;
assign LUT_2[50069] = 32'b11111111111111110101000010100100;
assign LUT_2[50070] = 32'b11111111111111111111000011000111;
assign LUT_2[50071] = 32'b11111111111111111011111011100000;
assign LUT_2[50072] = 32'b11111111111111110110011110000000;
assign LUT_2[50073] = 32'b11111111111111110011010110011001;
assign LUT_2[50074] = 32'b11111111111111111101010110111100;
assign LUT_2[50075] = 32'b11111111111111111010001111010101;
assign LUT_2[50076] = 32'b11111111111111110010111011101000;
assign LUT_2[50077] = 32'b11111111111111101111110100000001;
assign LUT_2[50078] = 32'b11111111111111111001110100100100;
assign LUT_2[50079] = 32'b11111111111111110110101100111101;
assign LUT_2[50080] = 32'b00000000000000000001100100000010;
assign LUT_2[50081] = 32'b11111111111111111110011100011011;
assign LUT_2[50082] = 32'b00000000000000001000011100111110;
assign LUT_2[50083] = 32'b00000000000000000101010101010111;
assign LUT_2[50084] = 32'b11111111111111111110000001101010;
assign LUT_2[50085] = 32'b11111111111111111010111010000011;
assign LUT_2[50086] = 32'b00000000000000000100111010100110;
assign LUT_2[50087] = 32'b00000000000000000001110010111111;
assign LUT_2[50088] = 32'b11111111111111111100010101011111;
assign LUT_2[50089] = 32'b11111111111111111001001101111000;
assign LUT_2[50090] = 32'b00000000000000000011001110011011;
assign LUT_2[50091] = 32'b00000000000000000000000110110100;
assign LUT_2[50092] = 32'b11111111111111111000110011000111;
assign LUT_2[50093] = 32'b11111111111111110101101011100000;
assign LUT_2[50094] = 32'b11111111111111111111101100000011;
assign LUT_2[50095] = 32'b11111111111111111100100100011100;
assign LUT_2[50096] = 32'b11111111111111111100001000001100;
assign LUT_2[50097] = 32'b11111111111111111001000000100101;
assign LUT_2[50098] = 32'b00000000000000000011000001001000;
assign LUT_2[50099] = 32'b11111111111111111111111001100001;
assign LUT_2[50100] = 32'b11111111111111111000100101110100;
assign LUT_2[50101] = 32'b11111111111111110101011110001101;
assign LUT_2[50102] = 32'b11111111111111111111011110110000;
assign LUT_2[50103] = 32'b11111111111111111100010111001001;
assign LUT_2[50104] = 32'b11111111111111110110111001101001;
assign LUT_2[50105] = 32'b11111111111111110011110010000010;
assign LUT_2[50106] = 32'b11111111111111111101110010100101;
assign LUT_2[50107] = 32'b11111111111111111010101010111110;
assign LUT_2[50108] = 32'b11111111111111110011010111010001;
assign LUT_2[50109] = 32'b11111111111111110000001111101010;
assign LUT_2[50110] = 32'b11111111111111111010010000001101;
assign LUT_2[50111] = 32'b11111111111111110111001000100110;
assign LUT_2[50112] = 32'b11111111111111111001010000111100;
assign LUT_2[50113] = 32'b11111111111111110110001001010101;
assign LUT_2[50114] = 32'b00000000000000000000001001111000;
assign LUT_2[50115] = 32'b11111111111111111101000010010001;
assign LUT_2[50116] = 32'b11111111111111110101101110100100;
assign LUT_2[50117] = 32'b11111111111111110010100110111101;
assign LUT_2[50118] = 32'b11111111111111111100100111100000;
assign LUT_2[50119] = 32'b11111111111111111001011111111001;
assign LUT_2[50120] = 32'b11111111111111110100000010011001;
assign LUT_2[50121] = 32'b11111111111111110000111010110010;
assign LUT_2[50122] = 32'b11111111111111111010111011010101;
assign LUT_2[50123] = 32'b11111111111111110111110011101110;
assign LUT_2[50124] = 32'b11111111111111110000100000000001;
assign LUT_2[50125] = 32'b11111111111111101101011000011010;
assign LUT_2[50126] = 32'b11111111111111110111011000111101;
assign LUT_2[50127] = 32'b11111111111111110100010001010110;
assign LUT_2[50128] = 32'b11111111111111110011110101000110;
assign LUT_2[50129] = 32'b11111111111111110000101101011111;
assign LUT_2[50130] = 32'b11111111111111111010101110000010;
assign LUT_2[50131] = 32'b11111111111111110111100110011011;
assign LUT_2[50132] = 32'b11111111111111110000010010101110;
assign LUT_2[50133] = 32'b11111111111111101101001011000111;
assign LUT_2[50134] = 32'b11111111111111110111001011101010;
assign LUT_2[50135] = 32'b11111111111111110100000100000011;
assign LUT_2[50136] = 32'b11111111111111101110100110100011;
assign LUT_2[50137] = 32'b11111111111111101011011110111100;
assign LUT_2[50138] = 32'b11111111111111110101011111011111;
assign LUT_2[50139] = 32'b11111111111111110010010111111000;
assign LUT_2[50140] = 32'b11111111111111101011000100001011;
assign LUT_2[50141] = 32'b11111111111111100111111100100100;
assign LUT_2[50142] = 32'b11111111111111110001111101000111;
assign LUT_2[50143] = 32'b11111111111111101110110101100000;
assign LUT_2[50144] = 32'b11111111111111111001101100100101;
assign LUT_2[50145] = 32'b11111111111111110110100100111110;
assign LUT_2[50146] = 32'b00000000000000000000100101100001;
assign LUT_2[50147] = 32'b11111111111111111101011101111010;
assign LUT_2[50148] = 32'b11111111111111110110001010001101;
assign LUT_2[50149] = 32'b11111111111111110011000010100110;
assign LUT_2[50150] = 32'b11111111111111111101000011001001;
assign LUT_2[50151] = 32'b11111111111111111001111011100010;
assign LUT_2[50152] = 32'b11111111111111110100011110000010;
assign LUT_2[50153] = 32'b11111111111111110001010110011011;
assign LUT_2[50154] = 32'b11111111111111111011010110111110;
assign LUT_2[50155] = 32'b11111111111111111000001111010111;
assign LUT_2[50156] = 32'b11111111111111110000111011101010;
assign LUT_2[50157] = 32'b11111111111111101101110100000011;
assign LUT_2[50158] = 32'b11111111111111110111110100100110;
assign LUT_2[50159] = 32'b11111111111111110100101100111111;
assign LUT_2[50160] = 32'b11111111111111110100010000101111;
assign LUT_2[50161] = 32'b11111111111111110001001001001000;
assign LUT_2[50162] = 32'b11111111111111111011001001101011;
assign LUT_2[50163] = 32'b11111111111111111000000010000100;
assign LUT_2[50164] = 32'b11111111111111110000101110010111;
assign LUT_2[50165] = 32'b11111111111111101101100110110000;
assign LUT_2[50166] = 32'b11111111111111110111100111010011;
assign LUT_2[50167] = 32'b11111111111111110100011111101100;
assign LUT_2[50168] = 32'b11111111111111101111000010001100;
assign LUT_2[50169] = 32'b11111111111111101011111010100101;
assign LUT_2[50170] = 32'b11111111111111110101111011001000;
assign LUT_2[50171] = 32'b11111111111111110010110011100001;
assign LUT_2[50172] = 32'b11111111111111101011011111110100;
assign LUT_2[50173] = 32'b11111111111111101000011000001101;
assign LUT_2[50174] = 32'b11111111111111110010011000110000;
assign LUT_2[50175] = 32'b11111111111111101111010001001001;
assign LUT_2[50176] = 32'b11111111111111111010101111110111;
assign LUT_2[50177] = 32'b11111111111111110111101000010000;
assign LUT_2[50178] = 32'b00000000000000000001101000110011;
assign LUT_2[50179] = 32'b11111111111111111110100001001100;
assign LUT_2[50180] = 32'b11111111111111110111001101011111;
assign LUT_2[50181] = 32'b11111111111111110100000101111000;
assign LUT_2[50182] = 32'b11111111111111111110000110011011;
assign LUT_2[50183] = 32'b11111111111111111010111110110100;
assign LUT_2[50184] = 32'b11111111111111110101100001010100;
assign LUT_2[50185] = 32'b11111111111111110010011001101101;
assign LUT_2[50186] = 32'b11111111111111111100011010010000;
assign LUT_2[50187] = 32'b11111111111111111001010010101001;
assign LUT_2[50188] = 32'b11111111111111110001111110111100;
assign LUT_2[50189] = 32'b11111111111111101110110111010101;
assign LUT_2[50190] = 32'b11111111111111111000110111111000;
assign LUT_2[50191] = 32'b11111111111111110101110000010001;
assign LUT_2[50192] = 32'b11111111111111110101010100000001;
assign LUT_2[50193] = 32'b11111111111111110010001100011010;
assign LUT_2[50194] = 32'b11111111111111111100001100111101;
assign LUT_2[50195] = 32'b11111111111111111001000101010110;
assign LUT_2[50196] = 32'b11111111111111110001110001101001;
assign LUT_2[50197] = 32'b11111111111111101110101010000010;
assign LUT_2[50198] = 32'b11111111111111111000101010100101;
assign LUT_2[50199] = 32'b11111111111111110101100010111110;
assign LUT_2[50200] = 32'b11111111111111110000000101011110;
assign LUT_2[50201] = 32'b11111111111111101100111101110111;
assign LUT_2[50202] = 32'b11111111111111110110111110011010;
assign LUT_2[50203] = 32'b11111111111111110011110110110011;
assign LUT_2[50204] = 32'b11111111111111101100100011000110;
assign LUT_2[50205] = 32'b11111111111111101001011011011111;
assign LUT_2[50206] = 32'b11111111111111110011011100000010;
assign LUT_2[50207] = 32'b11111111111111110000010100011011;
assign LUT_2[50208] = 32'b11111111111111111011001011100000;
assign LUT_2[50209] = 32'b11111111111111111000000011111001;
assign LUT_2[50210] = 32'b00000000000000000010000100011100;
assign LUT_2[50211] = 32'b11111111111111111110111100110101;
assign LUT_2[50212] = 32'b11111111111111110111101001001000;
assign LUT_2[50213] = 32'b11111111111111110100100001100001;
assign LUT_2[50214] = 32'b11111111111111111110100010000100;
assign LUT_2[50215] = 32'b11111111111111111011011010011101;
assign LUT_2[50216] = 32'b11111111111111110101111100111101;
assign LUT_2[50217] = 32'b11111111111111110010110101010110;
assign LUT_2[50218] = 32'b11111111111111111100110101111001;
assign LUT_2[50219] = 32'b11111111111111111001101110010010;
assign LUT_2[50220] = 32'b11111111111111110010011010100101;
assign LUT_2[50221] = 32'b11111111111111101111010010111110;
assign LUT_2[50222] = 32'b11111111111111111001010011100001;
assign LUT_2[50223] = 32'b11111111111111110110001011111010;
assign LUT_2[50224] = 32'b11111111111111110101101111101010;
assign LUT_2[50225] = 32'b11111111111111110010101000000011;
assign LUT_2[50226] = 32'b11111111111111111100101000100110;
assign LUT_2[50227] = 32'b11111111111111111001100000111111;
assign LUT_2[50228] = 32'b11111111111111110010001101010010;
assign LUT_2[50229] = 32'b11111111111111101111000101101011;
assign LUT_2[50230] = 32'b11111111111111111001000110001110;
assign LUT_2[50231] = 32'b11111111111111110101111110100111;
assign LUT_2[50232] = 32'b11111111111111110000100001000111;
assign LUT_2[50233] = 32'b11111111111111101101011001100000;
assign LUT_2[50234] = 32'b11111111111111110111011010000011;
assign LUT_2[50235] = 32'b11111111111111110100010010011100;
assign LUT_2[50236] = 32'b11111111111111101100111110101111;
assign LUT_2[50237] = 32'b11111111111111101001110111001000;
assign LUT_2[50238] = 32'b11111111111111110011110111101011;
assign LUT_2[50239] = 32'b11111111111111110000110000000100;
assign LUT_2[50240] = 32'b11111111111111110010111000011010;
assign LUT_2[50241] = 32'b11111111111111101111110000110011;
assign LUT_2[50242] = 32'b11111111111111111001110001010110;
assign LUT_2[50243] = 32'b11111111111111110110101001101111;
assign LUT_2[50244] = 32'b11111111111111101111010110000010;
assign LUT_2[50245] = 32'b11111111111111101100001110011011;
assign LUT_2[50246] = 32'b11111111111111110110001110111110;
assign LUT_2[50247] = 32'b11111111111111110011000111010111;
assign LUT_2[50248] = 32'b11111111111111101101101001110111;
assign LUT_2[50249] = 32'b11111111111111101010100010010000;
assign LUT_2[50250] = 32'b11111111111111110100100010110011;
assign LUT_2[50251] = 32'b11111111111111110001011011001100;
assign LUT_2[50252] = 32'b11111111111111101010000111011111;
assign LUT_2[50253] = 32'b11111111111111100110111111111000;
assign LUT_2[50254] = 32'b11111111111111110001000000011011;
assign LUT_2[50255] = 32'b11111111111111101101111000110100;
assign LUT_2[50256] = 32'b11111111111111101101011100100100;
assign LUT_2[50257] = 32'b11111111111111101010010100111101;
assign LUT_2[50258] = 32'b11111111111111110100010101100000;
assign LUT_2[50259] = 32'b11111111111111110001001101111001;
assign LUT_2[50260] = 32'b11111111111111101001111010001100;
assign LUT_2[50261] = 32'b11111111111111100110110010100101;
assign LUT_2[50262] = 32'b11111111111111110000110011001000;
assign LUT_2[50263] = 32'b11111111111111101101101011100001;
assign LUT_2[50264] = 32'b11111111111111101000001110000001;
assign LUT_2[50265] = 32'b11111111111111100101000110011010;
assign LUT_2[50266] = 32'b11111111111111101111000110111101;
assign LUT_2[50267] = 32'b11111111111111101011111111010110;
assign LUT_2[50268] = 32'b11111111111111100100101011101001;
assign LUT_2[50269] = 32'b11111111111111100001100100000010;
assign LUT_2[50270] = 32'b11111111111111101011100100100101;
assign LUT_2[50271] = 32'b11111111111111101000011100111110;
assign LUT_2[50272] = 32'b11111111111111110011010100000011;
assign LUT_2[50273] = 32'b11111111111111110000001100011100;
assign LUT_2[50274] = 32'b11111111111111111010001100111111;
assign LUT_2[50275] = 32'b11111111111111110111000101011000;
assign LUT_2[50276] = 32'b11111111111111101111110001101011;
assign LUT_2[50277] = 32'b11111111111111101100101010000100;
assign LUT_2[50278] = 32'b11111111111111110110101010100111;
assign LUT_2[50279] = 32'b11111111111111110011100011000000;
assign LUT_2[50280] = 32'b11111111111111101110000101100000;
assign LUT_2[50281] = 32'b11111111111111101010111101111001;
assign LUT_2[50282] = 32'b11111111111111110100111110011100;
assign LUT_2[50283] = 32'b11111111111111110001110110110101;
assign LUT_2[50284] = 32'b11111111111111101010100011001000;
assign LUT_2[50285] = 32'b11111111111111100111011011100001;
assign LUT_2[50286] = 32'b11111111111111110001011100000100;
assign LUT_2[50287] = 32'b11111111111111101110010100011101;
assign LUT_2[50288] = 32'b11111111111111101101111000001101;
assign LUT_2[50289] = 32'b11111111111111101010110000100110;
assign LUT_2[50290] = 32'b11111111111111110100110001001001;
assign LUT_2[50291] = 32'b11111111111111110001101001100010;
assign LUT_2[50292] = 32'b11111111111111101010010101110101;
assign LUT_2[50293] = 32'b11111111111111100111001110001110;
assign LUT_2[50294] = 32'b11111111111111110001001110110001;
assign LUT_2[50295] = 32'b11111111111111101110000111001010;
assign LUT_2[50296] = 32'b11111111111111101000101001101010;
assign LUT_2[50297] = 32'b11111111111111100101100010000011;
assign LUT_2[50298] = 32'b11111111111111101111100010100110;
assign LUT_2[50299] = 32'b11111111111111101100011010111111;
assign LUT_2[50300] = 32'b11111111111111100101000111010010;
assign LUT_2[50301] = 32'b11111111111111100001111111101011;
assign LUT_2[50302] = 32'b11111111111111101100000000001110;
assign LUT_2[50303] = 32'b11111111111111101000111000100111;
assign LUT_2[50304] = 32'b11111111111111111111000100000110;
assign LUT_2[50305] = 32'b11111111111111111011111100011111;
assign LUT_2[50306] = 32'b00000000000000000101111101000010;
assign LUT_2[50307] = 32'b00000000000000000010110101011011;
assign LUT_2[50308] = 32'b11111111111111111011100001101110;
assign LUT_2[50309] = 32'b11111111111111111000011010000111;
assign LUT_2[50310] = 32'b00000000000000000010011010101010;
assign LUT_2[50311] = 32'b11111111111111111111010011000011;
assign LUT_2[50312] = 32'b11111111111111111001110101100011;
assign LUT_2[50313] = 32'b11111111111111110110101101111100;
assign LUT_2[50314] = 32'b00000000000000000000101110011111;
assign LUT_2[50315] = 32'b11111111111111111101100110111000;
assign LUT_2[50316] = 32'b11111111111111110110010011001011;
assign LUT_2[50317] = 32'b11111111111111110011001011100100;
assign LUT_2[50318] = 32'b11111111111111111101001100000111;
assign LUT_2[50319] = 32'b11111111111111111010000100100000;
assign LUT_2[50320] = 32'b11111111111111111001101000010000;
assign LUT_2[50321] = 32'b11111111111111110110100000101001;
assign LUT_2[50322] = 32'b00000000000000000000100001001100;
assign LUT_2[50323] = 32'b11111111111111111101011001100101;
assign LUT_2[50324] = 32'b11111111111111110110000101111000;
assign LUT_2[50325] = 32'b11111111111111110010111110010001;
assign LUT_2[50326] = 32'b11111111111111111100111110110100;
assign LUT_2[50327] = 32'b11111111111111111001110111001101;
assign LUT_2[50328] = 32'b11111111111111110100011001101101;
assign LUT_2[50329] = 32'b11111111111111110001010010000110;
assign LUT_2[50330] = 32'b11111111111111111011010010101001;
assign LUT_2[50331] = 32'b11111111111111111000001011000010;
assign LUT_2[50332] = 32'b11111111111111110000110111010101;
assign LUT_2[50333] = 32'b11111111111111101101101111101110;
assign LUT_2[50334] = 32'b11111111111111110111110000010001;
assign LUT_2[50335] = 32'b11111111111111110100101000101010;
assign LUT_2[50336] = 32'b11111111111111111111011111101111;
assign LUT_2[50337] = 32'b11111111111111111100011000001000;
assign LUT_2[50338] = 32'b00000000000000000110011000101011;
assign LUT_2[50339] = 32'b00000000000000000011010001000100;
assign LUT_2[50340] = 32'b11111111111111111011111101010111;
assign LUT_2[50341] = 32'b11111111111111111000110101110000;
assign LUT_2[50342] = 32'b00000000000000000010110110010011;
assign LUT_2[50343] = 32'b11111111111111111111101110101100;
assign LUT_2[50344] = 32'b11111111111111111010010001001100;
assign LUT_2[50345] = 32'b11111111111111110111001001100101;
assign LUT_2[50346] = 32'b00000000000000000001001010001000;
assign LUT_2[50347] = 32'b11111111111111111110000010100001;
assign LUT_2[50348] = 32'b11111111111111110110101110110100;
assign LUT_2[50349] = 32'b11111111111111110011100111001101;
assign LUT_2[50350] = 32'b11111111111111111101100111110000;
assign LUT_2[50351] = 32'b11111111111111111010100000001001;
assign LUT_2[50352] = 32'b11111111111111111010000011111001;
assign LUT_2[50353] = 32'b11111111111111110110111100010010;
assign LUT_2[50354] = 32'b00000000000000000000111100110101;
assign LUT_2[50355] = 32'b11111111111111111101110101001110;
assign LUT_2[50356] = 32'b11111111111111110110100001100001;
assign LUT_2[50357] = 32'b11111111111111110011011001111010;
assign LUT_2[50358] = 32'b11111111111111111101011010011101;
assign LUT_2[50359] = 32'b11111111111111111010010010110110;
assign LUT_2[50360] = 32'b11111111111111110100110101010110;
assign LUT_2[50361] = 32'b11111111111111110001101101101111;
assign LUT_2[50362] = 32'b11111111111111111011101110010010;
assign LUT_2[50363] = 32'b11111111111111111000100110101011;
assign LUT_2[50364] = 32'b11111111111111110001010010111110;
assign LUT_2[50365] = 32'b11111111111111101110001011010111;
assign LUT_2[50366] = 32'b11111111111111111000001011111010;
assign LUT_2[50367] = 32'b11111111111111110101000100010011;
assign LUT_2[50368] = 32'b11111111111111110111001100101001;
assign LUT_2[50369] = 32'b11111111111111110100000101000010;
assign LUT_2[50370] = 32'b11111111111111111110000101100101;
assign LUT_2[50371] = 32'b11111111111111111010111101111110;
assign LUT_2[50372] = 32'b11111111111111110011101010010001;
assign LUT_2[50373] = 32'b11111111111111110000100010101010;
assign LUT_2[50374] = 32'b11111111111111111010100011001101;
assign LUT_2[50375] = 32'b11111111111111110111011011100110;
assign LUT_2[50376] = 32'b11111111111111110001111110000110;
assign LUT_2[50377] = 32'b11111111111111101110110110011111;
assign LUT_2[50378] = 32'b11111111111111111000110111000010;
assign LUT_2[50379] = 32'b11111111111111110101101111011011;
assign LUT_2[50380] = 32'b11111111111111101110011011101110;
assign LUT_2[50381] = 32'b11111111111111101011010100000111;
assign LUT_2[50382] = 32'b11111111111111110101010100101010;
assign LUT_2[50383] = 32'b11111111111111110010001101000011;
assign LUT_2[50384] = 32'b11111111111111110001110000110011;
assign LUT_2[50385] = 32'b11111111111111101110101001001100;
assign LUT_2[50386] = 32'b11111111111111111000101001101111;
assign LUT_2[50387] = 32'b11111111111111110101100010001000;
assign LUT_2[50388] = 32'b11111111111111101110001110011011;
assign LUT_2[50389] = 32'b11111111111111101011000110110100;
assign LUT_2[50390] = 32'b11111111111111110101000111010111;
assign LUT_2[50391] = 32'b11111111111111110001111111110000;
assign LUT_2[50392] = 32'b11111111111111101100100010010000;
assign LUT_2[50393] = 32'b11111111111111101001011010101001;
assign LUT_2[50394] = 32'b11111111111111110011011011001100;
assign LUT_2[50395] = 32'b11111111111111110000010011100101;
assign LUT_2[50396] = 32'b11111111111111101000111111111000;
assign LUT_2[50397] = 32'b11111111111111100101111000010001;
assign LUT_2[50398] = 32'b11111111111111101111111000110100;
assign LUT_2[50399] = 32'b11111111111111101100110001001101;
assign LUT_2[50400] = 32'b11111111111111110111101000010010;
assign LUT_2[50401] = 32'b11111111111111110100100000101011;
assign LUT_2[50402] = 32'b11111111111111111110100001001110;
assign LUT_2[50403] = 32'b11111111111111111011011001100111;
assign LUT_2[50404] = 32'b11111111111111110100000101111010;
assign LUT_2[50405] = 32'b11111111111111110000111110010011;
assign LUT_2[50406] = 32'b11111111111111111010111110110110;
assign LUT_2[50407] = 32'b11111111111111110111110111001111;
assign LUT_2[50408] = 32'b11111111111111110010011001101111;
assign LUT_2[50409] = 32'b11111111111111101111010010001000;
assign LUT_2[50410] = 32'b11111111111111111001010010101011;
assign LUT_2[50411] = 32'b11111111111111110110001011000100;
assign LUT_2[50412] = 32'b11111111111111101110110111010111;
assign LUT_2[50413] = 32'b11111111111111101011101111110000;
assign LUT_2[50414] = 32'b11111111111111110101110000010011;
assign LUT_2[50415] = 32'b11111111111111110010101000101100;
assign LUT_2[50416] = 32'b11111111111111110010001100011100;
assign LUT_2[50417] = 32'b11111111111111101111000100110101;
assign LUT_2[50418] = 32'b11111111111111111001000101011000;
assign LUT_2[50419] = 32'b11111111111111110101111101110001;
assign LUT_2[50420] = 32'b11111111111111101110101010000100;
assign LUT_2[50421] = 32'b11111111111111101011100010011101;
assign LUT_2[50422] = 32'b11111111111111110101100011000000;
assign LUT_2[50423] = 32'b11111111111111110010011011011001;
assign LUT_2[50424] = 32'b11111111111111101100111101111001;
assign LUT_2[50425] = 32'b11111111111111101001110110010010;
assign LUT_2[50426] = 32'b11111111111111110011110110110101;
assign LUT_2[50427] = 32'b11111111111111110000101111001110;
assign LUT_2[50428] = 32'b11111111111111101001011011100001;
assign LUT_2[50429] = 32'b11111111111111100110010011111010;
assign LUT_2[50430] = 32'b11111111111111110000010100011101;
assign LUT_2[50431] = 32'b11111111111111101101001100110110;
assign LUT_2[50432] = 32'b11111111111111111110101110011101;
assign LUT_2[50433] = 32'b11111111111111111011100110110110;
assign LUT_2[50434] = 32'b00000000000000000101100111011001;
assign LUT_2[50435] = 32'b00000000000000000010011111110010;
assign LUT_2[50436] = 32'b11111111111111111011001100000101;
assign LUT_2[50437] = 32'b11111111111111111000000100011110;
assign LUT_2[50438] = 32'b00000000000000000010000101000001;
assign LUT_2[50439] = 32'b11111111111111111110111101011010;
assign LUT_2[50440] = 32'b11111111111111111001011111111010;
assign LUT_2[50441] = 32'b11111111111111110110011000010011;
assign LUT_2[50442] = 32'b00000000000000000000011000110110;
assign LUT_2[50443] = 32'b11111111111111111101010001001111;
assign LUT_2[50444] = 32'b11111111111111110101111101100010;
assign LUT_2[50445] = 32'b11111111111111110010110101111011;
assign LUT_2[50446] = 32'b11111111111111111100110110011110;
assign LUT_2[50447] = 32'b11111111111111111001101110110111;
assign LUT_2[50448] = 32'b11111111111111111001010010100111;
assign LUT_2[50449] = 32'b11111111111111110110001011000000;
assign LUT_2[50450] = 32'b00000000000000000000001011100011;
assign LUT_2[50451] = 32'b11111111111111111101000011111100;
assign LUT_2[50452] = 32'b11111111111111110101110000001111;
assign LUT_2[50453] = 32'b11111111111111110010101000101000;
assign LUT_2[50454] = 32'b11111111111111111100101001001011;
assign LUT_2[50455] = 32'b11111111111111111001100001100100;
assign LUT_2[50456] = 32'b11111111111111110100000100000100;
assign LUT_2[50457] = 32'b11111111111111110000111100011101;
assign LUT_2[50458] = 32'b11111111111111111010111101000000;
assign LUT_2[50459] = 32'b11111111111111110111110101011001;
assign LUT_2[50460] = 32'b11111111111111110000100001101100;
assign LUT_2[50461] = 32'b11111111111111101101011010000101;
assign LUT_2[50462] = 32'b11111111111111110111011010101000;
assign LUT_2[50463] = 32'b11111111111111110100010011000001;
assign LUT_2[50464] = 32'b11111111111111111111001010000110;
assign LUT_2[50465] = 32'b11111111111111111100000010011111;
assign LUT_2[50466] = 32'b00000000000000000110000011000010;
assign LUT_2[50467] = 32'b00000000000000000010111011011011;
assign LUT_2[50468] = 32'b11111111111111111011100111101110;
assign LUT_2[50469] = 32'b11111111111111111000100000000111;
assign LUT_2[50470] = 32'b00000000000000000010100000101010;
assign LUT_2[50471] = 32'b11111111111111111111011001000011;
assign LUT_2[50472] = 32'b11111111111111111001111011100011;
assign LUT_2[50473] = 32'b11111111111111110110110011111100;
assign LUT_2[50474] = 32'b00000000000000000000110100011111;
assign LUT_2[50475] = 32'b11111111111111111101101100111000;
assign LUT_2[50476] = 32'b11111111111111110110011001001011;
assign LUT_2[50477] = 32'b11111111111111110011010001100100;
assign LUT_2[50478] = 32'b11111111111111111101010010000111;
assign LUT_2[50479] = 32'b11111111111111111010001010100000;
assign LUT_2[50480] = 32'b11111111111111111001101110010000;
assign LUT_2[50481] = 32'b11111111111111110110100110101001;
assign LUT_2[50482] = 32'b00000000000000000000100111001100;
assign LUT_2[50483] = 32'b11111111111111111101011111100101;
assign LUT_2[50484] = 32'b11111111111111110110001011111000;
assign LUT_2[50485] = 32'b11111111111111110011000100010001;
assign LUT_2[50486] = 32'b11111111111111111101000100110100;
assign LUT_2[50487] = 32'b11111111111111111001111101001101;
assign LUT_2[50488] = 32'b11111111111111110100011111101101;
assign LUT_2[50489] = 32'b11111111111111110001011000000110;
assign LUT_2[50490] = 32'b11111111111111111011011000101001;
assign LUT_2[50491] = 32'b11111111111111111000010001000010;
assign LUT_2[50492] = 32'b11111111111111110000111101010101;
assign LUT_2[50493] = 32'b11111111111111101101110101101110;
assign LUT_2[50494] = 32'b11111111111111110111110110010001;
assign LUT_2[50495] = 32'b11111111111111110100101110101010;
assign LUT_2[50496] = 32'b11111111111111110110110111000000;
assign LUT_2[50497] = 32'b11111111111111110011101111011001;
assign LUT_2[50498] = 32'b11111111111111111101101111111100;
assign LUT_2[50499] = 32'b11111111111111111010101000010101;
assign LUT_2[50500] = 32'b11111111111111110011010100101000;
assign LUT_2[50501] = 32'b11111111111111110000001101000001;
assign LUT_2[50502] = 32'b11111111111111111010001101100100;
assign LUT_2[50503] = 32'b11111111111111110111000101111101;
assign LUT_2[50504] = 32'b11111111111111110001101000011101;
assign LUT_2[50505] = 32'b11111111111111101110100000110110;
assign LUT_2[50506] = 32'b11111111111111111000100001011001;
assign LUT_2[50507] = 32'b11111111111111110101011001110010;
assign LUT_2[50508] = 32'b11111111111111101110000110000101;
assign LUT_2[50509] = 32'b11111111111111101010111110011110;
assign LUT_2[50510] = 32'b11111111111111110100111111000001;
assign LUT_2[50511] = 32'b11111111111111110001110111011010;
assign LUT_2[50512] = 32'b11111111111111110001011011001010;
assign LUT_2[50513] = 32'b11111111111111101110010011100011;
assign LUT_2[50514] = 32'b11111111111111111000010100000110;
assign LUT_2[50515] = 32'b11111111111111110101001100011111;
assign LUT_2[50516] = 32'b11111111111111101101111000110010;
assign LUT_2[50517] = 32'b11111111111111101010110001001011;
assign LUT_2[50518] = 32'b11111111111111110100110001101110;
assign LUT_2[50519] = 32'b11111111111111110001101010000111;
assign LUT_2[50520] = 32'b11111111111111101100001100100111;
assign LUT_2[50521] = 32'b11111111111111101001000101000000;
assign LUT_2[50522] = 32'b11111111111111110011000101100011;
assign LUT_2[50523] = 32'b11111111111111101111111101111100;
assign LUT_2[50524] = 32'b11111111111111101000101010001111;
assign LUT_2[50525] = 32'b11111111111111100101100010101000;
assign LUT_2[50526] = 32'b11111111111111101111100011001011;
assign LUT_2[50527] = 32'b11111111111111101100011011100100;
assign LUT_2[50528] = 32'b11111111111111110111010010101001;
assign LUT_2[50529] = 32'b11111111111111110100001011000010;
assign LUT_2[50530] = 32'b11111111111111111110001011100101;
assign LUT_2[50531] = 32'b11111111111111111011000011111110;
assign LUT_2[50532] = 32'b11111111111111110011110000010001;
assign LUT_2[50533] = 32'b11111111111111110000101000101010;
assign LUT_2[50534] = 32'b11111111111111111010101001001101;
assign LUT_2[50535] = 32'b11111111111111110111100001100110;
assign LUT_2[50536] = 32'b11111111111111110010000100000110;
assign LUT_2[50537] = 32'b11111111111111101110111100011111;
assign LUT_2[50538] = 32'b11111111111111111000111101000010;
assign LUT_2[50539] = 32'b11111111111111110101110101011011;
assign LUT_2[50540] = 32'b11111111111111101110100001101110;
assign LUT_2[50541] = 32'b11111111111111101011011010000111;
assign LUT_2[50542] = 32'b11111111111111110101011010101010;
assign LUT_2[50543] = 32'b11111111111111110010010011000011;
assign LUT_2[50544] = 32'b11111111111111110001110110110011;
assign LUT_2[50545] = 32'b11111111111111101110101111001100;
assign LUT_2[50546] = 32'b11111111111111111000101111101111;
assign LUT_2[50547] = 32'b11111111111111110101101000001000;
assign LUT_2[50548] = 32'b11111111111111101110010100011011;
assign LUT_2[50549] = 32'b11111111111111101011001100110100;
assign LUT_2[50550] = 32'b11111111111111110101001101010111;
assign LUT_2[50551] = 32'b11111111111111110010000101110000;
assign LUT_2[50552] = 32'b11111111111111101100101000010000;
assign LUT_2[50553] = 32'b11111111111111101001100000101001;
assign LUT_2[50554] = 32'b11111111111111110011100001001100;
assign LUT_2[50555] = 32'b11111111111111110000011001100101;
assign LUT_2[50556] = 32'b11111111111111101001000101111000;
assign LUT_2[50557] = 32'b11111111111111100101111110010001;
assign LUT_2[50558] = 32'b11111111111111101111111110110100;
assign LUT_2[50559] = 32'b11111111111111101100110111001101;
assign LUT_2[50560] = 32'b00000000000000000011000010101100;
assign LUT_2[50561] = 32'b11111111111111111111111011000101;
assign LUT_2[50562] = 32'b00000000000000001001111011101000;
assign LUT_2[50563] = 32'b00000000000000000110110100000001;
assign LUT_2[50564] = 32'b11111111111111111111100000010100;
assign LUT_2[50565] = 32'b11111111111111111100011000101101;
assign LUT_2[50566] = 32'b00000000000000000110011001010000;
assign LUT_2[50567] = 32'b00000000000000000011010001101001;
assign LUT_2[50568] = 32'b11111111111111111101110100001001;
assign LUT_2[50569] = 32'b11111111111111111010101100100010;
assign LUT_2[50570] = 32'b00000000000000000100101101000101;
assign LUT_2[50571] = 32'b00000000000000000001100101011110;
assign LUT_2[50572] = 32'b11111111111111111010010001110001;
assign LUT_2[50573] = 32'b11111111111111110111001010001010;
assign LUT_2[50574] = 32'b00000000000000000001001010101101;
assign LUT_2[50575] = 32'b11111111111111111110000011000110;
assign LUT_2[50576] = 32'b11111111111111111101100110110110;
assign LUT_2[50577] = 32'b11111111111111111010011111001111;
assign LUT_2[50578] = 32'b00000000000000000100011111110010;
assign LUT_2[50579] = 32'b00000000000000000001011000001011;
assign LUT_2[50580] = 32'b11111111111111111010000100011110;
assign LUT_2[50581] = 32'b11111111111111110110111100110111;
assign LUT_2[50582] = 32'b00000000000000000000111101011010;
assign LUT_2[50583] = 32'b11111111111111111101110101110011;
assign LUT_2[50584] = 32'b11111111111111111000011000010011;
assign LUT_2[50585] = 32'b11111111111111110101010000101100;
assign LUT_2[50586] = 32'b11111111111111111111010001001111;
assign LUT_2[50587] = 32'b11111111111111111100001001101000;
assign LUT_2[50588] = 32'b11111111111111110100110101111011;
assign LUT_2[50589] = 32'b11111111111111110001101110010100;
assign LUT_2[50590] = 32'b11111111111111111011101110110111;
assign LUT_2[50591] = 32'b11111111111111111000100111010000;
assign LUT_2[50592] = 32'b00000000000000000011011110010101;
assign LUT_2[50593] = 32'b00000000000000000000010110101110;
assign LUT_2[50594] = 32'b00000000000000001010010111010001;
assign LUT_2[50595] = 32'b00000000000000000111001111101010;
assign LUT_2[50596] = 32'b11111111111111111111111011111101;
assign LUT_2[50597] = 32'b11111111111111111100110100010110;
assign LUT_2[50598] = 32'b00000000000000000110110100111001;
assign LUT_2[50599] = 32'b00000000000000000011101101010010;
assign LUT_2[50600] = 32'b11111111111111111110001111110010;
assign LUT_2[50601] = 32'b11111111111111111011001000001011;
assign LUT_2[50602] = 32'b00000000000000000101001000101110;
assign LUT_2[50603] = 32'b00000000000000000010000001000111;
assign LUT_2[50604] = 32'b11111111111111111010101101011010;
assign LUT_2[50605] = 32'b11111111111111110111100101110011;
assign LUT_2[50606] = 32'b00000000000000000001100110010110;
assign LUT_2[50607] = 32'b11111111111111111110011110101111;
assign LUT_2[50608] = 32'b11111111111111111110000010011111;
assign LUT_2[50609] = 32'b11111111111111111010111010111000;
assign LUT_2[50610] = 32'b00000000000000000100111011011011;
assign LUT_2[50611] = 32'b00000000000000000001110011110100;
assign LUT_2[50612] = 32'b11111111111111111010100000000111;
assign LUT_2[50613] = 32'b11111111111111110111011000100000;
assign LUT_2[50614] = 32'b00000000000000000001011001000011;
assign LUT_2[50615] = 32'b11111111111111111110010001011100;
assign LUT_2[50616] = 32'b11111111111111111000110011111100;
assign LUT_2[50617] = 32'b11111111111111110101101100010101;
assign LUT_2[50618] = 32'b11111111111111111111101100111000;
assign LUT_2[50619] = 32'b11111111111111111100100101010001;
assign LUT_2[50620] = 32'b11111111111111110101010001100100;
assign LUT_2[50621] = 32'b11111111111111110010001001111101;
assign LUT_2[50622] = 32'b11111111111111111100001010100000;
assign LUT_2[50623] = 32'b11111111111111111001000010111001;
assign LUT_2[50624] = 32'b11111111111111111011001011001111;
assign LUT_2[50625] = 32'b11111111111111111000000011101000;
assign LUT_2[50626] = 32'b00000000000000000010000100001011;
assign LUT_2[50627] = 32'b11111111111111111110111100100100;
assign LUT_2[50628] = 32'b11111111111111110111101000110111;
assign LUT_2[50629] = 32'b11111111111111110100100001010000;
assign LUT_2[50630] = 32'b11111111111111111110100001110011;
assign LUT_2[50631] = 32'b11111111111111111011011010001100;
assign LUT_2[50632] = 32'b11111111111111110101111100101100;
assign LUT_2[50633] = 32'b11111111111111110010110101000101;
assign LUT_2[50634] = 32'b11111111111111111100110101101000;
assign LUT_2[50635] = 32'b11111111111111111001101110000001;
assign LUT_2[50636] = 32'b11111111111111110010011010010100;
assign LUT_2[50637] = 32'b11111111111111101111010010101101;
assign LUT_2[50638] = 32'b11111111111111111001010011010000;
assign LUT_2[50639] = 32'b11111111111111110110001011101001;
assign LUT_2[50640] = 32'b11111111111111110101101111011001;
assign LUT_2[50641] = 32'b11111111111111110010100111110010;
assign LUT_2[50642] = 32'b11111111111111111100101000010101;
assign LUT_2[50643] = 32'b11111111111111111001100000101110;
assign LUT_2[50644] = 32'b11111111111111110010001101000001;
assign LUT_2[50645] = 32'b11111111111111101111000101011010;
assign LUT_2[50646] = 32'b11111111111111111001000101111101;
assign LUT_2[50647] = 32'b11111111111111110101111110010110;
assign LUT_2[50648] = 32'b11111111111111110000100000110110;
assign LUT_2[50649] = 32'b11111111111111101101011001001111;
assign LUT_2[50650] = 32'b11111111111111110111011001110010;
assign LUT_2[50651] = 32'b11111111111111110100010010001011;
assign LUT_2[50652] = 32'b11111111111111101100111110011110;
assign LUT_2[50653] = 32'b11111111111111101001110110110111;
assign LUT_2[50654] = 32'b11111111111111110011110111011010;
assign LUT_2[50655] = 32'b11111111111111110000101111110011;
assign LUT_2[50656] = 32'b11111111111111111011100110111000;
assign LUT_2[50657] = 32'b11111111111111111000011111010001;
assign LUT_2[50658] = 32'b00000000000000000010011111110100;
assign LUT_2[50659] = 32'b11111111111111111111011000001101;
assign LUT_2[50660] = 32'b11111111111111111000000100100000;
assign LUT_2[50661] = 32'b11111111111111110100111100111001;
assign LUT_2[50662] = 32'b11111111111111111110111101011100;
assign LUT_2[50663] = 32'b11111111111111111011110101110101;
assign LUT_2[50664] = 32'b11111111111111110110011000010101;
assign LUT_2[50665] = 32'b11111111111111110011010000101110;
assign LUT_2[50666] = 32'b11111111111111111101010001010001;
assign LUT_2[50667] = 32'b11111111111111111010001001101010;
assign LUT_2[50668] = 32'b11111111111111110010110101111101;
assign LUT_2[50669] = 32'b11111111111111101111101110010110;
assign LUT_2[50670] = 32'b11111111111111111001101110111001;
assign LUT_2[50671] = 32'b11111111111111110110100111010010;
assign LUT_2[50672] = 32'b11111111111111110110001011000010;
assign LUT_2[50673] = 32'b11111111111111110011000011011011;
assign LUT_2[50674] = 32'b11111111111111111101000011111110;
assign LUT_2[50675] = 32'b11111111111111111001111100010111;
assign LUT_2[50676] = 32'b11111111111111110010101000101010;
assign LUT_2[50677] = 32'b11111111111111101111100001000011;
assign LUT_2[50678] = 32'b11111111111111111001100001100110;
assign LUT_2[50679] = 32'b11111111111111110110011001111111;
assign LUT_2[50680] = 32'b11111111111111110000111100011111;
assign LUT_2[50681] = 32'b11111111111111101101110100111000;
assign LUT_2[50682] = 32'b11111111111111110111110101011011;
assign LUT_2[50683] = 32'b11111111111111110100101101110100;
assign LUT_2[50684] = 32'b11111111111111101101011010000111;
assign LUT_2[50685] = 32'b11111111111111101010010010100000;
assign LUT_2[50686] = 32'b11111111111111110100010011000011;
assign LUT_2[50687] = 32'b11111111111111110001001011011100;
assign LUT_2[50688] = 32'b11111111111111111111100001101001;
assign LUT_2[50689] = 32'b11111111111111111100011010000010;
assign LUT_2[50690] = 32'b00000000000000000110011010100101;
assign LUT_2[50691] = 32'b00000000000000000011010010111110;
assign LUT_2[50692] = 32'b11111111111111111011111111010001;
assign LUT_2[50693] = 32'b11111111111111111000110111101010;
assign LUT_2[50694] = 32'b00000000000000000010111000001101;
assign LUT_2[50695] = 32'b11111111111111111111110000100110;
assign LUT_2[50696] = 32'b11111111111111111010010011000110;
assign LUT_2[50697] = 32'b11111111111111110111001011011111;
assign LUT_2[50698] = 32'b00000000000000000001001100000010;
assign LUT_2[50699] = 32'b11111111111111111110000100011011;
assign LUT_2[50700] = 32'b11111111111111110110110000101110;
assign LUT_2[50701] = 32'b11111111111111110011101001000111;
assign LUT_2[50702] = 32'b11111111111111111101101001101010;
assign LUT_2[50703] = 32'b11111111111111111010100010000011;
assign LUT_2[50704] = 32'b11111111111111111010000101110011;
assign LUT_2[50705] = 32'b11111111111111110110111110001100;
assign LUT_2[50706] = 32'b00000000000000000000111110101111;
assign LUT_2[50707] = 32'b11111111111111111101110111001000;
assign LUT_2[50708] = 32'b11111111111111110110100011011011;
assign LUT_2[50709] = 32'b11111111111111110011011011110100;
assign LUT_2[50710] = 32'b11111111111111111101011100010111;
assign LUT_2[50711] = 32'b11111111111111111010010100110000;
assign LUT_2[50712] = 32'b11111111111111110100110111010000;
assign LUT_2[50713] = 32'b11111111111111110001101111101001;
assign LUT_2[50714] = 32'b11111111111111111011110000001100;
assign LUT_2[50715] = 32'b11111111111111111000101000100101;
assign LUT_2[50716] = 32'b11111111111111110001010100111000;
assign LUT_2[50717] = 32'b11111111111111101110001101010001;
assign LUT_2[50718] = 32'b11111111111111111000001101110100;
assign LUT_2[50719] = 32'b11111111111111110101000110001101;
assign LUT_2[50720] = 32'b11111111111111111111111101010010;
assign LUT_2[50721] = 32'b11111111111111111100110101101011;
assign LUT_2[50722] = 32'b00000000000000000110110110001110;
assign LUT_2[50723] = 32'b00000000000000000011101110100111;
assign LUT_2[50724] = 32'b11111111111111111100011010111010;
assign LUT_2[50725] = 32'b11111111111111111001010011010011;
assign LUT_2[50726] = 32'b00000000000000000011010011110110;
assign LUT_2[50727] = 32'b00000000000000000000001100001111;
assign LUT_2[50728] = 32'b11111111111111111010101110101111;
assign LUT_2[50729] = 32'b11111111111111110111100111001000;
assign LUT_2[50730] = 32'b00000000000000000001100111101011;
assign LUT_2[50731] = 32'b11111111111111111110100000000100;
assign LUT_2[50732] = 32'b11111111111111110111001100010111;
assign LUT_2[50733] = 32'b11111111111111110100000100110000;
assign LUT_2[50734] = 32'b11111111111111111110000101010011;
assign LUT_2[50735] = 32'b11111111111111111010111101101100;
assign LUT_2[50736] = 32'b11111111111111111010100001011100;
assign LUT_2[50737] = 32'b11111111111111110111011001110101;
assign LUT_2[50738] = 32'b00000000000000000001011010011000;
assign LUT_2[50739] = 32'b11111111111111111110010010110001;
assign LUT_2[50740] = 32'b11111111111111110110111111000100;
assign LUT_2[50741] = 32'b11111111111111110011110111011101;
assign LUT_2[50742] = 32'b11111111111111111101111000000000;
assign LUT_2[50743] = 32'b11111111111111111010110000011001;
assign LUT_2[50744] = 32'b11111111111111110101010010111001;
assign LUT_2[50745] = 32'b11111111111111110010001011010010;
assign LUT_2[50746] = 32'b11111111111111111100001011110101;
assign LUT_2[50747] = 32'b11111111111111111001000100001110;
assign LUT_2[50748] = 32'b11111111111111110001110000100001;
assign LUT_2[50749] = 32'b11111111111111101110101000111010;
assign LUT_2[50750] = 32'b11111111111111111000101001011101;
assign LUT_2[50751] = 32'b11111111111111110101100001110110;
assign LUT_2[50752] = 32'b11111111111111110111101010001100;
assign LUT_2[50753] = 32'b11111111111111110100100010100101;
assign LUT_2[50754] = 32'b11111111111111111110100011001000;
assign LUT_2[50755] = 32'b11111111111111111011011011100001;
assign LUT_2[50756] = 32'b11111111111111110100000111110100;
assign LUT_2[50757] = 32'b11111111111111110001000000001101;
assign LUT_2[50758] = 32'b11111111111111111011000000110000;
assign LUT_2[50759] = 32'b11111111111111110111111001001001;
assign LUT_2[50760] = 32'b11111111111111110010011011101001;
assign LUT_2[50761] = 32'b11111111111111101111010100000010;
assign LUT_2[50762] = 32'b11111111111111111001010100100101;
assign LUT_2[50763] = 32'b11111111111111110110001100111110;
assign LUT_2[50764] = 32'b11111111111111101110111001010001;
assign LUT_2[50765] = 32'b11111111111111101011110001101010;
assign LUT_2[50766] = 32'b11111111111111110101110010001101;
assign LUT_2[50767] = 32'b11111111111111110010101010100110;
assign LUT_2[50768] = 32'b11111111111111110010001110010110;
assign LUT_2[50769] = 32'b11111111111111101111000110101111;
assign LUT_2[50770] = 32'b11111111111111111001000111010010;
assign LUT_2[50771] = 32'b11111111111111110101111111101011;
assign LUT_2[50772] = 32'b11111111111111101110101011111110;
assign LUT_2[50773] = 32'b11111111111111101011100100010111;
assign LUT_2[50774] = 32'b11111111111111110101100100111010;
assign LUT_2[50775] = 32'b11111111111111110010011101010011;
assign LUT_2[50776] = 32'b11111111111111101100111111110011;
assign LUT_2[50777] = 32'b11111111111111101001111000001100;
assign LUT_2[50778] = 32'b11111111111111110011111000101111;
assign LUT_2[50779] = 32'b11111111111111110000110001001000;
assign LUT_2[50780] = 32'b11111111111111101001011101011011;
assign LUT_2[50781] = 32'b11111111111111100110010101110100;
assign LUT_2[50782] = 32'b11111111111111110000010110010111;
assign LUT_2[50783] = 32'b11111111111111101101001110110000;
assign LUT_2[50784] = 32'b11111111111111111000000101110101;
assign LUT_2[50785] = 32'b11111111111111110100111110001110;
assign LUT_2[50786] = 32'b11111111111111111110111110110001;
assign LUT_2[50787] = 32'b11111111111111111011110111001010;
assign LUT_2[50788] = 32'b11111111111111110100100011011101;
assign LUT_2[50789] = 32'b11111111111111110001011011110110;
assign LUT_2[50790] = 32'b11111111111111111011011100011001;
assign LUT_2[50791] = 32'b11111111111111111000010100110010;
assign LUT_2[50792] = 32'b11111111111111110010110111010010;
assign LUT_2[50793] = 32'b11111111111111101111101111101011;
assign LUT_2[50794] = 32'b11111111111111111001110000001110;
assign LUT_2[50795] = 32'b11111111111111110110101000100111;
assign LUT_2[50796] = 32'b11111111111111101111010100111010;
assign LUT_2[50797] = 32'b11111111111111101100001101010011;
assign LUT_2[50798] = 32'b11111111111111110110001101110110;
assign LUT_2[50799] = 32'b11111111111111110011000110001111;
assign LUT_2[50800] = 32'b11111111111111110010101001111111;
assign LUT_2[50801] = 32'b11111111111111101111100010011000;
assign LUT_2[50802] = 32'b11111111111111111001100010111011;
assign LUT_2[50803] = 32'b11111111111111110110011011010100;
assign LUT_2[50804] = 32'b11111111111111101111000111100111;
assign LUT_2[50805] = 32'b11111111111111101100000000000000;
assign LUT_2[50806] = 32'b11111111111111110110000000100011;
assign LUT_2[50807] = 32'b11111111111111110010111000111100;
assign LUT_2[50808] = 32'b11111111111111101101011011011100;
assign LUT_2[50809] = 32'b11111111111111101010010011110101;
assign LUT_2[50810] = 32'b11111111111111110100010100011000;
assign LUT_2[50811] = 32'b11111111111111110001001100110001;
assign LUT_2[50812] = 32'b11111111111111101001111001000100;
assign LUT_2[50813] = 32'b11111111111111100110110001011101;
assign LUT_2[50814] = 32'b11111111111111110000110010000000;
assign LUT_2[50815] = 32'b11111111111111101101101010011001;
assign LUT_2[50816] = 32'b00000000000000000011110101111000;
assign LUT_2[50817] = 32'b00000000000000000000101110010001;
assign LUT_2[50818] = 32'b00000000000000001010101110110100;
assign LUT_2[50819] = 32'b00000000000000000111100111001101;
assign LUT_2[50820] = 32'b00000000000000000000010011100000;
assign LUT_2[50821] = 32'b11111111111111111101001011111001;
assign LUT_2[50822] = 32'b00000000000000000111001100011100;
assign LUT_2[50823] = 32'b00000000000000000100000100110101;
assign LUT_2[50824] = 32'b11111111111111111110100111010101;
assign LUT_2[50825] = 32'b11111111111111111011011111101110;
assign LUT_2[50826] = 32'b00000000000000000101100000010001;
assign LUT_2[50827] = 32'b00000000000000000010011000101010;
assign LUT_2[50828] = 32'b11111111111111111011000100111101;
assign LUT_2[50829] = 32'b11111111111111110111111101010110;
assign LUT_2[50830] = 32'b00000000000000000001111101111001;
assign LUT_2[50831] = 32'b11111111111111111110110110010010;
assign LUT_2[50832] = 32'b11111111111111111110011010000010;
assign LUT_2[50833] = 32'b11111111111111111011010010011011;
assign LUT_2[50834] = 32'b00000000000000000101010010111110;
assign LUT_2[50835] = 32'b00000000000000000010001011010111;
assign LUT_2[50836] = 32'b11111111111111111010110111101010;
assign LUT_2[50837] = 32'b11111111111111110111110000000011;
assign LUT_2[50838] = 32'b00000000000000000001110000100110;
assign LUT_2[50839] = 32'b11111111111111111110101000111111;
assign LUT_2[50840] = 32'b11111111111111111001001011011111;
assign LUT_2[50841] = 32'b11111111111111110110000011111000;
assign LUT_2[50842] = 32'b00000000000000000000000100011011;
assign LUT_2[50843] = 32'b11111111111111111100111100110100;
assign LUT_2[50844] = 32'b11111111111111110101101001000111;
assign LUT_2[50845] = 32'b11111111111111110010100001100000;
assign LUT_2[50846] = 32'b11111111111111111100100010000011;
assign LUT_2[50847] = 32'b11111111111111111001011010011100;
assign LUT_2[50848] = 32'b00000000000000000100010001100001;
assign LUT_2[50849] = 32'b00000000000000000001001001111010;
assign LUT_2[50850] = 32'b00000000000000001011001010011101;
assign LUT_2[50851] = 32'b00000000000000001000000010110110;
assign LUT_2[50852] = 32'b00000000000000000000101111001001;
assign LUT_2[50853] = 32'b11111111111111111101100111100010;
assign LUT_2[50854] = 32'b00000000000000000111101000000101;
assign LUT_2[50855] = 32'b00000000000000000100100000011110;
assign LUT_2[50856] = 32'b11111111111111111111000010111110;
assign LUT_2[50857] = 32'b11111111111111111011111011010111;
assign LUT_2[50858] = 32'b00000000000000000101111011111010;
assign LUT_2[50859] = 32'b00000000000000000010110100010011;
assign LUT_2[50860] = 32'b11111111111111111011100000100110;
assign LUT_2[50861] = 32'b11111111111111111000011000111111;
assign LUT_2[50862] = 32'b00000000000000000010011001100010;
assign LUT_2[50863] = 32'b11111111111111111111010001111011;
assign LUT_2[50864] = 32'b11111111111111111110110101101011;
assign LUT_2[50865] = 32'b11111111111111111011101110000100;
assign LUT_2[50866] = 32'b00000000000000000101101110100111;
assign LUT_2[50867] = 32'b00000000000000000010100111000000;
assign LUT_2[50868] = 32'b11111111111111111011010011010011;
assign LUT_2[50869] = 32'b11111111111111111000001011101100;
assign LUT_2[50870] = 32'b00000000000000000010001100001111;
assign LUT_2[50871] = 32'b11111111111111111111000100101000;
assign LUT_2[50872] = 32'b11111111111111111001100111001000;
assign LUT_2[50873] = 32'b11111111111111110110011111100001;
assign LUT_2[50874] = 32'b00000000000000000000100000000100;
assign LUT_2[50875] = 32'b11111111111111111101011000011101;
assign LUT_2[50876] = 32'b11111111111111110110000100110000;
assign LUT_2[50877] = 32'b11111111111111110010111101001001;
assign LUT_2[50878] = 32'b11111111111111111100111101101100;
assign LUT_2[50879] = 32'b11111111111111111001110110000101;
assign LUT_2[50880] = 32'b11111111111111111011111110011011;
assign LUT_2[50881] = 32'b11111111111111111000110110110100;
assign LUT_2[50882] = 32'b00000000000000000010110111010111;
assign LUT_2[50883] = 32'b11111111111111111111101111110000;
assign LUT_2[50884] = 32'b11111111111111111000011100000011;
assign LUT_2[50885] = 32'b11111111111111110101010100011100;
assign LUT_2[50886] = 32'b11111111111111111111010100111111;
assign LUT_2[50887] = 32'b11111111111111111100001101011000;
assign LUT_2[50888] = 32'b11111111111111110110101111111000;
assign LUT_2[50889] = 32'b11111111111111110011101000010001;
assign LUT_2[50890] = 32'b11111111111111111101101000110100;
assign LUT_2[50891] = 32'b11111111111111111010100001001101;
assign LUT_2[50892] = 32'b11111111111111110011001101100000;
assign LUT_2[50893] = 32'b11111111111111110000000101111001;
assign LUT_2[50894] = 32'b11111111111111111010000110011100;
assign LUT_2[50895] = 32'b11111111111111110110111110110101;
assign LUT_2[50896] = 32'b11111111111111110110100010100101;
assign LUT_2[50897] = 32'b11111111111111110011011010111110;
assign LUT_2[50898] = 32'b11111111111111111101011011100001;
assign LUT_2[50899] = 32'b11111111111111111010010011111010;
assign LUT_2[50900] = 32'b11111111111111110011000000001101;
assign LUT_2[50901] = 32'b11111111111111101111111000100110;
assign LUT_2[50902] = 32'b11111111111111111001111001001001;
assign LUT_2[50903] = 32'b11111111111111110110110001100010;
assign LUT_2[50904] = 32'b11111111111111110001010100000010;
assign LUT_2[50905] = 32'b11111111111111101110001100011011;
assign LUT_2[50906] = 32'b11111111111111111000001100111110;
assign LUT_2[50907] = 32'b11111111111111110101000101010111;
assign LUT_2[50908] = 32'b11111111111111101101110001101010;
assign LUT_2[50909] = 32'b11111111111111101010101010000011;
assign LUT_2[50910] = 32'b11111111111111110100101010100110;
assign LUT_2[50911] = 32'b11111111111111110001100010111111;
assign LUT_2[50912] = 32'b11111111111111111100011010000100;
assign LUT_2[50913] = 32'b11111111111111111001010010011101;
assign LUT_2[50914] = 32'b00000000000000000011010011000000;
assign LUT_2[50915] = 32'b00000000000000000000001011011001;
assign LUT_2[50916] = 32'b11111111111111111000110111101100;
assign LUT_2[50917] = 32'b11111111111111110101110000000101;
assign LUT_2[50918] = 32'b11111111111111111111110000101000;
assign LUT_2[50919] = 32'b11111111111111111100101001000001;
assign LUT_2[50920] = 32'b11111111111111110111001011100001;
assign LUT_2[50921] = 32'b11111111111111110100000011111010;
assign LUT_2[50922] = 32'b11111111111111111110000100011101;
assign LUT_2[50923] = 32'b11111111111111111010111100110110;
assign LUT_2[50924] = 32'b11111111111111110011101001001001;
assign LUT_2[50925] = 32'b11111111111111110000100001100010;
assign LUT_2[50926] = 32'b11111111111111111010100010000101;
assign LUT_2[50927] = 32'b11111111111111110111011010011110;
assign LUT_2[50928] = 32'b11111111111111110110111110001110;
assign LUT_2[50929] = 32'b11111111111111110011110110100111;
assign LUT_2[50930] = 32'b11111111111111111101110111001010;
assign LUT_2[50931] = 32'b11111111111111111010101111100011;
assign LUT_2[50932] = 32'b11111111111111110011011011110110;
assign LUT_2[50933] = 32'b11111111111111110000010100001111;
assign LUT_2[50934] = 32'b11111111111111111010010100110010;
assign LUT_2[50935] = 32'b11111111111111110111001101001011;
assign LUT_2[50936] = 32'b11111111111111110001101111101011;
assign LUT_2[50937] = 32'b11111111111111101110101000000100;
assign LUT_2[50938] = 32'b11111111111111111000101000100111;
assign LUT_2[50939] = 32'b11111111111111110101100001000000;
assign LUT_2[50940] = 32'b11111111111111101110001101010011;
assign LUT_2[50941] = 32'b11111111111111101011000101101100;
assign LUT_2[50942] = 32'b11111111111111110101000110001111;
assign LUT_2[50943] = 32'b11111111111111110001111110101000;
assign LUT_2[50944] = 32'b00000000000000000011100000001111;
assign LUT_2[50945] = 32'b00000000000000000000011000101000;
assign LUT_2[50946] = 32'b00000000000000001010011001001011;
assign LUT_2[50947] = 32'b00000000000000000111010001100100;
assign LUT_2[50948] = 32'b11111111111111111111111101110111;
assign LUT_2[50949] = 32'b11111111111111111100110110010000;
assign LUT_2[50950] = 32'b00000000000000000110110110110011;
assign LUT_2[50951] = 32'b00000000000000000011101111001100;
assign LUT_2[50952] = 32'b11111111111111111110010001101100;
assign LUT_2[50953] = 32'b11111111111111111011001010000101;
assign LUT_2[50954] = 32'b00000000000000000101001010101000;
assign LUT_2[50955] = 32'b00000000000000000010000011000001;
assign LUT_2[50956] = 32'b11111111111111111010101111010100;
assign LUT_2[50957] = 32'b11111111111111110111100111101101;
assign LUT_2[50958] = 32'b00000000000000000001101000010000;
assign LUT_2[50959] = 32'b11111111111111111110100000101001;
assign LUT_2[50960] = 32'b11111111111111111110000100011001;
assign LUT_2[50961] = 32'b11111111111111111010111100110010;
assign LUT_2[50962] = 32'b00000000000000000100111101010101;
assign LUT_2[50963] = 32'b00000000000000000001110101101110;
assign LUT_2[50964] = 32'b11111111111111111010100010000001;
assign LUT_2[50965] = 32'b11111111111111110111011010011010;
assign LUT_2[50966] = 32'b00000000000000000001011010111101;
assign LUT_2[50967] = 32'b11111111111111111110010011010110;
assign LUT_2[50968] = 32'b11111111111111111000110101110110;
assign LUT_2[50969] = 32'b11111111111111110101101110001111;
assign LUT_2[50970] = 32'b11111111111111111111101110110010;
assign LUT_2[50971] = 32'b11111111111111111100100111001011;
assign LUT_2[50972] = 32'b11111111111111110101010011011110;
assign LUT_2[50973] = 32'b11111111111111110010001011110111;
assign LUT_2[50974] = 32'b11111111111111111100001100011010;
assign LUT_2[50975] = 32'b11111111111111111001000100110011;
assign LUT_2[50976] = 32'b00000000000000000011111011111000;
assign LUT_2[50977] = 32'b00000000000000000000110100010001;
assign LUT_2[50978] = 32'b00000000000000001010110100110100;
assign LUT_2[50979] = 32'b00000000000000000111101101001101;
assign LUT_2[50980] = 32'b00000000000000000000011001100000;
assign LUT_2[50981] = 32'b11111111111111111101010001111001;
assign LUT_2[50982] = 32'b00000000000000000111010010011100;
assign LUT_2[50983] = 32'b00000000000000000100001010110101;
assign LUT_2[50984] = 32'b11111111111111111110101101010101;
assign LUT_2[50985] = 32'b11111111111111111011100101101110;
assign LUT_2[50986] = 32'b00000000000000000101100110010001;
assign LUT_2[50987] = 32'b00000000000000000010011110101010;
assign LUT_2[50988] = 32'b11111111111111111011001010111101;
assign LUT_2[50989] = 32'b11111111111111111000000011010110;
assign LUT_2[50990] = 32'b00000000000000000010000011111001;
assign LUT_2[50991] = 32'b11111111111111111110111100010010;
assign LUT_2[50992] = 32'b11111111111111111110100000000010;
assign LUT_2[50993] = 32'b11111111111111111011011000011011;
assign LUT_2[50994] = 32'b00000000000000000101011000111110;
assign LUT_2[50995] = 32'b00000000000000000010010001010111;
assign LUT_2[50996] = 32'b11111111111111111010111101101010;
assign LUT_2[50997] = 32'b11111111111111110111110110000011;
assign LUT_2[50998] = 32'b00000000000000000001110110100110;
assign LUT_2[50999] = 32'b11111111111111111110101110111111;
assign LUT_2[51000] = 32'b11111111111111111001010001011111;
assign LUT_2[51001] = 32'b11111111111111110110001001111000;
assign LUT_2[51002] = 32'b00000000000000000000001010011011;
assign LUT_2[51003] = 32'b11111111111111111101000010110100;
assign LUT_2[51004] = 32'b11111111111111110101101111000111;
assign LUT_2[51005] = 32'b11111111111111110010100111100000;
assign LUT_2[51006] = 32'b11111111111111111100101000000011;
assign LUT_2[51007] = 32'b11111111111111111001100000011100;
assign LUT_2[51008] = 32'b11111111111111111011101000110010;
assign LUT_2[51009] = 32'b11111111111111111000100001001011;
assign LUT_2[51010] = 32'b00000000000000000010100001101110;
assign LUT_2[51011] = 32'b11111111111111111111011010000111;
assign LUT_2[51012] = 32'b11111111111111111000000110011010;
assign LUT_2[51013] = 32'b11111111111111110100111110110011;
assign LUT_2[51014] = 32'b11111111111111111110111111010110;
assign LUT_2[51015] = 32'b11111111111111111011110111101111;
assign LUT_2[51016] = 32'b11111111111111110110011010001111;
assign LUT_2[51017] = 32'b11111111111111110011010010101000;
assign LUT_2[51018] = 32'b11111111111111111101010011001011;
assign LUT_2[51019] = 32'b11111111111111111010001011100100;
assign LUT_2[51020] = 32'b11111111111111110010110111110111;
assign LUT_2[51021] = 32'b11111111111111101111110000010000;
assign LUT_2[51022] = 32'b11111111111111111001110000110011;
assign LUT_2[51023] = 32'b11111111111111110110101001001100;
assign LUT_2[51024] = 32'b11111111111111110110001100111100;
assign LUT_2[51025] = 32'b11111111111111110011000101010101;
assign LUT_2[51026] = 32'b11111111111111111101000101111000;
assign LUT_2[51027] = 32'b11111111111111111001111110010001;
assign LUT_2[51028] = 32'b11111111111111110010101010100100;
assign LUT_2[51029] = 32'b11111111111111101111100010111101;
assign LUT_2[51030] = 32'b11111111111111111001100011100000;
assign LUT_2[51031] = 32'b11111111111111110110011011111001;
assign LUT_2[51032] = 32'b11111111111111110000111110011001;
assign LUT_2[51033] = 32'b11111111111111101101110110110010;
assign LUT_2[51034] = 32'b11111111111111110111110111010101;
assign LUT_2[51035] = 32'b11111111111111110100101111101110;
assign LUT_2[51036] = 32'b11111111111111101101011100000001;
assign LUT_2[51037] = 32'b11111111111111101010010100011010;
assign LUT_2[51038] = 32'b11111111111111110100010100111101;
assign LUT_2[51039] = 32'b11111111111111110001001101010110;
assign LUT_2[51040] = 32'b11111111111111111100000100011011;
assign LUT_2[51041] = 32'b11111111111111111000111100110100;
assign LUT_2[51042] = 32'b00000000000000000010111101010111;
assign LUT_2[51043] = 32'b11111111111111111111110101110000;
assign LUT_2[51044] = 32'b11111111111111111000100010000011;
assign LUT_2[51045] = 32'b11111111111111110101011010011100;
assign LUT_2[51046] = 32'b11111111111111111111011010111111;
assign LUT_2[51047] = 32'b11111111111111111100010011011000;
assign LUT_2[51048] = 32'b11111111111111110110110101111000;
assign LUT_2[51049] = 32'b11111111111111110011101110010001;
assign LUT_2[51050] = 32'b11111111111111111101101110110100;
assign LUT_2[51051] = 32'b11111111111111111010100111001101;
assign LUT_2[51052] = 32'b11111111111111110011010011100000;
assign LUT_2[51053] = 32'b11111111111111110000001011111001;
assign LUT_2[51054] = 32'b11111111111111111010001100011100;
assign LUT_2[51055] = 32'b11111111111111110111000100110101;
assign LUT_2[51056] = 32'b11111111111111110110101000100101;
assign LUT_2[51057] = 32'b11111111111111110011100000111110;
assign LUT_2[51058] = 32'b11111111111111111101100001100001;
assign LUT_2[51059] = 32'b11111111111111111010011001111010;
assign LUT_2[51060] = 32'b11111111111111110011000110001101;
assign LUT_2[51061] = 32'b11111111111111101111111110100110;
assign LUT_2[51062] = 32'b11111111111111111001111111001001;
assign LUT_2[51063] = 32'b11111111111111110110110111100010;
assign LUT_2[51064] = 32'b11111111111111110001011010000010;
assign LUT_2[51065] = 32'b11111111111111101110010010011011;
assign LUT_2[51066] = 32'b11111111111111111000010010111110;
assign LUT_2[51067] = 32'b11111111111111110101001011010111;
assign LUT_2[51068] = 32'b11111111111111101101110111101010;
assign LUT_2[51069] = 32'b11111111111111101010110000000011;
assign LUT_2[51070] = 32'b11111111111111110100110000100110;
assign LUT_2[51071] = 32'b11111111111111110001101000111111;
assign LUT_2[51072] = 32'b00000000000000000111110100011110;
assign LUT_2[51073] = 32'b00000000000000000100101100110111;
assign LUT_2[51074] = 32'b00000000000000001110101101011010;
assign LUT_2[51075] = 32'b00000000000000001011100101110011;
assign LUT_2[51076] = 32'b00000000000000000100010010000110;
assign LUT_2[51077] = 32'b00000000000000000001001010011111;
assign LUT_2[51078] = 32'b00000000000000001011001011000010;
assign LUT_2[51079] = 32'b00000000000000001000000011011011;
assign LUT_2[51080] = 32'b00000000000000000010100101111011;
assign LUT_2[51081] = 32'b11111111111111111111011110010100;
assign LUT_2[51082] = 32'b00000000000000001001011110110111;
assign LUT_2[51083] = 32'b00000000000000000110010111010000;
assign LUT_2[51084] = 32'b11111111111111111111000011100011;
assign LUT_2[51085] = 32'b11111111111111111011111011111100;
assign LUT_2[51086] = 32'b00000000000000000101111100011111;
assign LUT_2[51087] = 32'b00000000000000000010110100111000;
assign LUT_2[51088] = 32'b00000000000000000010011000101000;
assign LUT_2[51089] = 32'b11111111111111111111010001000001;
assign LUT_2[51090] = 32'b00000000000000001001010001100100;
assign LUT_2[51091] = 32'b00000000000000000110001001111101;
assign LUT_2[51092] = 32'b11111111111111111110110110010000;
assign LUT_2[51093] = 32'b11111111111111111011101110101001;
assign LUT_2[51094] = 32'b00000000000000000101101111001100;
assign LUT_2[51095] = 32'b00000000000000000010100111100101;
assign LUT_2[51096] = 32'b11111111111111111101001010000101;
assign LUT_2[51097] = 32'b11111111111111111010000010011110;
assign LUT_2[51098] = 32'b00000000000000000100000011000001;
assign LUT_2[51099] = 32'b00000000000000000000111011011010;
assign LUT_2[51100] = 32'b11111111111111111001100111101101;
assign LUT_2[51101] = 32'b11111111111111110110100000000110;
assign LUT_2[51102] = 32'b00000000000000000000100000101001;
assign LUT_2[51103] = 32'b11111111111111111101011001000010;
assign LUT_2[51104] = 32'b00000000000000001000010000000111;
assign LUT_2[51105] = 32'b00000000000000000101001000100000;
assign LUT_2[51106] = 32'b00000000000000001111001001000011;
assign LUT_2[51107] = 32'b00000000000000001100000001011100;
assign LUT_2[51108] = 32'b00000000000000000100101101101111;
assign LUT_2[51109] = 32'b00000000000000000001100110001000;
assign LUT_2[51110] = 32'b00000000000000001011100110101011;
assign LUT_2[51111] = 32'b00000000000000001000011111000100;
assign LUT_2[51112] = 32'b00000000000000000011000001100100;
assign LUT_2[51113] = 32'b11111111111111111111111001111101;
assign LUT_2[51114] = 32'b00000000000000001001111010100000;
assign LUT_2[51115] = 32'b00000000000000000110110010111001;
assign LUT_2[51116] = 32'b11111111111111111111011111001100;
assign LUT_2[51117] = 32'b11111111111111111100010111100101;
assign LUT_2[51118] = 32'b00000000000000000110011000001000;
assign LUT_2[51119] = 32'b00000000000000000011010000100001;
assign LUT_2[51120] = 32'b00000000000000000010110100010001;
assign LUT_2[51121] = 32'b11111111111111111111101100101010;
assign LUT_2[51122] = 32'b00000000000000001001101101001101;
assign LUT_2[51123] = 32'b00000000000000000110100101100110;
assign LUT_2[51124] = 32'b11111111111111111111010001111001;
assign LUT_2[51125] = 32'b11111111111111111100001010010010;
assign LUT_2[51126] = 32'b00000000000000000110001010110101;
assign LUT_2[51127] = 32'b00000000000000000011000011001110;
assign LUT_2[51128] = 32'b11111111111111111101100101101110;
assign LUT_2[51129] = 32'b11111111111111111010011110000111;
assign LUT_2[51130] = 32'b00000000000000000100011110101010;
assign LUT_2[51131] = 32'b00000000000000000001010111000011;
assign LUT_2[51132] = 32'b11111111111111111010000011010110;
assign LUT_2[51133] = 32'b11111111111111110110111011101111;
assign LUT_2[51134] = 32'b00000000000000000000111100010010;
assign LUT_2[51135] = 32'b11111111111111111101110100101011;
assign LUT_2[51136] = 32'b11111111111111111111111101000001;
assign LUT_2[51137] = 32'b11111111111111111100110101011010;
assign LUT_2[51138] = 32'b00000000000000000110110101111101;
assign LUT_2[51139] = 32'b00000000000000000011101110010110;
assign LUT_2[51140] = 32'b11111111111111111100011010101001;
assign LUT_2[51141] = 32'b11111111111111111001010011000010;
assign LUT_2[51142] = 32'b00000000000000000011010011100101;
assign LUT_2[51143] = 32'b00000000000000000000001011111110;
assign LUT_2[51144] = 32'b11111111111111111010101110011110;
assign LUT_2[51145] = 32'b11111111111111110111100110110111;
assign LUT_2[51146] = 32'b00000000000000000001100111011010;
assign LUT_2[51147] = 32'b11111111111111111110011111110011;
assign LUT_2[51148] = 32'b11111111111111110111001100000110;
assign LUT_2[51149] = 32'b11111111111111110100000100011111;
assign LUT_2[51150] = 32'b11111111111111111110000101000010;
assign LUT_2[51151] = 32'b11111111111111111010111101011011;
assign LUT_2[51152] = 32'b11111111111111111010100001001011;
assign LUT_2[51153] = 32'b11111111111111110111011001100100;
assign LUT_2[51154] = 32'b00000000000000000001011010000111;
assign LUT_2[51155] = 32'b11111111111111111110010010100000;
assign LUT_2[51156] = 32'b11111111111111110110111110110011;
assign LUT_2[51157] = 32'b11111111111111110011110111001100;
assign LUT_2[51158] = 32'b11111111111111111101110111101111;
assign LUT_2[51159] = 32'b11111111111111111010110000001000;
assign LUT_2[51160] = 32'b11111111111111110101010010101000;
assign LUT_2[51161] = 32'b11111111111111110010001011000001;
assign LUT_2[51162] = 32'b11111111111111111100001011100100;
assign LUT_2[51163] = 32'b11111111111111111001000011111101;
assign LUT_2[51164] = 32'b11111111111111110001110000010000;
assign LUT_2[51165] = 32'b11111111111111101110101000101001;
assign LUT_2[51166] = 32'b11111111111111111000101001001100;
assign LUT_2[51167] = 32'b11111111111111110101100001100101;
assign LUT_2[51168] = 32'b00000000000000000000011000101010;
assign LUT_2[51169] = 32'b11111111111111111101010001000011;
assign LUT_2[51170] = 32'b00000000000000000111010001100110;
assign LUT_2[51171] = 32'b00000000000000000100001001111111;
assign LUT_2[51172] = 32'b11111111111111111100110110010010;
assign LUT_2[51173] = 32'b11111111111111111001101110101011;
assign LUT_2[51174] = 32'b00000000000000000011101111001110;
assign LUT_2[51175] = 32'b00000000000000000000100111100111;
assign LUT_2[51176] = 32'b11111111111111111011001010000111;
assign LUT_2[51177] = 32'b11111111111111111000000010100000;
assign LUT_2[51178] = 32'b00000000000000000010000011000011;
assign LUT_2[51179] = 32'b11111111111111111110111011011100;
assign LUT_2[51180] = 32'b11111111111111110111100111101111;
assign LUT_2[51181] = 32'b11111111111111110100100000001000;
assign LUT_2[51182] = 32'b11111111111111111110100000101011;
assign LUT_2[51183] = 32'b11111111111111111011011001000100;
assign LUT_2[51184] = 32'b11111111111111111010111100110100;
assign LUT_2[51185] = 32'b11111111111111110111110101001101;
assign LUT_2[51186] = 32'b00000000000000000001110101110000;
assign LUT_2[51187] = 32'b11111111111111111110101110001001;
assign LUT_2[51188] = 32'b11111111111111110111011010011100;
assign LUT_2[51189] = 32'b11111111111111110100010010110101;
assign LUT_2[51190] = 32'b11111111111111111110010011011000;
assign LUT_2[51191] = 32'b11111111111111111011001011110001;
assign LUT_2[51192] = 32'b11111111111111110101101110010001;
assign LUT_2[51193] = 32'b11111111111111110010100110101010;
assign LUT_2[51194] = 32'b11111111111111111100100111001101;
assign LUT_2[51195] = 32'b11111111111111111001011111100110;
assign LUT_2[51196] = 32'b11111111111111110010001011111001;
assign LUT_2[51197] = 32'b11111111111111101111000100010010;
assign LUT_2[51198] = 32'b11111111111111111001000100110101;
assign LUT_2[51199] = 32'b11111111111111110101111101001110;
assign LUT_2[51200] = 32'b11111111111111101111111001101110;
assign LUT_2[51201] = 32'b11111111111111101100110010000111;
assign LUT_2[51202] = 32'b11111111111111110110110010101010;
assign LUT_2[51203] = 32'b11111111111111110011101011000011;
assign LUT_2[51204] = 32'b11111111111111101100010111010110;
assign LUT_2[51205] = 32'b11111111111111101001001111101111;
assign LUT_2[51206] = 32'b11111111111111110011010000010010;
assign LUT_2[51207] = 32'b11111111111111110000001000101011;
assign LUT_2[51208] = 32'b11111111111111101010101011001011;
assign LUT_2[51209] = 32'b11111111111111100111100011100100;
assign LUT_2[51210] = 32'b11111111111111110001100100000111;
assign LUT_2[51211] = 32'b11111111111111101110011100100000;
assign LUT_2[51212] = 32'b11111111111111100111001000110011;
assign LUT_2[51213] = 32'b11111111111111100100000001001100;
assign LUT_2[51214] = 32'b11111111111111101110000001101111;
assign LUT_2[51215] = 32'b11111111111111101010111010001000;
assign LUT_2[51216] = 32'b11111111111111101010011101111000;
assign LUT_2[51217] = 32'b11111111111111100111010110010001;
assign LUT_2[51218] = 32'b11111111111111110001010110110100;
assign LUT_2[51219] = 32'b11111111111111101110001111001101;
assign LUT_2[51220] = 32'b11111111111111100110111011100000;
assign LUT_2[51221] = 32'b11111111111111100011110011111001;
assign LUT_2[51222] = 32'b11111111111111101101110100011100;
assign LUT_2[51223] = 32'b11111111111111101010101100110101;
assign LUT_2[51224] = 32'b11111111111111100101001111010101;
assign LUT_2[51225] = 32'b11111111111111100010000111101110;
assign LUT_2[51226] = 32'b11111111111111101100001000010001;
assign LUT_2[51227] = 32'b11111111111111101001000000101010;
assign LUT_2[51228] = 32'b11111111111111100001101100111101;
assign LUT_2[51229] = 32'b11111111111111011110100101010110;
assign LUT_2[51230] = 32'b11111111111111101000100101111001;
assign LUT_2[51231] = 32'b11111111111111100101011110010010;
assign LUT_2[51232] = 32'b11111111111111110000010101010111;
assign LUT_2[51233] = 32'b11111111111111101101001101110000;
assign LUT_2[51234] = 32'b11111111111111110111001110010011;
assign LUT_2[51235] = 32'b11111111111111110100000110101100;
assign LUT_2[51236] = 32'b11111111111111101100110010111111;
assign LUT_2[51237] = 32'b11111111111111101001101011011000;
assign LUT_2[51238] = 32'b11111111111111110011101011111011;
assign LUT_2[51239] = 32'b11111111111111110000100100010100;
assign LUT_2[51240] = 32'b11111111111111101011000110110100;
assign LUT_2[51241] = 32'b11111111111111100111111111001101;
assign LUT_2[51242] = 32'b11111111111111110001111111110000;
assign LUT_2[51243] = 32'b11111111111111101110111000001001;
assign LUT_2[51244] = 32'b11111111111111100111100100011100;
assign LUT_2[51245] = 32'b11111111111111100100011100110101;
assign LUT_2[51246] = 32'b11111111111111101110011101011000;
assign LUT_2[51247] = 32'b11111111111111101011010101110001;
assign LUT_2[51248] = 32'b11111111111111101010111001100001;
assign LUT_2[51249] = 32'b11111111111111100111110001111010;
assign LUT_2[51250] = 32'b11111111111111110001110010011101;
assign LUT_2[51251] = 32'b11111111111111101110101010110110;
assign LUT_2[51252] = 32'b11111111111111100111010111001001;
assign LUT_2[51253] = 32'b11111111111111100100001111100010;
assign LUT_2[51254] = 32'b11111111111111101110010000000101;
assign LUT_2[51255] = 32'b11111111111111101011001000011110;
assign LUT_2[51256] = 32'b11111111111111100101101010111110;
assign LUT_2[51257] = 32'b11111111111111100010100011010111;
assign LUT_2[51258] = 32'b11111111111111101100100011111010;
assign LUT_2[51259] = 32'b11111111111111101001011100010011;
assign LUT_2[51260] = 32'b11111111111111100010001000100110;
assign LUT_2[51261] = 32'b11111111111111011111000000111111;
assign LUT_2[51262] = 32'b11111111111111101001000001100010;
assign LUT_2[51263] = 32'b11111111111111100101111001111011;
assign LUT_2[51264] = 32'b11111111111111101000000010010001;
assign LUT_2[51265] = 32'b11111111111111100100111010101010;
assign LUT_2[51266] = 32'b11111111111111101110111011001101;
assign LUT_2[51267] = 32'b11111111111111101011110011100110;
assign LUT_2[51268] = 32'b11111111111111100100011111111001;
assign LUT_2[51269] = 32'b11111111111111100001011000010010;
assign LUT_2[51270] = 32'b11111111111111101011011000110101;
assign LUT_2[51271] = 32'b11111111111111101000010001001110;
assign LUT_2[51272] = 32'b11111111111111100010110011101110;
assign LUT_2[51273] = 32'b11111111111111011111101100000111;
assign LUT_2[51274] = 32'b11111111111111101001101100101010;
assign LUT_2[51275] = 32'b11111111111111100110100101000011;
assign LUT_2[51276] = 32'b11111111111111011111010001010110;
assign LUT_2[51277] = 32'b11111111111111011100001001101111;
assign LUT_2[51278] = 32'b11111111111111100110001010010010;
assign LUT_2[51279] = 32'b11111111111111100011000010101011;
assign LUT_2[51280] = 32'b11111111111111100010100110011011;
assign LUT_2[51281] = 32'b11111111111111011111011110110100;
assign LUT_2[51282] = 32'b11111111111111101001011111010111;
assign LUT_2[51283] = 32'b11111111111111100110010111110000;
assign LUT_2[51284] = 32'b11111111111111011111000100000011;
assign LUT_2[51285] = 32'b11111111111111011011111100011100;
assign LUT_2[51286] = 32'b11111111111111100101111100111111;
assign LUT_2[51287] = 32'b11111111111111100010110101011000;
assign LUT_2[51288] = 32'b11111111111111011101010111111000;
assign LUT_2[51289] = 32'b11111111111111011010010000010001;
assign LUT_2[51290] = 32'b11111111111111100100010000110100;
assign LUT_2[51291] = 32'b11111111111111100001001001001101;
assign LUT_2[51292] = 32'b11111111111111011001110101100000;
assign LUT_2[51293] = 32'b11111111111111010110101101111001;
assign LUT_2[51294] = 32'b11111111111111100000101110011100;
assign LUT_2[51295] = 32'b11111111111111011101100110110101;
assign LUT_2[51296] = 32'b11111111111111101000011101111010;
assign LUT_2[51297] = 32'b11111111111111100101010110010011;
assign LUT_2[51298] = 32'b11111111111111101111010110110110;
assign LUT_2[51299] = 32'b11111111111111101100001111001111;
assign LUT_2[51300] = 32'b11111111111111100100111011100010;
assign LUT_2[51301] = 32'b11111111111111100001110011111011;
assign LUT_2[51302] = 32'b11111111111111101011110100011110;
assign LUT_2[51303] = 32'b11111111111111101000101100110111;
assign LUT_2[51304] = 32'b11111111111111100011001111010111;
assign LUT_2[51305] = 32'b11111111111111100000000111110000;
assign LUT_2[51306] = 32'b11111111111111101010001000010011;
assign LUT_2[51307] = 32'b11111111111111100111000000101100;
assign LUT_2[51308] = 32'b11111111111111011111101100111111;
assign LUT_2[51309] = 32'b11111111111111011100100101011000;
assign LUT_2[51310] = 32'b11111111111111100110100101111011;
assign LUT_2[51311] = 32'b11111111111111100011011110010100;
assign LUT_2[51312] = 32'b11111111111111100011000010000100;
assign LUT_2[51313] = 32'b11111111111111011111111010011101;
assign LUT_2[51314] = 32'b11111111111111101001111011000000;
assign LUT_2[51315] = 32'b11111111111111100110110011011001;
assign LUT_2[51316] = 32'b11111111111111011111011111101100;
assign LUT_2[51317] = 32'b11111111111111011100011000000101;
assign LUT_2[51318] = 32'b11111111111111100110011000101000;
assign LUT_2[51319] = 32'b11111111111111100011010001000001;
assign LUT_2[51320] = 32'b11111111111111011101110011100001;
assign LUT_2[51321] = 32'b11111111111111011010101011111010;
assign LUT_2[51322] = 32'b11111111111111100100101100011101;
assign LUT_2[51323] = 32'b11111111111111100001100100110110;
assign LUT_2[51324] = 32'b11111111111111011010010001001001;
assign LUT_2[51325] = 32'b11111111111111010111001001100010;
assign LUT_2[51326] = 32'b11111111111111100001001010000101;
assign LUT_2[51327] = 32'b11111111111111011110000010011110;
assign LUT_2[51328] = 32'b11111111111111110100001101111101;
assign LUT_2[51329] = 32'b11111111111111110001000110010110;
assign LUT_2[51330] = 32'b11111111111111111011000110111001;
assign LUT_2[51331] = 32'b11111111111111110111111111010010;
assign LUT_2[51332] = 32'b11111111111111110000101011100101;
assign LUT_2[51333] = 32'b11111111111111101101100011111110;
assign LUT_2[51334] = 32'b11111111111111110111100100100001;
assign LUT_2[51335] = 32'b11111111111111110100011100111010;
assign LUT_2[51336] = 32'b11111111111111101110111111011010;
assign LUT_2[51337] = 32'b11111111111111101011110111110011;
assign LUT_2[51338] = 32'b11111111111111110101111000010110;
assign LUT_2[51339] = 32'b11111111111111110010110000101111;
assign LUT_2[51340] = 32'b11111111111111101011011101000010;
assign LUT_2[51341] = 32'b11111111111111101000010101011011;
assign LUT_2[51342] = 32'b11111111111111110010010101111110;
assign LUT_2[51343] = 32'b11111111111111101111001110010111;
assign LUT_2[51344] = 32'b11111111111111101110110010000111;
assign LUT_2[51345] = 32'b11111111111111101011101010100000;
assign LUT_2[51346] = 32'b11111111111111110101101011000011;
assign LUT_2[51347] = 32'b11111111111111110010100011011100;
assign LUT_2[51348] = 32'b11111111111111101011001111101111;
assign LUT_2[51349] = 32'b11111111111111101000001000001000;
assign LUT_2[51350] = 32'b11111111111111110010001000101011;
assign LUT_2[51351] = 32'b11111111111111101111000001000100;
assign LUT_2[51352] = 32'b11111111111111101001100011100100;
assign LUT_2[51353] = 32'b11111111111111100110011011111101;
assign LUT_2[51354] = 32'b11111111111111110000011100100000;
assign LUT_2[51355] = 32'b11111111111111101101010100111001;
assign LUT_2[51356] = 32'b11111111111111100110000001001100;
assign LUT_2[51357] = 32'b11111111111111100010111001100101;
assign LUT_2[51358] = 32'b11111111111111101100111010001000;
assign LUT_2[51359] = 32'b11111111111111101001110010100001;
assign LUT_2[51360] = 32'b11111111111111110100101001100110;
assign LUT_2[51361] = 32'b11111111111111110001100001111111;
assign LUT_2[51362] = 32'b11111111111111111011100010100010;
assign LUT_2[51363] = 32'b11111111111111111000011010111011;
assign LUT_2[51364] = 32'b11111111111111110001000111001110;
assign LUT_2[51365] = 32'b11111111111111101101111111100111;
assign LUT_2[51366] = 32'b11111111111111111000000000001010;
assign LUT_2[51367] = 32'b11111111111111110100111000100011;
assign LUT_2[51368] = 32'b11111111111111101111011011000011;
assign LUT_2[51369] = 32'b11111111111111101100010011011100;
assign LUT_2[51370] = 32'b11111111111111110110010011111111;
assign LUT_2[51371] = 32'b11111111111111110011001100011000;
assign LUT_2[51372] = 32'b11111111111111101011111000101011;
assign LUT_2[51373] = 32'b11111111111111101000110001000100;
assign LUT_2[51374] = 32'b11111111111111110010110001100111;
assign LUT_2[51375] = 32'b11111111111111101111101010000000;
assign LUT_2[51376] = 32'b11111111111111101111001101110000;
assign LUT_2[51377] = 32'b11111111111111101100000110001001;
assign LUT_2[51378] = 32'b11111111111111110110000110101100;
assign LUT_2[51379] = 32'b11111111111111110010111111000101;
assign LUT_2[51380] = 32'b11111111111111101011101011011000;
assign LUT_2[51381] = 32'b11111111111111101000100011110001;
assign LUT_2[51382] = 32'b11111111111111110010100100010100;
assign LUT_2[51383] = 32'b11111111111111101111011100101101;
assign LUT_2[51384] = 32'b11111111111111101001111111001101;
assign LUT_2[51385] = 32'b11111111111111100110110111100110;
assign LUT_2[51386] = 32'b11111111111111110000111000001001;
assign LUT_2[51387] = 32'b11111111111111101101110000100010;
assign LUT_2[51388] = 32'b11111111111111100110011100110101;
assign LUT_2[51389] = 32'b11111111111111100011010101001110;
assign LUT_2[51390] = 32'b11111111111111101101010101110001;
assign LUT_2[51391] = 32'b11111111111111101010001110001010;
assign LUT_2[51392] = 32'b11111111111111101100010110100000;
assign LUT_2[51393] = 32'b11111111111111101001001110111001;
assign LUT_2[51394] = 32'b11111111111111110011001111011100;
assign LUT_2[51395] = 32'b11111111111111110000000111110101;
assign LUT_2[51396] = 32'b11111111111111101000110100001000;
assign LUT_2[51397] = 32'b11111111111111100101101100100001;
assign LUT_2[51398] = 32'b11111111111111101111101101000100;
assign LUT_2[51399] = 32'b11111111111111101100100101011101;
assign LUT_2[51400] = 32'b11111111111111100111000111111101;
assign LUT_2[51401] = 32'b11111111111111100100000000010110;
assign LUT_2[51402] = 32'b11111111111111101110000000111001;
assign LUT_2[51403] = 32'b11111111111111101010111001010010;
assign LUT_2[51404] = 32'b11111111111111100011100101100101;
assign LUT_2[51405] = 32'b11111111111111100000011101111110;
assign LUT_2[51406] = 32'b11111111111111101010011110100001;
assign LUT_2[51407] = 32'b11111111111111100111010110111010;
assign LUT_2[51408] = 32'b11111111111111100110111010101010;
assign LUT_2[51409] = 32'b11111111111111100011110011000011;
assign LUT_2[51410] = 32'b11111111111111101101110011100110;
assign LUT_2[51411] = 32'b11111111111111101010101011111111;
assign LUT_2[51412] = 32'b11111111111111100011011000010010;
assign LUT_2[51413] = 32'b11111111111111100000010000101011;
assign LUT_2[51414] = 32'b11111111111111101010010001001110;
assign LUT_2[51415] = 32'b11111111111111100111001001100111;
assign LUT_2[51416] = 32'b11111111111111100001101100000111;
assign LUT_2[51417] = 32'b11111111111111011110100100100000;
assign LUT_2[51418] = 32'b11111111111111101000100101000011;
assign LUT_2[51419] = 32'b11111111111111100101011101011100;
assign LUT_2[51420] = 32'b11111111111111011110001001101111;
assign LUT_2[51421] = 32'b11111111111111011011000010001000;
assign LUT_2[51422] = 32'b11111111111111100101000010101011;
assign LUT_2[51423] = 32'b11111111111111100001111011000100;
assign LUT_2[51424] = 32'b11111111111111101100110010001001;
assign LUT_2[51425] = 32'b11111111111111101001101010100010;
assign LUT_2[51426] = 32'b11111111111111110011101011000101;
assign LUT_2[51427] = 32'b11111111111111110000100011011110;
assign LUT_2[51428] = 32'b11111111111111101001001111110001;
assign LUT_2[51429] = 32'b11111111111111100110001000001010;
assign LUT_2[51430] = 32'b11111111111111110000001000101101;
assign LUT_2[51431] = 32'b11111111111111101101000001000110;
assign LUT_2[51432] = 32'b11111111111111100111100011100110;
assign LUT_2[51433] = 32'b11111111111111100100011011111111;
assign LUT_2[51434] = 32'b11111111111111101110011100100010;
assign LUT_2[51435] = 32'b11111111111111101011010100111011;
assign LUT_2[51436] = 32'b11111111111111100100000001001110;
assign LUT_2[51437] = 32'b11111111111111100000111001100111;
assign LUT_2[51438] = 32'b11111111111111101010111010001010;
assign LUT_2[51439] = 32'b11111111111111100111110010100011;
assign LUT_2[51440] = 32'b11111111111111100111010110010011;
assign LUT_2[51441] = 32'b11111111111111100100001110101100;
assign LUT_2[51442] = 32'b11111111111111101110001111001111;
assign LUT_2[51443] = 32'b11111111111111101011000111101000;
assign LUT_2[51444] = 32'b11111111111111100011110011111011;
assign LUT_2[51445] = 32'b11111111111111100000101100010100;
assign LUT_2[51446] = 32'b11111111111111101010101100110111;
assign LUT_2[51447] = 32'b11111111111111100111100101010000;
assign LUT_2[51448] = 32'b11111111111111100010000111110000;
assign LUT_2[51449] = 32'b11111111111111011111000000001001;
assign LUT_2[51450] = 32'b11111111111111101001000000101100;
assign LUT_2[51451] = 32'b11111111111111100101111001000101;
assign LUT_2[51452] = 32'b11111111111111011110100101011000;
assign LUT_2[51453] = 32'b11111111111111011011011101110001;
assign LUT_2[51454] = 32'b11111111111111100101011110010100;
assign LUT_2[51455] = 32'b11111111111111100010010110101101;
assign LUT_2[51456] = 32'b11111111111111110011111000010100;
assign LUT_2[51457] = 32'b11111111111111110000110000101101;
assign LUT_2[51458] = 32'b11111111111111111010110001010000;
assign LUT_2[51459] = 32'b11111111111111110111101001101001;
assign LUT_2[51460] = 32'b11111111111111110000010101111100;
assign LUT_2[51461] = 32'b11111111111111101101001110010101;
assign LUT_2[51462] = 32'b11111111111111110111001110111000;
assign LUT_2[51463] = 32'b11111111111111110100000111010001;
assign LUT_2[51464] = 32'b11111111111111101110101001110001;
assign LUT_2[51465] = 32'b11111111111111101011100010001010;
assign LUT_2[51466] = 32'b11111111111111110101100010101101;
assign LUT_2[51467] = 32'b11111111111111110010011011000110;
assign LUT_2[51468] = 32'b11111111111111101011000111011001;
assign LUT_2[51469] = 32'b11111111111111100111111111110010;
assign LUT_2[51470] = 32'b11111111111111110010000000010101;
assign LUT_2[51471] = 32'b11111111111111101110111000101110;
assign LUT_2[51472] = 32'b11111111111111101110011100011110;
assign LUT_2[51473] = 32'b11111111111111101011010100110111;
assign LUT_2[51474] = 32'b11111111111111110101010101011010;
assign LUT_2[51475] = 32'b11111111111111110010001101110011;
assign LUT_2[51476] = 32'b11111111111111101010111010000110;
assign LUT_2[51477] = 32'b11111111111111100111110010011111;
assign LUT_2[51478] = 32'b11111111111111110001110011000010;
assign LUT_2[51479] = 32'b11111111111111101110101011011011;
assign LUT_2[51480] = 32'b11111111111111101001001101111011;
assign LUT_2[51481] = 32'b11111111111111100110000110010100;
assign LUT_2[51482] = 32'b11111111111111110000000110110111;
assign LUT_2[51483] = 32'b11111111111111101100111111010000;
assign LUT_2[51484] = 32'b11111111111111100101101011100011;
assign LUT_2[51485] = 32'b11111111111111100010100011111100;
assign LUT_2[51486] = 32'b11111111111111101100100100011111;
assign LUT_2[51487] = 32'b11111111111111101001011100111000;
assign LUT_2[51488] = 32'b11111111111111110100010011111101;
assign LUT_2[51489] = 32'b11111111111111110001001100010110;
assign LUT_2[51490] = 32'b11111111111111111011001100111001;
assign LUT_2[51491] = 32'b11111111111111111000000101010010;
assign LUT_2[51492] = 32'b11111111111111110000110001100101;
assign LUT_2[51493] = 32'b11111111111111101101101001111110;
assign LUT_2[51494] = 32'b11111111111111110111101010100001;
assign LUT_2[51495] = 32'b11111111111111110100100010111010;
assign LUT_2[51496] = 32'b11111111111111101111000101011010;
assign LUT_2[51497] = 32'b11111111111111101011111101110011;
assign LUT_2[51498] = 32'b11111111111111110101111110010110;
assign LUT_2[51499] = 32'b11111111111111110010110110101111;
assign LUT_2[51500] = 32'b11111111111111101011100011000010;
assign LUT_2[51501] = 32'b11111111111111101000011011011011;
assign LUT_2[51502] = 32'b11111111111111110010011011111110;
assign LUT_2[51503] = 32'b11111111111111101111010100010111;
assign LUT_2[51504] = 32'b11111111111111101110111000000111;
assign LUT_2[51505] = 32'b11111111111111101011110000100000;
assign LUT_2[51506] = 32'b11111111111111110101110001000011;
assign LUT_2[51507] = 32'b11111111111111110010101001011100;
assign LUT_2[51508] = 32'b11111111111111101011010101101111;
assign LUT_2[51509] = 32'b11111111111111101000001110001000;
assign LUT_2[51510] = 32'b11111111111111110010001110101011;
assign LUT_2[51511] = 32'b11111111111111101111000111000100;
assign LUT_2[51512] = 32'b11111111111111101001101001100100;
assign LUT_2[51513] = 32'b11111111111111100110100001111101;
assign LUT_2[51514] = 32'b11111111111111110000100010100000;
assign LUT_2[51515] = 32'b11111111111111101101011010111001;
assign LUT_2[51516] = 32'b11111111111111100110000111001100;
assign LUT_2[51517] = 32'b11111111111111100010111111100101;
assign LUT_2[51518] = 32'b11111111111111101101000000001000;
assign LUT_2[51519] = 32'b11111111111111101001111000100001;
assign LUT_2[51520] = 32'b11111111111111101100000000110111;
assign LUT_2[51521] = 32'b11111111111111101000111001010000;
assign LUT_2[51522] = 32'b11111111111111110010111001110011;
assign LUT_2[51523] = 32'b11111111111111101111110010001100;
assign LUT_2[51524] = 32'b11111111111111101000011110011111;
assign LUT_2[51525] = 32'b11111111111111100101010110111000;
assign LUT_2[51526] = 32'b11111111111111101111010111011011;
assign LUT_2[51527] = 32'b11111111111111101100001111110100;
assign LUT_2[51528] = 32'b11111111111111100110110010010100;
assign LUT_2[51529] = 32'b11111111111111100011101010101101;
assign LUT_2[51530] = 32'b11111111111111101101101011010000;
assign LUT_2[51531] = 32'b11111111111111101010100011101001;
assign LUT_2[51532] = 32'b11111111111111100011001111111100;
assign LUT_2[51533] = 32'b11111111111111100000001000010101;
assign LUT_2[51534] = 32'b11111111111111101010001000111000;
assign LUT_2[51535] = 32'b11111111111111100111000001010001;
assign LUT_2[51536] = 32'b11111111111111100110100101000001;
assign LUT_2[51537] = 32'b11111111111111100011011101011010;
assign LUT_2[51538] = 32'b11111111111111101101011101111101;
assign LUT_2[51539] = 32'b11111111111111101010010110010110;
assign LUT_2[51540] = 32'b11111111111111100011000010101001;
assign LUT_2[51541] = 32'b11111111111111011111111011000010;
assign LUT_2[51542] = 32'b11111111111111101001111011100101;
assign LUT_2[51543] = 32'b11111111111111100110110011111110;
assign LUT_2[51544] = 32'b11111111111111100001010110011110;
assign LUT_2[51545] = 32'b11111111111111011110001110110111;
assign LUT_2[51546] = 32'b11111111111111101000001111011010;
assign LUT_2[51547] = 32'b11111111111111100101000111110011;
assign LUT_2[51548] = 32'b11111111111111011101110100000110;
assign LUT_2[51549] = 32'b11111111111111011010101100011111;
assign LUT_2[51550] = 32'b11111111111111100100101101000010;
assign LUT_2[51551] = 32'b11111111111111100001100101011011;
assign LUT_2[51552] = 32'b11111111111111101100011100100000;
assign LUT_2[51553] = 32'b11111111111111101001010100111001;
assign LUT_2[51554] = 32'b11111111111111110011010101011100;
assign LUT_2[51555] = 32'b11111111111111110000001101110101;
assign LUT_2[51556] = 32'b11111111111111101000111010001000;
assign LUT_2[51557] = 32'b11111111111111100101110010100001;
assign LUT_2[51558] = 32'b11111111111111101111110011000100;
assign LUT_2[51559] = 32'b11111111111111101100101011011101;
assign LUT_2[51560] = 32'b11111111111111100111001101111101;
assign LUT_2[51561] = 32'b11111111111111100100000110010110;
assign LUT_2[51562] = 32'b11111111111111101110000110111001;
assign LUT_2[51563] = 32'b11111111111111101010111111010010;
assign LUT_2[51564] = 32'b11111111111111100011101011100101;
assign LUT_2[51565] = 32'b11111111111111100000100011111110;
assign LUT_2[51566] = 32'b11111111111111101010100100100001;
assign LUT_2[51567] = 32'b11111111111111100111011100111010;
assign LUT_2[51568] = 32'b11111111111111100111000000101010;
assign LUT_2[51569] = 32'b11111111111111100011111001000011;
assign LUT_2[51570] = 32'b11111111111111101101111001100110;
assign LUT_2[51571] = 32'b11111111111111101010110001111111;
assign LUT_2[51572] = 32'b11111111111111100011011110010010;
assign LUT_2[51573] = 32'b11111111111111100000010110101011;
assign LUT_2[51574] = 32'b11111111111111101010010111001110;
assign LUT_2[51575] = 32'b11111111111111100111001111100111;
assign LUT_2[51576] = 32'b11111111111111100001110010000111;
assign LUT_2[51577] = 32'b11111111111111011110101010100000;
assign LUT_2[51578] = 32'b11111111111111101000101011000011;
assign LUT_2[51579] = 32'b11111111111111100101100011011100;
assign LUT_2[51580] = 32'b11111111111111011110001111101111;
assign LUT_2[51581] = 32'b11111111111111011011001000001000;
assign LUT_2[51582] = 32'b11111111111111100101001000101011;
assign LUT_2[51583] = 32'b11111111111111100010000001000100;
assign LUT_2[51584] = 32'b11111111111111111000001100100011;
assign LUT_2[51585] = 32'b11111111111111110101000100111100;
assign LUT_2[51586] = 32'b11111111111111111111000101011111;
assign LUT_2[51587] = 32'b11111111111111111011111101111000;
assign LUT_2[51588] = 32'b11111111111111110100101010001011;
assign LUT_2[51589] = 32'b11111111111111110001100010100100;
assign LUT_2[51590] = 32'b11111111111111111011100011000111;
assign LUT_2[51591] = 32'b11111111111111111000011011100000;
assign LUT_2[51592] = 32'b11111111111111110010111110000000;
assign LUT_2[51593] = 32'b11111111111111101111110110011001;
assign LUT_2[51594] = 32'b11111111111111111001110110111100;
assign LUT_2[51595] = 32'b11111111111111110110101111010101;
assign LUT_2[51596] = 32'b11111111111111101111011011101000;
assign LUT_2[51597] = 32'b11111111111111101100010100000001;
assign LUT_2[51598] = 32'b11111111111111110110010100100100;
assign LUT_2[51599] = 32'b11111111111111110011001100111101;
assign LUT_2[51600] = 32'b11111111111111110010110000101101;
assign LUT_2[51601] = 32'b11111111111111101111101001000110;
assign LUT_2[51602] = 32'b11111111111111111001101001101001;
assign LUT_2[51603] = 32'b11111111111111110110100010000010;
assign LUT_2[51604] = 32'b11111111111111101111001110010101;
assign LUT_2[51605] = 32'b11111111111111101100000110101110;
assign LUT_2[51606] = 32'b11111111111111110110000111010001;
assign LUT_2[51607] = 32'b11111111111111110010111111101010;
assign LUT_2[51608] = 32'b11111111111111101101100010001010;
assign LUT_2[51609] = 32'b11111111111111101010011010100011;
assign LUT_2[51610] = 32'b11111111111111110100011011000110;
assign LUT_2[51611] = 32'b11111111111111110001010011011111;
assign LUT_2[51612] = 32'b11111111111111101001111111110010;
assign LUT_2[51613] = 32'b11111111111111100110111000001011;
assign LUT_2[51614] = 32'b11111111111111110000111000101110;
assign LUT_2[51615] = 32'b11111111111111101101110001000111;
assign LUT_2[51616] = 32'b11111111111111111000101000001100;
assign LUT_2[51617] = 32'b11111111111111110101100000100101;
assign LUT_2[51618] = 32'b11111111111111111111100001001000;
assign LUT_2[51619] = 32'b11111111111111111100011001100001;
assign LUT_2[51620] = 32'b11111111111111110101000101110100;
assign LUT_2[51621] = 32'b11111111111111110001111110001101;
assign LUT_2[51622] = 32'b11111111111111111011111110110000;
assign LUT_2[51623] = 32'b11111111111111111000110111001001;
assign LUT_2[51624] = 32'b11111111111111110011011001101001;
assign LUT_2[51625] = 32'b11111111111111110000010010000010;
assign LUT_2[51626] = 32'b11111111111111111010010010100101;
assign LUT_2[51627] = 32'b11111111111111110111001010111110;
assign LUT_2[51628] = 32'b11111111111111101111110111010001;
assign LUT_2[51629] = 32'b11111111111111101100101111101010;
assign LUT_2[51630] = 32'b11111111111111110110110000001101;
assign LUT_2[51631] = 32'b11111111111111110011101000100110;
assign LUT_2[51632] = 32'b11111111111111110011001100010110;
assign LUT_2[51633] = 32'b11111111111111110000000100101111;
assign LUT_2[51634] = 32'b11111111111111111010000101010010;
assign LUT_2[51635] = 32'b11111111111111110110111101101011;
assign LUT_2[51636] = 32'b11111111111111101111101001111110;
assign LUT_2[51637] = 32'b11111111111111101100100010010111;
assign LUT_2[51638] = 32'b11111111111111110110100010111010;
assign LUT_2[51639] = 32'b11111111111111110011011011010011;
assign LUT_2[51640] = 32'b11111111111111101101111101110011;
assign LUT_2[51641] = 32'b11111111111111101010110110001100;
assign LUT_2[51642] = 32'b11111111111111110100110110101111;
assign LUT_2[51643] = 32'b11111111111111110001101111001000;
assign LUT_2[51644] = 32'b11111111111111101010011011011011;
assign LUT_2[51645] = 32'b11111111111111100111010011110100;
assign LUT_2[51646] = 32'b11111111111111110001010100010111;
assign LUT_2[51647] = 32'b11111111111111101110001100110000;
assign LUT_2[51648] = 32'b11111111111111110000010101000110;
assign LUT_2[51649] = 32'b11111111111111101101001101011111;
assign LUT_2[51650] = 32'b11111111111111110111001110000010;
assign LUT_2[51651] = 32'b11111111111111110100000110011011;
assign LUT_2[51652] = 32'b11111111111111101100110010101110;
assign LUT_2[51653] = 32'b11111111111111101001101011000111;
assign LUT_2[51654] = 32'b11111111111111110011101011101010;
assign LUT_2[51655] = 32'b11111111111111110000100100000011;
assign LUT_2[51656] = 32'b11111111111111101011000110100011;
assign LUT_2[51657] = 32'b11111111111111100111111110111100;
assign LUT_2[51658] = 32'b11111111111111110001111111011111;
assign LUT_2[51659] = 32'b11111111111111101110110111111000;
assign LUT_2[51660] = 32'b11111111111111100111100100001011;
assign LUT_2[51661] = 32'b11111111111111100100011100100100;
assign LUT_2[51662] = 32'b11111111111111101110011101000111;
assign LUT_2[51663] = 32'b11111111111111101011010101100000;
assign LUT_2[51664] = 32'b11111111111111101010111001010000;
assign LUT_2[51665] = 32'b11111111111111100111110001101001;
assign LUT_2[51666] = 32'b11111111111111110001110010001100;
assign LUT_2[51667] = 32'b11111111111111101110101010100101;
assign LUT_2[51668] = 32'b11111111111111100111010110111000;
assign LUT_2[51669] = 32'b11111111111111100100001111010001;
assign LUT_2[51670] = 32'b11111111111111101110001111110100;
assign LUT_2[51671] = 32'b11111111111111101011001000001101;
assign LUT_2[51672] = 32'b11111111111111100101101010101101;
assign LUT_2[51673] = 32'b11111111111111100010100011000110;
assign LUT_2[51674] = 32'b11111111111111101100100011101001;
assign LUT_2[51675] = 32'b11111111111111101001011100000010;
assign LUT_2[51676] = 32'b11111111111111100010001000010101;
assign LUT_2[51677] = 32'b11111111111111011111000000101110;
assign LUT_2[51678] = 32'b11111111111111101001000001010001;
assign LUT_2[51679] = 32'b11111111111111100101111001101010;
assign LUT_2[51680] = 32'b11111111111111110000110000101111;
assign LUT_2[51681] = 32'b11111111111111101101101001001000;
assign LUT_2[51682] = 32'b11111111111111110111101001101011;
assign LUT_2[51683] = 32'b11111111111111110100100010000100;
assign LUT_2[51684] = 32'b11111111111111101101001110010111;
assign LUT_2[51685] = 32'b11111111111111101010000110110000;
assign LUT_2[51686] = 32'b11111111111111110100000111010011;
assign LUT_2[51687] = 32'b11111111111111110000111111101100;
assign LUT_2[51688] = 32'b11111111111111101011100010001100;
assign LUT_2[51689] = 32'b11111111111111101000011010100101;
assign LUT_2[51690] = 32'b11111111111111110010011011001000;
assign LUT_2[51691] = 32'b11111111111111101111010011100001;
assign LUT_2[51692] = 32'b11111111111111100111111111110100;
assign LUT_2[51693] = 32'b11111111111111100100111000001101;
assign LUT_2[51694] = 32'b11111111111111101110111000110000;
assign LUT_2[51695] = 32'b11111111111111101011110001001001;
assign LUT_2[51696] = 32'b11111111111111101011010100111001;
assign LUT_2[51697] = 32'b11111111111111101000001101010010;
assign LUT_2[51698] = 32'b11111111111111110010001101110101;
assign LUT_2[51699] = 32'b11111111111111101111000110001110;
assign LUT_2[51700] = 32'b11111111111111100111110010100001;
assign LUT_2[51701] = 32'b11111111111111100100101010111010;
assign LUT_2[51702] = 32'b11111111111111101110101011011101;
assign LUT_2[51703] = 32'b11111111111111101011100011110110;
assign LUT_2[51704] = 32'b11111111111111100110000110010110;
assign LUT_2[51705] = 32'b11111111111111100010111110101111;
assign LUT_2[51706] = 32'b11111111111111101100111111010010;
assign LUT_2[51707] = 32'b11111111111111101001110111101011;
assign LUT_2[51708] = 32'b11111111111111100010100011111110;
assign LUT_2[51709] = 32'b11111111111111011111011100010111;
assign LUT_2[51710] = 32'b11111111111111101001011100111010;
assign LUT_2[51711] = 32'b11111111111111100110010101010011;
assign LUT_2[51712] = 32'b11111111111111110100101011100000;
assign LUT_2[51713] = 32'b11111111111111110001100011111001;
assign LUT_2[51714] = 32'b11111111111111111011100100011100;
assign LUT_2[51715] = 32'b11111111111111111000011100110101;
assign LUT_2[51716] = 32'b11111111111111110001001001001000;
assign LUT_2[51717] = 32'b11111111111111101110000001100001;
assign LUT_2[51718] = 32'b11111111111111111000000010000100;
assign LUT_2[51719] = 32'b11111111111111110100111010011101;
assign LUT_2[51720] = 32'b11111111111111101111011100111101;
assign LUT_2[51721] = 32'b11111111111111101100010101010110;
assign LUT_2[51722] = 32'b11111111111111110110010101111001;
assign LUT_2[51723] = 32'b11111111111111110011001110010010;
assign LUT_2[51724] = 32'b11111111111111101011111010100101;
assign LUT_2[51725] = 32'b11111111111111101000110010111110;
assign LUT_2[51726] = 32'b11111111111111110010110011100001;
assign LUT_2[51727] = 32'b11111111111111101111101011111010;
assign LUT_2[51728] = 32'b11111111111111101111001111101010;
assign LUT_2[51729] = 32'b11111111111111101100001000000011;
assign LUT_2[51730] = 32'b11111111111111110110001000100110;
assign LUT_2[51731] = 32'b11111111111111110011000000111111;
assign LUT_2[51732] = 32'b11111111111111101011101101010010;
assign LUT_2[51733] = 32'b11111111111111101000100101101011;
assign LUT_2[51734] = 32'b11111111111111110010100110001110;
assign LUT_2[51735] = 32'b11111111111111101111011110100111;
assign LUT_2[51736] = 32'b11111111111111101010000001000111;
assign LUT_2[51737] = 32'b11111111111111100110111001100000;
assign LUT_2[51738] = 32'b11111111111111110000111010000011;
assign LUT_2[51739] = 32'b11111111111111101101110010011100;
assign LUT_2[51740] = 32'b11111111111111100110011110101111;
assign LUT_2[51741] = 32'b11111111111111100011010111001000;
assign LUT_2[51742] = 32'b11111111111111101101010111101011;
assign LUT_2[51743] = 32'b11111111111111101010010000000100;
assign LUT_2[51744] = 32'b11111111111111110101000111001001;
assign LUT_2[51745] = 32'b11111111111111110001111111100010;
assign LUT_2[51746] = 32'b11111111111111111100000000000101;
assign LUT_2[51747] = 32'b11111111111111111000111000011110;
assign LUT_2[51748] = 32'b11111111111111110001100100110001;
assign LUT_2[51749] = 32'b11111111111111101110011101001010;
assign LUT_2[51750] = 32'b11111111111111111000011101101101;
assign LUT_2[51751] = 32'b11111111111111110101010110000110;
assign LUT_2[51752] = 32'b11111111111111101111111000100110;
assign LUT_2[51753] = 32'b11111111111111101100110000111111;
assign LUT_2[51754] = 32'b11111111111111110110110001100010;
assign LUT_2[51755] = 32'b11111111111111110011101001111011;
assign LUT_2[51756] = 32'b11111111111111101100010110001110;
assign LUT_2[51757] = 32'b11111111111111101001001110100111;
assign LUT_2[51758] = 32'b11111111111111110011001111001010;
assign LUT_2[51759] = 32'b11111111111111110000000111100011;
assign LUT_2[51760] = 32'b11111111111111101111101011010011;
assign LUT_2[51761] = 32'b11111111111111101100100011101100;
assign LUT_2[51762] = 32'b11111111111111110110100100001111;
assign LUT_2[51763] = 32'b11111111111111110011011100101000;
assign LUT_2[51764] = 32'b11111111111111101100001000111011;
assign LUT_2[51765] = 32'b11111111111111101001000001010100;
assign LUT_2[51766] = 32'b11111111111111110011000001110111;
assign LUT_2[51767] = 32'b11111111111111101111111010010000;
assign LUT_2[51768] = 32'b11111111111111101010011100110000;
assign LUT_2[51769] = 32'b11111111111111100111010101001001;
assign LUT_2[51770] = 32'b11111111111111110001010101101100;
assign LUT_2[51771] = 32'b11111111111111101110001110000101;
assign LUT_2[51772] = 32'b11111111111111100110111010011000;
assign LUT_2[51773] = 32'b11111111111111100011110010110001;
assign LUT_2[51774] = 32'b11111111111111101101110011010100;
assign LUT_2[51775] = 32'b11111111111111101010101011101101;
assign LUT_2[51776] = 32'b11111111111111101100110100000011;
assign LUT_2[51777] = 32'b11111111111111101001101100011100;
assign LUT_2[51778] = 32'b11111111111111110011101100111111;
assign LUT_2[51779] = 32'b11111111111111110000100101011000;
assign LUT_2[51780] = 32'b11111111111111101001010001101011;
assign LUT_2[51781] = 32'b11111111111111100110001010000100;
assign LUT_2[51782] = 32'b11111111111111110000001010100111;
assign LUT_2[51783] = 32'b11111111111111101101000011000000;
assign LUT_2[51784] = 32'b11111111111111100111100101100000;
assign LUT_2[51785] = 32'b11111111111111100100011101111001;
assign LUT_2[51786] = 32'b11111111111111101110011110011100;
assign LUT_2[51787] = 32'b11111111111111101011010110110101;
assign LUT_2[51788] = 32'b11111111111111100100000011001000;
assign LUT_2[51789] = 32'b11111111111111100000111011100001;
assign LUT_2[51790] = 32'b11111111111111101010111100000100;
assign LUT_2[51791] = 32'b11111111111111100111110100011101;
assign LUT_2[51792] = 32'b11111111111111100111011000001101;
assign LUT_2[51793] = 32'b11111111111111100100010000100110;
assign LUT_2[51794] = 32'b11111111111111101110010001001001;
assign LUT_2[51795] = 32'b11111111111111101011001001100010;
assign LUT_2[51796] = 32'b11111111111111100011110101110101;
assign LUT_2[51797] = 32'b11111111111111100000101110001110;
assign LUT_2[51798] = 32'b11111111111111101010101110110001;
assign LUT_2[51799] = 32'b11111111111111100111100111001010;
assign LUT_2[51800] = 32'b11111111111111100010001001101010;
assign LUT_2[51801] = 32'b11111111111111011111000010000011;
assign LUT_2[51802] = 32'b11111111111111101001000010100110;
assign LUT_2[51803] = 32'b11111111111111100101111010111111;
assign LUT_2[51804] = 32'b11111111111111011110100111010010;
assign LUT_2[51805] = 32'b11111111111111011011011111101011;
assign LUT_2[51806] = 32'b11111111111111100101100000001110;
assign LUT_2[51807] = 32'b11111111111111100010011000100111;
assign LUT_2[51808] = 32'b11111111111111101101001111101100;
assign LUT_2[51809] = 32'b11111111111111101010001000000101;
assign LUT_2[51810] = 32'b11111111111111110100001000101000;
assign LUT_2[51811] = 32'b11111111111111110001000001000001;
assign LUT_2[51812] = 32'b11111111111111101001101101010100;
assign LUT_2[51813] = 32'b11111111111111100110100101101101;
assign LUT_2[51814] = 32'b11111111111111110000100110010000;
assign LUT_2[51815] = 32'b11111111111111101101011110101001;
assign LUT_2[51816] = 32'b11111111111111101000000001001001;
assign LUT_2[51817] = 32'b11111111111111100100111001100010;
assign LUT_2[51818] = 32'b11111111111111101110111010000101;
assign LUT_2[51819] = 32'b11111111111111101011110010011110;
assign LUT_2[51820] = 32'b11111111111111100100011110110001;
assign LUT_2[51821] = 32'b11111111111111100001010111001010;
assign LUT_2[51822] = 32'b11111111111111101011010111101101;
assign LUT_2[51823] = 32'b11111111111111101000010000000110;
assign LUT_2[51824] = 32'b11111111111111100111110011110110;
assign LUT_2[51825] = 32'b11111111111111100100101100001111;
assign LUT_2[51826] = 32'b11111111111111101110101100110010;
assign LUT_2[51827] = 32'b11111111111111101011100101001011;
assign LUT_2[51828] = 32'b11111111111111100100010001011110;
assign LUT_2[51829] = 32'b11111111111111100001001001110111;
assign LUT_2[51830] = 32'b11111111111111101011001010011010;
assign LUT_2[51831] = 32'b11111111111111101000000010110011;
assign LUT_2[51832] = 32'b11111111111111100010100101010011;
assign LUT_2[51833] = 32'b11111111111111011111011101101100;
assign LUT_2[51834] = 32'b11111111111111101001011110001111;
assign LUT_2[51835] = 32'b11111111111111100110010110101000;
assign LUT_2[51836] = 32'b11111111111111011111000010111011;
assign LUT_2[51837] = 32'b11111111111111011011111011010100;
assign LUT_2[51838] = 32'b11111111111111100101111011110111;
assign LUT_2[51839] = 32'b11111111111111100010110100010000;
assign LUT_2[51840] = 32'b11111111111111111000111111101111;
assign LUT_2[51841] = 32'b11111111111111110101111000001000;
assign LUT_2[51842] = 32'b11111111111111111111111000101011;
assign LUT_2[51843] = 32'b11111111111111111100110001000100;
assign LUT_2[51844] = 32'b11111111111111110101011101010111;
assign LUT_2[51845] = 32'b11111111111111110010010101110000;
assign LUT_2[51846] = 32'b11111111111111111100010110010011;
assign LUT_2[51847] = 32'b11111111111111111001001110101100;
assign LUT_2[51848] = 32'b11111111111111110011110001001100;
assign LUT_2[51849] = 32'b11111111111111110000101001100101;
assign LUT_2[51850] = 32'b11111111111111111010101010001000;
assign LUT_2[51851] = 32'b11111111111111110111100010100001;
assign LUT_2[51852] = 32'b11111111111111110000001110110100;
assign LUT_2[51853] = 32'b11111111111111101101000111001101;
assign LUT_2[51854] = 32'b11111111111111110111000111110000;
assign LUT_2[51855] = 32'b11111111111111110100000000001001;
assign LUT_2[51856] = 32'b11111111111111110011100011111001;
assign LUT_2[51857] = 32'b11111111111111110000011100010010;
assign LUT_2[51858] = 32'b11111111111111111010011100110101;
assign LUT_2[51859] = 32'b11111111111111110111010101001110;
assign LUT_2[51860] = 32'b11111111111111110000000001100001;
assign LUT_2[51861] = 32'b11111111111111101100111001111010;
assign LUT_2[51862] = 32'b11111111111111110110111010011101;
assign LUT_2[51863] = 32'b11111111111111110011110010110110;
assign LUT_2[51864] = 32'b11111111111111101110010101010110;
assign LUT_2[51865] = 32'b11111111111111101011001101101111;
assign LUT_2[51866] = 32'b11111111111111110101001110010010;
assign LUT_2[51867] = 32'b11111111111111110010000110101011;
assign LUT_2[51868] = 32'b11111111111111101010110010111110;
assign LUT_2[51869] = 32'b11111111111111100111101011010111;
assign LUT_2[51870] = 32'b11111111111111110001101011111010;
assign LUT_2[51871] = 32'b11111111111111101110100100010011;
assign LUT_2[51872] = 32'b11111111111111111001011011011000;
assign LUT_2[51873] = 32'b11111111111111110110010011110001;
assign LUT_2[51874] = 32'b00000000000000000000010100010100;
assign LUT_2[51875] = 32'b11111111111111111101001100101101;
assign LUT_2[51876] = 32'b11111111111111110101111001000000;
assign LUT_2[51877] = 32'b11111111111111110010110001011001;
assign LUT_2[51878] = 32'b11111111111111111100110001111100;
assign LUT_2[51879] = 32'b11111111111111111001101010010101;
assign LUT_2[51880] = 32'b11111111111111110100001100110101;
assign LUT_2[51881] = 32'b11111111111111110001000101001110;
assign LUT_2[51882] = 32'b11111111111111111011000101110001;
assign LUT_2[51883] = 32'b11111111111111110111111110001010;
assign LUT_2[51884] = 32'b11111111111111110000101010011101;
assign LUT_2[51885] = 32'b11111111111111101101100010110110;
assign LUT_2[51886] = 32'b11111111111111110111100011011001;
assign LUT_2[51887] = 32'b11111111111111110100011011110010;
assign LUT_2[51888] = 32'b11111111111111110011111111100010;
assign LUT_2[51889] = 32'b11111111111111110000110111111011;
assign LUT_2[51890] = 32'b11111111111111111010111000011110;
assign LUT_2[51891] = 32'b11111111111111110111110000110111;
assign LUT_2[51892] = 32'b11111111111111110000011101001010;
assign LUT_2[51893] = 32'b11111111111111101101010101100011;
assign LUT_2[51894] = 32'b11111111111111110111010110000110;
assign LUT_2[51895] = 32'b11111111111111110100001110011111;
assign LUT_2[51896] = 32'b11111111111111101110110000111111;
assign LUT_2[51897] = 32'b11111111111111101011101001011000;
assign LUT_2[51898] = 32'b11111111111111110101101001111011;
assign LUT_2[51899] = 32'b11111111111111110010100010010100;
assign LUT_2[51900] = 32'b11111111111111101011001110100111;
assign LUT_2[51901] = 32'b11111111111111101000000111000000;
assign LUT_2[51902] = 32'b11111111111111110010000111100011;
assign LUT_2[51903] = 32'b11111111111111101110111111111100;
assign LUT_2[51904] = 32'b11111111111111110001001000010010;
assign LUT_2[51905] = 32'b11111111111111101110000000101011;
assign LUT_2[51906] = 32'b11111111111111111000000001001110;
assign LUT_2[51907] = 32'b11111111111111110100111001100111;
assign LUT_2[51908] = 32'b11111111111111101101100101111010;
assign LUT_2[51909] = 32'b11111111111111101010011110010011;
assign LUT_2[51910] = 32'b11111111111111110100011110110110;
assign LUT_2[51911] = 32'b11111111111111110001010111001111;
assign LUT_2[51912] = 32'b11111111111111101011111001101111;
assign LUT_2[51913] = 32'b11111111111111101000110010001000;
assign LUT_2[51914] = 32'b11111111111111110010110010101011;
assign LUT_2[51915] = 32'b11111111111111101111101011000100;
assign LUT_2[51916] = 32'b11111111111111101000010111010111;
assign LUT_2[51917] = 32'b11111111111111100101001111110000;
assign LUT_2[51918] = 32'b11111111111111101111010000010011;
assign LUT_2[51919] = 32'b11111111111111101100001000101100;
assign LUT_2[51920] = 32'b11111111111111101011101100011100;
assign LUT_2[51921] = 32'b11111111111111101000100100110101;
assign LUT_2[51922] = 32'b11111111111111110010100101011000;
assign LUT_2[51923] = 32'b11111111111111101111011101110001;
assign LUT_2[51924] = 32'b11111111111111101000001010000100;
assign LUT_2[51925] = 32'b11111111111111100101000010011101;
assign LUT_2[51926] = 32'b11111111111111101111000011000000;
assign LUT_2[51927] = 32'b11111111111111101011111011011001;
assign LUT_2[51928] = 32'b11111111111111100110011101111001;
assign LUT_2[51929] = 32'b11111111111111100011010110010010;
assign LUT_2[51930] = 32'b11111111111111101101010110110101;
assign LUT_2[51931] = 32'b11111111111111101010001111001110;
assign LUT_2[51932] = 32'b11111111111111100010111011100001;
assign LUT_2[51933] = 32'b11111111111111011111110011111010;
assign LUT_2[51934] = 32'b11111111111111101001110100011101;
assign LUT_2[51935] = 32'b11111111111111100110101100110110;
assign LUT_2[51936] = 32'b11111111111111110001100011111011;
assign LUT_2[51937] = 32'b11111111111111101110011100010100;
assign LUT_2[51938] = 32'b11111111111111111000011100110111;
assign LUT_2[51939] = 32'b11111111111111110101010101010000;
assign LUT_2[51940] = 32'b11111111111111101110000001100011;
assign LUT_2[51941] = 32'b11111111111111101010111001111100;
assign LUT_2[51942] = 32'b11111111111111110100111010011111;
assign LUT_2[51943] = 32'b11111111111111110001110010111000;
assign LUT_2[51944] = 32'b11111111111111101100010101011000;
assign LUT_2[51945] = 32'b11111111111111101001001101110001;
assign LUT_2[51946] = 32'b11111111111111110011001110010100;
assign LUT_2[51947] = 32'b11111111111111110000000110101101;
assign LUT_2[51948] = 32'b11111111111111101000110011000000;
assign LUT_2[51949] = 32'b11111111111111100101101011011001;
assign LUT_2[51950] = 32'b11111111111111101111101011111100;
assign LUT_2[51951] = 32'b11111111111111101100100100010101;
assign LUT_2[51952] = 32'b11111111111111101100001000000101;
assign LUT_2[51953] = 32'b11111111111111101001000000011110;
assign LUT_2[51954] = 32'b11111111111111110011000001000001;
assign LUT_2[51955] = 32'b11111111111111101111111001011010;
assign LUT_2[51956] = 32'b11111111111111101000100101101101;
assign LUT_2[51957] = 32'b11111111111111100101011110000110;
assign LUT_2[51958] = 32'b11111111111111101111011110101001;
assign LUT_2[51959] = 32'b11111111111111101100010111000010;
assign LUT_2[51960] = 32'b11111111111111100110111001100010;
assign LUT_2[51961] = 32'b11111111111111100011110001111011;
assign LUT_2[51962] = 32'b11111111111111101101110010011110;
assign LUT_2[51963] = 32'b11111111111111101010101010110111;
assign LUT_2[51964] = 32'b11111111111111100011010111001010;
assign LUT_2[51965] = 32'b11111111111111100000001111100011;
assign LUT_2[51966] = 32'b11111111111111101010010000000110;
assign LUT_2[51967] = 32'b11111111111111100111001000011111;
assign LUT_2[51968] = 32'b11111111111111111000101010000110;
assign LUT_2[51969] = 32'b11111111111111110101100010011111;
assign LUT_2[51970] = 32'b11111111111111111111100011000010;
assign LUT_2[51971] = 32'b11111111111111111100011011011011;
assign LUT_2[51972] = 32'b11111111111111110101000111101110;
assign LUT_2[51973] = 32'b11111111111111110010000000000111;
assign LUT_2[51974] = 32'b11111111111111111100000000101010;
assign LUT_2[51975] = 32'b11111111111111111000111001000011;
assign LUT_2[51976] = 32'b11111111111111110011011011100011;
assign LUT_2[51977] = 32'b11111111111111110000010011111100;
assign LUT_2[51978] = 32'b11111111111111111010010100011111;
assign LUT_2[51979] = 32'b11111111111111110111001100111000;
assign LUT_2[51980] = 32'b11111111111111101111111001001011;
assign LUT_2[51981] = 32'b11111111111111101100110001100100;
assign LUT_2[51982] = 32'b11111111111111110110110010000111;
assign LUT_2[51983] = 32'b11111111111111110011101010100000;
assign LUT_2[51984] = 32'b11111111111111110011001110010000;
assign LUT_2[51985] = 32'b11111111111111110000000110101001;
assign LUT_2[51986] = 32'b11111111111111111010000111001100;
assign LUT_2[51987] = 32'b11111111111111110110111111100101;
assign LUT_2[51988] = 32'b11111111111111101111101011111000;
assign LUT_2[51989] = 32'b11111111111111101100100100010001;
assign LUT_2[51990] = 32'b11111111111111110110100100110100;
assign LUT_2[51991] = 32'b11111111111111110011011101001101;
assign LUT_2[51992] = 32'b11111111111111101101111111101101;
assign LUT_2[51993] = 32'b11111111111111101010111000000110;
assign LUT_2[51994] = 32'b11111111111111110100111000101001;
assign LUT_2[51995] = 32'b11111111111111110001110001000010;
assign LUT_2[51996] = 32'b11111111111111101010011101010101;
assign LUT_2[51997] = 32'b11111111111111100111010101101110;
assign LUT_2[51998] = 32'b11111111111111110001010110010001;
assign LUT_2[51999] = 32'b11111111111111101110001110101010;
assign LUT_2[52000] = 32'b11111111111111111001000101101111;
assign LUT_2[52001] = 32'b11111111111111110101111110001000;
assign LUT_2[52002] = 32'b11111111111111111111111110101011;
assign LUT_2[52003] = 32'b11111111111111111100110111000100;
assign LUT_2[52004] = 32'b11111111111111110101100011010111;
assign LUT_2[52005] = 32'b11111111111111110010011011110000;
assign LUT_2[52006] = 32'b11111111111111111100011100010011;
assign LUT_2[52007] = 32'b11111111111111111001010100101100;
assign LUT_2[52008] = 32'b11111111111111110011110111001100;
assign LUT_2[52009] = 32'b11111111111111110000101111100101;
assign LUT_2[52010] = 32'b11111111111111111010110000001000;
assign LUT_2[52011] = 32'b11111111111111110111101000100001;
assign LUT_2[52012] = 32'b11111111111111110000010100110100;
assign LUT_2[52013] = 32'b11111111111111101101001101001101;
assign LUT_2[52014] = 32'b11111111111111110111001101110000;
assign LUT_2[52015] = 32'b11111111111111110100000110001001;
assign LUT_2[52016] = 32'b11111111111111110011101001111001;
assign LUT_2[52017] = 32'b11111111111111110000100010010010;
assign LUT_2[52018] = 32'b11111111111111111010100010110101;
assign LUT_2[52019] = 32'b11111111111111110111011011001110;
assign LUT_2[52020] = 32'b11111111111111110000000111100001;
assign LUT_2[52021] = 32'b11111111111111101100111111111010;
assign LUT_2[52022] = 32'b11111111111111110111000000011101;
assign LUT_2[52023] = 32'b11111111111111110011111000110110;
assign LUT_2[52024] = 32'b11111111111111101110011011010110;
assign LUT_2[52025] = 32'b11111111111111101011010011101111;
assign LUT_2[52026] = 32'b11111111111111110101010100010010;
assign LUT_2[52027] = 32'b11111111111111110010001100101011;
assign LUT_2[52028] = 32'b11111111111111101010111000111110;
assign LUT_2[52029] = 32'b11111111111111100111110001010111;
assign LUT_2[52030] = 32'b11111111111111110001110001111010;
assign LUT_2[52031] = 32'b11111111111111101110101010010011;
assign LUT_2[52032] = 32'b11111111111111110000110010101001;
assign LUT_2[52033] = 32'b11111111111111101101101011000010;
assign LUT_2[52034] = 32'b11111111111111110111101011100101;
assign LUT_2[52035] = 32'b11111111111111110100100011111110;
assign LUT_2[52036] = 32'b11111111111111101101010000010001;
assign LUT_2[52037] = 32'b11111111111111101010001000101010;
assign LUT_2[52038] = 32'b11111111111111110100001001001101;
assign LUT_2[52039] = 32'b11111111111111110001000001100110;
assign LUT_2[52040] = 32'b11111111111111101011100100000110;
assign LUT_2[52041] = 32'b11111111111111101000011100011111;
assign LUT_2[52042] = 32'b11111111111111110010011101000010;
assign LUT_2[52043] = 32'b11111111111111101111010101011011;
assign LUT_2[52044] = 32'b11111111111111101000000001101110;
assign LUT_2[52045] = 32'b11111111111111100100111010000111;
assign LUT_2[52046] = 32'b11111111111111101110111010101010;
assign LUT_2[52047] = 32'b11111111111111101011110011000011;
assign LUT_2[52048] = 32'b11111111111111101011010110110011;
assign LUT_2[52049] = 32'b11111111111111101000001111001100;
assign LUT_2[52050] = 32'b11111111111111110010001111101111;
assign LUT_2[52051] = 32'b11111111111111101111001000001000;
assign LUT_2[52052] = 32'b11111111111111100111110100011011;
assign LUT_2[52053] = 32'b11111111111111100100101100110100;
assign LUT_2[52054] = 32'b11111111111111101110101101010111;
assign LUT_2[52055] = 32'b11111111111111101011100101110000;
assign LUT_2[52056] = 32'b11111111111111100110001000010000;
assign LUT_2[52057] = 32'b11111111111111100011000000101001;
assign LUT_2[52058] = 32'b11111111111111101101000001001100;
assign LUT_2[52059] = 32'b11111111111111101001111001100101;
assign LUT_2[52060] = 32'b11111111111111100010100101111000;
assign LUT_2[52061] = 32'b11111111111111011111011110010001;
assign LUT_2[52062] = 32'b11111111111111101001011110110100;
assign LUT_2[52063] = 32'b11111111111111100110010111001101;
assign LUT_2[52064] = 32'b11111111111111110001001110010010;
assign LUT_2[52065] = 32'b11111111111111101110000110101011;
assign LUT_2[52066] = 32'b11111111111111111000000111001110;
assign LUT_2[52067] = 32'b11111111111111110100111111100111;
assign LUT_2[52068] = 32'b11111111111111101101101011111010;
assign LUT_2[52069] = 32'b11111111111111101010100100010011;
assign LUT_2[52070] = 32'b11111111111111110100100100110110;
assign LUT_2[52071] = 32'b11111111111111110001011101001111;
assign LUT_2[52072] = 32'b11111111111111101011111111101111;
assign LUT_2[52073] = 32'b11111111111111101000111000001000;
assign LUT_2[52074] = 32'b11111111111111110010111000101011;
assign LUT_2[52075] = 32'b11111111111111101111110001000100;
assign LUT_2[52076] = 32'b11111111111111101000011101010111;
assign LUT_2[52077] = 32'b11111111111111100101010101110000;
assign LUT_2[52078] = 32'b11111111111111101111010110010011;
assign LUT_2[52079] = 32'b11111111111111101100001110101100;
assign LUT_2[52080] = 32'b11111111111111101011110010011100;
assign LUT_2[52081] = 32'b11111111111111101000101010110101;
assign LUT_2[52082] = 32'b11111111111111110010101011011000;
assign LUT_2[52083] = 32'b11111111111111101111100011110001;
assign LUT_2[52084] = 32'b11111111111111101000010000000100;
assign LUT_2[52085] = 32'b11111111111111100101001000011101;
assign LUT_2[52086] = 32'b11111111111111101111001001000000;
assign LUT_2[52087] = 32'b11111111111111101100000001011001;
assign LUT_2[52088] = 32'b11111111111111100110100011111001;
assign LUT_2[52089] = 32'b11111111111111100011011100010010;
assign LUT_2[52090] = 32'b11111111111111101101011100110101;
assign LUT_2[52091] = 32'b11111111111111101010010101001110;
assign LUT_2[52092] = 32'b11111111111111100011000001100001;
assign LUT_2[52093] = 32'b11111111111111011111111001111010;
assign LUT_2[52094] = 32'b11111111111111101001111010011101;
assign LUT_2[52095] = 32'b11111111111111100110110010110110;
assign LUT_2[52096] = 32'b11111111111111111100111110010101;
assign LUT_2[52097] = 32'b11111111111111111001110110101110;
assign LUT_2[52098] = 32'b00000000000000000011110111010001;
assign LUT_2[52099] = 32'b00000000000000000000101111101010;
assign LUT_2[52100] = 32'b11111111111111111001011011111101;
assign LUT_2[52101] = 32'b11111111111111110110010100010110;
assign LUT_2[52102] = 32'b00000000000000000000010100111001;
assign LUT_2[52103] = 32'b11111111111111111101001101010010;
assign LUT_2[52104] = 32'b11111111111111110111101111110010;
assign LUT_2[52105] = 32'b11111111111111110100101000001011;
assign LUT_2[52106] = 32'b11111111111111111110101000101110;
assign LUT_2[52107] = 32'b11111111111111111011100001000111;
assign LUT_2[52108] = 32'b11111111111111110100001101011010;
assign LUT_2[52109] = 32'b11111111111111110001000101110011;
assign LUT_2[52110] = 32'b11111111111111111011000110010110;
assign LUT_2[52111] = 32'b11111111111111110111111110101111;
assign LUT_2[52112] = 32'b11111111111111110111100010011111;
assign LUT_2[52113] = 32'b11111111111111110100011010111000;
assign LUT_2[52114] = 32'b11111111111111111110011011011011;
assign LUT_2[52115] = 32'b11111111111111111011010011110100;
assign LUT_2[52116] = 32'b11111111111111110100000000000111;
assign LUT_2[52117] = 32'b11111111111111110000111000100000;
assign LUT_2[52118] = 32'b11111111111111111010111001000011;
assign LUT_2[52119] = 32'b11111111111111110111110001011100;
assign LUT_2[52120] = 32'b11111111111111110010010011111100;
assign LUT_2[52121] = 32'b11111111111111101111001100010101;
assign LUT_2[52122] = 32'b11111111111111111001001100111000;
assign LUT_2[52123] = 32'b11111111111111110110000101010001;
assign LUT_2[52124] = 32'b11111111111111101110110001100100;
assign LUT_2[52125] = 32'b11111111111111101011101001111101;
assign LUT_2[52126] = 32'b11111111111111110101101010100000;
assign LUT_2[52127] = 32'b11111111111111110010100010111001;
assign LUT_2[52128] = 32'b11111111111111111101011001111110;
assign LUT_2[52129] = 32'b11111111111111111010010010010111;
assign LUT_2[52130] = 32'b00000000000000000100010010111010;
assign LUT_2[52131] = 32'b00000000000000000001001011010011;
assign LUT_2[52132] = 32'b11111111111111111001110111100110;
assign LUT_2[52133] = 32'b11111111111111110110101111111111;
assign LUT_2[52134] = 32'b00000000000000000000110000100010;
assign LUT_2[52135] = 32'b11111111111111111101101000111011;
assign LUT_2[52136] = 32'b11111111111111111000001011011011;
assign LUT_2[52137] = 32'b11111111111111110101000011110100;
assign LUT_2[52138] = 32'b11111111111111111111000100010111;
assign LUT_2[52139] = 32'b11111111111111111011111100110000;
assign LUT_2[52140] = 32'b11111111111111110100101001000011;
assign LUT_2[52141] = 32'b11111111111111110001100001011100;
assign LUT_2[52142] = 32'b11111111111111111011100001111111;
assign LUT_2[52143] = 32'b11111111111111111000011010011000;
assign LUT_2[52144] = 32'b11111111111111110111111110001000;
assign LUT_2[52145] = 32'b11111111111111110100110110100001;
assign LUT_2[52146] = 32'b11111111111111111110110111000100;
assign LUT_2[52147] = 32'b11111111111111111011101111011101;
assign LUT_2[52148] = 32'b11111111111111110100011011110000;
assign LUT_2[52149] = 32'b11111111111111110001010100001001;
assign LUT_2[52150] = 32'b11111111111111111011010100101100;
assign LUT_2[52151] = 32'b11111111111111111000001101000101;
assign LUT_2[52152] = 32'b11111111111111110010101111100101;
assign LUT_2[52153] = 32'b11111111111111101111100111111110;
assign LUT_2[52154] = 32'b11111111111111111001101000100001;
assign LUT_2[52155] = 32'b11111111111111110110100000111010;
assign LUT_2[52156] = 32'b11111111111111101111001101001101;
assign LUT_2[52157] = 32'b11111111111111101100000101100110;
assign LUT_2[52158] = 32'b11111111111111110110000110001001;
assign LUT_2[52159] = 32'b11111111111111110010111110100010;
assign LUT_2[52160] = 32'b11111111111111110101000110111000;
assign LUT_2[52161] = 32'b11111111111111110001111111010001;
assign LUT_2[52162] = 32'b11111111111111111011111111110100;
assign LUT_2[52163] = 32'b11111111111111111000111000001101;
assign LUT_2[52164] = 32'b11111111111111110001100100100000;
assign LUT_2[52165] = 32'b11111111111111101110011100111001;
assign LUT_2[52166] = 32'b11111111111111111000011101011100;
assign LUT_2[52167] = 32'b11111111111111110101010101110101;
assign LUT_2[52168] = 32'b11111111111111101111111000010101;
assign LUT_2[52169] = 32'b11111111111111101100110000101110;
assign LUT_2[52170] = 32'b11111111111111110110110001010001;
assign LUT_2[52171] = 32'b11111111111111110011101001101010;
assign LUT_2[52172] = 32'b11111111111111101100010101111101;
assign LUT_2[52173] = 32'b11111111111111101001001110010110;
assign LUT_2[52174] = 32'b11111111111111110011001110111001;
assign LUT_2[52175] = 32'b11111111111111110000000111010010;
assign LUT_2[52176] = 32'b11111111111111101111101011000010;
assign LUT_2[52177] = 32'b11111111111111101100100011011011;
assign LUT_2[52178] = 32'b11111111111111110110100011111110;
assign LUT_2[52179] = 32'b11111111111111110011011100010111;
assign LUT_2[52180] = 32'b11111111111111101100001000101010;
assign LUT_2[52181] = 32'b11111111111111101001000001000011;
assign LUT_2[52182] = 32'b11111111111111110011000001100110;
assign LUT_2[52183] = 32'b11111111111111101111111001111111;
assign LUT_2[52184] = 32'b11111111111111101010011100011111;
assign LUT_2[52185] = 32'b11111111111111100111010100111000;
assign LUT_2[52186] = 32'b11111111111111110001010101011011;
assign LUT_2[52187] = 32'b11111111111111101110001101110100;
assign LUT_2[52188] = 32'b11111111111111100110111010000111;
assign LUT_2[52189] = 32'b11111111111111100011110010100000;
assign LUT_2[52190] = 32'b11111111111111101101110011000011;
assign LUT_2[52191] = 32'b11111111111111101010101011011100;
assign LUT_2[52192] = 32'b11111111111111110101100010100001;
assign LUT_2[52193] = 32'b11111111111111110010011010111010;
assign LUT_2[52194] = 32'b11111111111111111100011011011101;
assign LUT_2[52195] = 32'b11111111111111111001010011110110;
assign LUT_2[52196] = 32'b11111111111111110010000000001001;
assign LUT_2[52197] = 32'b11111111111111101110111000100010;
assign LUT_2[52198] = 32'b11111111111111111000111001000101;
assign LUT_2[52199] = 32'b11111111111111110101110001011110;
assign LUT_2[52200] = 32'b11111111111111110000010011111110;
assign LUT_2[52201] = 32'b11111111111111101101001100010111;
assign LUT_2[52202] = 32'b11111111111111110111001100111010;
assign LUT_2[52203] = 32'b11111111111111110100000101010011;
assign LUT_2[52204] = 32'b11111111111111101100110001100110;
assign LUT_2[52205] = 32'b11111111111111101001101001111111;
assign LUT_2[52206] = 32'b11111111111111110011101010100010;
assign LUT_2[52207] = 32'b11111111111111110000100010111011;
assign LUT_2[52208] = 32'b11111111111111110000000110101011;
assign LUT_2[52209] = 32'b11111111111111101100111111000100;
assign LUT_2[52210] = 32'b11111111111111110110111111100111;
assign LUT_2[52211] = 32'b11111111111111110011111000000000;
assign LUT_2[52212] = 32'b11111111111111101100100100010011;
assign LUT_2[52213] = 32'b11111111111111101001011100101100;
assign LUT_2[52214] = 32'b11111111111111110011011101001111;
assign LUT_2[52215] = 32'b11111111111111110000010101101000;
assign LUT_2[52216] = 32'b11111111111111101010111000001000;
assign LUT_2[52217] = 32'b11111111111111100111110000100001;
assign LUT_2[52218] = 32'b11111111111111110001110001000100;
assign LUT_2[52219] = 32'b11111111111111101110101001011101;
assign LUT_2[52220] = 32'b11111111111111100111010101110000;
assign LUT_2[52221] = 32'b11111111111111100100001110001001;
assign LUT_2[52222] = 32'b11111111111111101110001110101100;
assign LUT_2[52223] = 32'b11111111111111101011000111000101;
assign LUT_2[52224] = 32'b11111111111111110110100101110011;
assign LUT_2[52225] = 32'b11111111111111110011011110001100;
assign LUT_2[52226] = 32'b11111111111111111101011110101111;
assign LUT_2[52227] = 32'b11111111111111111010010111001000;
assign LUT_2[52228] = 32'b11111111111111110011000011011011;
assign LUT_2[52229] = 32'b11111111111111101111111011110100;
assign LUT_2[52230] = 32'b11111111111111111001111100010111;
assign LUT_2[52231] = 32'b11111111111111110110110100110000;
assign LUT_2[52232] = 32'b11111111111111110001010111010000;
assign LUT_2[52233] = 32'b11111111111111101110001111101001;
assign LUT_2[52234] = 32'b11111111111111111000010000001100;
assign LUT_2[52235] = 32'b11111111111111110101001000100101;
assign LUT_2[52236] = 32'b11111111111111101101110100111000;
assign LUT_2[52237] = 32'b11111111111111101010101101010001;
assign LUT_2[52238] = 32'b11111111111111110100101101110100;
assign LUT_2[52239] = 32'b11111111111111110001100110001101;
assign LUT_2[52240] = 32'b11111111111111110001001001111101;
assign LUT_2[52241] = 32'b11111111111111101110000010010110;
assign LUT_2[52242] = 32'b11111111111111111000000010111001;
assign LUT_2[52243] = 32'b11111111111111110100111011010010;
assign LUT_2[52244] = 32'b11111111111111101101100111100101;
assign LUT_2[52245] = 32'b11111111111111101010011111111110;
assign LUT_2[52246] = 32'b11111111111111110100100000100001;
assign LUT_2[52247] = 32'b11111111111111110001011000111010;
assign LUT_2[52248] = 32'b11111111111111101011111011011010;
assign LUT_2[52249] = 32'b11111111111111101000110011110011;
assign LUT_2[52250] = 32'b11111111111111110010110100010110;
assign LUT_2[52251] = 32'b11111111111111101111101100101111;
assign LUT_2[52252] = 32'b11111111111111101000011001000010;
assign LUT_2[52253] = 32'b11111111111111100101010001011011;
assign LUT_2[52254] = 32'b11111111111111101111010001111110;
assign LUT_2[52255] = 32'b11111111111111101100001010010111;
assign LUT_2[52256] = 32'b11111111111111110111000001011100;
assign LUT_2[52257] = 32'b11111111111111110011111001110101;
assign LUT_2[52258] = 32'b11111111111111111101111010011000;
assign LUT_2[52259] = 32'b11111111111111111010110010110001;
assign LUT_2[52260] = 32'b11111111111111110011011111000100;
assign LUT_2[52261] = 32'b11111111111111110000010111011101;
assign LUT_2[52262] = 32'b11111111111111111010011000000000;
assign LUT_2[52263] = 32'b11111111111111110111010000011001;
assign LUT_2[52264] = 32'b11111111111111110001110010111001;
assign LUT_2[52265] = 32'b11111111111111101110101011010010;
assign LUT_2[52266] = 32'b11111111111111111000101011110101;
assign LUT_2[52267] = 32'b11111111111111110101100100001110;
assign LUT_2[52268] = 32'b11111111111111101110010000100001;
assign LUT_2[52269] = 32'b11111111111111101011001000111010;
assign LUT_2[52270] = 32'b11111111111111110101001001011101;
assign LUT_2[52271] = 32'b11111111111111110010000001110110;
assign LUT_2[52272] = 32'b11111111111111110001100101100110;
assign LUT_2[52273] = 32'b11111111111111101110011101111111;
assign LUT_2[52274] = 32'b11111111111111111000011110100010;
assign LUT_2[52275] = 32'b11111111111111110101010110111011;
assign LUT_2[52276] = 32'b11111111111111101110000011001110;
assign LUT_2[52277] = 32'b11111111111111101010111011100111;
assign LUT_2[52278] = 32'b11111111111111110100111100001010;
assign LUT_2[52279] = 32'b11111111111111110001110100100011;
assign LUT_2[52280] = 32'b11111111111111101100010111000011;
assign LUT_2[52281] = 32'b11111111111111101001001111011100;
assign LUT_2[52282] = 32'b11111111111111110011001111111111;
assign LUT_2[52283] = 32'b11111111111111110000001000011000;
assign LUT_2[52284] = 32'b11111111111111101000110100101011;
assign LUT_2[52285] = 32'b11111111111111100101101101000100;
assign LUT_2[52286] = 32'b11111111111111101111101101100111;
assign LUT_2[52287] = 32'b11111111111111101100100110000000;
assign LUT_2[52288] = 32'b11111111111111101110101110010110;
assign LUT_2[52289] = 32'b11111111111111101011100110101111;
assign LUT_2[52290] = 32'b11111111111111110101100111010010;
assign LUT_2[52291] = 32'b11111111111111110010011111101011;
assign LUT_2[52292] = 32'b11111111111111101011001011111110;
assign LUT_2[52293] = 32'b11111111111111101000000100010111;
assign LUT_2[52294] = 32'b11111111111111110010000100111010;
assign LUT_2[52295] = 32'b11111111111111101110111101010011;
assign LUT_2[52296] = 32'b11111111111111101001011111110011;
assign LUT_2[52297] = 32'b11111111111111100110011000001100;
assign LUT_2[52298] = 32'b11111111111111110000011000101111;
assign LUT_2[52299] = 32'b11111111111111101101010001001000;
assign LUT_2[52300] = 32'b11111111111111100101111101011011;
assign LUT_2[52301] = 32'b11111111111111100010110101110100;
assign LUT_2[52302] = 32'b11111111111111101100110110010111;
assign LUT_2[52303] = 32'b11111111111111101001101110110000;
assign LUT_2[52304] = 32'b11111111111111101001010010100000;
assign LUT_2[52305] = 32'b11111111111111100110001010111001;
assign LUT_2[52306] = 32'b11111111111111110000001011011100;
assign LUT_2[52307] = 32'b11111111111111101101000011110101;
assign LUT_2[52308] = 32'b11111111111111100101110000001000;
assign LUT_2[52309] = 32'b11111111111111100010101000100001;
assign LUT_2[52310] = 32'b11111111111111101100101001000100;
assign LUT_2[52311] = 32'b11111111111111101001100001011101;
assign LUT_2[52312] = 32'b11111111111111100100000011111101;
assign LUT_2[52313] = 32'b11111111111111100000111100010110;
assign LUT_2[52314] = 32'b11111111111111101010111100111001;
assign LUT_2[52315] = 32'b11111111111111100111110101010010;
assign LUT_2[52316] = 32'b11111111111111100000100001100101;
assign LUT_2[52317] = 32'b11111111111111011101011001111110;
assign LUT_2[52318] = 32'b11111111111111100111011010100001;
assign LUT_2[52319] = 32'b11111111111111100100010010111010;
assign LUT_2[52320] = 32'b11111111111111101111001001111111;
assign LUT_2[52321] = 32'b11111111111111101100000010011000;
assign LUT_2[52322] = 32'b11111111111111110110000010111011;
assign LUT_2[52323] = 32'b11111111111111110010111011010100;
assign LUT_2[52324] = 32'b11111111111111101011100111100111;
assign LUT_2[52325] = 32'b11111111111111101000100000000000;
assign LUT_2[52326] = 32'b11111111111111110010100000100011;
assign LUT_2[52327] = 32'b11111111111111101111011000111100;
assign LUT_2[52328] = 32'b11111111111111101001111011011100;
assign LUT_2[52329] = 32'b11111111111111100110110011110101;
assign LUT_2[52330] = 32'b11111111111111110000110100011000;
assign LUT_2[52331] = 32'b11111111111111101101101100110001;
assign LUT_2[52332] = 32'b11111111111111100110011001000100;
assign LUT_2[52333] = 32'b11111111111111100011010001011101;
assign LUT_2[52334] = 32'b11111111111111101101010010000000;
assign LUT_2[52335] = 32'b11111111111111101010001010011001;
assign LUT_2[52336] = 32'b11111111111111101001101110001001;
assign LUT_2[52337] = 32'b11111111111111100110100110100010;
assign LUT_2[52338] = 32'b11111111111111110000100111000101;
assign LUT_2[52339] = 32'b11111111111111101101011111011110;
assign LUT_2[52340] = 32'b11111111111111100110001011110001;
assign LUT_2[52341] = 32'b11111111111111100011000100001010;
assign LUT_2[52342] = 32'b11111111111111101101000100101101;
assign LUT_2[52343] = 32'b11111111111111101001111101000110;
assign LUT_2[52344] = 32'b11111111111111100100011111100110;
assign LUT_2[52345] = 32'b11111111111111100001010111111111;
assign LUT_2[52346] = 32'b11111111111111101011011000100010;
assign LUT_2[52347] = 32'b11111111111111101000010000111011;
assign LUT_2[52348] = 32'b11111111111111100000111101001110;
assign LUT_2[52349] = 32'b11111111111111011101110101100111;
assign LUT_2[52350] = 32'b11111111111111100111110110001010;
assign LUT_2[52351] = 32'b11111111111111100100101110100011;
assign LUT_2[52352] = 32'b11111111111111111010111010000010;
assign LUT_2[52353] = 32'b11111111111111110111110010011011;
assign LUT_2[52354] = 32'b00000000000000000001110010111110;
assign LUT_2[52355] = 32'b11111111111111111110101011010111;
assign LUT_2[52356] = 32'b11111111111111110111010111101010;
assign LUT_2[52357] = 32'b11111111111111110100010000000011;
assign LUT_2[52358] = 32'b11111111111111111110010000100110;
assign LUT_2[52359] = 32'b11111111111111111011001000111111;
assign LUT_2[52360] = 32'b11111111111111110101101011011111;
assign LUT_2[52361] = 32'b11111111111111110010100011111000;
assign LUT_2[52362] = 32'b11111111111111111100100100011011;
assign LUT_2[52363] = 32'b11111111111111111001011100110100;
assign LUT_2[52364] = 32'b11111111111111110010001001000111;
assign LUT_2[52365] = 32'b11111111111111101111000001100000;
assign LUT_2[52366] = 32'b11111111111111111001000010000011;
assign LUT_2[52367] = 32'b11111111111111110101111010011100;
assign LUT_2[52368] = 32'b11111111111111110101011110001100;
assign LUT_2[52369] = 32'b11111111111111110010010110100101;
assign LUT_2[52370] = 32'b11111111111111111100010111001000;
assign LUT_2[52371] = 32'b11111111111111111001001111100001;
assign LUT_2[52372] = 32'b11111111111111110001111011110100;
assign LUT_2[52373] = 32'b11111111111111101110110100001101;
assign LUT_2[52374] = 32'b11111111111111111000110100110000;
assign LUT_2[52375] = 32'b11111111111111110101101101001001;
assign LUT_2[52376] = 32'b11111111111111110000001111101001;
assign LUT_2[52377] = 32'b11111111111111101101001000000010;
assign LUT_2[52378] = 32'b11111111111111110111001000100101;
assign LUT_2[52379] = 32'b11111111111111110100000000111110;
assign LUT_2[52380] = 32'b11111111111111101100101101010001;
assign LUT_2[52381] = 32'b11111111111111101001100101101010;
assign LUT_2[52382] = 32'b11111111111111110011100110001101;
assign LUT_2[52383] = 32'b11111111111111110000011110100110;
assign LUT_2[52384] = 32'b11111111111111111011010101101011;
assign LUT_2[52385] = 32'b11111111111111111000001110000100;
assign LUT_2[52386] = 32'b00000000000000000010001110100111;
assign LUT_2[52387] = 32'b11111111111111111111000111000000;
assign LUT_2[52388] = 32'b11111111111111110111110011010011;
assign LUT_2[52389] = 32'b11111111111111110100101011101100;
assign LUT_2[52390] = 32'b11111111111111111110101100001111;
assign LUT_2[52391] = 32'b11111111111111111011100100101000;
assign LUT_2[52392] = 32'b11111111111111110110000111001000;
assign LUT_2[52393] = 32'b11111111111111110010111111100001;
assign LUT_2[52394] = 32'b11111111111111111101000000000100;
assign LUT_2[52395] = 32'b11111111111111111001111000011101;
assign LUT_2[52396] = 32'b11111111111111110010100100110000;
assign LUT_2[52397] = 32'b11111111111111101111011101001001;
assign LUT_2[52398] = 32'b11111111111111111001011101101100;
assign LUT_2[52399] = 32'b11111111111111110110010110000101;
assign LUT_2[52400] = 32'b11111111111111110101111001110101;
assign LUT_2[52401] = 32'b11111111111111110010110010001110;
assign LUT_2[52402] = 32'b11111111111111111100110010110001;
assign LUT_2[52403] = 32'b11111111111111111001101011001010;
assign LUT_2[52404] = 32'b11111111111111110010010111011101;
assign LUT_2[52405] = 32'b11111111111111101111001111110110;
assign LUT_2[52406] = 32'b11111111111111111001010000011001;
assign LUT_2[52407] = 32'b11111111111111110110001000110010;
assign LUT_2[52408] = 32'b11111111111111110000101011010010;
assign LUT_2[52409] = 32'b11111111111111101101100011101011;
assign LUT_2[52410] = 32'b11111111111111110111100100001110;
assign LUT_2[52411] = 32'b11111111111111110100011100100111;
assign LUT_2[52412] = 32'b11111111111111101101001000111010;
assign LUT_2[52413] = 32'b11111111111111101010000001010011;
assign LUT_2[52414] = 32'b11111111111111110100000001110110;
assign LUT_2[52415] = 32'b11111111111111110000111010001111;
assign LUT_2[52416] = 32'b11111111111111110011000010100101;
assign LUT_2[52417] = 32'b11111111111111101111111010111110;
assign LUT_2[52418] = 32'b11111111111111111001111011100001;
assign LUT_2[52419] = 32'b11111111111111110110110011111010;
assign LUT_2[52420] = 32'b11111111111111101111100000001101;
assign LUT_2[52421] = 32'b11111111111111101100011000100110;
assign LUT_2[52422] = 32'b11111111111111110110011001001001;
assign LUT_2[52423] = 32'b11111111111111110011010001100010;
assign LUT_2[52424] = 32'b11111111111111101101110100000010;
assign LUT_2[52425] = 32'b11111111111111101010101100011011;
assign LUT_2[52426] = 32'b11111111111111110100101100111110;
assign LUT_2[52427] = 32'b11111111111111110001100101010111;
assign LUT_2[52428] = 32'b11111111111111101010010001101010;
assign LUT_2[52429] = 32'b11111111111111100111001010000011;
assign LUT_2[52430] = 32'b11111111111111110001001010100110;
assign LUT_2[52431] = 32'b11111111111111101110000010111111;
assign LUT_2[52432] = 32'b11111111111111101101100110101111;
assign LUT_2[52433] = 32'b11111111111111101010011111001000;
assign LUT_2[52434] = 32'b11111111111111110100011111101011;
assign LUT_2[52435] = 32'b11111111111111110001011000000100;
assign LUT_2[52436] = 32'b11111111111111101010000100010111;
assign LUT_2[52437] = 32'b11111111111111100110111100110000;
assign LUT_2[52438] = 32'b11111111111111110000111101010011;
assign LUT_2[52439] = 32'b11111111111111101101110101101100;
assign LUT_2[52440] = 32'b11111111111111101000011000001100;
assign LUT_2[52441] = 32'b11111111111111100101010000100101;
assign LUT_2[52442] = 32'b11111111111111101111010001001000;
assign LUT_2[52443] = 32'b11111111111111101100001001100001;
assign LUT_2[52444] = 32'b11111111111111100100110101110100;
assign LUT_2[52445] = 32'b11111111111111100001101110001101;
assign LUT_2[52446] = 32'b11111111111111101011101110110000;
assign LUT_2[52447] = 32'b11111111111111101000100111001001;
assign LUT_2[52448] = 32'b11111111111111110011011110001110;
assign LUT_2[52449] = 32'b11111111111111110000010110100111;
assign LUT_2[52450] = 32'b11111111111111111010010111001010;
assign LUT_2[52451] = 32'b11111111111111110111001111100011;
assign LUT_2[52452] = 32'b11111111111111101111111011110110;
assign LUT_2[52453] = 32'b11111111111111101100110100001111;
assign LUT_2[52454] = 32'b11111111111111110110110100110010;
assign LUT_2[52455] = 32'b11111111111111110011101101001011;
assign LUT_2[52456] = 32'b11111111111111101110001111101011;
assign LUT_2[52457] = 32'b11111111111111101011001000000100;
assign LUT_2[52458] = 32'b11111111111111110101001000100111;
assign LUT_2[52459] = 32'b11111111111111110010000001000000;
assign LUT_2[52460] = 32'b11111111111111101010101101010011;
assign LUT_2[52461] = 32'b11111111111111100111100101101100;
assign LUT_2[52462] = 32'b11111111111111110001100110001111;
assign LUT_2[52463] = 32'b11111111111111101110011110101000;
assign LUT_2[52464] = 32'b11111111111111101110000010011000;
assign LUT_2[52465] = 32'b11111111111111101010111010110001;
assign LUT_2[52466] = 32'b11111111111111110100111011010100;
assign LUT_2[52467] = 32'b11111111111111110001110011101101;
assign LUT_2[52468] = 32'b11111111111111101010100000000000;
assign LUT_2[52469] = 32'b11111111111111100111011000011001;
assign LUT_2[52470] = 32'b11111111111111110001011000111100;
assign LUT_2[52471] = 32'b11111111111111101110010001010101;
assign LUT_2[52472] = 32'b11111111111111101000110011110101;
assign LUT_2[52473] = 32'b11111111111111100101101100001110;
assign LUT_2[52474] = 32'b11111111111111101111101100110001;
assign LUT_2[52475] = 32'b11111111111111101100100101001010;
assign LUT_2[52476] = 32'b11111111111111100101010001011101;
assign LUT_2[52477] = 32'b11111111111111100010001001110110;
assign LUT_2[52478] = 32'b11111111111111101100001010011001;
assign LUT_2[52479] = 32'b11111111111111101001000010110010;
assign LUT_2[52480] = 32'b11111111111111111010100100011001;
assign LUT_2[52481] = 32'b11111111111111110111011100110010;
assign LUT_2[52482] = 32'b00000000000000000001011101010101;
assign LUT_2[52483] = 32'b11111111111111111110010101101110;
assign LUT_2[52484] = 32'b11111111111111110111000010000001;
assign LUT_2[52485] = 32'b11111111111111110011111010011010;
assign LUT_2[52486] = 32'b11111111111111111101111010111101;
assign LUT_2[52487] = 32'b11111111111111111010110011010110;
assign LUT_2[52488] = 32'b11111111111111110101010101110110;
assign LUT_2[52489] = 32'b11111111111111110010001110001111;
assign LUT_2[52490] = 32'b11111111111111111100001110110010;
assign LUT_2[52491] = 32'b11111111111111111001000111001011;
assign LUT_2[52492] = 32'b11111111111111110001110011011110;
assign LUT_2[52493] = 32'b11111111111111101110101011110111;
assign LUT_2[52494] = 32'b11111111111111111000101100011010;
assign LUT_2[52495] = 32'b11111111111111110101100100110011;
assign LUT_2[52496] = 32'b11111111111111110101001000100011;
assign LUT_2[52497] = 32'b11111111111111110010000000111100;
assign LUT_2[52498] = 32'b11111111111111111100000001011111;
assign LUT_2[52499] = 32'b11111111111111111000111001111000;
assign LUT_2[52500] = 32'b11111111111111110001100110001011;
assign LUT_2[52501] = 32'b11111111111111101110011110100100;
assign LUT_2[52502] = 32'b11111111111111111000011111000111;
assign LUT_2[52503] = 32'b11111111111111110101010111100000;
assign LUT_2[52504] = 32'b11111111111111101111111010000000;
assign LUT_2[52505] = 32'b11111111111111101100110010011001;
assign LUT_2[52506] = 32'b11111111111111110110110010111100;
assign LUT_2[52507] = 32'b11111111111111110011101011010101;
assign LUT_2[52508] = 32'b11111111111111101100010111101000;
assign LUT_2[52509] = 32'b11111111111111101001010000000001;
assign LUT_2[52510] = 32'b11111111111111110011010000100100;
assign LUT_2[52511] = 32'b11111111111111110000001000111101;
assign LUT_2[52512] = 32'b11111111111111111011000000000010;
assign LUT_2[52513] = 32'b11111111111111110111111000011011;
assign LUT_2[52514] = 32'b00000000000000000001111000111110;
assign LUT_2[52515] = 32'b11111111111111111110110001010111;
assign LUT_2[52516] = 32'b11111111111111110111011101101010;
assign LUT_2[52517] = 32'b11111111111111110100010110000011;
assign LUT_2[52518] = 32'b11111111111111111110010110100110;
assign LUT_2[52519] = 32'b11111111111111111011001110111111;
assign LUT_2[52520] = 32'b11111111111111110101110001011111;
assign LUT_2[52521] = 32'b11111111111111110010101001111000;
assign LUT_2[52522] = 32'b11111111111111111100101010011011;
assign LUT_2[52523] = 32'b11111111111111111001100010110100;
assign LUT_2[52524] = 32'b11111111111111110010001111000111;
assign LUT_2[52525] = 32'b11111111111111101111000111100000;
assign LUT_2[52526] = 32'b11111111111111111001001000000011;
assign LUT_2[52527] = 32'b11111111111111110110000000011100;
assign LUT_2[52528] = 32'b11111111111111110101100100001100;
assign LUT_2[52529] = 32'b11111111111111110010011100100101;
assign LUT_2[52530] = 32'b11111111111111111100011101001000;
assign LUT_2[52531] = 32'b11111111111111111001010101100001;
assign LUT_2[52532] = 32'b11111111111111110010000001110100;
assign LUT_2[52533] = 32'b11111111111111101110111010001101;
assign LUT_2[52534] = 32'b11111111111111111000111010110000;
assign LUT_2[52535] = 32'b11111111111111110101110011001001;
assign LUT_2[52536] = 32'b11111111111111110000010101101001;
assign LUT_2[52537] = 32'b11111111111111101101001110000010;
assign LUT_2[52538] = 32'b11111111111111110111001110100101;
assign LUT_2[52539] = 32'b11111111111111110100000110111110;
assign LUT_2[52540] = 32'b11111111111111101100110011010001;
assign LUT_2[52541] = 32'b11111111111111101001101011101010;
assign LUT_2[52542] = 32'b11111111111111110011101100001101;
assign LUT_2[52543] = 32'b11111111111111110000100100100110;
assign LUT_2[52544] = 32'b11111111111111110010101100111100;
assign LUT_2[52545] = 32'b11111111111111101111100101010101;
assign LUT_2[52546] = 32'b11111111111111111001100101111000;
assign LUT_2[52547] = 32'b11111111111111110110011110010001;
assign LUT_2[52548] = 32'b11111111111111101111001010100100;
assign LUT_2[52549] = 32'b11111111111111101100000010111101;
assign LUT_2[52550] = 32'b11111111111111110110000011100000;
assign LUT_2[52551] = 32'b11111111111111110010111011111001;
assign LUT_2[52552] = 32'b11111111111111101101011110011001;
assign LUT_2[52553] = 32'b11111111111111101010010110110010;
assign LUT_2[52554] = 32'b11111111111111110100010111010101;
assign LUT_2[52555] = 32'b11111111111111110001001111101110;
assign LUT_2[52556] = 32'b11111111111111101001111100000001;
assign LUT_2[52557] = 32'b11111111111111100110110100011010;
assign LUT_2[52558] = 32'b11111111111111110000110100111101;
assign LUT_2[52559] = 32'b11111111111111101101101101010110;
assign LUT_2[52560] = 32'b11111111111111101101010001000110;
assign LUT_2[52561] = 32'b11111111111111101010001001011111;
assign LUT_2[52562] = 32'b11111111111111110100001010000010;
assign LUT_2[52563] = 32'b11111111111111110001000010011011;
assign LUT_2[52564] = 32'b11111111111111101001101110101110;
assign LUT_2[52565] = 32'b11111111111111100110100111000111;
assign LUT_2[52566] = 32'b11111111111111110000100111101010;
assign LUT_2[52567] = 32'b11111111111111101101100000000011;
assign LUT_2[52568] = 32'b11111111111111101000000010100011;
assign LUT_2[52569] = 32'b11111111111111100100111010111100;
assign LUT_2[52570] = 32'b11111111111111101110111011011111;
assign LUT_2[52571] = 32'b11111111111111101011110011111000;
assign LUT_2[52572] = 32'b11111111111111100100100000001011;
assign LUT_2[52573] = 32'b11111111111111100001011000100100;
assign LUT_2[52574] = 32'b11111111111111101011011001000111;
assign LUT_2[52575] = 32'b11111111111111101000010001100000;
assign LUT_2[52576] = 32'b11111111111111110011001000100101;
assign LUT_2[52577] = 32'b11111111111111110000000000111110;
assign LUT_2[52578] = 32'b11111111111111111010000001100001;
assign LUT_2[52579] = 32'b11111111111111110110111001111010;
assign LUT_2[52580] = 32'b11111111111111101111100110001101;
assign LUT_2[52581] = 32'b11111111111111101100011110100110;
assign LUT_2[52582] = 32'b11111111111111110110011111001001;
assign LUT_2[52583] = 32'b11111111111111110011010111100010;
assign LUT_2[52584] = 32'b11111111111111101101111010000010;
assign LUT_2[52585] = 32'b11111111111111101010110010011011;
assign LUT_2[52586] = 32'b11111111111111110100110010111110;
assign LUT_2[52587] = 32'b11111111111111110001101011010111;
assign LUT_2[52588] = 32'b11111111111111101010010111101010;
assign LUT_2[52589] = 32'b11111111111111100111010000000011;
assign LUT_2[52590] = 32'b11111111111111110001010000100110;
assign LUT_2[52591] = 32'b11111111111111101110001000111111;
assign LUT_2[52592] = 32'b11111111111111101101101100101111;
assign LUT_2[52593] = 32'b11111111111111101010100101001000;
assign LUT_2[52594] = 32'b11111111111111110100100101101011;
assign LUT_2[52595] = 32'b11111111111111110001011110000100;
assign LUT_2[52596] = 32'b11111111111111101010001010010111;
assign LUT_2[52597] = 32'b11111111111111100111000010110000;
assign LUT_2[52598] = 32'b11111111111111110001000011010011;
assign LUT_2[52599] = 32'b11111111111111101101111011101100;
assign LUT_2[52600] = 32'b11111111111111101000011110001100;
assign LUT_2[52601] = 32'b11111111111111100101010110100101;
assign LUT_2[52602] = 32'b11111111111111101111010111001000;
assign LUT_2[52603] = 32'b11111111111111101100001111100001;
assign LUT_2[52604] = 32'b11111111111111100100111011110100;
assign LUT_2[52605] = 32'b11111111111111100001110100001101;
assign LUT_2[52606] = 32'b11111111111111101011110100110000;
assign LUT_2[52607] = 32'b11111111111111101000101101001001;
assign LUT_2[52608] = 32'b11111111111111111110111000101000;
assign LUT_2[52609] = 32'b11111111111111111011110001000001;
assign LUT_2[52610] = 32'b00000000000000000101110001100100;
assign LUT_2[52611] = 32'b00000000000000000010101001111101;
assign LUT_2[52612] = 32'b11111111111111111011010110010000;
assign LUT_2[52613] = 32'b11111111111111111000001110101001;
assign LUT_2[52614] = 32'b00000000000000000010001111001100;
assign LUT_2[52615] = 32'b11111111111111111111000111100101;
assign LUT_2[52616] = 32'b11111111111111111001101010000101;
assign LUT_2[52617] = 32'b11111111111111110110100010011110;
assign LUT_2[52618] = 32'b00000000000000000000100011000001;
assign LUT_2[52619] = 32'b11111111111111111101011011011010;
assign LUT_2[52620] = 32'b11111111111111110110000111101101;
assign LUT_2[52621] = 32'b11111111111111110011000000000110;
assign LUT_2[52622] = 32'b11111111111111111101000000101001;
assign LUT_2[52623] = 32'b11111111111111111001111001000010;
assign LUT_2[52624] = 32'b11111111111111111001011100110010;
assign LUT_2[52625] = 32'b11111111111111110110010101001011;
assign LUT_2[52626] = 32'b00000000000000000000010101101110;
assign LUT_2[52627] = 32'b11111111111111111101001110000111;
assign LUT_2[52628] = 32'b11111111111111110101111010011010;
assign LUT_2[52629] = 32'b11111111111111110010110010110011;
assign LUT_2[52630] = 32'b11111111111111111100110011010110;
assign LUT_2[52631] = 32'b11111111111111111001101011101111;
assign LUT_2[52632] = 32'b11111111111111110100001110001111;
assign LUT_2[52633] = 32'b11111111111111110001000110101000;
assign LUT_2[52634] = 32'b11111111111111111011000111001011;
assign LUT_2[52635] = 32'b11111111111111110111111111100100;
assign LUT_2[52636] = 32'b11111111111111110000101011110111;
assign LUT_2[52637] = 32'b11111111111111101101100100010000;
assign LUT_2[52638] = 32'b11111111111111110111100100110011;
assign LUT_2[52639] = 32'b11111111111111110100011101001100;
assign LUT_2[52640] = 32'b11111111111111111111010100010001;
assign LUT_2[52641] = 32'b11111111111111111100001100101010;
assign LUT_2[52642] = 32'b00000000000000000110001101001101;
assign LUT_2[52643] = 32'b00000000000000000011000101100110;
assign LUT_2[52644] = 32'b11111111111111111011110001111001;
assign LUT_2[52645] = 32'b11111111111111111000101010010010;
assign LUT_2[52646] = 32'b00000000000000000010101010110101;
assign LUT_2[52647] = 32'b11111111111111111111100011001110;
assign LUT_2[52648] = 32'b11111111111111111010000101101110;
assign LUT_2[52649] = 32'b11111111111111110110111110000111;
assign LUT_2[52650] = 32'b00000000000000000000111110101010;
assign LUT_2[52651] = 32'b11111111111111111101110111000011;
assign LUT_2[52652] = 32'b11111111111111110110100011010110;
assign LUT_2[52653] = 32'b11111111111111110011011011101111;
assign LUT_2[52654] = 32'b11111111111111111101011100010010;
assign LUT_2[52655] = 32'b11111111111111111010010100101011;
assign LUT_2[52656] = 32'b11111111111111111001111000011011;
assign LUT_2[52657] = 32'b11111111111111110110110000110100;
assign LUT_2[52658] = 32'b00000000000000000000110001010111;
assign LUT_2[52659] = 32'b11111111111111111101101001110000;
assign LUT_2[52660] = 32'b11111111111111110110010110000011;
assign LUT_2[52661] = 32'b11111111111111110011001110011100;
assign LUT_2[52662] = 32'b11111111111111111101001110111111;
assign LUT_2[52663] = 32'b11111111111111111010000111011000;
assign LUT_2[52664] = 32'b11111111111111110100101001111000;
assign LUT_2[52665] = 32'b11111111111111110001100010010001;
assign LUT_2[52666] = 32'b11111111111111111011100010110100;
assign LUT_2[52667] = 32'b11111111111111111000011011001101;
assign LUT_2[52668] = 32'b11111111111111110001000111100000;
assign LUT_2[52669] = 32'b11111111111111101101111111111001;
assign LUT_2[52670] = 32'b11111111111111111000000000011100;
assign LUT_2[52671] = 32'b11111111111111110100111000110101;
assign LUT_2[52672] = 32'b11111111111111110111000001001011;
assign LUT_2[52673] = 32'b11111111111111110011111001100100;
assign LUT_2[52674] = 32'b11111111111111111101111010000111;
assign LUT_2[52675] = 32'b11111111111111111010110010100000;
assign LUT_2[52676] = 32'b11111111111111110011011110110011;
assign LUT_2[52677] = 32'b11111111111111110000010111001100;
assign LUT_2[52678] = 32'b11111111111111111010010111101111;
assign LUT_2[52679] = 32'b11111111111111110111010000001000;
assign LUT_2[52680] = 32'b11111111111111110001110010101000;
assign LUT_2[52681] = 32'b11111111111111101110101011000001;
assign LUT_2[52682] = 32'b11111111111111111000101011100100;
assign LUT_2[52683] = 32'b11111111111111110101100011111101;
assign LUT_2[52684] = 32'b11111111111111101110010000010000;
assign LUT_2[52685] = 32'b11111111111111101011001000101001;
assign LUT_2[52686] = 32'b11111111111111110101001001001100;
assign LUT_2[52687] = 32'b11111111111111110010000001100101;
assign LUT_2[52688] = 32'b11111111111111110001100101010101;
assign LUT_2[52689] = 32'b11111111111111101110011101101110;
assign LUT_2[52690] = 32'b11111111111111111000011110010001;
assign LUT_2[52691] = 32'b11111111111111110101010110101010;
assign LUT_2[52692] = 32'b11111111111111101110000010111101;
assign LUT_2[52693] = 32'b11111111111111101010111011010110;
assign LUT_2[52694] = 32'b11111111111111110100111011111001;
assign LUT_2[52695] = 32'b11111111111111110001110100010010;
assign LUT_2[52696] = 32'b11111111111111101100010110110010;
assign LUT_2[52697] = 32'b11111111111111101001001111001011;
assign LUT_2[52698] = 32'b11111111111111110011001111101110;
assign LUT_2[52699] = 32'b11111111111111110000001000000111;
assign LUT_2[52700] = 32'b11111111111111101000110100011010;
assign LUT_2[52701] = 32'b11111111111111100101101100110011;
assign LUT_2[52702] = 32'b11111111111111101111101101010110;
assign LUT_2[52703] = 32'b11111111111111101100100101101111;
assign LUT_2[52704] = 32'b11111111111111110111011100110100;
assign LUT_2[52705] = 32'b11111111111111110100010101001101;
assign LUT_2[52706] = 32'b11111111111111111110010101110000;
assign LUT_2[52707] = 32'b11111111111111111011001110001001;
assign LUT_2[52708] = 32'b11111111111111110011111010011100;
assign LUT_2[52709] = 32'b11111111111111110000110010110101;
assign LUT_2[52710] = 32'b11111111111111111010110011011000;
assign LUT_2[52711] = 32'b11111111111111110111101011110001;
assign LUT_2[52712] = 32'b11111111111111110010001110010001;
assign LUT_2[52713] = 32'b11111111111111101111000110101010;
assign LUT_2[52714] = 32'b11111111111111111001000111001101;
assign LUT_2[52715] = 32'b11111111111111110101111111100110;
assign LUT_2[52716] = 32'b11111111111111101110101011111001;
assign LUT_2[52717] = 32'b11111111111111101011100100010010;
assign LUT_2[52718] = 32'b11111111111111110101100100110101;
assign LUT_2[52719] = 32'b11111111111111110010011101001110;
assign LUT_2[52720] = 32'b11111111111111110010000000111110;
assign LUT_2[52721] = 32'b11111111111111101110111001010111;
assign LUT_2[52722] = 32'b11111111111111111000111001111010;
assign LUT_2[52723] = 32'b11111111111111110101110010010011;
assign LUT_2[52724] = 32'b11111111111111101110011110100110;
assign LUT_2[52725] = 32'b11111111111111101011010110111111;
assign LUT_2[52726] = 32'b11111111111111110101010111100010;
assign LUT_2[52727] = 32'b11111111111111110010001111111011;
assign LUT_2[52728] = 32'b11111111111111101100110010011011;
assign LUT_2[52729] = 32'b11111111111111101001101010110100;
assign LUT_2[52730] = 32'b11111111111111110011101011010111;
assign LUT_2[52731] = 32'b11111111111111110000100011110000;
assign LUT_2[52732] = 32'b11111111111111101001010000000011;
assign LUT_2[52733] = 32'b11111111111111100110001000011100;
assign LUT_2[52734] = 32'b11111111111111110000001000111111;
assign LUT_2[52735] = 32'b11111111111111101101000001011000;
assign LUT_2[52736] = 32'b11111111111111111011010111100101;
assign LUT_2[52737] = 32'b11111111111111111000001111111110;
assign LUT_2[52738] = 32'b00000000000000000010010000100001;
assign LUT_2[52739] = 32'b11111111111111111111001000111010;
assign LUT_2[52740] = 32'b11111111111111110111110101001101;
assign LUT_2[52741] = 32'b11111111111111110100101101100110;
assign LUT_2[52742] = 32'b11111111111111111110101110001001;
assign LUT_2[52743] = 32'b11111111111111111011100110100010;
assign LUT_2[52744] = 32'b11111111111111110110001001000010;
assign LUT_2[52745] = 32'b11111111111111110011000001011011;
assign LUT_2[52746] = 32'b11111111111111111101000001111110;
assign LUT_2[52747] = 32'b11111111111111111001111010010111;
assign LUT_2[52748] = 32'b11111111111111110010100110101010;
assign LUT_2[52749] = 32'b11111111111111101111011111000011;
assign LUT_2[52750] = 32'b11111111111111111001011111100110;
assign LUT_2[52751] = 32'b11111111111111110110010111111111;
assign LUT_2[52752] = 32'b11111111111111110101111011101111;
assign LUT_2[52753] = 32'b11111111111111110010110100001000;
assign LUT_2[52754] = 32'b11111111111111111100110100101011;
assign LUT_2[52755] = 32'b11111111111111111001101101000100;
assign LUT_2[52756] = 32'b11111111111111110010011001010111;
assign LUT_2[52757] = 32'b11111111111111101111010001110000;
assign LUT_2[52758] = 32'b11111111111111111001010010010011;
assign LUT_2[52759] = 32'b11111111111111110110001010101100;
assign LUT_2[52760] = 32'b11111111111111110000101101001100;
assign LUT_2[52761] = 32'b11111111111111101101100101100101;
assign LUT_2[52762] = 32'b11111111111111110111100110001000;
assign LUT_2[52763] = 32'b11111111111111110100011110100001;
assign LUT_2[52764] = 32'b11111111111111101101001010110100;
assign LUT_2[52765] = 32'b11111111111111101010000011001101;
assign LUT_2[52766] = 32'b11111111111111110100000011110000;
assign LUT_2[52767] = 32'b11111111111111110000111100001001;
assign LUT_2[52768] = 32'b11111111111111111011110011001110;
assign LUT_2[52769] = 32'b11111111111111111000101011100111;
assign LUT_2[52770] = 32'b00000000000000000010101100001010;
assign LUT_2[52771] = 32'b11111111111111111111100100100011;
assign LUT_2[52772] = 32'b11111111111111111000010000110110;
assign LUT_2[52773] = 32'b11111111111111110101001001001111;
assign LUT_2[52774] = 32'b11111111111111111111001001110010;
assign LUT_2[52775] = 32'b11111111111111111100000010001011;
assign LUT_2[52776] = 32'b11111111111111110110100100101011;
assign LUT_2[52777] = 32'b11111111111111110011011101000100;
assign LUT_2[52778] = 32'b11111111111111111101011101100111;
assign LUT_2[52779] = 32'b11111111111111111010010110000000;
assign LUT_2[52780] = 32'b11111111111111110011000010010011;
assign LUT_2[52781] = 32'b11111111111111101111111010101100;
assign LUT_2[52782] = 32'b11111111111111111001111011001111;
assign LUT_2[52783] = 32'b11111111111111110110110011101000;
assign LUT_2[52784] = 32'b11111111111111110110010111011000;
assign LUT_2[52785] = 32'b11111111111111110011001111110001;
assign LUT_2[52786] = 32'b11111111111111111101010000010100;
assign LUT_2[52787] = 32'b11111111111111111010001000101101;
assign LUT_2[52788] = 32'b11111111111111110010110101000000;
assign LUT_2[52789] = 32'b11111111111111101111101101011001;
assign LUT_2[52790] = 32'b11111111111111111001101101111100;
assign LUT_2[52791] = 32'b11111111111111110110100110010101;
assign LUT_2[52792] = 32'b11111111111111110001001000110101;
assign LUT_2[52793] = 32'b11111111111111101110000001001110;
assign LUT_2[52794] = 32'b11111111111111111000000001110001;
assign LUT_2[52795] = 32'b11111111111111110100111010001010;
assign LUT_2[52796] = 32'b11111111111111101101100110011101;
assign LUT_2[52797] = 32'b11111111111111101010011110110110;
assign LUT_2[52798] = 32'b11111111111111110100011111011001;
assign LUT_2[52799] = 32'b11111111111111110001010111110010;
assign LUT_2[52800] = 32'b11111111111111110011100000001000;
assign LUT_2[52801] = 32'b11111111111111110000011000100001;
assign LUT_2[52802] = 32'b11111111111111111010011001000100;
assign LUT_2[52803] = 32'b11111111111111110111010001011101;
assign LUT_2[52804] = 32'b11111111111111101111111101110000;
assign LUT_2[52805] = 32'b11111111111111101100110110001001;
assign LUT_2[52806] = 32'b11111111111111110110110110101100;
assign LUT_2[52807] = 32'b11111111111111110011101111000101;
assign LUT_2[52808] = 32'b11111111111111101110010001100101;
assign LUT_2[52809] = 32'b11111111111111101011001001111110;
assign LUT_2[52810] = 32'b11111111111111110101001010100001;
assign LUT_2[52811] = 32'b11111111111111110010000010111010;
assign LUT_2[52812] = 32'b11111111111111101010101111001101;
assign LUT_2[52813] = 32'b11111111111111100111100111100110;
assign LUT_2[52814] = 32'b11111111111111110001101000001001;
assign LUT_2[52815] = 32'b11111111111111101110100000100010;
assign LUT_2[52816] = 32'b11111111111111101110000100010010;
assign LUT_2[52817] = 32'b11111111111111101010111100101011;
assign LUT_2[52818] = 32'b11111111111111110100111101001110;
assign LUT_2[52819] = 32'b11111111111111110001110101100111;
assign LUT_2[52820] = 32'b11111111111111101010100001111010;
assign LUT_2[52821] = 32'b11111111111111100111011010010011;
assign LUT_2[52822] = 32'b11111111111111110001011010110110;
assign LUT_2[52823] = 32'b11111111111111101110010011001111;
assign LUT_2[52824] = 32'b11111111111111101000110101101111;
assign LUT_2[52825] = 32'b11111111111111100101101110001000;
assign LUT_2[52826] = 32'b11111111111111101111101110101011;
assign LUT_2[52827] = 32'b11111111111111101100100111000100;
assign LUT_2[52828] = 32'b11111111111111100101010011010111;
assign LUT_2[52829] = 32'b11111111111111100010001011110000;
assign LUT_2[52830] = 32'b11111111111111101100001100010011;
assign LUT_2[52831] = 32'b11111111111111101001000100101100;
assign LUT_2[52832] = 32'b11111111111111110011111011110001;
assign LUT_2[52833] = 32'b11111111111111110000110100001010;
assign LUT_2[52834] = 32'b11111111111111111010110100101101;
assign LUT_2[52835] = 32'b11111111111111110111101101000110;
assign LUT_2[52836] = 32'b11111111111111110000011001011001;
assign LUT_2[52837] = 32'b11111111111111101101010001110010;
assign LUT_2[52838] = 32'b11111111111111110111010010010101;
assign LUT_2[52839] = 32'b11111111111111110100001010101110;
assign LUT_2[52840] = 32'b11111111111111101110101101001110;
assign LUT_2[52841] = 32'b11111111111111101011100101100111;
assign LUT_2[52842] = 32'b11111111111111110101100110001010;
assign LUT_2[52843] = 32'b11111111111111110010011110100011;
assign LUT_2[52844] = 32'b11111111111111101011001010110110;
assign LUT_2[52845] = 32'b11111111111111101000000011001111;
assign LUT_2[52846] = 32'b11111111111111110010000011110010;
assign LUT_2[52847] = 32'b11111111111111101110111100001011;
assign LUT_2[52848] = 32'b11111111111111101110011111111011;
assign LUT_2[52849] = 32'b11111111111111101011011000010100;
assign LUT_2[52850] = 32'b11111111111111110101011000110111;
assign LUT_2[52851] = 32'b11111111111111110010010001010000;
assign LUT_2[52852] = 32'b11111111111111101010111101100011;
assign LUT_2[52853] = 32'b11111111111111100111110101111100;
assign LUT_2[52854] = 32'b11111111111111110001110110011111;
assign LUT_2[52855] = 32'b11111111111111101110101110111000;
assign LUT_2[52856] = 32'b11111111111111101001010001011000;
assign LUT_2[52857] = 32'b11111111111111100110001001110001;
assign LUT_2[52858] = 32'b11111111111111110000001010010100;
assign LUT_2[52859] = 32'b11111111111111101101000010101101;
assign LUT_2[52860] = 32'b11111111111111100101101111000000;
assign LUT_2[52861] = 32'b11111111111111100010100111011001;
assign LUT_2[52862] = 32'b11111111111111101100100111111100;
assign LUT_2[52863] = 32'b11111111111111101001100000010101;
assign LUT_2[52864] = 32'b11111111111111111111101011110100;
assign LUT_2[52865] = 32'b11111111111111111100100100001101;
assign LUT_2[52866] = 32'b00000000000000000110100100110000;
assign LUT_2[52867] = 32'b00000000000000000011011101001001;
assign LUT_2[52868] = 32'b11111111111111111100001001011100;
assign LUT_2[52869] = 32'b11111111111111111001000001110101;
assign LUT_2[52870] = 32'b00000000000000000011000010011000;
assign LUT_2[52871] = 32'b11111111111111111111111010110001;
assign LUT_2[52872] = 32'b11111111111111111010011101010001;
assign LUT_2[52873] = 32'b11111111111111110111010101101010;
assign LUT_2[52874] = 32'b00000000000000000001010110001101;
assign LUT_2[52875] = 32'b11111111111111111110001110100110;
assign LUT_2[52876] = 32'b11111111111111110110111010111001;
assign LUT_2[52877] = 32'b11111111111111110011110011010010;
assign LUT_2[52878] = 32'b11111111111111111101110011110101;
assign LUT_2[52879] = 32'b11111111111111111010101100001110;
assign LUT_2[52880] = 32'b11111111111111111010001111111110;
assign LUT_2[52881] = 32'b11111111111111110111001000010111;
assign LUT_2[52882] = 32'b00000000000000000001001000111010;
assign LUT_2[52883] = 32'b11111111111111111110000001010011;
assign LUT_2[52884] = 32'b11111111111111110110101101100110;
assign LUT_2[52885] = 32'b11111111111111110011100101111111;
assign LUT_2[52886] = 32'b11111111111111111101100110100010;
assign LUT_2[52887] = 32'b11111111111111111010011110111011;
assign LUT_2[52888] = 32'b11111111111111110101000001011011;
assign LUT_2[52889] = 32'b11111111111111110001111001110100;
assign LUT_2[52890] = 32'b11111111111111111011111010010111;
assign LUT_2[52891] = 32'b11111111111111111000110010110000;
assign LUT_2[52892] = 32'b11111111111111110001011111000011;
assign LUT_2[52893] = 32'b11111111111111101110010111011100;
assign LUT_2[52894] = 32'b11111111111111111000010111111111;
assign LUT_2[52895] = 32'b11111111111111110101010000011000;
assign LUT_2[52896] = 32'b00000000000000000000000111011101;
assign LUT_2[52897] = 32'b11111111111111111100111111110110;
assign LUT_2[52898] = 32'b00000000000000000111000000011001;
assign LUT_2[52899] = 32'b00000000000000000011111000110010;
assign LUT_2[52900] = 32'b11111111111111111100100101000101;
assign LUT_2[52901] = 32'b11111111111111111001011101011110;
assign LUT_2[52902] = 32'b00000000000000000011011110000001;
assign LUT_2[52903] = 32'b00000000000000000000010110011010;
assign LUT_2[52904] = 32'b11111111111111111010111000111010;
assign LUT_2[52905] = 32'b11111111111111110111110001010011;
assign LUT_2[52906] = 32'b00000000000000000001110001110110;
assign LUT_2[52907] = 32'b11111111111111111110101010001111;
assign LUT_2[52908] = 32'b11111111111111110111010110100010;
assign LUT_2[52909] = 32'b11111111111111110100001110111011;
assign LUT_2[52910] = 32'b11111111111111111110001111011110;
assign LUT_2[52911] = 32'b11111111111111111011000111110111;
assign LUT_2[52912] = 32'b11111111111111111010101011100111;
assign LUT_2[52913] = 32'b11111111111111110111100100000000;
assign LUT_2[52914] = 32'b00000000000000000001100100100011;
assign LUT_2[52915] = 32'b11111111111111111110011100111100;
assign LUT_2[52916] = 32'b11111111111111110111001001001111;
assign LUT_2[52917] = 32'b11111111111111110100000001101000;
assign LUT_2[52918] = 32'b11111111111111111110000010001011;
assign LUT_2[52919] = 32'b11111111111111111010111010100100;
assign LUT_2[52920] = 32'b11111111111111110101011101000100;
assign LUT_2[52921] = 32'b11111111111111110010010101011101;
assign LUT_2[52922] = 32'b11111111111111111100010110000000;
assign LUT_2[52923] = 32'b11111111111111111001001110011001;
assign LUT_2[52924] = 32'b11111111111111110001111010101100;
assign LUT_2[52925] = 32'b11111111111111101110110011000101;
assign LUT_2[52926] = 32'b11111111111111111000110011101000;
assign LUT_2[52927] = 32'b11111111111111110101101100000001;
assign LUT_2[52928] = 32'b11111111111111110111110100010111;
assign LUT_2[52929] = 32'b11111111111111110100101100110000;
assign LUT_2[52930] = 32'b11111111111111111110101101010011;
assign LUT_2[52931] = 32'b11111111111111111011100101101100;
assign LUT_2[52932] = 32'b11111111111111110100010001111111;
assign LUT_2[52933] = 32'b11111111111111110001001010011000;
assign LUT_2[52934] = 32'b11111111111111111011001010111011;
assign LUT_2[52935] = 32'b11111111111111111000000011010100;
assign LUT_2[52936] = 32'b11111111111111110010100101110100;
assign LUT_2[52937] = 32'b11111111111111101111011110001101;
assign LUT_2[52938] = 32'b11111111111111111001011110110000;
assign LUT_2[52939] = 32'b11111111111111110110010111001001;
assign LUT_2[52940] = 32'b11111111111111101111000011011100;
assign LUT_2[52941] = 32'b11111111111111101011111011110101;
assign LUT_2[52942] = 32'b11111111111111110101111100011000;
assign LUT_2[52943] = 32'b11111111111111110010110100110001;
assign LUT_2[52944] = 32'b11111111111111110010011000100001;
assign LUT_2[52945] = 32'b11111111111111101111010000111010;
assign LUT_2[52946] = 32'b11111111111111111001010001011101;
assign LUT_2[52947] = 32'b11111111111111110110001001110110;
assign LUT_2[52948] = 32'b11111111111111101110110110001001;
assign LUT_2[52949] = 32'b11111111111111101011101110100010;
assign LUT_2[52950] = 32'b11111111111111110101101111000101;
assign LUT_2[52951] = 32'b11111111111111110010100111011110;
assign LUT_2[52952] = 32'b11111111111111101101001001111110;
assign LUT_2[52953] = 32'b11111111111111101010000010010111;
assign LUT_2[52954] = 32'b11111111111111110100000010111010;
assign LUT_2[52955] = 32'b11111111111111110000111011010011;
assign LUT_2[52956] = 32'b11111111111111101001100111100110;
assign LUT_2[52957] = 32'b11111111111111100110011111111111;
assign LUT_2[52958] = 32'b11111111111111110000100000100010;
assign LUT_2[52959] = 32'b11111111111111101101011000111011;
assign LUT_2[52960] = 32'b11111111111111111000010000000000;
assign LUT_2[52961] = 32'b11111111111111110101001000011001;
assign LUT_2[52962] = 32'b11111111111111111111001000111100;
assign LUT_2[52963] = 32'b11111111111111111100000001010101;
assign LUT_2[52964] = 32'b11111111111111110100101101101000;
assign LUT_2[52965] = 32'b11111111111111110001100110000001;
assign LUT_2[52966] = 32'b11111111111111111011100110100100;
assign LUT_2[52967] = 32'b11111111111111111000011110111101;
assign LUT_2[52968] = 32'b11111111111111110011000001011101;
assign LUT_2[52969] = 32'b11111111111111101111111001110110;
assign LUT_2[52970] = 32'b11111111111111111001111010011001;
assign LUT_2[52971] = 32'b11111111111111110110110010110010;
assign LUT_2[52972] = 32'b11111111111111101111011111000101;
assign LUT_2[52973] = 32'b11111111111111101100010111011110;
assign LUT_2[52974] = 32'b11111111111111110110011000000001;
assign LUT_2[52975] = 32'b11111111111111110011010000011010;
assign LUT_2[52976] = 32'b11111111111111110010110100001010;
assign LUT_2[52977] = 32'b11111111111111101111101100100011;
assign LUT_2[52978] = 32'b11111111111111111001101101000110;
assign LUT_2[52979] = 32'b11111111111111110110100101011111;
assign LUT_2[52980] = 32'b11111111111111101111010001110010;
assign LUT_2[52981] = 32'b11111111111111101100001010001011;
assign LUT_2[52982] = 32'b11111111111111110110001010101110;
assign LUT_2[52983] = 32'b11111111111111110011000011000111;
assign LUT_2[52984] = 32'b11111111111111101101100101100111;
assign LUT_2[52985] = 32'b11111111111111101010011110000000;
assign LUT_2[52986] = 32'b11111111111111110100011110100011;
assign LUT_2[52987] = 32'b11111111111111110001010110111100;
assign LUT_2[52988] = 32'b11111111111111101010000011001111;
assign LUT_2[52989] = 32'b11111111111111100110111011101000;
assign LUT_2[52990] = 32'b11111111111111110000111100001011;
assign LUT_2[52991] = 32'b11111111111111101101110100100100;
assign LUT_2[52992] = 32'b11111111111111111111010110001011;
assign LUT_2[52993] = 32'b11111111111111111100001110100100;
assign LUT_2[52994] = 32'b00000000000000000110001111000111;
assign LUT_2[52995] = 32'b00000000000000000011000111100000;
assign LUT_2[52996] = 32'b11111111111111111011110011110011;
assign LUT_2[52997] = 32'b11111111111111111000101100001100;
assign LUT_2[52998] = 32'b00000000000000000010101100101111;
assign LUT_2[52999] = 32'b11111111111111111111100101001000;
assign LUT_2[53000] = 32'b11111111111111111010000111101000;
assign LUT_2[53001] = 32'b11111111111111110111000000000001;
assign LUT_2[53002] = 32'b00000000000000000001000000100100;
assign LUT_2[53003] = 32'b11111111111111111101111000111101;
assign LUT_2[53004] = 32'b11111111111111110110100101010000;
assign LUT_2[53005] = 32'b11111111111111110011011101101001;
assign LUT_2[53006] = 32'b11111111111111111101011110001100;
assign LUT_2[53007] = 32'b11111111111111111010010110100101;
assign LUT_2[53008] = 32'b11111111111111111001111010010101;
assign LUT_2[53009] = 32'b11111111111111110110110010101110;
assign LUT_2[53010] = 32'b00000000000000000000110011010001;
assign LUT_2[53011] = 32'b11111111111111111101101011101010;
assign LUT_2[53012] = 32'b11111111111111110110010111111101;
assign LUT_2[53013] = 32'b11111111111111110011010000010110;
assign LUT_2[53014] = 32'b11111111111111111101010000111001;
assign LUT_2[53015] = 32'b11111111111111111010001001010010;
assign LUT_2[53016] = 32'b11111111111111110100101011110010;
assign LUT_2[53017] = 32'b11111111111111110001100100001011;
assign LUT_2[53018] = 32'b11111111111111111011100100101110;
assign LUT_2[53019] = 32'b11111111111111111000011101000111;
assign LUT_2[53020] = 32'b11111111111111110001001001011010;
assign LUT_2[53021] = 32'b11111111111111101110000001110011;
assign LUT_2[53022] = 32'b11111111111111111000000010010110;
assign LUT_2[53023] = 32'b11111111111111110100111010101111;
assign LUT_2[53024] = 32'b11111111111111111111110001110100;
assign LUT_2[53025] = 32'b11111111111111111100101010001101;
assign LUT_2[53026] = 32'b00000000000000000110101010110000;
assign LUT_2[53027] = 32'b00000000000000000011100011001001;
assign LUT_2[53028] = 32'b11111111111111111100001111011100;
assign LUT_2[53029] = 32'b11111111111111111001000111110101;
assign LUT_2[53030] = 32'b00000000000000000011001000011000;
assign LUT_2[53031] = 32'b00000000000000000000000000110001;
assign LUT_2[53032] = 32'b11111111111111111010100011010001;
assign LUT_2[53033] = 32'b11111111111111110111011011101010;
assign LUT_2[53034] = 32'b00000000000000000001011100001101;
assign LUT_2[53035] = 32'b11111111111111111110010100100110;
assign LUT_2[53036] = 32'b11111111111111110111000000111001;
assign LUT_2[53037] = 32'b11111111111111110011111001010010;
assign LUT_2[53038] = 32'b11111111111111111101111001110101;
assign LUT_2[53039] = 32'b11111111111111111010110010001110;
assign LUT_2[53040] = 32'b11111111111111111010010101111110;
assign LUT_2[53041] = 32'b11111111111111110111001110010111;
assign LUT_2[53042] = 32'b00000000000000000001001110111010;
assign LUT_2[53043] = 32'b11111111111111111110000111010011;
assign LUT_2[53044] = 32'b11111111111111110110110011100110;
assign LUT_2[53045] = 32'b11111111111111110011101011111111;
assign LUT_2[53046] = 32'b11111111111111111101101100100010;
assign LUT_2[53047] = 32'b11111111111111111010100100111011;
assign LUT_2[53048] = 32'b11111111111111110101000111011011;
assign LUT_2[53049] = 32'b11111111111111110001111111110100;
assign LUT_2[53050] = 32'b11111111111111111100000000010111;
assign LUT_2[53051] = 32'b11111111111111111000111000110000;
assign LUT_2[53052] = 32'b11111111111111110001100101000011;
assign LUT_2[53053] = 32'b11111111111111101110011101011100;
assign LUT_2[53054] = 32'b11111111111111111000011101111111;
assign LUT_2[53055] = 32'b11111111111111110101010110011000;
assign LUT_2[53056] = 32'b11111111111111110111011110101110;
assign LUT_2[53057] = 32'b11111111111111110100010111000111;
assign LUT_2[53058] = 32'b11111111111111111110010111101010;
assign LUT_2[53059] = 32'b11111111111111111011010000000011;
assign LUT_2[53060] = 32'b11111111111111110011111100010110;
assign LUT_2[53061] = 32'b11111111111111110000110100101111;
assign LUT_2[53062] = 32'b11111111111111111010110101010010;
assign LUT_2[53063] = 32'b11111111111111110111101101101011;
assign LUT_2[53064] = 32'b11111111111111110010010000001011;
assign LUT_2[53065] = 32'b11111111111111101111001000100100;
assign LUT_2[53066] = 32'b11111111111111111001001001000111;
assign LUT_2[53067] = 32'b11111111111111110110000001100000;
assign LUT_2[53068] = 32'b11111111111111101110101101110011;
assign LUT_2[53069] = 32'b11111111111111101011100110001100;
assign LUT_2[53070] = 32'b11111111111111110101100110101111;
assign LUT_2[53071] = 32'b11111111111111110010011111001000;
assign LUT_2[53072] = 32'b11111111111111110010000010111000;
assign LUT_2[53073] = 32'b11111111111111101110111011010001;
assign LUT_2[53074] = 32'b11111111111111111000111011110100;
assign LUT_2[53075] = 32'b11111111111111110101110100001101;
assign LUT_2[53076] = 32'b11111111111111101110100000100000;
assign LUT_2[53077] = 32'b11111111111111101011011000111001;
assign LUT_2[53078] = 32'b11111111111111110101011001011100;
assign LUT_2[53079] = 32'b11111111111111110010010001110101;
assign LUT_2[53080] = 32'b11111111111111101100110100010101;
assign LUT_2[53081] = 32'b11111111111111101001101100101110;
assign LUT_2[53082] = 32'b11111111111111110011101101010001;
assign LUT_2[53083] = 32'b11111111111111110000100101101010;
assign LUT_2[53084] = 32'b11111111111111101001010001111101;
assign LUT_2[53085] = 32'b11111111111111100110001010010110;
assign LUT_2[53086] = 32'b11111111111111110000001010111001;
assign LUT_2[53087] = 32'b11111111111111101101000011010010;
assign LUT_2[53088] = 32'b11111111111111110111111010010111;
assign LUT_2[53089] = 32'b11111111111111110100110010110000;
assign LUT_2[53090] = 32'b11111111111111111110110011010011;
assign LUT_2[53091] = 32'b11111111111111111011101011101100;
assign LUT_2[53092] = 32'b11111111111111110100010111111111;
assign LUT_2[53093] = 32'b11111111111111110001010000011000;
assign LUT_2[53094] = 32'b11111111111111111011010000111011;
assign LUT_2[53095] = 32'b11111111111111111000001001010100;
assign LUT_2[53096] = 32'b11111111111111110010101011110100;
assign LUT_2[53097] = 32'b11111111111111101111100100001101;
assign LUT_2[53098] = 32'b11111111111111111001100100110000;
assign LUT_2[53099] = 32'b11111111111111110110011101001001;
assign LUT_2[53100] = 32'b11111111111111101111001001011100;
assign LUT_2[53101] = 32'b11111111111111101100000001110101;
assign LUT_2[53102] = 32'b11111111111111110110000010011000;
assign LUT_2[53103] = 32'b11111111111111110010111010110001;
assign LUT_2[53104] = 32'b11111111111111110010011110100001;
assign LUT_2[53105] = 32'b11111111111111101111010110111010;
assign LUT_2[53106] = 32'b11111111111111111001010111011101;
assign LUT_2[53107] = 32'b11111111111111110110001111110110;
assign LUT_2[53108] = 32'b11111111111111101110111100001001;
assign LUT_2[53109] = 32'b11111111111111101011110100100010;
assign LUT_2[53110] = 32'b11111111111111110101110101000101;
assign LUT_2[53111] = 32'b11111111111111110010101101011110;
assign LUT_2[53112] = 32'b11111111111111101101001111111110;
assign LUT_2[53113] = 32'b11111111111111101010001000010111;
assign LUT_2[53114] = 32'b11111111111111110100001000111010;
assign LUT_2[53115] = 32'b11111111111111110001000001010011;
assign LUT_2[53116] = 32'b11111111111111101001101101100110;
assign LUT_2[53117] = 32'b11111111111111100110100101111111;
assign LUT_2[53118] = 32'b11111111111111110000100110100010;
assign LUT_2[53119] = 32'b11111111111111101101011110111011;
assign LUT_2[53120] = 32'b00000000000000000011101010011010;
assign LUT_2[53121] = 32'b00000000000000000000100010110011;
assign LUT_2[53122] = 32'b00000000000000001010100011010110;
assign LUT_2[53123] = 32'b00000000000000000111011011101111;
assign LUT_2[53124] = 32'b00000000000000000000001000000010;
assign LUT_2[53125] = 32'b11111111111111111101000000011011;
assign LUT_2[53126] = 32'b00000000000000000111000000111110;
assign LUT_2[53127] = 32'b00000000000000000011111001010111;
assign LUT_2[53128] = 32'b11111111111111111110011011110111;
assign LUT_2[53129] = 32'b11111111111111111011010100010000;
assign LUT_2[53130] = 32'b00000000000000000101010100110011;
assign LUT_2[53131] = 32'b00000000000000000010001101001100;
assign LUT_2[53132] = 32'b11111111111111111010111001011111;
assign LUT_2[53133] = 32'b11111111111111110111110001111000;
assign LUT_2[53134] = 32'b00000000000000000001110010011011;
assign LUT_2[53135] = 32'b11111111111111111110101010110100;
assign LUT_2[53136] = 32'b11111111111111111110001110100100;
assign LUT_2[53137] = 32'b11111111111111111011000110111101;
assign LUT_2[53138] = 32'b00000000000000000101000111100000;
assign LUT_2[53139] = 32'b00000000000000000001111111111001;
assign LUT_2[53140] = 32'b11111111111111111010101100001100;
assign LUT_2[53141] = 32'b11111111111111110111100100100101;
assign LUT_2[53142] = 32'b00000000000000000001100101001000;
assign LUT_2[53143] = 32'b11111111111111111110011101100001;
assign LUT_2[53144] = 32'b11111111111111111001000000000001;
assign LUT_2[53145] = 32'b11111111111111110101111000011010;
assign LUT_2[53146] = 32'b11111111111111111111111000111101;
assign LUT_2[53147] = 32'b11111111111111111100110001010110;
assign LUT_2[53148] = 32'b11111111111111110101011101101001;
assign LUT_2[53149] = 32'b11111111111111110010010110000010;
assign LUT_2[53150] = 32'b11111111111111111100010110100101;
assign LUT_2[53151] = 32'b11111111111111111001001110111110;
assign LUT_2[53152] = 32'b00000000000000000100000110000011;
assign LUT_2[53153] = 32'b00000000000000000000111110011100;
assign LUT_2[53154] = 32'b00000000000000001010111110111111;
assign LUT_2[53155] = 32'b00000000000000000111110111011000;
assign LUT_2[53156] = 32'b00000000000000000000100011101011;
assign LUT_2[53157] = 32'b11111111111111111101011100000100;
assign LUT_2[53158] = 32'b00000000000000000111011100100111;
assign LUT_2[53159] = 32'b00000000000000000100010101000000;
assign LUT_2[53160] = 32'b11111111111111111110110111100000;
assign LUT_2[53161] = 32'b11111111111111111011101111111001;
assign LUT_2[53162] = 32'b00000000000000000101110000011100;
assign LUT_2[53163] = 32'b00000000000000000010101000110101;
assign LUT_2[53164] = 32'b11111111111111111011010101001000;
assign LUT_2[53165] = 32'b11111111111111111000001101100001;
assign LUT_2[53166] = 32'b00000000000000000010001110000100;
assign LUT_2[53167] = 32'b11111111111111111111000110011101;
assign LUT_2[53168] = 32'b11111111111111111110101010001101;
assign LUT_2[53169] = 32'b11111111111111111011100010100110;
assign LUT_2[53170] = 32'b00000000000000000101100011001001;
assign LUT_2[53171] = 32'b00000000000000000010011011100010;
assign LUT_2[53172] = 32'b11111111111111111011000111110101;
assign LUT_2[53173] = 32'b11111111111111111000000000001110;
assign LUT_2[53174] = 32'b00000000000000000010000000110001;
assign LUT_2[53175] = 32'b11111111111111111110111001001010;
assign LUT_2[53176] = 32'b11111111111111111001011011101010;
assign LUT_2[53177] = 32'b11111111111111110110010100000011;
assign LUT_2[53178] = 32'b00000000000000000000010100100110;
assign LUT_2[53179] = 32'b11111111111111111101001100111111;
assign LUT_2[53180] = 32'b11111111111111110101111001010010;
assign LUT_2[53181] = 32'b11111111111111110010110001101011;
assign LUT_2[53182] = 32'b11111111111111111100110010001110;
assign LUT_2[53183] = 32'b11111111111111111001101010100111;
assign LUT_2[53184] = 32'b11111111111111111011110010111101;
assign LUT_2[53185] = 32'b11111111111111111000101011010110;
assign LUT_2[53186] = 32'b00000000000000000010101011111001;
assign LUT_2[53187] = 32'b11111111111111111111100100010010;
assign LUT_2[53188] = 32'b11111111111111111000010000100101;
assign LUT_2[53189] = 32'b11111111111111110101001000111110;
assign LUT_2[53190] = 32'b11111111111111111111001001100001;
assign LUT_2[53191] = 32'b11111111111111111100000001111010;
assign LUT_2[53192] = 32'b11111111111111110110100100011010;
assign LUT_2[53193] = 32'b11111111111111110011011100110011;
assign LUT_2[53194] = 32'b11111111111111111101011101010110;
assign LUT_2[53195] = 32'b11111111111111111010010101101111;
assign LUT_2[53196] = 32'b11111111111111110011000010000010;
assign LUT_2[53197] = 32'b11111111111111101111111010011011;
assign LUT_2[53198] = 32'b11111111111111111001111010111110;
assign LUT_2[53199] = 32'b11111111111111110110110011010111;
assign LUT_2[53200] = 32'b11111111111111110110010111000111;
assign LUT_2[53201] = 32'b11111111111111110011001111100000;
assign LUT_2[53202] = 32'b11111111111111111101010000000011;
assign LUT_2[53203] = 32'b11111111111111111010001000011100;
assign LUT_2[53204] = 32'b11111111111111110010110100101111;
assign LUT_2[53205] = 32'b11111111111111101111101101001000;
assign LUT_2[53206] = 32'b11111111111111111001101101101011;
assign LUT_2[53207] = 32'b11111111111111110110100110000100;
assign LUT_2[53208] = 32'b11111111111111110001001000100100;
assign LUT_2[53209] = 32'b11111111111111101110000000111101;
assign LUT_2[53210] = 32'b11111111111111111000000001100000;
assign LUT_2[53211] = 32'b11111111111111110100111001111001;
assign LUT_2[53212] = 32'b11111111111111101101100110001100;
assign LUT_2[53213] = 32'b11111111111111101010011110100101;
assign LUT_2[53214] = 32'b11111111111111110100011111001000;
assign LUT_2[53215] = 32'b11111111111111110001010111100001;
assign LUT_2[53216] = 32'b11111111111111111100001110100110;
assign LUT_2[53217] = 32'b11111111111111111001000110111111;
assign LUT_2[53218] = 32'b00000000000000000011000111100010;
assign LUT_2[53219] = 32'b11111111111111111111111111111011;
assign LUT_2[53220] = 32'b11111111111111111000101100001110;
assign LUT_2[53221] = 32'b11111111111111110101100100100111;
assign LUT_2[53222] = 32'b11111111111111111111100101001010;
assign LUT_2[53223] = 32'b11111111111111111100011101100011;
assign LUT_2[53224] = 32'b11111111111111110111000000000011;
assign LUT_2[53225] = 32'b11111111111111110011111000011100;
assign LUT_2[53226] = 32'b11111111111111111101111000111111;
assign LUT_2[53227] = 32'b11111111111111111010110001011000;
assign LUT_2[53228] = 32'b11111111111111110011011101101011;
assign LUT_2[53229] = 32'b11111111111111110000010110000100;
assign LUT_2[53230] = 32'b11111111111111111010010110100111;
assign LUT_2[53231] = 32'b11111111111111110111001111000000;
assign LUT_2[53232] = 32'b11111111111111110110110010110000;
assign LUT_2[53233] = 32'b11111111111111110011101011001001;
assign LUT_2[53234] = 32'b11111111111111111101101011101100;
assign LUT_2[53235] = 32'b11111111111111111010100100000101;
assign LUT_2[53236] = 32'b11111111111111110011010000011000;
assign LUT_2[53237] = 32'b11111111111111110000001000110001;
assign LUT_2[53238] = 32'b11111111111111111010001001010100;
assign LUT_2[53239] = 32'b11111111111111110111000001101101;
assign LUT_2[53240] = 32'b11111111111111110001100100001101;
assign LUT_2[53241] = 32'b11111111111111101110011100100110;
assign LUT_2[53242] = 32'b11111111111111111000011101001001;
assign LUT_2[53243] = 32'b11111111111111110101010101100010;
assign LUT_2[53244] = 32'b11111111111111101110000001110101;
assign LUT_2[53245] = 32'b11111111111111101010111010001110;
assign LUT_2[53246] = 32'b11111111111111110100111010110001;
assign LUT_2[53247] = 32'b11111111111111110001110011001010;
assign LUT_2[53248] = 32'b11111111111111110011000111111101;
assign LUT_2[53249] = 32'b11111111111111110000000000010110;
assign LUT_2[53250] = 32'b11111111111111111010000000111001;
assign LUT_2[53251] = 32'b11111111111111110110111001010010;
assign LUT_2[53252] = 32'b11111111111111101111100101100101;
assign LUT_2[53253] = 32'b11111111111111101100011101111110;
assign LUT_2[53254] = 32'b11111111111111110110011110100001;
assign LUT_2[53255] = 32'b11111111111111110011010110111010;
assign LUT_2[53256] = 32'b11111111111111101101111001011010;
assign LUT_2[53257] = 32'b11111111111111101010110001110011;
assign LUT_2[53258] = 32'b11111111111111110100110010010110;
assign LUT_2[53259] = 32'b11111111111111110001101010101111;
assign LUT_2[53260] = 32'b11111111111111101010010111000010;
assign LUT_2[53261] = 32'b11111111111111100111001111011011;
assign LUT_2[53262] = 32'b11111111111111110001001111111110;
assign LUT_2[53263] = 32'b11111111111111101110001000010111;
assign LUT_2[53264] = 32'b11111111111111101101101100000111;
assign LUT_2[53265] = 32'b11111111111111101010100100100000;
assign LUT_2[53266] = 32'b11111111111111110100100101000011;
assign LUT_2[53267] = 32'b11111111111111110001011101011100;
assign LUT_2[53268] = 32'b11111111111111101010001001101111;
assign LUT_2[53269] = 32'b11111111111111100111000010001000;
assign LUT_2[53270] = 32'b11111111111111110001000010101011;
assign LUT_2[53271] = 32'b11111111111111101101111011000100;
assign LUT_2[53272] = 32'b11111111111111101000011101100100;
assign LUT_2[53273] = 32'b11111111111111100101010101111101;
assign LUT_2[53274] = 32'b11111111111111101111010110100000;
assign LUT_2[53275] = 32'b11111111111111101100001110111001;
assign LUT_2[53276] = 32'b11111111111111100100111011001100;
assign LUT_2[53277] = 32'b11111111111111100001110011100101;
assign LUT_2[53278] = 32'b11111111111111101011110100001000;
assign LUT_2[53279] = 32'b11111111111111101000101100100001;
assign LUT_2[53280] = 32'b11111111111111110011100011100110;
assign LUT_2[53281] = 32'b11111111111111110000011011111111;
assign LUT_2[53282] = 32'b11111111111111111010011100100010;
assign LUT_2[53283] = 32'b11111111111111110111010100111011;
assign LUT_2[53284] = 32'b11111111111111110000000001001110;
assign LUT_2[53285] = 32'b11111111111111101100111001100111;
assign LUT_2[53286] = 32'b11111111111111110110111010001010;
assign LUT_2[53287] = 32'b11111111111111110011110010100011;
assign LUT_2[53288] = 32'b11111111111111101110010101000011;
assign LUT_2[53289] = 32'b11111111111111101011001101011100;
assign LUT_2[53290] = 32'b11111111111111110101001101111111;
assign LUT_2[53291] = 32'b11111111111111110010000110011000;
assign LUT_2[53292] = 32'b11111111111111101010110010101011;
assign LUT_2[53293] = 32'b11111111111111100111101011000100;
assign LUT_2[53294] = 32'b11111111111111110001101011100111;
assign LUT_2[53295] = 32'b11111111111111101110100100000000;
assign LUT_2[53296] = 32'b11111111111111101110000111110000;
assign LUT_2[53297] = 32'b11111111111111101011000000001001;
assign LUT_2[53298] = 32'b11111111111111110101000000101100;
assign LUT_2[53299] = 32'b11111111111111110001111001000101;
assign LUT_2[53300] = 32'b11111111111111101010100101011000;
assign LUT_2[53301] = 32'b11111111111111100111011101110001;
assign LUT_2[53302] = 32'b11111111111111110001011110010100;
assign LUT_2[53303] = 32'b11111111111111101110010110101101;
assign LUT_2[53304] = 32'b11111111111111101000111001001101;
assign LUT_2[53305] = 32'b11111111111111100101110001100110;
assign LUT_2[53306] = 32'b11111111111111101111110010001001;
assign LUT_2[53307] = 32'b11111111111111101100101010100010;
assign LUT_2[53308] = 32'b11111111111111100101010110110101;
assign LUT_2[53309] = 32'b11111111111111100010001111001110;
assign LUT_2[53310] = 32'b11111111111111101100001111110001;
assign LUT_2[53311] = 32'b11111111111111101001001000001010;
assign LUT_2[53312] = 32'b11111111111111101011010000100000;
assign LUT_2[53313] = 32'b11111111111111101000001000111001;
assign LUT_2[53314] = 32'b11111111111111110010001001011100;
assign LUT_2[53315] = 32'b11111111111111101111000001110101;
assign LUT_2[53316] = 32'b11111111111111100111101110001000;
assign LUT_2[53317] = 32'b11111111111111100100100110100001;
assign LUT_2[53318] = 32'b11111111111111101110100111000100;
assign LUT_2[53319] = 32'b11111111111111101011011111011101;
assign LUT_2[53320] = 32'b11111111111111100110000001111101;
assign LUT_2[53321] = 32'b11111111111111100010111010010110;
assign LUT_2[53322] = 32'b11111111111111101100111010111001;
assign LUT_2[53323] = 32'b11111111111111101001110011010010;
assign LUT_2[53324] = 32'b11111111111111100010011111100101;
assign LUT_2[53325] = 32'b11111111111111011111010111111110;
assign LUT_2[53326] = 32'b11111111111111101001011000100001;
assign LUT_2[53327] = 32'b11111111111111100110010000111010;
assign LUT_2[53328] = 32'b11111111111111100101110100101010;
assign LUT_2[53329] = 32'b11111111111111100010101101000011;
assign LUT_2[53330] = 32'b11111111111111101100101101100110;
assign LUT_2[53331] = 32'b11111111111111101001100101111111;
assign LUT_2[53332] = 32'b11111111111111100010010010010010;
assign LUT_2[53333] = 32'b11111111111111011111001010101011;
assign LUT_2[53334] = 32'b11111111111111101001001011001110;
assign LUT_2[53335] = 32'b11111111111111100110000011100111;
assign LUT_2[53336] = 32'b11111111111111100000100110000111;
assign LUT_2[53337] = 32'b11111111111111011101011110100000;
assign LUT_2[53338] = 32'b11111111111111100111011111000011;
assign LUT_2[53339] = 32'b11111111111111100100010111011100;
assign LUT_2[53340] = 32'b11111111111111011101000011101111;
assign LUT_2[53341] = 32'b11111111111111011001111100001000;
assign LUT_2[53342] = 32'b11111111111111100011111100101011;
assign LUT_2[53343] = 32'b11111111111111100000110101000100;
assign LUT_2[53344] = 32'b11111111111111101011101100001001;
assign LUT_2[53345] = 32'b11111111111111101000100100100010;
assign LUT_2[53346] = 32'b11111111111111110010100101000101;
assign LUT_2[53347] = 32'b11111111111111101111011101011110;
assign LUT_2[53348] = 32'b11111111111111101000001001110001;
assign LUT_2[53349] = 32'b11111111111111100101000010001010;
assign LUT_2[53350] = 32'b11111111111111101111000010101101;
assign LUT_2[53351] = 32'b11111111111111101011111011000110;
assign LUT_2[53352] = 32'b11111111111111100110011101100110;
assign LUT_2[53353] = 32'b11111111111111100011010101111111;
assign LUT_2[53354] = 32'b11111111111111101101010110100010;
assign LUT_2[53355] = 32'b11111111111111101010001110111011;
assign LUT_2[53356] = 32'b11111111111111100010111011001110;
assign LUT_2[53357] = 32'b11111111111111011111110011100111;
assign LUT_2[53358] = 32'b11111111111111101001110100001010;
assign LUT_2[53359] = 32'b11111111111111100110101100100011;
assign LUT_2[53360] = 32'b11111111111111100110010000010011;
assign LUT_2[53361] = 32'b11111111111111100011001000101100;
assign LUT_2[53362] = 32'b11111111111111101101001001001111;
assign LUT_2[53363] = 32'b11111111111111101010000001101000;
assign LUT_2[53364] = 32'b11111111111111100010101101111011;
assign LUT_2[53365] = 32'b11111111111111011111100110010100;
assign LUT_2[53366] = 32'b11111111111111101001100110110111;
assign LUT_2[53367] = 32'b11111111111111100110011111010000;
assign LUT_2[53368] = 32'b11111111111111100001000001110000;
assign LUT_2[53369] = 32'b11111111111111011101111010001001;
assign LUT_2[53370] = 32'b11111111111111100111111010101100;
assign LUT_2[53371] = 32'b11111111111111100100110011000101;
assign LUT_2[53372] = 32'b11111111111111011101011111011000;
assign LUT_2[53373] = 32'b11111111111111011010010111110001;
assign LUT_2[53374] = 32'b11111111111111100100011000010100;
assign LUT_2[53375] = 32'b11111111111111100001010000101101;
assign LUT_2[53376] = 32'b11111111111111110111011100001100;
assign LUT_2[53377] = 32'b11111111111111110100010100100101;
assign LUT_2[53378] = 32'b11111111111111111110010101001000;
assign LUT_2[53379] = 32'b11111111111111111011001101100001;
assign LUT_2[53380] = 32'b11111111111111110011111001110100;
assign LUT_2[53381] = 32'b11111111111111110000110010001101;
assign LUT_2[53382] = 32'b11111111111111111010110010110000;
assign LUT_2[53383] = 32'b11111111111111110111101011001001;
assign LUT_2[53384] = 32'b11111111111111110010001101101001;
assign LUT_2[53385] = 32'b11111111111111101111000110000010;
assign LUT_2[53386] = 32'b11111111111111111001000110100101;
assign LUT_2[53387] = 32'b11111111111111110101111110111110;
assign LUT_2[53388] = 32'b11111111111111101110101011010001;
assign LUT_2[53389] = 32'b11111111111111101011100011101010;
assign LUT_2[53390] = 32'b11111111111111110101100100001101;
assign LUT_2[53391] = 32'b11111111111111110010011100100110;
assign LUT_2[53392] = 32'b11111111111111110010000000010110;
assign LUT_2[53393] = 32'b11111111111111101110111000101111;
assign LUT_2[53394] = 32'b11111111111111111000111001010010;
assign LUT_2[53395] = 32'b11111111111111110101110001101011;
assign LUT_2[53396] = 32'b11111111111111101110011101111110;
assign LUT_2[53397] = 32'b11111111111111101011010110010111;
assign LUT_2[53398] = 32'b11111111111111110101010110111010;
assign LUT_2[53399] = 32'b11111111111111110010001111010011;
assign LUT_2[53400] = 32'b11111111111111101100110001110011;
assign LUT_2[53401] = 32'b11111111111111101001101010001100;
assign LUT_2[53402] = 32'b11111111111111110011101010101111;
assign LUT_2[53403] = 32'b11111111111111110000100011001000;
assign LUT_2[53404] = 32'b11111111111111101001001111011011;
assign LUT_2[53405] = 32'b11111111111111100110000111110100;
assign LUT_2[53406] = 32'b11111111111111110000001000010111;
assign LUT_2[53407] = 32'b11111111111111101101000000110000;
assign LUT_2[53408] = 32'b11111111111111110111110111110101;
assign LUT_2[53409] = 32'b11111111111111110100110000001110;
assign LUT_2[53410] = 32'b11111111111111111110110000110001;
assign LUT_2[53411] = 32'b11111111111111111011101001001010;
assign LUT_2[53412] = 32'b11111111111111110100010101011101;
assign LUT_2[53413] = 32'b11111111111111110001001101110110;
assign LUT_2[53414] = 32'b11111111111111111011001110011001;
assign LUT_2[53415] = 32'b11111111111111111000000110110010;
assign LUT_2[53416] = 32'b11111111111111110010101001010010;
assign LUT_2[53417] = 32'b11111111111111101111100001101011;
assign LUT_2[53418] = 32'b11111111111111111001100010001110;
assign LUT_2[53419] = 32'b11111111111111110110011010100111;
assign LUT_2[53420] = 32'b11111111111111101111000110111010;
assign LUT_2[53421] = 32'b11111111111111101011111111010011;
assign LUT_2[53422] = 32'b11111111111111110101111111110110;
assign LUT_2[53423] = 32'b11111111111111110010111000001111;
assign LUT_2[53424] = 32'b11111111111111110010011011111111;
assign LUT_2[53425] = 32'b11111111111111101111010100011000;
assign LUT_2[53426] = 32'b11111111111111111001010100111011;
assign LUT_2[53427] = 32'b11111111111111110110001101010100;
assign LUT_2[53428] = 32'b11111111111111101110111001100111;
assign LUT_2[53429] = 32'b11111111111111101011110010000000;
assign LUT_2[53430] = 32'b11111111111111110101110010100011;
assign LUT_2[53431] = 32'b11111111111111110010101010111100;
assign LUT_2[53432] = 32'b11111111111111101101001101011100;
assign LUT_2[53433] = 32'b11111111111111101010000101110101;
assign LUT_2[53434] = 32'b11111111111111110100000110011000;
assign LUT_2[53435] = 32'b11111111111111110000111110110001;
assign LUT_2[53436] = 32'b11111111111111101001101011000100;
assign LUT_2[53437] = 32'b11111111111111100110100011011101;
assign LUT_2[53438] = 32'b11111111111111110000100100000000;
assign LUT_2[53439] = 32'b11111111111111101101011100011001;
assign LUT_2[53440] = 32'b11111111111111101111100100101111;
assign LUT_2[53441] = 32'b11111111111111101100011101001000;
assign LUT_2[53442] = 32'b11111111111111110110011101101011;
assign LUT_2[53443] = 32'b11111111111111110011010110000100;
assign LUT_2[53444] = 32'b11111111111111101100000010010111;
assign LUT_2[53445] = 32'b11111111111111101000111010110000;
assign LUT_2[53446] = 32'b11111111111111110010111011010011;
assign LUT_2[53447] = 32'b11111111111111101111110011101100;
assign LUT_2[53448] = 32'b11111111111111101010010110001100;
assign LUT_2[53449] = 32'b11111111111111100111001110100101;
assign LUT_2[53450] = 32'b11111111111111110001001111001000;
assign LUT_2[53451] = 32'b11111111111111101110000111100001;
assign LUT_2[53452] = 32'b11111111111111100110110011110100;
assign LUT_2[53453] = 32'b11111111111111100011101100001101;
assign LUT_2[53454] = 32'b11111111111111101101101100110000;
assign LUT_2[53455] = 32'b11111111111111101010100101001001;
assign LUT_2[53456] = 32'b11111111111111101010001000111001;
assign LUT_2[53457] = 32'b11111111111111100111000001010010;
assign LUT_2[53458] = 32'b11111111111111110001000001110101;
assign LUT_2[53459] = 32'b11111111111111101101111010001110;
assign LUT_2[53460] = 32'b11111111111111100110100110100001;
assign LUT_2[53461] = 32'b11111111111111100011011110111010;
assign LUT_2[53462] = 32'b11111111111111101101011111011101;
assign LUT_2[53463] = 32'b11111111111111101010010111110110;
assign LUT_2[53464] = 32'b11111111111111100100111010010110;
assign LUT_2[53465] = 32'b11111111111111100001110010101111;
assign LUT_2[53466] = 32'b11111111111111101011110011010010;
assign LUT_2[53467] = 32'b11111111111111101000101011101011;
assign LUT_2[53468] = 32'b11111111111111100001010111111110;
assign LUT_2[53469] = 32'b11111111111111011110010000010111;
assign LUT_2[53470] = 32'b11111111111111101000010000111010;
assign LUT_2[53471] = 32'b11111111111111100101001001010011;
assign LUT_2[53472] = 32'b11111111111111110000000000011000;
assign LUT_2[53473] = 32'b11111111111111101100111000110001;
assign LUT_2[53474] = 32'b11111111111111110110111001010100;
assign LUT_2[53475] = 32'b11111111111111110011110001101101;
assign LUT_2[53476] = 32'b11111111111111101100011110000000;
assign LUT_2[53477] = 32'b11111111111111101001010110011001;
assign LUT_2[53478] = 32'b11111111111111110011010110111100;
assign LUT_2[53479] = 32'b11111111111111110000001111010101;
assign LUT_2[53480] = 32'b11111111111111101010110001110101;
assign LUT_2[53481] = 32'b11111111111111100111101010001110;
assign LUT_2[53482] = 32'b11111111111111110001101010110001;
assign LUT_2[53483] = 32'b11111111111111101110100011001010;
assign LUT_2[53484] = 32'b11111111111111100111001111011101;
assign LUT_2[53485] = 32'b11111111111111100100000111110110;
assign LUT_2[53486] = 32'b11111111111111101110001000011001;
assign LUT_2[53487] = 32'b11111111111111101011000000110010;
assign LUT_2[53488] = 32'b11111111111111101010100100100010;
assign LUT_2[53489] = 32'b11111111111111100111011100111011;
assign LUT_2[53490] = 32'b11111111111111110001011101011110;
assign LUT_2[53491] = 32'b11111111111111101110010101110111;
assign LUT_2[53492] = 32'b11111111111111100111000010001010;
assign LUT_2[53493] = 32'b11111111111111100011111010100011;
assign LUT_2[53494] = 32'b11111111111111101101111011000110;
assign LUT_2[53495] = 32'b11111111111111101010110011011111;
assign LUT_2[53496] = 32'b11111111111111100101010101111111;
assign LUT_2[53497] = 32'b11111111111111100010001110011000;
assign LUT_2[53498] = 32'b11111111111111101100001110111011;
assign LUT_2[53499] = 32'b11111111111111101001000111010100;
assign LUT_2[53500] = 32'b11111111111111100001110011100111;
assign LUT_2[53501] = 32'b11111111111111011110101100000000;
assign LUT_2[53502] = 32'b11111111111111101000101100100011;
assign LUT_2[53503] = 32'b11111111111111100101100100111100;
assign LUT_2[53504] = 32'b11111111111111110111000110100011;
assign LUT_2[53505] = 32'b11111111111111110011111110111100;
assign LUT_2[53506] = 32'b11111111111111111101111111011111;
assign LUT_2[53507] = 32'b11111111111111111010110111111000;
assign LUT_2[53508] = 32'b11111111111111110011100100001011;
assign LUT_2[53509] = 32'b11111111111111110000011100100100;
assign LUT_2[53510] = 32'b11111111111111111010011101000111;
assign LUT_2[53511] = 32'b11111111111111110111010101100000;
assign LUT_2[53512] = 32'b11111111111111110001111000000000;
assign LUT_2[53513] = 32'b11111111111111101110110000011001;
assign LUT_2[53514] = 32'b11111111111111111000110000111100;
assign LUT_2[53515] = 32'b11111111111111110101101001010101;
assign LUT_2[53516] = 32'b11111111111111101110010101101000;
assign LUT_2[53517] = 32'b11111111111111101011001110000001;
assign LUT_2[53518] = 32'b11111111111111110101001110100100;
assign LUT_2[53519] = 32'b11111111111111110010000110111101;
assign LUT_2[53520] = 32'b11111111111111110001101010101101;
assign LUT_2[53521] = 32'b11111111111111101110100011000110;
assign LUT_2[53522] = 32'b11111111111111111000100011101001;
assign LUT_2[53523] = 32'b11111111111111110101011100000010;
assign LUT_2[53524] = 32'b11111111111111101110001000010101;
assign LUT_2[53525] = 32'b11111111111111101011000000101110;
assign LUT_2[53526] = 32'b11111111111111110101000001010001;
assign LUT_2[53527] = 32'b11111111111111110001111001101010;
assign LUT_2[53528] = 32'b11111111111111101100011100001010;
assign LUT_2[53529] = 32'b11111111111111101001010100100011;
assign LUT_2[53530] = 32'b11111111111111110011010101000110;
assign LUT_2[53531] = 32'b11111111111111110000001101011111;
assign LUT_2[53532] = 32'b11111111111111101000111001110010;
assign LUT_2[53533] = 32'b11111111111111100101110010001011;
assign LUT_2[53534] = 32'b11111111111111101111110010101110;
assign LUT_2[53535] = 32'b11111111111111101100101011000111;
assign LUT_2[53536] = 32'b11111111111111110111100010001100;
assign LUT_2[53537] = 32'b11111111111111110100011010100101;
assign LUT_2[53538] = 32'b11111111111111111110011011001000;
assign LUT_2[53539] = 32'b11111111111111111011010011100001;
assign LUT_2[53540] = 32'b11111111111111110011111111110100;
assign LUT_2[53541] = 32'b11111111111111110000111000001101;
assign LUT_2[53542] = 32'b11111111111111111010111000110000;
assign LUT_2[53543] = 32'b11111111111111110111110001001001;
assign LUT_2[53544] = 32'b11111111111111110010010011101001;
assign LUT_2[53545] = 32'b11111111111111101111001100000010;
assign LUT_2[53546] = 32'b11111111111111111001001100100101;
assign LUT_2[53547] = 32'b11111111111111110110000100111110;
assign LUT_2[53548] = 32'b11111111111111101110110001010001;
assign LUT_2[53549] = 32'b11111111111111101011101001101010;
assign LUT_2[53550] = 32'b11111111111111110101101010001101;
assign LUT_2[53551] = 32'b11111111111111110010100010100110;
assign LUT_2[53552] = 32'b11111111111111110010000110010110;
assign LUT_2[53553] = 32'b11111111111111101110111110101111;
assign LUT_2[53554] = 32'b11111111111111111000111111010010;
assign LUT_2[53555] = 32'b11111111111111110101110111101011;
assign LUT_2[53556] = 32'b11111111111111101110100011111110;
assign LUT_2[53557] = 32'b11111111111111101011011100010111;
assign LUT_2[53558] = 32'b11111111111111110101011100111010;
assign LUT_2[53559] = 32'b11111111111111110010010101010011;
assign LUT_2[53560] = 32'b11111111111111101100110111110011;
assign LUT_2[53561] = 32'b11111111111111101001110000001100;
assign LUT_2[53562] = 32'b11111111111111110011110000101111;
assign LUT_2[53563] = 32'b11111111111111110000101001001000;
assign LUT_2[53564] = 32'b11111111111111101001010101011011;
assign LUT_2[53565] = 32'b11111111111111100110001101110100;
assign LUT_2[53566] = 32'b11111111111111110000001110010111;
assign LUT_2[53567] = 32'b11111111111111101101000110110000;
assign LUT_2[53568] = 32'b11111111111111101111001111000110;
assign LUT_2[53569] = 32'b11111111111111101100000111011111;
assign LUT_2[53570] = 32'b11111111111111110110001000000010;
assign LUT_2[53571] = 32'b11111111111111110011000000011011;
assign LUT_2[53572] = 32'b11111111111111101011101100101110;
assign LUT_2[53573] = 32'b11111111111111101000100101000111;
assign LUT_2[53574] = 32'b11111111111111110010100101101010;
assign LUT_2[53575] = 32'b11111111111111101111011110000011;
assign LUT_2[53576] = 32'b11111111111111101010000000100011;
assign LUT_2[53577] = 32'b11111111111111100110111000111100;
assign LUT_2[53578] = 32'b11111111111111110000111001011111;
assign LUT_2[53579] = 32'b11111111111111101101110001111000;
assign LUT_2[53580] = 32'b11111111111111100110011110001011;
assign LUT_2[53581] = 32'b11111111111111100011010110100100;
assign LUT_2[53582] = 32'b11111111111111101101010111000111;
assign LUT_2[53583] = 32'b11111111111111101010001111100000;
assign LUT_2[53584] = 32'b11111111111111101001110011010000;
assign LUT_2[53585] = 32'b11111111111111100110101011101001;
assign LUT_2[53586] = 32'b11111111111111110000101100001100;
assign LUT_2[53587] = 32'b11111111111111101101100100100101;
assign LUT_2[53588] = 32'b11111111111111100110010000111000;
assign LUT_2[53589] = 32'b11111111111111100011001001010001;
assign LUT_2[53590] = 32'b11111111111111101101001001110100;
assign LUT_2[53591] = 32'b11111111111111101010000010001101;
assign LUT_2[53592] = 32'b11111111111111100100100100101101;
assign LUT_2[53593] = 32'b11111111111111100001011101000110;
assign LUT_2[53594] = 32'b11111111111111101011011101101001;
assign LUT_2[53595] = 32'b11111111111111101000010110000010;
assign LUT_2[53596] = 32'b11111111111111100001000010010101;
assign LUT_2[53597] = 32'b11111111111111011101111010101110;
assign LUT_2[53598] = 32'b11111111111111100111111011010001;
assign LUT_2[53599] = 32'b11111111111111100100110011101010;
assign LUT_2[53600] = 32'b11111111111111101111101010101111;
assign LUT_2[53601] = 32'b11111111111111101100100011001000;
assign LUT_2[53602] = 32'b11111111111111110110100011101011;
assign LUT_2[53603] = 32'b11111111111111110011011100000100;
assign LUT_2[53604] = 32'b11111111111111101100001000010111;
assign LUT_2[53605] = 32'b11111111111111101001000000110000;
assign LUT_2[53606] = 32'b11111111111111110011000001010011;
assign LUT_2[53607] = 32'b11111111111111101111111001101100;
assign LUT_2[53608] = 32'b11111111111111101010011100001100;
assign LUT_2[53609] = 32'b11111111111111100111010100100101;
assign LUT_2[53610] = 32'b11111111111111110001010101001000;
assign LUT_2[53611] = 32'b11111111111111101110001101100001;
assign LUT_2[53612] = 32'b11111111111111100110111001110100;
assign LUT_2[53613] = 32'b11111111111111100011110010001101;
assign LUT_2[53614] = 32'b11111111111111101101110010110000;
assign LUT_2[53615] = 32'b11111111111111101010101011001001;
assign LUT_2[53616] = 32'b11111111111111101010001110111001;
assign LUT_2[53617] = 32'b11111111111111100111000111010010;
assign LUT_2[53618] = 32'b11111111111111110001000111110101;
assign LUT_2[53619] = 32'b11111111111111101110000000001110;
assign LUT_2[53620] = 32'b11111111111111100110101100100001;
assign LUT_2[53621] = 32'b11111111111111100011100100111010;
assign LUT_2[53622] = 32'b11111111111111101101100101011101;
assign LUT_2[53623] = 32'b11111111111111101010011101110110;
assign LUT_2[53624] = 32'b11111111111111100101000000010110;
assign LUT_2[53625] = 32'b11111111111111100001111000101111;
assign LUT_2[53626] = 32'b11111111111111101011111001010010;
assign LUT_2[53627] = 32'b11111111111111101000110001101011;
assign LUT_2[53628] = 32'b11111111111111100001011101111110;
assign LUT_2[53629] = 32'b11111111111111011110010110010111;
assign LUT_2[53630] = 32'b11111111111111101000010110111010;
assign LUT_2[53631] = 32'b11111111111111100101001111010011;
assign LUT_2[53632] = 32'b11111111111111111011011010110010;
assign LUT_2[53633] = 32'b11111111111111111000010011001011;
assign LUT_2[53634] = 32'b00000000000000000010010011101110;
assign LUT_2[53635] = 32'b11111111111111111111001100000111;
assign LUT_2[53636] = 32'b11111111111111110111111000011010;
assign LUT_2[53637] = 32'b11111111111111110100110000110011;
assign LUT_2[53638] = 32'b11111111111111111110110001010110;
assign LUT_2[53639] = 32'b11111111111111111011101001101111;
assign LUT_2[53640] = 32'b11111111111111110110001100001111;
assign LUT_2[53641] = 32'b11111111111111110011000100101000;
assign LUT_2[53642] = 32'b11111111111111111101000101001011;
assign LUT_2[53643] = 32'b11111111111111111001111101100100;
assign LUT_2[53644] = 32'b11111111111111110010101001110111;
assign LUT_2[53645] = 32'b11111111111111101111100010010000;
assign LUT_2[53646] = 32'b11111111111111111001100010110011;
assign LUT_2[53647] = 32'b11111111111111110110011011001100;
assign LUT_2[53648] = 32'b11111111111111110101111110111100;
assign LUT_2[53649] = 32'b11111111111111110010110111010101;
assign LUT_2[53650] = 32'b11111111111111111100110111111000;
assign LUT_2[53651] = 32'b11111111111111111001110000010001;
assign LUT_2[53652] = 32'b11111111111111110010011100100100;
assign LUT_2[53653] = 32'b11111111111111101111010100111101;
assign LUT_2[53654] = 32'b11111111111111111001010101100000;
assign LUT_2[53655] = 32'b11111111111111110110001101111001;
assign LUT_2[53656] = 32'b11111111111111110000110000011001;
assign LUT_2[53657] = 32'b11111111111111101101101000110010;
assign LUT_2[53658] = 32'b11111111111111110111101001010101;
assign LUT_2[53659] = 32'b11111111111111110100100001101110;
assign LUT_2[53660] = 32'b11111111111111101101001110000001;
assign LUT_2[53661] = 32'b11111111111111101010000110011010;
assign LUT_2[53662] = 32'b11111111111111110100000110111101;
assign LUT_2[53663] = 32'b11111111111111110000111111010110;
assign LUT_2[53664] = 32'b11111111111111111011110110011011;
assign LUT_2[53665] = 32'b11111111111111111000101110110100;
assign LUT_2[53666] = 32'b00000000000000000010101111010111;
assign LUT_2[53667] = 32'b11111111111111111111100111110000;
assign LUT_2[53668] = 32'b11111111111111111000010100000011;
assign LUT_2[53669] = 32'b11111111111111110101001100011100;
assign LUT_2[53670] = 32'b11111111111111111111001100111111;
assign LUT_2[53671] = 32'b11111111111111111100000101011000;
assign LUT_2[53672] = 32'b11111111111111110110100111111000;
assign LUT_2[53673] = 32'b11111111111111110011100000010001;
assign LUT_2[53674] = 32'b11111111111111111101100000110100;
assign LUT_2[53675] = 32'b11111111111111111010011001001101;
assign LUT_2[53676] = 32'b11111111111111110011000101100000;
assign LUT_2[53677] = 32'b11111111111111101111111101111001;
assign LUT_2[53678] = 32'b11111111111111111001111110011100;
assign LUT_2[53679] = 32'b11111111111111110110110110110101;
assign LUT_2[53680] = 32'b11111111111111110110011010100101;
assign LUT_2[53681] = 32'b11111111111111110011010010111110;
assign LUT_2[53682] = 32'b11111111111111111101010011100001;
assign LUT_2[53683] = 32'b11111111111111111010001011111010;
assign LUT_2[53684] = 32'b11111111111111110010111000001101;
assign LUT_2[53685] = 32'b11111111111111101111110000100110;
assign LUT_2[53686] = 32'b11111111111111111001110001001001;
assign LUT_2[53687] = 32'b11111111111111110110101001100010;
assign LUT_2[53688] = 32'b11111111111111110001001100000010;
assign LUT_2[53689] = 32'b11111111111111101110000100011011;
assign LUT_2[53690] = 32'b11111111111111111000000100111110;
assign LUT_2[53691] = 32'b11111111111111110100111101010111;
assign LUT_2[53692] = 32'b11111111111111101101101001101010;
assign LUT_2[53693] = 32'b11111111111111101010100010000011;
assign LUT_2[53694] = 32'b11111111111111110100100010100110;
assign LUT_2[53695] = 32'b11111111111111110001011010111111;
assign LUT_2[53696] = 32'b11111111111111110011100011010101;
assign LUT_2[53697] = 32'b11111111111111110000011011101110;
assign LUT_2[53698] = 32'b11111111111111111010011100010001;
assign LUT_2[53699] = 32'b11111111111111110111010100101010;
assign LUT_2[53700] = 32'b11111111111111110000000000111101;
assign LUT_2[53701] = 32'b11111111111111101100111001010110;
assign LUT_2[53702] = 32'b11111111111111110110111001111001;
assign LUT_2[53703] = 32'b11111111111111110011110010010010;
assign LUT_2[53704] = 32'b11111111111111101110010100110010;
assign LUT_2[53705] = 32'b11111111111111101011001101001011;
assign LUT_2[53706] = 32'b11111111111111110101001101101110;
assign LUT_2[53707] = 32'b11111111111111110010000110000111;
assign LUT_2[53708] = 32'b11111111111111101010110010011010;
assign LUT_2[53709] = 32'b11111111111111100111101010110011;
assign LUT_2[53710] = 32'b11111111111111110001101011010110;
assign LUT_2[53711] = 32'b11111111111111101110100011101111;
assign LUT_2[53712] = 32'b11111111111111101110000111011111;
assign LUT_2[53713] = 32'b11111111111111101010111111111000;
assign LUT_2[53714] = 32'b11111111111111110101000000011011;
assign LUT_2[53715] = 32'b11111111111111110001111000110100;
assign LUT_2[53716] = 32'b11111111111111101010100101000111;
assign LUT_2[53717] = 32'b11111111111111100111011101100000;
assign LUT_2[53718] = 32'b11111111111111110001011110000011;
assign LUT_2[53719] = 32'b11111111111111101110010110011100;
assign LUT_2[53720] = 32'b11111111111111101000111000111100;
assign LUT_2[53721] = 32'b11111111111111100101110001010101;
assign LUT_2[53722] = 32'b11111111111111101111110001111000;
assign LUT_2[53723] = 32'b11111111111111101100101010010001;
assign LUT_2[53724] = 32'b11111111111111100101010110100100;
assign LUT_2[53725] = 32'b11111111111111100010001110111101;
assign LUT_2[53726] = 32'b11111111111111101100001111100000;
assign LUT_2[53727] = 32'b11111111111111101001000111111001;
assign LUT_2[53728] = 32'b11111111111111110011111110111110;
assign LUT_2[53729] = 32'b11111111111111110000110111010111;
assign LUT_2[53730] = 32'b11111111111111111010110111111010;
assign LUT_2[53731] = 32'b11111111111111110111110000010011;
assign LUT_2[53732] = 32'b11111111111111110000011100100110;
assign LUT_2[53733] = 32'b11111111111111101101010100111111;
assign LUT_2[53734] = 32'b11111111111111110111010101100010;
assign LUT_2[53735] = 32'b11111111111111110100001101111011;
assign LUT_2[53736] = 32'b11111111111111101110110000011011;
assign LUT_2[53737] = 32'b11111111111111101011101000110100;
assign LUT_2[53738] = 32'b11111111111111110101101001010111;
assign LUT_2[53739] = 32'b11111111111111110010100001110000;
assign LUT_2[53740] = 32'b11111111111111101011001110000011;
assign LUT_2[53741] = 32'b11111111111111101000000110011100;
assign LUT_2[53742] = 32'b11111111111111110010000110111111;
assign LUT_2[53743] = 32'b11111111111111101110111111011000;
assign LUT_2[53744] = 32'b11111111111111101110100011001000;
assign LUT_2[53745] = 32'b11111111111111101011011011100001;
assign LUT_2[53746] = 32'b11111111111111110101011100000100;
assign LUT_2[53747] = 32'b11111111111111110010010100011101;
assign LUT_2[53748] = 32'b11111111111111101011000000110000;
assign LUT_2[53749] = 32'b11111111111111100111111001001001;
assign LUT_2[53750] = 32'b11111111111111110001111001101100;
assign LUT_2[53751] = 32'b11111111111111101110110010000101;
assign LUT_2[53752] = 32'b11111111111111101001010100100101;
assign LUT_2[53753] = 32'b11111111111111100110001100111110;
assign LUT_2[53754] = 32'b11111111111111110000001101100001;
assign LUT_2[53755] = 32'b11111111111111101101000101111010;
assign LUT_2[53756] = 32'b11111111111111100101110010001101;
assign LUT_2[53757] = 32'b11111111111111100010101010100110;
assign LUT_2[53758] = 32'b11111111111111101100101011001001;
assign LUT_2[53759] = 32'b11111111111111101001100011100010;
assign LUT_2[53760] = 32'b11111111111111110111111001101111;
assign LUT_2[53761] = 32'b11111111111111110100110010001000;
assign LUT_2[53762] = 32'b11111111111111111110110010101011;
assign LUT_2[53763] = 32'b11111111111111111011101011000100;
assign LUT_2[53764] = 32'b11111111111111110100010111010111;
assign LUT_2[53765] = 32'b11111111111111110001001111110000;
assign LUT_2[53766] = 32'b11111111111111111011010000010011;
assign LUT_2[53767] = 32'b11111111111111111000001000101100;
assign LUT_2[53768] = 32'b11111111111111110010101011001100;
assign LUT_2[53769] = 32'b11111111111111101111100011100101;
assign LUT_2[53770] = 32'b11111111111111111001100100001000;
assign LUT_2[53771] = 32'b11111111111111110110011100100001;
assign LUT_2[53772] = 32'b11111111111111101111001000110100;
assign LUT_2[53773] = 32'b11111111111111101100000001001101;
assign LUT_2[53774] = 32'b11111111111111110110000001110000;
assign LUT_2[53775] = 32'b11111111111111110010111010001001;
assign LUT_2[53776] = 32'b11111111111111110010011101111001;
assign LUT_2[53777] = 32'b11111111111111101111010110010010;
assign LUT_2[53778] = 32'b11111111111111111001010110110101;
assign LUT_2[53779] = 32'b11111111111111110110001111001110;
assign LUT_2[53780] = 32'b11111111111111101110111011100001;
assign LUT_2[53781] = 32'b11111111111111101011110011111010;
assign LUT_2[53782] = 32'b11111111111111110101110100011101;
assign LUT_2[53783] = 32'b11111111111111110010101100110110;
assign LUT_2[53784] = 32'b11111111111111101101001111010110;
assign LUT_2[53785] = 32'b11111111111111101010000111101111;
assign LUT_2[53786] = 32'b11111111111111110100001000010010;
assign LUT_2[53787] = 32'b11111111111111110001000000101011;
assign LUT_2[53788] = 32'b11111111111111101001101100111110;
assign LUT_2[53789] = 32'b11111111111111100110100101010111;
assign LUT_2[53790] = 32'b11111111111111110000100101111010;
assign LUT_2[53791] = 32'b11111111111111101101011110010011;
assign LUT_2[53792] = 32'b11111111111111111000010101011000;
assign LUT_2[53793] = 32'b11111111111111110101001101110001;
assign LUT_2[53794] = 32'b11111111111111111111001110010100;
assign LUT_2[53795] = 32'b11111111111111111100000110101101;
assign LUT_2[53796] = 32'b11111111111111110100110011000000;
assign LUT_2[53797] = 32'b11111111111111110001101011011001;
assign LUT_2[53798] = 32'b11111111111111111011101011111100;
assign LUT_2[53799] = 32'b11111111111111111000100100010101;
assign LUT_2[53800] = 32'b11111111111111110011000110110101;
assign LUT_2[53801] = 32'b11111111111111101111111111001110;
assign LUT_2[53802] = 32'b11111111111111111001111111110001;
assign LUT_2[53803] = 32'b11111111111111110110111000001010;
assign LUT_2[53804] = 32'b11111111111111101111100100011101;
assign LUT_2[53805] = 32'b11111111111111101100011100110110;
assign LUT_2[53806] = 32'b11111111111111110110011101011001;
assign LUT_2[53807] = 32'b11111111111111110011010101110010;
assign LUT_2[53808] = 32'b11111111111111110010111001100010;
assign LUT_2[53809] = 32'b11111111111111101111110001111011;
assign LUT_2[53810] = 32'b11111111111111111001110010011110;
assign LUT_2[53811] = 32'b11111111111111110110101010110111;
assign LUT_2[53812] = 32'b11111111111111101111010111001010;
assign LUT_2[53813] = 32'b11111111111111101100001111100011;
assign LUT_2[53814] = 32'b11111111111111110110010000000110;
assign LUT_2[53815] = 32'b11111111111111110011001000011111;
assign LUT_2[53816] = 32'b11111111111111101101101010111111;
assign LUT_2[53817] = 32'b11111111111111101010100011011000;
assign LUT_2[53818] = 32'b11111111111111110100100011111011;
assign LUT_2[53819] = 32'b11111111111111110001011100010100;
assign LUT_2[53820] = 32'b11111111111111101010001000100111;
assign LUT_2[53821] = 32'b11111111111111100111000001000000;
assign LUT_2[53822] = 32'b11111111111111110001000001100011;
assign LUT_2[53823] = 32'b11111111111111101101111001111100;
assign LUT_2[53824] = 32'b11111111111111110000000010010010;
assign LUT_2[53825] = 32'b11111111111111101100111010101011;
assign LUT_2[53826] = 32'b11111111111111110110111011001110;
assign LUT_2[53827] = 32'b11111111111111110011110011100111;
assign LUT_2[53828] = 32'b11111111111111101100011111111010;
assign LUT_2[53829] = 32'b11111111111111101001011000010011;
assign LUT_2[53830] = 32'b11111111111111110011011000110110;
assign LUT_2[53831] = 32'b11111111111111110000010001001111;
assign LUT_2[53832] = 32'b11111111111111101010110011101111;
assign LUT_2[53833] = 32'b11111111111111100111101100001000;
assign LUT_2[53834] = 32'b11111111111111110001101100101011;
assign LUT_2[53835] = 32'b11111111111111101110100101000100;
assign LUT_2[53836] = 32'b11111111111111100111010001010111;
assign LUT_2[53837] = 32'b11111111111111100100001001110000;
assign LUT_2[53838] = 32'b11111111111111101110001010010011;
assign LUT_2[53839] = 32'b11111111111111101011000010101100;
assign LUT_2[53840] = 32'b11111111111111101010100110011100;
assign LUT_2[53841] = 32'b11111111111111100111011110110101;
assign LUT_2[53842] = 32'b11111111111111110001011111011000;
assign LUT_2[53843] = 32'b11111111111111101110010111110001;
assign LUT_2[53844] = 32'b11111111111111100111000100000100;
assign LUT_2[53845] = 32'b11111111111111100011111100011101;
assign LUT_2[53846] = 32'b11111111111111101101111101000000;
assign LUT_2[53847] = 32'b11111111111111101010110101011001;
assign LUT_2[53848] = 32'b11111111111111100101010111111001;
assign LUT_2[53849] = 32'b11111111111111100010010000010010;
assign LUT_2[53850] = 32'b11111111111111101100010000110101;
assign LUT_2[53851] = 32'b11111111111111101001001001001110;
assign LUT_2[53852] = 32'b11111111111111100001110101100001;
assign LUT_2[53853] = 32'b11111111111111011110101101111010;
assign LUT_2[53854] = 32'b11111111111111101000101110011101;
assign LUT_2[53855] = 32'b11111111111111100101100110110110;
assign LUT_2[53856] = 32'b11111111111111110000011101111011;
assign LUT_2[53857] = 32'b11111111111111101101010110010100;
assign LUT_2[53858] = 32'b11111111111111110111010110110111;
assign LUT_2[53859] = 32'b11111111111111110100001111010000;
assign LUT_2[53860] = 32'b11111111111111101100111011100011;
assign LUT_2[53861] = 32'b11111111111111101001110011111100;
assign LUT_2[53862] = 32'b11111111111111110011110100011111;
assign LUT_2[53863] = 32'b11111111111111110000101100111000;
assign LUT_2[53864] = 32'b11111111111111101011001111011000;
assign LUT_2[53865] = 32'b11111111111111101000000111110001;
assign LUT_2[53866] = 32'b11111111111111110010001000010100;
assign LUT_2[53867] = 32'b11111111111111101111000000101101;
assign LUT_2[53868] = 32'b11111111111111100111101101000000;
assign LUT_2[53869] = 32'b11111111111111100100100101011001;
assign LUT_2[53870] = 32'b11111111111111101110100101111100;
assign LUT_2[53871] = 32'b11111111111111101011011110010101;
assign LUT_2[53872] = 32'b11111111111111101011000010000101;
assign LUT_2[53873] = 32'b11111111111111100111111010011110;
assign LUT_2[53874] = 32'b11111111111111110001111011000001;
assign LUT_2[53875] = 32'b11111111111111101110110011011010;
assign LUT_2[53876] = 32'b11111111111111100111011111101101;
assign LUT_2[53877] = 32'b11111111111111100100011000000110;
assign LUT_2[53878] = 32'b11111111111111101110011000101001;
assign LUT_2[53879] = 32'b11111111111111101011010001000010;
assign LUT_2[53880] = 32'b11111111111111100101110011100010;
assign LUT_2[53881] = 32'b11111111111111100010101011111011;
assign LUT_2[53882] = 32'b11111111111111101100101100011110;
assign LUT_2[53883] = 32'b11111111111111101001100100110111;
assign LUT_2[53884] = 32'b11111111111111100010010001001010;
assign LUT_2[53885] = 32'b11111111111111011111001001100011;
assign LUT_2[53886] = 32'b11111111111111101001001010000110;
assign LUT_2[53887] = 32'b11111111111111100110000010011111;
assign LUT_2[53888] = 32'b11111111111111111100001101111110;
assign LUT_2[53889] = 32'b11111111111111111001000110010111;
assign LUT_2[53890] = 32'b00000000000000000011000110111010;
assign LUT_2[53891] = 32'b11111111111111111111111111010011;
assign LUT_2[53892] = 32'b11111111111111111000101011100110;
assign LUT_2[53893] = 32'b11111111111111110101100011111111;
assign LUT_2[53894] = 32'b11111111111111111111100100100010;
assign LUT_2[53895] = 32'b11111111111111111100011100111011;
assign LUT_2[53896] = 32'b11111111111111110110111111011011;
assign LUT_2[53897] = 32'b11111111111111110011110111110100;
assign LUT_2[53898] = 32'b11111111111111111101111000010111;
assign LUT_2[53899] = 32'b11111111111111111010110000110000;
assign LUT_2[53900] = 32'b11111111111111110011011101000011;
assign LUT_2[53901] = 32'b11111111111111110000010101011100;
assign LUT_2[53902] = 32'b11111111111111111010010101111111;
assign LUT_2[53903] = 32'b11111111111111110111001110011000;
assign LUT_2[53904] = 32'b11111111111111110110110010001000;
assign LUT_2[53905] = 32'b11111111111111110011101010100001;
assign LUT_2[53906] = 32'b11111111111111111101101011000100;
assign LUT_2[53907] = 32'b11111111111111111010100011011101;
assign LUT_2[53908] = 32'b11111111111111110011001111110000;
assign LUT_2[53909] = 32'b11111111111111110000001000001001;
assign LUT_2[53910] = 32'b11111111111111111010001000101100;
assign LUT_2[53911] = 32'b11111111111111110111000001000101;
assign LUT_2[53912] = 32'b11111111111111110001100011100101;
assign LUT_2[53913] = 32'b11111111111111101110011011111110;
assign LUT_2[53914] = 32'b11111111111111111000011100100001;
assign LUT_2[53915] = 32'b11111111111111110101010100111010;
assign LUT_2[53916] = 32'b11111111111111101110000001001101;
assign LUT_2[53917] = 32'b11111111111111101010111001100110;
assign LUT_2[53918] = 32'b11111111111111110100111010001001;
assign LUT_2[53919] = 32'b11111111111111110001110010100010;
assign LUT_2[53920] = 32'b11111111111111111100101001100111;
assign LUT_2[53921] = 32'b11111111111111111001100010000000;
assign LUT_2[53922] = 32'b00000000000000000011100010100011;
assign LUT_2[53923] = 32'b00000000000000000000011010111100;
assign LUT_2[53924] = 32'b11111111111111111001000111001111;
assign LUT_2[53925] = 32'b11111111111111110101111111101000;
assign LUT_2[53926] = 32'b00000000000000000000000000001011;
assign LUT_2[53927] = 32'b11111111111111111100111000100100;
assign LUT_2[53928] = 32'b11111111111111110111011011000100;
assign LUT_2[53929] = 32'b11111111111111110100010011011101;
assign LUT_2[53930] = 32'b11111111111111111110010100000000;
assign LUT_2[53931] = 32'b11111111111111111011001100011001;
assign LUT_2[53932] = 32'b11111111111111110011111000101100;
assign LUT_2[53933] = 32'b11111111111111110000110001000101;
assign LUT_2[53934] = 32'b11111111111111111010110001101000;
assign LUT_2[53935] = 32'b11111111111111110111101010000001;
assign LUT_2[53936] = 32'b11111111111111110111001101110001;
assign LUT_2[53937] = 32'b11111111111111110100000110001010;
assign LUT_2[53938] = 32'b11111111111111111110000110101101;
assign LUT_2[53939] = 32'b11111111111111111010111111000110;
assign LUT_2[53940] = 32'b11111111111111110011101011011001;
assign LUT_2[53941] = 32'b11111111111111110000100011110010;
assign LUT_2[53942] = 32'b11111111111111111010100100010101;
assign LUT_2[53943] = 32'b11111111111111110111011100101110;
assign LUT_2[53944] = 32'b11111111111111110001111111001110;
assign LUT_2[53945] = 32'b11111111111111101110110111100111;
assign LUT_2[53946] = 32'b11111111111111111000111000001010;
assign LUT_2[53947] = 32'b11111111111111110101110000100011;
assign LUT_2[53948] = 32'b11111111111111101110011100110110;
assign LUT_2[53949] = 32'b11111111111111101011010101001111;
assign LUT_2[53950] = 32'b11111111111111110101010101110010;
assign LUT_2[53951] = 32'b11111111111111110010001110001011;
assign LUT_2[53952] = 32'b11111111111111110100010110100001;
assign LUT_2[53953] = 32'b11111111111111110001001110111010;
assign LUT_2[53954] = 32'b11111111111111111011001111011101;
assign LUT_2[53955] = 32'b11111111111111111000000111110110;
assign LUT_2[53956] = 32'b11111111111111110000110100001001;
assign LUT_2[53957] = 32'b11111111111111101101101100100010;
assign LUT_2[53958] = 32'b11111111111111110111101101000101;
assign LUT_2[53959] = 32'b11111111111111110100100101011110;
assign LUT_2[53960] = 32'b11111111111111101111000111111110;
assign LUT_2[53961] = 32'b11111111111111101100000000010111;
assign LUT_2[53962] = 32'b11111111111111110110000000111010;
assign LUT_2[53963] = 32'b11111111111111110010111001010011;
assign LUT_2[53964] = 32'b11111111111111101011100101100110;
assign LUT_2[53965] = 32'b11111111111111101000011101111111;
assign LUT_2[53966] = 32'b11111111111111110010011110100010;
assign LUT_2[53967] = 32'b11111111111111101111010110111011;
assign LUT_2[53968] = 32'b11111111111111101110111010101011;
assign LUT_2[53969] = 32'b11111111111111101011110011000100;
assign LUT_2[53970] = 32'b11111111111111110101110011100111;
assign LUT_2[53971] = 32'b11111111111111110010101100000000;
assign LUT_2[53972] = 32'b11111111111111101011011000010011;
assign LUT_2[53973] = 32'b11111111111111101000010000101100;
assign LUT_2[53974] = 32'b11111111111111110010010001001111;
assign LUT_2[53975] = 32'b11111111111111101111001001101000;
assign LUT_2[53976] = 32'b11111111111111101001101100001000;
assign LUT_2[53977] = 32'b11111111111111100110100100100001;
assign LUT_2[53978] = 32'b11111111111111110000100101000100;
assign LUT_2[53979] = 32'b11111111111111101101011101011101;
assign LUT_2[53980] = 32'b11111111111111100110001001110000;
assign LUT_2[53981] = 32'b11111111111111100011000010001001;
assign LUT_2[53982] = 32'b11111111111111101101000010101100;
assign LUT_2[53983] = 32'b11111111111111101001111011000101;
assign LUT_2[53984] = 32'b11111111111111110100110010001010;
assign LUT_2[53985] = 32'b11111111111111110001101010100011;
assign LUT_2[53986] = 32'b11111111111111111011101011000110;
assign LUT_2[53987] = 32'b11111111111111111000100011011111;
assign LUT_2[53988] = 32'b11111111111111110001001111110010;
assign LUT_2[53989] = 32'b11111111111111101110001000001011;
assign LUT_2[53990] = 32'b11111111111111111000001000101110;
assign LUT_2[53991] = 32'b11111111111111110101000001000111;
assign LUT_2[53992] = 32'b11111111111111101111100011100111;
assign LUT_2[53993] = 32'b11111111111111101100011100000000;
assign LUT_2[53994] = 32'b11111111111111110110011100100011;
assign LUT_2[53995] = 32'b11111111111111110011010100111100;
assign LUT_2[53996] = 32'b11111111111111101100000001001111;
assign LUT_2[53997] = 32'b11111111111111101000111001101000;
assign LUT_2[53998] = 32'b11111111111111110010111010001011;
assign LUT_2[53999] = 32'b11111111111111101111110010100100;
assign LUT_2[54000] = 32'b11111111111111101111010110010100;
assign LUT_2[54001] = 32'b11111111111111101100001110101101;
assign LUT_2[54002] = 32'b11111111111111110110001111010000;
assign LUT_2[54003] = 32'b11111111111111110011000111101001;
assign LUT_2[54004] = 32'b11111111111111101011110011111100;
assign LUT_2[54005] = 32'b11111111111111101000101100010101;
assign LUT_2[54006] = 32'b11111111111111110010101100111000;
assign LUT_2[54007] = 32'b11111111111111101111100101010001;
assign LUT_2[54008] = 32'b11111111111111101010000111110001;
assign LUT_2[54009] = 32'b11111111111111100111000000001010;
assign LUT_2[54010] = 32'b11111111111111110001000000101101;
assign LUT_2[54011] = 32'b11111111111111101101111001000110;
assign LUT_2[54012] = 32'b11111111111111100110100101011001;
assign LUT_2[54013] = 32'b11111111111111100011011101110010;
assign LUT_2[54014] = 32'b11111111111111101101011110010101;
assign LUT_2[54015] = 32'b11111111111111101010010110101110;
assign LUT_2[54016] = 32'b11111111111111111011111000010101;
assign LUT_2[54017] = 32'b11111111111111111000110000101110;
assign LUT_2[54018] = 32'b00000000000000000010110001010001;
assign LUT_2[54019] = 32'b11111111111111111111101001101010;
assign LUT_2[54020] = 32'b11111111111111111000010101111101;
assign LUT_2[54021] = 32'b11111111111111110101001110010110;
assign LUT_2[54022] = 32'b11111111111111111111001110111001;
assign LUT_2[54023] = 32'b11111111111111111100000111010010;
assign LUT_2[54024] = 32'b11111111111111110110101001110010;
assign LUT_2[54025] = 32'b11111111111111110011100010001011;
assign LUT_2[54026] = 32'b11111111111111111101100010101110;
assign LUT_2[54027] = 32'b11111111111111111010011011000111;
assign LUT_2[54028] = 32'b11111111111111110011000111011010;
assign LUT_2[54029] = 32'b11111111111111101111111111110011;
assign LUT_2[54030] = 32'b11111111111111111010000000010110;
assign LUT_2[54031] = 32'b11111111111111110110111000101111;
assign LUT_2[54032] = 32'b11111111111111110110011100011111;
assign LUT_2[54033] = 32'b11111111111111110011010100111000;
assign LUT_2[54034] = 32'b11111111111111111101010101011011;
assign LUT_2[54035] = 32'b11111111111111111010001101110100;
assign LUT_2[54036] = 32'b11111111111111110010111010000111;
assign LUT_2[54037] = 32'b11111111111111101111110010100000;
assign LUT_2[54038] = 32'b11111111111111111001110011000011;
assign LUT_2[54039] = 32'b11111111111111110110101011011100;
assign LUT_2[54040] = 32'b11111111111111110001001101111100;
assign LUT_2[54041] = 32'b11111111111111101110000110010101;
assign LUT_2[54042] = 32'b11111111111111111000000110111000;
assign LUT_2[54043] = 32'b11111111111111110100111111010001;
assign LUT_2[54044] = 32'b11111111111111101101101011100100;
assign LUT_2[54045] = 32'b11111111111111101010100011111101;
assign LUT_2[54046] = 32'b11111111111111110100100100100000;
assign LUT_2[54047] = 32'b11111111111111110001011100111001;
assign LUT_2[54048] = 32'b11111111111111111100010011111110;
assign LUT_2[54049] = 32'b11111111111111111001001100010111;
assign LUT_2[54050] = 32'b00000000000000000011001100111010;
assign LUT_2[54051] = 32'b00000000000000000000000101010011;
assign LUT_2[54052] = 32'b11111111111111111000110001100110;
assign LUT_2[54053] = 32'b11111111111111110101101001111111;
assign LUT_2[54054] = 32'b11111111111111111111101010100010;
assign LUT_2[54055] = 32'b11111111111111111100100010111011;
assign LUT_2[54056] = 32'b11111111111111110111000101011011;
assign LUT_2[54057] = 32'b11111111111111110011111101110100;
assign LUT_2[54058] = 32'b11111111111111111101111110010111;
assign LUT_2[54059] = 32'b11111111111111111010110110110000;
assign LUT_2[54060] = 32'b11111111111111110011100011000011;
assign LUT_2[54061] = 32'b11111111111111110000011011011100;
assign LUT_2[54062] = 32'b11111111111111111010011011111111;
assign LUT_2[54063] = 32'b11111111111111110111010100011000;
assign LUT_2[54064] = 32'b11111111111111110110111000001000;
assign LUT_2[54065] = 32'b11111111111111110011110000100001;
assign LUT_2[54066] = 32'b11111111111111111101110001000100;
assign LUT_2[54067] = 32'b11111111111111111010101001011101;
assign LUT_2[54068] = 32'b11111111111111110011010101110000;
assign LUT_2[54069] = 32'b11111111111111110000001110001001;
assign LUT_2[54070] = 32'b11111111111111111010001110101100;
assign LUT_2[54071] = 32'b11111111111111110111000111000101;
assign LUT_2[54072] = 32'b11111111111111110001101001100101;
assign LUT_2[54073] = 32'b11111111111111101110100001111110;
assign LUT_2[54074] = 32'b11111111111111111000100010100001;
assign LUT_2[54075] = 32'b11111111111111110101011010111010;
assign LUT_2[54076] = 32'b11111111111111101110000111001101;
assign LUT_2[54077] = 32'b11111111111111101010111111100110;
assign LUT_2[54078] = 32'b11111111111111110101000000001001;
assign LUT_2[54079] = 32'b11111111111111110001111000100010;
assign LUT_2[54080] = 32'b11111111111111110100000000111000;
assign LUT_2[54081] = 32'b11111111111111110000111001010001;
assign LUT_2[54082] = 32'b11111111111111111010111001110100;
assign LUT_2[54083] = 32'b11111111111111110111110010001101;
assign LUT_2[54084] = 32'b11111111111111110000011110100000;
assign LUT_2[54085] = 32'b11111111111111101101010110111001;
assign LUT_2[54086] = 32'b11111111111111110111010111011100;
assign LUT_2[54087] = 32'b11111111111111110100001111110101;
assign LUT_2[54088] = 32'b11111111111111101110110010010101;
assign LUT_2[54089] = 32'b11111111111111101011101010101110;
assign LUT_2[54090] = 32'b11111111111111110101101011010001;
assign LUT_2[54091] = 32'b11111111111111110010100011101010;
assign LUT_2[54092] = 32'b11111111111111101011001111111101;
assign LUT_2[54093] = 32'b11111111111111101000001000010110;
assign LUT_2[54094] = 32'b11111111111111110010001000111001;
assign LUT_2[54095] = 32'b11111111111111101111000001010010;
assign LUT_2[54096] = 32'b11111111111111101110100101000010;
assign LUT_2[54097] = 32'b11111111111111101011011101011011;
assign LUT_2[54098] = 32'b11111111111111110101011101111110;
assign LUT_2[54099] = 32'b11111111111111110010010110010111;
assign LUT_2[54100] = 32'b11111111111111101011000010101010;
assign LUT_2[54101] = 32'b11111111111111100111111011000011;
assign LUT_2[54102] = 32'b11111111111111110001111011100110;
assign LUT_2[54103] = 32'b11111111111111101110110011111111;
assign LUT_2[54104] = 32'b11111111111111101001010110011111;
assign LUT_2[54105] = 32'b11111111111111100110001110111000;
assign LUT_2[54106] = 32'b11111111111111110000001111011011;
assign LUT_2[54107] = 32'b11111111111111101101000111110100;
assign LUT_2[54108] = 32'b11111111111111100101110100000111;
assign LUT_2[54109] = 32'b11111111111111100010101100100000;
assign LUT_2[54110] = 32'b11111111111111101100101101000011;
assign LUT_2[54111] = 32'b11111111111111101001100101011100;
assign LUT_2[54112] = 32'b11111111111111110100011100100001;
assign LUT_2[54113] = 32'b11111111111111110001010100111010;
assign LUT_2[54114] = 32'b11111111111111111011010101011101;
assign LUT_2[54115] = 32'b11111111111111111000001101110110;
assign LUT_2[54116] = 32'b11111111111111110000111010001001;
assign LUT_2[54117] = 32'b11111111111111101101110010100010;
assign LUT_2[54118] = 32'b11111111111111110111110011000101;
assign LUT_2[54119] = 32'b11111111111111110100101011011110;
assign LUT_2[54120] = 32'b11111111111111101111001101111110;
assign LUT_2[54121] = 32'b11111111111111101100000110010111;
assign LUT_2[54122] = 32'b11111111111111110110000110111010;
assign LUT_2[54123] = 32'b11111111111111110010111111010011;
assign LUT_2[54124] = 32'b11111111111111101011101011100110;
assign LUT_2[54125] = 32'b11111111111111101000100011111111;
assign LUT_2[54126] = 32'b11111111111111110010100100100010;
assign LUT_2[54127] = 32'b11111111111111101111011100111011;
assign LUT_2[54128] = 32'b11111111111111101111000000101011;
assign LUT_2[54129] = 32'b11111111111111101011111001000100;
assign LUT_2[54130] = 32'b11111111111111110101111001100111;
assign LUT_2[54131] = 32'b11111111111111110010110010000000;
assign LUT_2[54132] = 32'b11111111111111101011011110010011;
assign LUT_2[54133] = 32'b11111111111111101000010110101100;
assign LUT_2[54134] = 32'b11111111111111110010010111001111;
assign LUT_2[54135] = 32'b11111111111111101111001111101000;
assign LUT_2[54136] = 32'b11111111111111101001110010001000;
assign LUT_2[54137] = 32'b11111111111111100110101010100001;
assign LUT_2[54138] = 32'b11111111111111110000101011000100;
assign LUT_2[54139] = 32'b11111111111111101101100011011101;
assign LUT_2[54140] = 32'b11111111111111100110001111110000;
assign LUT_2[54141] = 32'b11111111111111100011001000001001;
assign LUT_2[54142] = 32'b11111111111111101101001000101100;
assign LUT_2[54143] = 32'b11111111111111101010000001000101;
assign LUT_2[54144] = 32'b00000000000000000000001100100100;
assign LUT_2[54145] = 32'b11111111111111111101000100111101;
assign LUT_2[54146] = 32'b00000000000000000111000101100000;
assign LUT_2[54147] = 32'b00000000000000000011111101111001;
assign LUT_2[54148] = 32'b11111111111111111100101010001100;
assign LUT_2[54149] = 32'b11111111111111111001100010100101;
assign LUT_2[54150] = 32'b00000000000000000011100011001000;
assign LUT_2[54151] = 32'b00000000000000000000011011100001;
assign LUT_2[54152] = 32'b11111111111111111010111110000001;
assign LUT_2[54153] = 32'b11111111111111110111110110011010;
assign LUT_2[54154] = 32'b00000000000000000001110110111101;
assign LUT_2[54155] = 32'b11111111111111111110101111010110;
assign LUT_2[54156] = 32'b11111111111111110111011011101001;
assign LUT_2[54157] = 32'b11111111111111110100010100000010;
assign LUT_2[54158] = 32'b11111111111111111110010100100101;
assign LUT_2[54159] = 32'b11111111111111111011001100111110;
assign LUT_2[54160] = 32'b11111111111111111010110000101110;
assign LUT_2[54161] = 32'b11111111111111110111101001000111;
assign LUT_2[54162] = 32'b00000000000000000001101001101010;
assign LUT_2[54163] = 32'b11111111111111111110100010000011;
assign LUT_2[54164] = 32'b11111111111111110111001110010110;
assign LUT_2[54165] = 32'b11111111111111110100000110101111;
assign LUT_2[54166] = 32'b11111111111111111110000111010010;
assign LUT_2[54167] = 32'b11111111111111111010111111101011;
assign LUT_2[54168] = 32'b11111111111111110101100010001011;
assign LUT_2[54169] = 32'b11111111111111110010011010100100;
assign LUT_2[54170] = 32'b11111111111111111100011011000111;
assign LUT_2[54171] = 32'b11111111111111111001010011100000;
assign LUT_2[54172] = 32'b11111111111111110001111111110011;
assign LUT_2[54173] = 32'b11111111111111101110111000001100;
assign LUT_2[54174] = 32'b11111111111111111000111000101111;
assign LUT_2[54175] = 32'b11111111111111110101110001001000;
assign LUT_2[54176] = 32'b00000000000000000000101000001101;
assign LUT_2[54177] = 32'b11111111111111111101100000100110;
assign LUT_2[54178] = 32'b00000000000000000111100001001001;
assign LUT_2[54179] = 32'b00000000000000000100011001100010;
assign LUT_2[54180] = 32'b11111111111111111101000101110101;
assign LUT_2[54181] = 32'b11111111111111111001111110001110;
assign LUT_2[54182] = 32'b00000000000000000011111110110001;
assign LUT_2[54183] = 32'b00000000000000000000110111001010;
assign LUT_2[54184] = 32'b11111111111111111011011001101010;
assign LUT_2[54185] = 32'b11111111111111111000010010000011;
assign LUT_2[54186] = 32'b00000000000000000010010010100110;
assign LUT_2[54187] = 32'b11111111111111111111001010111111;
assign LUT_2[54188] = 32'b11111111111111110111110111010010;
assign LUT_2[54189] = 32'b11111111111111110100101111101011;
assign LUT_2[54190] = 32'b11111111111111111110110000001110;
assign LUT_2[54191] = 32'b11111111111111111011101000100111;
assign LUT_2[54192] = 32'b11111111111111111011001100010111;
assign LUT_2[54193] = 32'b11111111111111111000000100110000;
assign LUT_2[54194] = 32'b00000000000000000010000101010011;
assign LUT_2[54195] = 32'b11111111111111111110111101101100;
assign LUT_2[54196] = 32'b11111111111111110111101001111111;
assign LUT_2[54197] = 32'b11111111111111110100100010011000;
assign LUT_2[54198] = 32'b11111111111111111110100010111011;
assign LUT_2[54199] = 32'b11111111111111111011011011010100;
assign LUT_2[54200] = 32'b11111111111111110101111101110100;
assign LUT_2[54201] = 32'b11111111111111110010110110001101;
assign LUT_2[54202] = 32'b11111111111111111100110110110000;
assign LUT_2[54203] = 32'b11111111111111111001101111001001;
assign LUT_2[54204] = 32'b11111111111111110010011011011100;
assign LUT_2[54205] = 32'b11111111111111101111010011110101;
assign LUT_2[54206] = 32'b11111111111111111001010100011000;
assign LUT_2[54207] = 32'b11111111111111110110001100110001;
assign LUT_2[54208] = 32'b11111111111111111000010101000111;
assign LUT_2[54209] = 32'b11111111111111110101001101100000;
assign LUT_2[54210] = 32'b11111111111111111111001110000011;
assign LUT_2[54211] = 32'b11111111111111111100000110011100;
assign LUT_2[54212] = 32'b11111111111111110100110010101111;
assign LUT_2[54213] = 32'b11111111111111110001101011001000;
assign LUT_2[54214] = 32'b11111111111111111011101011101011;
assign LUT_2[54215] = 32'b11111111111111111000100100000100;
assign LUT_2[54216] = 32'b11111111111111110011000110100100;
assign LUT_2[54217] = 32'b11111111111111101111111110111101;
assign LUT_2[54218] = 32'b11111111111111111001111111100000;
assign LUT_2[54219] = 32'b11111111111111110110110111111001;
assign LUT_2[54220] = 32'b11111111111111101111100100001100;
assign LUT_2[54221] = 32'b11111111111111101100011100100101;
assign LUT_2[54222] = 32'b11111111111111110110011101001000;
assign LUT_2[54223] = 32'b11111111111111110011010101100001;
assign LUT_2[54224] = 32'b11111111111111110010111001010001;
assign LUT_2[54225] = 32'b11111111111111101111110001101010;
assign LUT_2[54226] = 32'b11111111111111111001110010001101;
assign LUT_2[54227] = 32'b11111111111111110110101010100110;
assign LUT_2[54228] = 32'b11111111111111101111010110111001;
assign LUT_2[54229] = 32'b11111111111111101100001111010010;
assign LUT_2[54230] = 32'b11111111111111110110001111110101;
assign LUT_2[54231] = 32'b11111111111111110011001000001110;
assign LUT_2[54232] = 32'b11111111111111101101101010101110;
assign LUT_2[54233] = 32'b11111111111111101010100011000111;
assign LUT_2[54234] = 32'b11111111111111110100100011101010;
assign LUT_2[54235] = 32'b11111111111111110001011100000011;
assign LUT_2[54236] = 32'b11111111111111101010001000010110;
assign LUT_2[54237] = 32'b11111111111111100111000000101111;
assign LUT_2[54238] = 32'b11111111111111110001000001010010;
assign LUT_2[54239] = 32'b11111111111111101101111001101011;
assign LUT_2[54240] = 32'b11111111111111111000110000110000;
assign LUT_2[54241] = 32'b11111111111111110101101001001001;
assign LUT_2[54242] = 32'b11111111111111111111101001101100;
assign LUT_2[54243] = 32'b11111111111111111100100010000101;
assign LUT_2[54244] = 32'b11111111111111110101001110011000;
assign LUT_2[54245] = 32'b11111111111111110010000110110001;
assign LUT_2[54246] = 32'b11111111111111111100000111010100;
assign LUT_2[54247] = 32'b11111111111111111000111111101101;
assign LUT_2[54248] = 32'b11111111111111110011100010001101;
assign LUT_2[54249] = 32'b11111111111111110000011010100110;
assign LUT_2[54250] = 32'b11111111111111111010011011001001;
assign LUT_2[54251] = 32'b11111111111111110111010011100010;
assign LUT_2[54252] = 32'b11111111111111101111111111110101;
assign LUT_2[54253] = 32'b11111111111111101100111000001110;
assign LUT_2[54254] = 32'b11111111111111110110111000110001;
assign LUT_2[54255] = 32'b11111111111111110011110001001010;
assign LUT_2[54256] = 32'b11111111111111110011010100111010;
assign LUT_2[54257] = 32'b11111111111111110000001101010011;
assign LUT_2[54258] = 32'b11111111111111111010001101110110;
assign LUT_2[54259] = 32'b11111111111111110111000110001111;
assign LUT_2[54260] = 32'b11111111111111101111110010100010;
assign LUT_2[54261] = 32'b11111111111111101100101010111011;
assign LUT_2[54262] = 32'b11111111111111110110101011011110;
assign LUT_2[54263] = 32'b11111111111111110011100011110111;
assign LUT_2[54264] = 32'b11111111111111101110000110010111;
assign LUT_2[54265] = 32'b11111111111111101010111110110000;
assign LUT_2[54266] = 32'b11111111111111110100111111010011;
assign LUT_2[54267] = 32'b11111111111111110001110111101100;
assign LUT_2[54268] = 32'b11111111111111101010100011111111;
assign LUT_2[54269] = 32'b11111111111111100111011100011000;
assign LUT_2[54270] = 32'b11111111111111110001011100111011;
assign LUT_2[54271] = 32'b11111111111111101110010101010100;
assign LUT_2[54272] = 32'b11111111111111111001110100000010;
assign LUT_2[54273] = 32'b11111111111111110110101100011011;
assign LUT_2[54274] = 32'b00000000000000000000101100111110;
assign LUT_2[54275] = 32'b11111111111111111101100101010111;
assign LUT_2[54276] = 32'b11111111111111110110010001101010;
assign LUT_2[54277] = 32'b11111111111111110011001010000011;
assign LUT_2[54278] = 32'b11111111111111111101001010100110;
assign LUT_2[54279] = 32'b11111111111111111010000010111111;
assign LUT_2[54280] = 32'b11111111111111110100100101011111;
assign LUT_2[54281] = 32'b11111111111111110001011101111000;
assign LUT_2[54282] = 32'b11111111111111111011011110011011;
assign LUT_2[54283] = 32'b11111111111111111000010110110100;
assign LUT_2[54284] = 32'b11111111111111110001000011000111;
assign LUT_2[54285] = 32'b11111111111111101101111011100000;
assign LUT_2[54286] = 32'b11111111111111110111111100000011;
assign LUT_2[54287] = 32'b11111111111111110100110100011100;
assign LUT_2[54288] = 32'b11111111111111110100011000001100;
assign LUT_2[54289] = 32'b11111111111111110001010000100101;
assign LUT_2[54290] = 32'b11111111111111111011010001001000;
assign LUT_2[54291] = 32'b11111111111111111000001001100001;
assign LUT_2[54292] = 32'b11111111111111110000110101110100;
assign LUT_2[54293] = 32'b11111111111111101101101110001101;
assign LUT_2[54294] = 32'b11111111111111110111101110110000;
assign LUT_2[54295] = 32'b11111111111111110100100111001001;
assign LUT_2[54296] = 32'b11111111111111101111001001101001;
assign LUT_2[54297] = 32'b11111111111111101100000010000010;
assign LUT_2[54298] = 32'b11111111111111110110000010100101;
assign LUT_2[54299] = 32'b11111111111111110010111010111110;
assign LUT_2[54300] = 32'b11111111111111101011100111010001;
assign LUT_2[54301] = 32'b11111111111111101000011111101010;
assign LUT_2[54302] = 32'b11111111111111110010100000001101;
assign LUT_2[54303] = 32'b11111111111111101111011000100110;
assign LUT_2[54304] = 32'b11111111111111111010001111101011;
assign LUT_2[54305] = 32'b11111111111111110111001000000100;
assign LUT_2[54306] = 32'b00000000000000000001001000100111;
assign LUT_2[54307] = 32'b11111111111111111110000001000000;
assign LUT_2[54308] = 32'b11111111111111110110101101010011;
assign LUT_2[54309] = 32'b11111111111111110011100101101100;
assign LUT_2[54310] = 32'b11111111111111111101100110001111;
assign LUT_2[54311] = 32'b11111111111111111010011110101000;
assign LUT_2[54312] = 32'b11111111111111110101000001001000;
assign LUT_2[54313] = 32'b11111111111111110001111001100001;
assign LUT_2[54314] = 32'b11111111111111111011111010000100;
assign LUT_2[54315] = 32'b11111111111111111000110010011101;
assign LUT_2[54316] = 32'b11111111111111110001011110110000;
assign LUT_2[54317] = 32'b11111111111111101110010111001001;
assign LUT_2[54318] = 32'b11111111111111111000010111101100;
assign LUT_2[54319] = 32'b11111111111111110101010000000101;
assign LUT_2[54320] = 32'b11111111111111110100110011110101;
assign LUT_2[54321] = 32'b11111111111111110001101100001110;
assign LUT_2[54322] = 32'b11111111111111111011101100110001;
assign LUT_2[54323] = 32'b11111111111111111000100101001010;
assign LUT_2[54324] = 32'b11111111111111110001010001011101;
assign LUT_2[54325] = 32'b11111111111111101110001001110110;
assign LUT_2[54326] = 32'b11111111111111111000001010011001;
assign LUT_2[54327] = 32'b11111111111111110101000010110010;
assign LUT_2[54328] = 32'b11111111111111101111100101010010;
assign LUT_2[54329] = 32'b11111111111111101100011101101011;
assign LUT_2[54330] = 32'b11111111111111110110011110001110;
assign LUT_2[54331] = 32'b11111111111111110011010110100111;
assign LUT_2[54332] = 32'b11111111111111101100000010111010;
assign LUT_2[54333] = 32'b11111111111111101000111011010011;
assign LUT_2[54334] = 32'b11111111111111110010111011110110;
assign LUT_2[54335] = 32'b11111111111111101111110100001111;
assign LUT_2[54336] = 32'b11111111111111110001111100100101;
assign LUT_2[54337] = 32'b11111111111111101110110100111110;
assign LUT_2[54338] = 32'b11111111111111111000110101100001;
assign LUT_2[54339] = 32'b11111111111111110101101101111010;
assign LUT_2[54340] = 32'b11111111111111101110011010001101;
assign LUT_2[54341] = 32'b11111111111111101011010010100110;
assign LUT_2[54342] = 32'b11111111111111110101010011001001;
assign LUT_2[54343] = 32'b11111111111111110010001011100010;
assign LUT_2[54344] = 32'b11111111111111101100101110000010;
assign LUT_2[54345] = 32'b11111111111111101001100110011011;
assign LUT_2[54346] = 32'b11111111111111110011100110111110;
assign LUT_2[54347] = 32'b11111111111111110000011111010111;
assign LUT_2[54348] = 32'b11111111111111101001001011101010;
assign LUT_2[54349] = 32'b11111111111111100110000100000011;
assign LUT_2[54350] = 32'b11111111111111110000000100100110;
assign LUT_2[54351] = 32'b11111111111111101100111100111111;
assign LUT_2[54352] = 32'b11111111111111101100100000101111;
assign LUT_2[54353] = 32'b11111111111111101001011001001000;
assign LUT_2[54354] = 32'b11111111111111110011011001101011;
assign LUT_2[54355] = 32'b11111111111111110000010010000100;
assign LUT_2[54356] = 32'b11111111111111101000111110010111;
assign LUT_2[54357] = 32'b11111111111111100101110110110000;
assign LUT_2[54358] = 32'b11111111111111101111110111010011;
assign LUT_2[54359] = 32'b11111111111111101100101111101100;
assign LUT_2[54360] = 32'b11111111111111100111010010001100;
assign LUT_2[54361] = 32'b11111111111111100100001010100101;
assign LUT_2[54362] = 32'b11111111111111101110001011001000;
assign LUT_2[54363] = 32'b11111111111111101011000011100001;
assign LUT_2[54364] = 32'b11111111111111100011101111110100;
assign LUT_2[54365] = 32'b11111111111111100000101000001101;
assign LUT_2[54366] = 32'b11111111111111101010101000110000;
assign LUT_2[54367] = 32'b11111111111111100111100001001001;
assign LUT_2[54368] = 32'b11111111111111110010011000001110;
assign LUT_2[54369] = 32'b11111111111111101111010000100111;
assign LUT_2[54370] = 32'b11111111111111111001010001001010;
assign LUT_2[54371] = 32'b11111111111111110110001001100011;
assign LUT_2[54372] = 32'b11111111111111101110110101110110;
assign LUT_2[54373] = 32'b11111111111111101011101110001111;
assign LUT_2[54374] = 32'b11111111111111110101101110110010;
assign LUT_2[54375] = 32'b11111111111111110010100111001011;
assign LUT_2[54376] = 32'b11111111111111101101001001101011;
assign LUT_2[54377] = 32'b11111111111111101010000010000100;
assign LUT_2[54378] = 32'b11111111111111110100000010100111;
assign LUT_2[54379] = 32'b11111111111111110000111011000000;
assign LUT_2[54380] = 32'b11111111111111101001100111010011;
assign LUT_2[54381] = 32'b11111111111111100110011111101100;
assign LUT_2[54382] = 32'b11111111111111110000100000001111;
assign LUT_2[54383] = 32'b11111111111111101101011000101000;
assign LUT_2[54384] = 32'b11111111111111101100111100011000;
assign LUT_2[54385] = 32'b11111111111111101001110100110001;
assign LUT_2[54386] = 32'b11111111111111110011110101010100;
assign LUT_2[54387] = 32'b11111111111111110000101101101101;
assign LUT_2[54388] = 32'b11111111111111101001011010000000;
assign LUT_2[54389] = 32'b11111111111111100110010010011001;
assign LUT_2[54390] = 32'b11111111111111110000010010111100;
assign LUT_2[54391] = 32'b11111111111111101101001011010101;
assign LUT_2[54392] = 32'b11111111111111100111101101110101;
assign LUT_2[54393] = 32'b11111111111111100100100110001110;
assign LUT_2[54394] = 32'b11111111111111101110100110110001;
assign LUT_2[54395] = 32'b11111111111111101011011111001010;
assign LUT_2[54396] = 32'b11111111111111100100001011011101;
assign LUT_2[54397] = 32'b11111111111111100001000011110110;
assign LUT_2[54398] = 32'b11111111111111101011000100011001;
assign LUT_2[54399] = 32'b11111111111111100111111100110010;
assign LUT_2[54400] = 32'b11111111111111111110001000010001;
assign LUT_2[54401] = 32'b11111111111111111011000000101010;
assign LUT_2[54402] = 32'b00000000000000000101000001001101;
assign LUT_2[54403] = 32'b00000000000000000001111001100110;
assign LUT_2[54404] = 32'b11111111111111111010100101111001;
assign LUT_2[54405] = 32'b11111111111111110111011110010010;
assign LUT_2[54406] = 32'b00000000000000000001011110110101;
assign LUT_2[54407] = 32'b11111111111111111110010111001110;
assign LUT_2[54408] = 32'b11111111111111111000111001101110;
assign LUT_2[54409] = 32'b11111111111111110101110010000111;
assign LUT_2[54410] = 32'b11111111111111111111110010101010;
assign LUT_2[54411] = 32'b11111111111111111100101011000011;
assign LUT_2[54412] = 32'b11111111111111110101010111010110;
assign LUT_2[54413] = 32'b11111111111111110010001111101111;
assign LUT_2[54414] = 32'b11111111111111111100010000010010;
assign LUT_2[54415] = 32'b11111111111111111001001000101011;
assign LUT_2[54416] = 32'b11111111111111111000101100011011;
assign LUT_2[54417] = 32'b11111111111111110101100100110100;
assign LUT_2[54418] = 32'b11111111111111111111100101010111;
assign LUT_2[54419] = 32'b11111111111111111100011101110000;
assign LUT_2[54420] = 32'b11111111111111110101001010000011;
assign LUT_2[54421] = 32'b11111111111111110010000010011100;
assign LUT_2[54422] = 32'b11111111111111111100000010111111;
assign LUT_2[54423] = 32'b11111111111111111000111011011000;
assign LUT_2[54424] = 32'b11111111111111110011011101111000;
assign LUT_2[54425] = 32'b11111111111111110000010110010001;
assign LUT_2[54426] = 32'b11111111111111111010010110110100;
assign LUT_2[54427] = 32'b11111111111111110111001111001101;
assign LUT_2[54428] = 32'b11111111111111101111111011100000;
assign LUT_2[54429] = 32'b11111111111111101100110011111001;
assign LUT_2[54430] = 32'b11111111111111110110110100011100;
assign LUT_2[54431] = 32'b11111111111111110011101100110101;
assign LUT_2[54432] = 32'b11111111111111111110100011111010;
assign LUT_2[54433] = 32'b11111111111111111011011100010011;
assign LUT_2[54434] = 32'b00000000000000000101011100110110;
assign LUT_2[54435] = 32'b00000000000000000010010101001111;
assign LUT_2[54436] = 32'b11111111111111111011000001100010;
assign LUT_2[54437] = 32'b11111111111111110111111001111011;
assign LUT_2[54438] = 32'b00000000000000000001111010011110;
assign LUT_2[54439] = 32'b11111111111111111110110010110111;
assign LUT_2[54440] = 32'b11111111111111111001010101010111;
assign LUT_2[54441] = 32'b11111111111111110110001101110000;
assign LUT_2[54442] = 32'b00000000000000000000001110010011;
assign LUT_2[54443] = 32'b11111111111111111101000110101100;
assign LUT_2[54444] = 32'b11111111111111110101110010111111;
assign LUT_2[54445] = 32'b11111111111111110010101011011000;
assign LUT_2[54446] = 32'b11111111111111111100101011111011;
assign LUT_2[54447] = 32'b11111111111111111001100100010100;
assign LUT_2[54448] = 32'b11111111111111111001001000000100;
assign LUT_2[54449] = 32'b11111111111111110110000000011101;
assign LUT_2[54450] = 32'b00000000000000000000000001000000;
assign LUT_2[54451] = 32'b11111111111111111100111001011001;
assign LUT_2[54452] = 32'b11111111111111110101100101101100;
assign LUT_2[54453] = 32'b11111111111111110010011110000101;
assign LUT_2[54454] = 32'b11111111111111111100011110101000;
assign LUT_2[54455] = 32'b11111111111111111001010111000001;
assign LUT_2[54456] = 32'b11111111111111110011111001100001;
assign LUT_2[54457] = 32'b11111111111111110000110001111010;
assign LUT_2[54458] = 32'b11111111111111111010110010011101;
assign LUT_2[54459] = 32'b11111111111111110111101010110110;
assign LUT_2[54460] = 32'b11111111111111110000010111001001;
assign LUT_2[54461] = 32'b11111111111111101101001111100010;
assign LUT_2[54462] = 32'b11111111111111110111010000000101;
assign LUT_2[54463] = 32'b11111111111111110100001000011110;
assign LUT_2[54464] = 32'b11111111111111110110010000110100;
assign LUT_2[54465] = 32'b11111111111111110011001001001101;
assign LUT_2[54466] = 32'b11111111111111111101001001110000;
assign LUT_2[54467] = 32'b11111111111111111010000010001001;
assign LUT_2[54468] = 32'b11111111111111110010101110011100;
assign LUT_2[54469] = 32'b11111111111111101111100110110101;
assign LUT_2[54470] = 32'b11111111111111111001100111011000;
assign LUT_2[54471] = 32'b11111111111111110110011111110001;
assign LUT_2[54472] = 32'b11111111111111110001000010010001;
assign LUT_2[54473] = 32'b11111111111111101101111010101010;
assign LUT_2[54474] = 32'b11111111111111110111111011001101;
assign LUT_2[54475] = 32'b11111111111111110100110011100110;
assign LUT_2[54476] = 32'b11111111111111101101011111111001;
assign LUT_2[54477] = 32'b11111111111111101010011000010010;
assign LUT_2[54478] = 32'b11111111111111110100011000110101;
assign LUT_2[54479] = 32'b11111111111111110001010001001110;
assign LUT_2[54480] = 32'b11111111111111110000110100111110;
assign LUT_2[54481] = 32'b11111111111111101101101101010111;
assign LUT_2[54482] = 32'b11111111111111110111101101111010;
assign LUT_2[54483] = 32'b11111111111111110100100110010011;
assign LUT_2[54484] = 32'b11111111111111101101010010100110;
assign LUT_2[54485] = 32'b11111111111111101010001010111111;
assign LUT_2[54486] = 32'b11111111111111110100001011100010;
assign LUT_2[54487] = 32'b11111111111111110001000011111011;
assign LUT_2[54488] = 32'b11111111111111101011100110011011;
assign LUT_2[54489] = 32'b11111111111111101000011110110100;
assign LUT_2[54490] = 32'b11111111111111110010011111010111;
assign LUT_2[54491] = 32'b11111111111111101111010111110000;
assign LUT_2[54492] = 32'b11111111111111101000000100000011;
assign LUT_2[54493] = 32'b11111111111111100100111100011100;
assign LUT_2[54494] = 32'b11111111111111101110111100111111;
assign LUT_2[54495] = 32'b11111111111111101011110101011000;
assign LUT_2[54496] = 32'b11111111111111110110101100011101;
assign LUT_2[54497] = 32'b11111111111111110011100100110110;
assign LUT_2[54498] = 32'b11111111111111111101100101011001;
assign LUT_2[54499] = 32'b11111111111111111010011101110010;
assign LUT_2[54500] = 32'b11111111111111110011001010000101;
assign LUT_2[54501] = 32'b11111111111111110000000010011110;
assign LUT_2[54502] = 32'b11111111111111111010000011000001;
assign LUT_2[54503] = 32'b11111111111111110110111011011010;
assign LUT_2[54504] = 32'b11111111111111110001011101111010;
assign LUT_2[54505] = 32'b11111111111111101110010110010011;
assign LUT_2[54506] = 32'b11111111111111111000010110110110;
assign LUT_2[54507] = 32'b11111111111111110101001111001111;
assign LUT_2[54508] = 32'b11111111111111101101111011100010;
assign LUT_2[54509] = 32'b11111111111111101010110011111011;
assign LUT_2[54510] = 32'b11111111111111110100110100011110;
assign LUT_2[54511] = 32'b11111111111111110001101100110111;
assign LUT_2[54512] = 32'b11111111111111110001010000100111;
assign LUT_2[54513] = 32'b11111111111111101110001001000000;
assign LUT_2[54514] = 32'b11111111111111111000001001100011;
assign LUT_2[54515] = 32'b11111111111111110101000001111100;
assign LUT_2[54516] = 32'b11111111111111101101101110001111;
assign LUT_2[54517] = 32'b11111111111111101010100110101000;
assign LUT_2[54518] = 32'b11111111111111110100100111001011;
assign LUT_2[54519] = 32'b11111111111111110001011111100100;
assign LUT_2[54520] = 32'b11111111111111101100000010000100;
assign LUT_2[54521] = 32'b11111111111111101000111010011101;
assign LUT_2[54522] = 32'b11111111111111110010111011000000;
assign LUT_2[54523] = 32'b11111111111111101111110011011001;
assign LUT_2[54524] = 32'b11111111111111101000011111101100;
assign LUT_2[54525] = 32'b11111111111111100101011000000101;
assign LUT_2[54526] = 32'b11111111111111101111011000101000;
assign LUT_2[54527] = 32'b11111111111111101100010001000001;
assign LUT_2[54528] = 32'b11111111111111111101110010101000;
assign LUT_2[54529] = 32'b11111111111111111010101011000001;
assign LUT_2[54530] = 32'b00000000000000000100101011100100;
assign LUT_2[54531] = 32'b00000000000000000001100011111101;
assign LUT_2[54532] = 32'b11111111111111111010010000010000;
assign LUT_2[54533] = 32'b11111111111111110111001000101001;
assign LUT_2[54534] = 32'b00000000000000000001001001001100;
assign LUT_2[54535] = 32'b11111111111111111110000001100101;
assign LUT_2[54536] = 32'b11111111111111111000100100000101;
assign LUT_2[54537] = 32'b11111111111111110101011100011110;
assign LUT_2[54538] = 32'b11111111111111111111011101000001;
assign LUT_2[54539] = 32'b11111111111111111100010101011010;
assign LUT_2[54540] = 32'b11111111111111110101000001101101;
assign LUT_2[54541] = 32'b11111111111111110001111010000110;
assign LUT_2[54542] = 32'b11111111111111111011111010101001;
assign LUT_2[54543] = 32'b11111111111111111000110011000010;
assign LUT_2[54544] = 32'b11111111111111111000010110110010;
assign LUT_2[54545] = 32'b11111111111111110101001111001011;
assign LUT_2[54546] = 32'b11111111111111111111001111101110;
assign LUT_2[54547] = 32'b11111111111111111100001000000111;
assign LUT_2[54548] = 32'b11111111111111110100110100011010;
assign LUT_2[54549] = 32'b11111111111111110001101100110011;
assign LUT_2[54550] = 32'b11111111111111111011101101010110;
assign LUT_2[54551] = 32'b11111111111111111000100101101111;
assign LUT_2[54552] = 32'b11111111111111110011001000001111;
assign LUT_2[54553] = 32'b11111111111111110000000000101000;
assign LUT_2[54554] = 32'b11111111111111111010000001001011;
assign LUT_2[54555] = 32'b11111111111111110110111001100100;
assign LUT_2[54556] = 32'b11111111111111101111100101110111;
assign LUT_2[54557] = 32'b11111111111111101100011110010000;
assign LUT_2[54558] = 32'b11111111111111110110011110110011;
assign LUT_2[54559] = 32'b11111111111111110011010111001100;
assign LUT_2[54560] = 32'b11111111111111111110001110010001;
assign LUT_2[54561] = 32'b11111111111111111011000110101010;
assign LUT_2[54562] = 32'b00000000000000000101000111001101;
assign LUT_2[54563] = 32'b00000000000000000001111111100110;
assign LUT_2[54564] = 32'b11111111111111111010101011111001;
assign LUT_2[54565] = 32'b11111111111111110111100100010010;
assign LUT_2[54566] = 32'b00000000000000000001100100110101;
assign LUT_2[54567] = 32'b11111111111111111110011101001110;
assign LUT_2[54568] = 32'b11111111111111111000111111101110;
assign LUT_2[54569] = 32'b11111111111111110101111000000111;
assign LUT_2[54570] = 32'b11111111111111111111111000101010;
assign LUT_2[54571] = 32'b11111111111111111100110001000011;
assign LUT_2[54572] = 32'b11111111111111110101011101010110;
assign LUT_2[54573] = 32'b11111111111111110010010101101111;
assign LUT_2[54574] = 32'b11111111111111111100010110010010;
assign LUT_2[54575] = 32'b11111111111111111001001110101011;
assign LUT_2[54576] = 32'b11111111111111111000110010011011;
assign LUT_2[54577] = 32'b11111111111111110101101010110100;
assign LUT_2[54578] = 32'b11111111111111111111101011010111;
assign LUT_2[54579] = 32'b11111111111111111100100011110000;
assign LUT_2[54580] = 32'b11111111111111110101010000000011;
assign LUT_2[54581] = 32'b11111111111111110010001000011100;
assign LUT_2[54582] = 32'b11111111111111111100001000111111;
assign LUT_2[54583] = 32'b11111111111111111001000001011000;
assign LUT_2[54584] = 32'b11111111111111110011100011111000;
assign LUT_2[54585] = 32'b11111111111111110000011100010001;
assign LUT_2[54586] = 32'b11111111111111111010011100110100;
assign LUT_2[54587] = 32'b11111111111111110111010101001101;
assign LUT_2[54588] = 32'b11111111111111110000000001100000;
assign LUT_2[54589] = 32'b11111111111111101100111001111001;
assign LUT_2[54590] = 32'b11111111111111110110111010011100;
assign LUT_2[54591] = 32'b11111111111111110011110010110101;
assign LUT_2[54592] = 32'b11111111111111110101111011001011;
assign LUT_2[54593] = 32'b11111111111111110010110011100100;
assign LUT_2[54594] = 32'b11111111111111111100110100000111;
assign LUT_2[54595] = 32'b11111111111111111001101100100000;
assign LUT_2[54596] = 32'b11111111111111110010011000110011;
assign LUT_2[54597] = 32'b11111111111111101111010001001100;
assign LUT_2[54598] = 32'b11111111111111111001010001101111;
assign LUT_2[54599] = 32'b11111111111111110110001010001000;
assign LUT_2[54600] = 32'b11111111111111110000101100101000;
assign LUT_2[54601] = 32'b11111111111111101101100101000001;
assign LUT_2[54602] = 32'b11111111111111110111100101100100;
assign LUT_2[54603] = 32'b11111111111111110100011101111101;
assign LUT_2[54604] = 32'b11111111111111101101001010010000;
assign LUT_2[54605] = 32'b11111111111111101010000010101001;
assign LUT_2[54606] = 32'b11111111111111110100000011001100;
assign LUT_2[54607] = 32'b11111111111111110000111011100101;
assign LUT_2[54608] = 32'b11111111111111110000011111010101;
assign LUT_2[54609] = 32'b11111111111111101101010111101110;
assign LUT_2[54610] = 32'b11111111111111110111011000010001;
assign LUT_2[54611] = 32'b11111111111111110100010000101010;
assign LUT_2[54612] = 32'b11111111111111101100111100111101;
assign LUT_2[54613] = 32'b11111111111111101001110101010110;
assign LUT_2[54614] = 32'b11111111111111110011110101111001;
assign LUT_2[54615] = 32'b11111111111111110000101110010010;
assign LUT_2[54616] = 32'b11111111111111101011010000110010;
assign LUT_2[54617] = 32'b11111111111111101000001001001011;
assign LUT_2[54618] = 32'b11111111111111110010001001101110;
assign LUT_2[54619] = 32'b11111111111111101111000010000111;
assign LUT_2[54620] = 32'b11111111111111100111101110011010;
assign LUT_2[54621] = 32'b11111111111111100100100110110011;
assign LUT_2[54622] = 32'b11111111111111101110100111010110;
assign LUT_2[54623] = 32'b11111111111111101011011111101111;
assign LUT_2[54624] = 32'b11111111111111110110010110110100;
assign LUT_2[54625] = 32'b11111111111111110011001111001101;
assign LUT_2[54626] = 32'b11111111111111111101001111110000;
assign LUT_2[54627] = 32'b11111111111111111010001000001001;
assign LUT_2[54628] = 32'b11111111111111110010110100011100;
assign LUT_2[54629] = 32'b11111111111111101111101100110101;
assign LUT_2[54630] = 32'b11111111111111111001101101011000;
assign LUT_2[54631] = 32'b11111111111111110110100101110001;
assign LUT_2[54632] = 32'b11111111111111110001001000010001;
assign LUT_2[54633] = 32'b11111111111111101110000000101010;
assign LUT_2[54634] = 32'b11111111111111111000000001001101;
assign LUT_2[54635] = 32'b11111111111111110100111001100110;
assign LUT_2[54636] = 32'b11111111111111101101100101111001;
assign LUT_2[54637] = 32'b11111111111111101010011110010010;
assign LUT_2[54638] = 32'b11111111111111110100011110110101;
assign LUT_2[54639] = 32'b11111111111111110001010111001110;
assign LUT_2[54640] = 32'b11111111111111110000111010111110;
assign LUT_2[54641] = 32'b11111111111111101101110011010111;
assign LUT_2[54642] = 32'b11111111111111110111110011111010;
assign LUT_2[54643] = 32'b11111111111111110100101100010011;
assign LUT_2[54644] = 32'b11111111111111101101011000100110;
assign LUT_2[54645] = 32'b11111111111111101010010000111111;
assign LUT_2[54646] = 32'b11111111111111110100010001100010;
assign LUT_2[54647] = 32'b11111111111111110001001001111011;
assign LUT_2[54648] = 32'b11111111111111101011101100011011;
assign LUT_2[54649] = 32'b11111111111111101000100100110100;
assign LUT_2[54650] = 32'b11111111111111110010100101010111;
assign LUT_2[54651] = 32'b11111111111111101111011101110000;
assign LUT_2[54652] = 32'b11111111111111101000001010000011;
assign LUT_2[54653] = 32'b11111111111111100101000010011100;
assign LUT_2[54654] = 32'b11111111111111101111000010111111;
assign LUT_2[54655] = 32'b11111111111111101011111011011000;
assign LUT_2[54656] = 32'b00000000000000000010000110110111;
assign LUT_2[54657] = 32'b11111111111111111110111111010000;
assign LUT_2[54658] = 32'b00000000000000001000111111110011;
assign LUT_2[54659] = 32'b00000000000000000101111000001100;
assign LUT_2[54660] = 32'b11111111111111111110100100011111;
assign LUT_2[54661] = 32'b11111111111111111011011100111000;
assign LUT_2[54662] = 32'b00000000000000000101011101011011;
assign LUT_2[54663] = 32'b00000000000000000010010101110100;
assign LUT_2[54664] = 32'b11111111111111111100111000010100;
assign LUT_2[54665] = 32'b11111111111111111001110000101101;
assign LUT_2[54666] = 32'b00000000000000000011110001010000;
assign LUT_2[54667] = 32'b00000000000000000000101001101001;
assign LUT_2[54668] = 32'b11111111111111111001010101111100;
assign LUT_2[54669] = 32'b11111111111111110110001110010101;
assign LUT_2[54670] = 32'b00000000000000000000001110111000;
assign LUT_2[54671] = 32'b11111111111111111101000111010001;
assign LUT_2[54672] = 32'b11111111111111111100101011000001;
assign LUT_2[54673] = 32'b11111111111111111001100011011010;
assign LUT_2[54674] = 32'b00000000000000000011100011111101;
assign LUT_2[54675] = 32'b00000000000000000000011100010110;
assign LUT_2[54676] = 32'b11111111111111111001001000101001;
assign LUT_2[54677] = 32'b11111111111111110110000001000010;
assign LUT_2[54678] = 32'b00000000000000000000000001100101;
assign LUT_2[54679] = 32'b11111111111111111100111001111110;
assign LUT_2[54680] = 32'b11111111111111110111011100011110;
assign LUT_2[54681] = 32'b11111111111111110100010100110111;
assign LUT_2[54682] = 32'b11111111111111111110010101011010;
assign LUT_2[54683] = 32'b11111111111111111011001101110011;
assign LUT_2[54684] = 32'b11111111111111110011111010000110;
assign LUT_2[54685] = 32'b11111111111111110000110010011111;
assign LUT_2[54686] = 32'b11111111111111111010110011000010;
assign LUT_2[54687] = 32'b11111111111111110111101011011011;
assign LUT_2[54688] = 32'b00000000000000000010100010100000;
assign LUT_2[54689] = 32'b11111111111111111111011010111001;
assign LUT_2[54690] = 32'b00000000000000001001011011011100;
assign LUT_2[54691] = 32'b00000000000000000110010011110101;
assign LUT_2[54692] = 32'b11111111111111111111000000001000;
assign LUT_2[54693] = 32'b11111111111111111011111000100001;
assign LUT_2[54694] = 32'b00000000000000000101111001000100;
assign LUT_2[54695] = 32'b00000000000000000010110001011101;
assign LUT_2[54696] = 32'b11111111111111111101010011111101;
assign LUT_2[54697] = 32'b11111111111111111010001100010110;
assign LUT_2[54698] = 32'b00000000000000000100001100111001;
assign LUT_2[54699] = 32'b00000000000000000001000101010010;
assign LUT_2[54700] = 32'b11111111111111111001110001100101;
assign LUT_2[54701] = 32'b11111111111111110110101001111110;
assign LUT_2[54702] = 32'b00000000000000000000101010100001;
assign LUT_2[54703] = 32'b11111111111111111101100010111010;
assign LUT_2[54704] = 32'b11111111111111111101000110101010;
assign LUT_2[54705] = 32'b11111111111111111001111111000011;
assign LUT_2[54706] = 32'b00000000000000000011111111100110;
assign LUT_2[54707] = 32'b00000000000000000000110111111111;
assign LUT_2[54708] = 32'b11111111111111111001100100010010;
assign LUT_2[54709] = 32'b11111111111111110110011100101011;
assign LUT_2[54710] = 32'b00000000000000000000011101001110;
assign LUT_2[54711] = 32'b11111111111111111101010101100111;
assign LUT_2[54712] = 32'b11111111111111110111111000000111;
assign LUT_2[54713] = 32'b11111111111111110100110000100000;
assign LUT_2[54714] = 32'b11111111111111111110110001000011;
assign LUT_2[54715] = 32'b11111111111111111011101001011100;
assign LUT_2[54716] = 32'b11111111111111110100010101101111;
assign LUT_2[54717] = 32'b11111111111111110001001110001000;
assign LUT_2[54718] = 32'b11111111111111111011001110101011;
assign LUT_2[54719] = 32'b11111111111111111000000111000100;
assign LUT_2[54720] = 32'b11111111111111111010001111011010;
assign LUT_2[54721] = 32'b11111111111111110111000111110011;
assign LUT_2[54722] = 32'b00000000000000000001001000010110;
assign LUT_2[54723] = 32'b11111111111111111110000000101111;
assign LUT_2[54724] = 32'b11111111111111110110101101000010;
assign LUT_2[54725] = 32'b11111111111111110011100101011011;
assign LUT_2[54726] = 32'b11111111111111111101100101111110;
assign LUT_2[54727] = 32'b11111111111111111010011110010111;
assign LUT_2[54728] = 32'b11111111111111110101000000110111;
assign LUT_2[54729] = 32'b11111111111111110001111001010000;
assign LUT_2[54730] = 32'b11111111111111111011111001110011;
assign LUT_2[54731] = 32'b11111111111111111000110010001100;
assign LUT_2[54732] = 32'b11111111111111110001011110011111;
assign LUT_2[54733] = 32'b11111111111111101110010110111000;
assign LUT_2[54734] = 32'b11111111111111111000010111011011;
assign LUT_2[54735] = 32'b11111111111111110101001111110100;
assign LUT_2[54736] = 32'b11111111111111110100110011100100;
assign LUT_2[54737] = 32'b11111111111111110001101011111101;
assign LUT_2[54738] = 32'b11111111111111111011101100100000;
assign LUT_2[54739] = 32'b11111111111111111000100100111001;
assign LUT_2[54740] = 32'b11111111111111110001010001001100;
assign LUT_2[54741] = 32'b11111111111111101110001001100101;
assign LUT_2[54742] = 32'b11111111111111111000001010001000;
assign LUT_2[54743] = 32'b11111111111111110101000010100001;
assign LUT_2[54744] = 32'b11111111111111101111100101000001;
assign LUT_2[54745] = 32'b11111111111111101100011101011010;
assign LUT_2[54746] = 32'b11111111111111110110011101111101;
assign LUT_2[54747] = 32'b11111111111111110011010110010110;
assign LUT_2[54748] = 32'b11111111111111101100000010101001;
assign LUT_2[54749] = 32'b11111111111111101000111011000010;
assign LUT_2[54750] = 32'b11111111111111110010111011100101;
assign LUT_2[54751] = 32'b11111111111111101111110011111110;
assign LUT_2[54752] = 32'b11111111111111111010101011000011;
assign LUT_2[54753] = 32'b11111111111111110111100011011100;
assign LUT_2[54754] = 32'b00000000000000000001100011111111;
assign LUT_2[54755] = 32'b11111111111111111110011100011000;
assign LUT_2[54756] = 32'b11111111111111110111001000101011;
assign LUT_2[54757] = 32'b11111111111111110100000001000100;
assign LUT_2[54758] = 32'b11111111111111111110000001100111;
assign LUT_2[54759] = 32'b11111111111111111010111010000000;
assign LUT_2[54760] = 32'b11111111111111110101011100100000;
assign LUT_2[54761] = 32'b11111111111111110010010100111001;
assign LUT_2[54762] = 32'b11111111111111111100010101011100;
assign LUT_2[54763] = 32'b11111111111111111001001101110101;
assign LUT_2[54764] = 32'b11111111111111110001111010001000;
assign LUT_2[54765] = 32'b11111111111111101110110010100001;
assign LUT_2[54766] = 32'b11111111111111111000110011000100;
assign LUT_2[54767] = 32'b11111111111111110101101011011101;
assign LUT_2[54768] = 32'b11111111111111110101001111001101;
assign LUT_2[54769] = 32'b11111111111111110010000111100110;
assign LUT_2[54770] = 32'b11111111111111111100001000001001;
assign LUT_2[54771] = 32'b11111111111111111001000000100010;
assign LUT_2[54772] = 32'b11111111111111110001101100110101;
assign LUT_2[54773] = 32'b11111111111111101110100101001110;
assign LUT_2[54774] = 32'b11111111111111111000100101110001;
assign LUT_2[54775] = 32'b11111111111111110101011110001010;
assign LUT_2[54776] = 32'b11111111111111110000000000101010;
assign LUT_2[54777] = 32'b11111111111111101100111001000011;
assign LUT_2[54778] = 32'b11111111111111110110111001100110;
assign LUT_2[54779] = 32'b11111111111111110011110001111111;
assign LUT_2[54780] = 32'b11111111111111101100011110010010;
assign LUT_2[54781] = 32'b11111111111111101001010110101011;
assign LUT_2[54782] = 32'b11111111111111110011010111001110;
assign LUT_2[54783] = 32'b11111111111111110000001111100111;
assign LUT_2[54784] = 32'b11111111111111111110100101110100;
assign LUT_2[54785] = 32'b11111111111111111011011110001101;
assign LUT_2[54786] = 32'b00000000000000000101011110110000;
assign LUT_2[54787] = 32'b00000000000000000010010111001001;
assign LUT_2[54788] = 32'b11111111111111111011000011011100;
assign LUT_2[54789] = 32'b11111111111111110111111011110101;
assign LUT_2[54790] = 32'b00000000000000000001111100011000;
assign LUT_2[54791] = 32'b11111111111111111110110100110001;
assign LUT_2[54792] = 32'b11111111111111111001010111010001;
assign LUT_2[54793] = 32'b11111111111111110110001111101010;
assign LUT_2[54794] = 32'b00000000000000000000010000001101;
assign LUT_2[54795] = 32'b11111111111111111101001000100110;
assign LUT_2[54796] = 32'b11111111111111110101110100111001;
assign LUT_2[54797] = 32'b11111111111111110010101101010010;
assign LUT_2[54798] = 32'b11111111111111111100101101110101;
assign LUT_2[54799] = 32'b11111111111111111001100110001110;
assign LUT_2[54800] = 32'b11111111111111111001001001111110;
assign LUT_2[54801] = 32'b11111111111111110110000010010111;
assign LUT_2[54802] = 32'b00000000000000000000000010111010;
assign LUT_2[54803] = 32'b11111111111111111100111011010011;
assign LUT_2[54804] = 32'b11111111111111110101100111100110;
assign LUT_2[54805] = 32'b11111111111111110010011111111111;
assign LUT_2[54806] = 32'b11111111111111111100100000100010;
assign LUT_2[54807] = 32'b11111111111111111001011000111011;
assign LUT_2[54808] = 32'b11111111111111110011111011011011;
assign LUT_2[54809] = 32'b11111111111111110000110011110100;
assign LUT_2[54810] = 32'b11111111111111111010110100010111;
assign LUT_2[54811] = 32'b11111111111111110111101100110000;
assign LUT_2[54812] = 32'b11111111111111110000011001000011;
assign LUT_2[54813] = 32'b11111111111111101101010001011100;
assign LUT_2[54814] = 32'b11111111111111110111010001111111;
assign LUT_2[54815] = 32'b11111111111111110100001010011000;
assign LUT_2[54816] = 32'b11111111111111111111000001011101;
assign LUT_2[54817] = 32'b11111111111111111011111001110110;
assign LUT_2[54818] = 32'b00000000000000000101111010011001;
assign LUT_2[54819] = 32'b00000000000000000010110010110010;
assign LUT_2[54820] = 32'b11111111111111111011011111000101;
assign LUT_2[54821] = 32'b11111111111111111000010111011110;
assign LUT_2[54822] = 32'b00000000000000000010011000000001;
assign LUT_2[54823] = 32'b11111111111111111111010000011010;
assign LUT_2[54824] = 32'b11111111111111111001110010111010;
assign LUT_2[54825] = 32'b11111111111111110110101011010011;
assign LUT_2[54826] = 32'b00000000000000000000101011110110;
assign LUT_2[54827] = 32'b11111111111111111101100100001111;
assign LUT_2[54828] = 32'b11111111111111110110010000100010;
assign LUT_2[54829] = 32'b11111111111111110011001000111011;
assign LUT_2[54830] = 32'b11111111111111111101001001011110;
assign LUT_2[54831] = 32'b11111111111111111010000001110111;
assign LUT_2[54832] = 32'b11111111111111111001100101100111;
assign LUT_2[54833] = 32'b11111111111111110110011110000000;
assign LUT_2[54834] = 32'b00000000000000000000011110100011;
assign LUT_2[54835] = 32'b11111111111111111101010110111100;
assign LUT_2[54836] = 32'b11111111111111110110000011001111;
assign LUT_2[54837] = 32'b11111111111111110010111011101000;
assign LUT_2[54838] = 32'b11111111111111111100111100001011;
assign LUT_2[54839] = 32'b11111111111111111001110100100100;
assign LUT_2[54840] = 32'b11111111111111110100010111000100;
assign LUT_2[54841] = 32'b11111111111111110001001111011101;
assign LUT_2[54842] = 32'b11111111111111111011010000000000;
assign LUT_2[54843] = 32'b11111111111111111000001000011001;
assign LUT_2[54844] = 32'b11111111111111110000110100101100;
assign LUT_2[54845] = 32'b11111111111111101101101101000101;
assign LUT_2[54846] = 32'b11111111111111110111101101101000;
assign LUT_2[54847] = 32'b11111111111111110100100110000001;
assign LUT_2[54848] = 32'b11111111111111110110101110010111;
assign LUT_2[54849] = 32'b11111111111111110011100110110000;
assign LUT_2[54850] = 32'b11111111111111111101100111010011;
assign LUT_2[54851] = 32'b11111111111111111010011111101100;
assign LUT_2[54852] = 32'b11111111111111110011001011111111;
assign LUT_2[54853] = 32'b11111111111111110000000100011000;
assign LUT_2[54854] = 32'b11111111111111111010000100111011;
assign LUT_2[54855] = 32'b11111111111111110110111101010100;
assign LUT_2[54856] = 32'b11111111111111110001011111110100;
assign LUT_2[54857] = 32'b11111111111111101110011000001101;
assign LUT_2[54858] = 32'b11111111111111111000011000110000;
assign LUT_2[54859] = 32'b11111111111111110101010001001001;
assign LUT_2[54860] = 32'b11111111111111101101111101011100;
assign LUT_2[54861] = 32'b11111111111111101010110101110101;
assign LUT_2[54862] = 32'b11111111111111110100110110011000;
assign LUT_2[54863] = 32'b11111111111111110001101110110001;
assign LUT_2[54864] = 32'b11111111111111110001010010100001;
assign LUT_2[54865] = 32'b11111111111111101110001010111010;
assign LUT_2[54866] = 32'b11111111111111111000001011011101;
assign LUT_2[54867] = 32'b11111111111111110101000011110110;
assign LUT_2[54868] = 32'b11111111111111101101110000001001;
assign LUT_2[54869] = 32'b11111111111111101010101000100010;
assign LUT_2[54870] = 32'b11111111111111110100101001000101;
assign LUT_2[54871] = 32'b11111111111111110001100001011110;
assign LUT_2[54872] = 32'b11111111111111101100000011111110;
assign LUT_2[54873] = 32'b11111111111111101000111100010111;
assign LUT_2[54874] = 32'b11111111111111110010111100111010;
assign LUT_2[54875] = 32'b11111111111111101111110101010011;
assign LUT_2[54876] = 32'b11111111111111101000100001100110;
assign LUT_2[54877] = 32'b11111111111111100101011001111111;
assign LUT_2[54878] = 32'b11111111111111101111011010100010;
assign LUT_2[54879] = 32'b11111111111111101100010010111011;
assign LUT_2[54880] = 32'b11111111111111110111001010000000;
assign LUT_2[54881] = 32'b11111111111111110100000010011001;
assign LUT_2[54882] = 32'b11111111111111111110000010111100;
assign LUT_2[54883] = 32'b11111111111111111010111011010101;
assign LUT_2[54884] = 32'b11111111111111110011100111101000;
assign LUT_2[54885] = 32'b11111111111111110000100000000001;
assign LUT_2[54886] = 32'b11111111111111111010100000100100;
assign LUT_2[54887] = 32'b11111111111111110111011000111101;
assign LUT_2[54888] = 32'b11111111111111110001111011011101;
assign LUT_2[54889] = 32'b11111111111111101110110011110110;
assign LUT_2[54890] = 32'b11111111111111111000110100011001;
assign LUT_2[54891] = 32'b11111111111111110101101100110010;
assign LUT_2[54892] = 32'b11111111111111101110011001000101;
assign LUT_2[54893] = 32'b11111111111111101011010001011110;
assign LUT_2[54894] = 32'b11111111111111110101010010000001;
assign LUT_2[54895] = 32'b11111111111111110010001010011010;
assign LUT_2[54896] = 32'b11111111111111110001101110001010;
assign LUT_2[54897] = 32'b11111111111111101110100110100011;
assign LUT_2[54898] = 32'b11111111111111111000100111000110;
assign LUT_2[54899] = 32'b11111111111111110101011111011111;
assign LUT_2[54900] = 32'b11111111111111101110001011110010;
assign LUT_2[54901] = 32'b11111111111111101011000100001011;
assign LUT_2[54902] = 32'b11111111111111110101000100101110;
assign LUT_2[54903] = 32'b11111111111111110001111101000111;
assign LUT_2[54904] = 32'b11111111111111101100011111100111;
assign LUT_2[54905] = 32'b11111111111111101001011000000000;
assign LUT_2[54906] = 32'b11111111111111110011011000100011;
assign LUT_2[54907] = 32'b11111111111111110000010000111100;
assign LUT_2[54908] = 32'b11111111111111101000111101001111;
assign LUT_2[54909] = 32'b11111111111111100101110101101000;
assign LUT_2[54910] = 32'b11111111111111101111110110001011;
assign LUT_2[54911] = 32'b11111111111111101100101110100100;
assign LUT_2[54912] = 32'b00000000000000000010111010000011;
assign LUT_2[54913] = 32'b11111111111111111111110010011100;
assign LUT_2[54914] = 32'b00000000000000001001110010111111;
assign LUT_2[54915] = 32'b00000000000000000110101011011000;
assign LUT_2[54916] = 32'b11111111111111111111010111101011;
assign LUT_2[54917] = 32'b11111111111111111100010000000100;
assign LUT_2[54918] = 32'b00000000000000000110010000100111;
assign LUT_2[54919] = 32'b00000000000000000011001001000000;
assign LUT_2[54920] = 32'b11111111111111111101101011100000;
assign LUT_2[54921] = 32'b11111111111111111010100011111001;
assign LUT_2[54922] = 32'b00000000000000000100100100011100;
assign LUT_2[54923] = 32'b00000000000000000001011100110101;
assign LUT_2[54924] = 32'b11111111111111111010001001001000;
assign LUT_2[54925] = 32'b11111111111111110111000001100001;
assign LUT_2[54926] = 32'b00000000000000000001000010000100;
assign LUT_2[54927] = 32'b11111111111111111101111010011101;
assign LUT_2[54928] = 32'b11111111111111111101011110001101;
assign LUT_2[54929] = 32'b11111111111111111010010110100110;
assign LUT_2[54930] = 32'b00000000000000000100010111001001;
assign LUT_2[54931] = 32'b00000000000000000001001111100010;
assign LUT_2[54932] = 32'b11111111111111111001111011110101;
assign LUT_2[54933] = 32'b11111111111111110110110100001110;
assign LUT_2[54934] = 32'b00000000000000000000110100110001;
assign LUT_2[54935] = 32'b11111111111111111101101101001010;
assign LUT_2[54936] = 32'b11111111111111111000001111101010;
assign LUT_2[54937] = 32'b11111111111111110101001000000011;
assign LUT_2[54938] = 32'b11111111111111111111001000100110;
assign LUT_2[54939] = 32'b11111111111111111100000000111111;
assign LUT_2[54940] = 32'b11111111111111110100101101010010;
assign LUT_2[54941] = 32'b11111111111111110001100101101011;
assign LUT_2[54942] = 32'b11111111111111111011100110001110;
assign LUT_2[54943] = 32'b11111111111111111000011110100111;
assign LUT_2[54944] = 32'b00000000000000000011010101101100;
assign LUT_2[54945] = 32'b00000000000000000000001110000101;
assign LUT_2[54946] = 32'b00000000000000001010001110101000;
assign LUT_2[54947] = 32'b00000000000000000111000111000001;
assign LUT_2[54948] = 32'b11111111111111111111110011010100;
assign LUT_2[54949] = 32'b11111111111111111100101011101101;
assign LUT_2[54950] = 32'b00000000000000000110101100010000;
assign LUT_2[54951] = 32'b00000000000000000011100100101001;
assign LUT_2[54952] = 32'b11111111111111111110000111001001;
assign LUT_2[54953] = 32'b11111111111111111010111111100010;
assign LUT_2[54954] = 32'b00000000000000000101000000000101;
assign LUT_2[54955] = 32'b00000000000000000001111000011110;
assign LUT_2[54956] = 32'b11111111111111111010100100110001;
assign LUT_2[54957] = 32'b11111111111111110111011101001010;
assign LUT_2[54958] = 32'b00000000000000000001011101101101;
assign LUT_2[54959] = 32'b11111111111111111110010110000110;
assign LUT_2[54960] = 32'b11111111111111111101111001110110;
assign LUT_2[54961] = 32'b11111111111111111010110010001111;
assign LUT_2[54962] = 32'b00000000000000000100110010110010;
assign LUT_2[54963] = 32'b00000000000000000001101011001011;
assign LUT_2[54964] = 32'b11111111111111111010010111011110;
assign LUT_2[54965] = 32'b11111111111111110111001111110111;
assign LUT_2[54966] = 32'b00000000000000000001010000011010;
assign LUT_2[54967] = 32'b11111111111111111110001000110011;
assign LUT_2[54968] = 32'b11111111111111111000101011010011;
assign LUT_2[54969] = 32'b11111111111111110101100011101100;
assign LUT_2[54970] = 32'b11111111111111111111100100001111;
assign LUT_2[54971] = 32'b11111111111111111100011100101000;
assign LUT_2[54972] = 32'b11111111111111110101001000111011;
assign LUT_2[54973] = 32'b11111111111111110010000001010100;
assign LUT_2[54974] = 32'b11111111111111111100000001110111;
assign LUT_2[54975] = 32'b11111111111111111000111010010000;
assign LUT_2[54976] = 32'b11111111111111111011000010100110;
assign LUT_2[54977] = 32'b11111111111111110111111010111111;
assign LUT_2[54978] = 32'b00000000000000000001111011100010;
assign LUT_2[54979] = 32'b11111111111111111110110011111011;
assign LUT_2[54980] = 32'b11111111111111110111100000001110;
assign LUT_2[54981] = 32'b11111111111111110100011000100111;
assign LUT_2[54982] = 32'b11111111111111111110011001001010;
assign LUT_2[54983] = 32'b11111111111111111011010001100011;
assign LUT_2[54984] = 32'b11111111111111110101110100000011;
assign LUT_2[54985] = 32'b11111111111111110010101100011100;
assign LUT_2[54986] = 32'b11111111111111111100101100111111;
assign LUT_2[54987] = 32'b11111111111111111001100101011000;
assign LUT_2[54988] = 32'b11111111111111110010010001101011;
assign LUT_2[54989] = 32'b11111111111111101111001010000100;
assign LUT_2[54990] = 32'b11111111111111111001001010100111;
assign LUT_2[54991] = 32'b11111111111111110110000011000000;
assign LUT_2[54992] = 32'b11111111111111110101100110110000;
assign LUT_2[54993] = 32'b11111111111111110010011111001001;
assign LUT_2[54994] = 32'b11111111111111111100011111101100;
assign LUT_2[54995] = 32'b11111111111111111001011000000101;
assign LUT_2[54996] = 32'b11111111111111110010000100011000;
assign LUT_2[54997] = 32'b11111111111111101110111100110001;
assign LUT_2[54998] = 32'b11111111111111111000111101010100;
assign LUT_2[54999] = 32'b11111111111111110101110101101101;
assign LUT_2[55000] = 32'b11111111111111110000011000001101;
assign LUT_2[55001] = 32'b11111111111111101101010000100110;
assign LUT_2[55002] = 32'b11111111111111110111010001001001;
assign LUT_2[55003] = 32'b11111111111111110100001001100010;
assign LUT_2[55004] = 32'b11111111111111101100110101110101;
assign LUT_2[55005] = 32'b11111111111111101001101110001110;
assign LUT_2[55006] = 32'b11111111111111110011101110110001;
assign LUT_2[55007] = 32'b11111111111111110000100111001010;
assign LUT_2[55008] = 32'b11111111111111111011011110001111;
assign LUT_2[55009] = 32'b11111111111111111000010110101000;
assign LUT_2[55010] = 32'b00000000000000000010010111001011;
assign LUT_2[55011] = 32'b11111111111111111111001111100100;
assign LUT_2[55012] = 32'b11111111111111110111111011110111;
assign LUT_2[55013] = 32'b11111111111111110100110100010000;
assign LUT_2[55014] = 32'b11111111111111111110110100110011;
assign LUT_2[55015] = 32'b11111111111111111011101101001100;
assign LUT_2[55016] = 32'b11111111111111110110001111101100;
assign LUT_2[55017] = 32'b11111111111111110011001000000101;
assign LUT_2[55018] = 32'b11111111111111111101001000101000;
assign LUT_2[55019] = 32'b11111111111111111010000001000001;
assign LUT_2[55020] = 32'b11111111111111110010101101010100;
assign LUT_2[55021] = 32'b11111111111111101111100101101101;
assign LUT_2[55022] = 32'b11111111111111111001100110010000;
assign LUT_2[55023] = 32'b11111111111111110110011110101001;
assign LUT_2[55024] = 32'b11111111111111110110000010011001;
assign LUT_2[55025] = 32'b11111111111111110010111010110010;
assign LUT_2[55026] = 32'b11111111111111111100111011010101;
assign LUT_2[55027] = 32'b11111111111111111001110011101110;
assign LUT_2[55028] = 32'b11111111111111110010100000000001;
assign LUT_2[55029] = 32'b11111111111111101111011000011010;
assign LUT_2[55030] = 32'b11111111111111111001011000111101;
assign LUT_2[55031] = 32'b11111111111111110110010001010110;
assign LUT_2[55032] = 32'b11111111111111110000110011110110;
assign LUT_2[55033] = 32'b11111111111111101101101100001111;
assign LUT_2[55034] = 32'b11111111111111110111101100110010;
assign LUT_2[55035] = 32'b11111111111111110100100101001011;
assign LUT_2[55036] = 32'b11111111111111101101010001011110;
assign LUT_2[55037] = 32'b11111111111111101010001001110111;
assign LUT_2[55038] = 32'b11111111111111110100001010011010;
assign LUT_2[55039] = 32'b11111111111111110001000010110011;
assign LUT_2[55040] = 32'b00000000000000000010100100011010;
assign LUT_2[55041] = 32'b11111111111111111111011100110011;
assign LUT_2[55042] = 32'b00000000000000001001011101010110;
assign LUT_2[55043] = 32'b00000000000000000110010101101111;
assign LUT_2[55044] = 32'b11111111111111111111000010000010;
assign LUT_2[55045] = 32'b11111111111111111011111010011011;
assign LUT_2[55046] = 32'b00000000000000000101111010111110;
assign LUT_2[55047] = 32'b00000000000000000010110011010111;
assign LUT_2[55048] = 32'b11111111111111111101010101110111;
assign LUT_2[55049] = 32'b11111111111111111010001110010000;
assign LUT_2[55050] = 32'b00000000000000000100001110110011;
assign LUT_2[55051] = 32'b00000000000000000001000111001100;
assign LUT_2[55052] = 32'b11111111111111111001110011011111;
assign LUT_2[55053] = 32'b11111111111111110110101011111000;
assign LUT_2[55054] = 32'b00000000000000000000101100011011;
assign LUT_2[55055] = 32'b11111111111111111101100100110100;
assign LUT_2[55056] = 32'b11111111111111111101001000100100;
assign LUT_2[55057] = 32'b11111111111111111010000000111101;
assign LUT_2[55058] = 32'b00000000000000000100000001100000;
assign LUT_2[55059] = 32'b00000000000000000000111001111001;
assign LUT_2[55060] = 32'b11111111111111111001100110001100;
assign LUT_2[55061] = 32'b11111111111111110110011110100101;
assign LUT_2[55062] = 32'b00000000000000000000011111001000;
assign LUT_2[55063] = 32'b11111111111111111101010111100001;
assign LUT_2[55064] = 32'b11111111111111110111111010000001;
assign LUT_2[55065] = 32'b11111111111111110100110010011010;
assign LUT_2[55066] = 32'b11111111111111111110110010111101;
assign LUT_2[55067] = 32'b11111111111111111011101011010110;
assign LUT_2[55068] = 32'b11111111111111110100010111101001;
assign LUT_2[55069] = 32'b11111111111111110001010000000010;
assign LUT_2[55070] = 32'b11111111111111111011010000100101;
assign LUT_2[55071] = 32'b11111111111111111000001000111110;
assign LUT_2[55072] = 32'b00000000000000000011000000000011;
assign LUT_2[55073] = 32'b11111111111111111111111000011100;
assign LUT_2[55074] = 32'b00000000000000001001111000111111;
assign LUT_2[55075] = 32'b00000000000000000110110001011000;
assign LUT_2[55076] = 32'b11111111111111111111011101101011;
assign LUT_2[55077] = 32'b11111111111111111100010110000100;
assign LUT_2[55078] = 32'b00000000000000000110010110100111;
assign LUT_2[55079] = 32'b00000000000000000011001111000000;
assign LUT_2[55080] = 32'b11111111111111111101110001100000;
assign LUT_2[55081] = 32'b11111111111111111010101001111001;
assign LUT_2[55082] = 32'b00000000000000000100101010011100;
assign LUT_2[55083] = 32'b00000000000000000001100010110101;
assign LUT_2[55084] = 32'b11111111111111111010001111001000;
assign LUT_2[55085] = 32'b11111111111111110111000111100001;
assign LUT_2[55086] = 32'b00000000000000000001001000000100;
assign LUT_2[55087] = 32'b11111111111111111110000000011101;
assign LUT_2[55088] = 32'b11111111111111111101100100001101;
assign LUT_2[55089] = 32'b11111111111111111010011100100110;
assign LUT_2[55090] = 32'b00000000000000000100011101001001;
assign LUT_2[55091] = 32'b00000000000000000001010101100010;
assign LUT_2[55092] = 32'b11111111111111111010000001110101;
assign LUT_2[55093] = 32'b11111111111111110110111010001110;
assign LUT_2[55094] = 32'b00000000000000000000111010110001;
assign LUT_2[55095] = 32'b11111111111111111101110011001010;
assign LUT_2[55096] = 32'b11111111111111111000010101101010;
assign LUT_2[55097] = 32'b11111111111111110101001110000011;
assign LUT_2[55098] = 32'b11111111111111111111001110100110;
assign LUT_2[55099] = 32'b11111111111111111100000110111111;
assign LUT_2[55100] = 32'b11111111111111110100110011010010;
assign LUT_2[55101] = 32'b11111111111111110001101011101011;
assign LUT_2[55102] = 32'b11111111111111111011101100001110;
assign LUT_2[55103] = 32'b11111111111111111000100100100111;
assign LUT_2[55104] = 32'b11111111111111111010101100111101;
assign LUT_2[55105] = 32'b11111111111111110111100101010110;
assign LUT_2[55106] = 32'b00000000000000000001100101111001;
assign LUT_2[55107] = 32'b11111111111111111110011110010010;
assign LUT_2[55108] = 32'b11111111111111110111001010100101;
assign LUT_2[55109] = 32'b11111111111111110100000010111110;
assign LUT_2[55110] = 32'b11111111111111111110000011100001;
assign LUT_2[55111] = 32'b11111111111111111010111011111010;
assign LUT_2[55112] = 32'b11111111111111110101011110011010;
assign LUT_2[55113] = 32'b11111111111111110010010110110011;
assign LUT_2[55114] = 32'b11111111111111111100010111010110;
assign LUT_2[55115] = 32'b11111111111111111001001111101111;
assign LUT_2[55116] = 32'b11111111111111110001111100000010;
assign LUT_2[55117] = 32'b11111111111111101110110100011011;
assign LUT_2[55118] = 32'b11111111111111111000110100111110;
assign LUT_2[55119] = 32'b11111111111111110101101101010111;
assign LUT_2[55120] = 32'b11111111111111110101010001000111;
assign LUT_2[55121] = 32'b11111111111111110010001001100000;
assign LUT_2[55122] = 32'b11111111111111111100001010000011;
assign LUT_2[55123] = 32'b11111111111111111001000010011100;
assign LUT_2[55124] = 32'b11111111111111110001101110101111;
assign LUT_2[55125] = 32'b11111111111111101110100111001000;
assign LUT_2[55126] = 32'b11111111111111111000100111101011;
assign LUT_2[55127] = 32'b11111111111111110101100000000100;
assign LUT_2[55128] = 32'b11111111111111110000000010100100;
assign LUT_2[55129] = 32'b11111111111111101100111010111101;
assign LUT_2[55130] = 32'b11111111111111110110111011100000;
assign LUT_2[55131] = 32'b11111111111111110011110011111001;
assign LUT_2[55132] = 32'b11111111111111101100100000001100;
assign LUT_2[55133] = 32'b11111111111111101001011000100101;
assign LUT_2[55134] = 32'b11111111111111110011011001001000;
assign LUT_2[55135] = 32'b11111111111111110000010001100001;
assign LUT_2[55136] = 32'b11111111111111111011001000100110;
assign LUT_2[55137] = 32'b11111111111111111000000000111111;
assign LUT_2[55138] = 32'b00000000000000000010000001100010;
assign LUT_2[55139] = 32'b11111111111111111110111001111011;
assign LUT_2[55140] = 32'b11111111111111110111100110001110;
assign LUT_2[55141] = 32'b11111111111111110100011110100111;
assign LUT_2[55142] = 32'b11111111111111111110011111001010;
assign LUT_2[55143] = 32'b11111111111111111011010111100011;
assign LUT_2[55144] = 32'b11111111111111110101111010000011;
assign LUT_2[55145] = 32'b11111111111111110010110010011100;
assign LUT_2[55146] = 32'b11111111111111111100110010111111;
assign LUT_2[55147] = 32'b11111111111111111001101011011000;
assign LUT_2[55148] = 32'b11111111111111110010010111101011;
assign LUT_2[55149] = 32'b11111111111111101111010000000100;
assign LUT_2[55150] = 32'b11111111111111111001010000100111;
assign LUT_2[55151] = 32'b11111111111111110110001001000000;
assign LUT_2[55152] = 32'b11111111111111110101101100110000;
assign LUT_2[55153] = 32'b11111111111111110010100101001001;
assign LUT_2[55154] = 32'b11111111111111111100100101101100;
assign LUT_2[55155] = 32'b11111111111111111001011110000101;
assign LUT_2[55156] = 32'b11111111111111110010001010011000;
assign LUT_2[55157] = 32'b11111111111111101111000010110001;
assign LUT_2[55158] = 32'b11111111111111111001000011010100;
assign LUT_2[55159] = 32'b11111111111111110101111011101101;
assign LUT_2[55160] = 32'b11111111111111110000011110001101;
assign LUT_2[55161] = 32'b11111111111111101101010110100110;
assign LUT_2[55162] = 32'b11111111111111110111010111001001;
assign LUT_2[55163] = 32'b11111111111111110100001111100010;
assign LUT_2[55164] = 32'b11111111111111101100111011110101;
assign LUT_2[55165] = 32'b11111111111111101001110100001110;
assign LUT_2[55166] = 32'b11111111111111110011110100110001;
assign LUT_2[55167] = 32'b11111111111111110000101101001010;
assign LUT_2[55168] = 32'b00000000000000000110111000101001;
assign LUT_2[55169] = 32'b00000000000000000011110001000010;
assign LUT_2[55170] = 32'b00000000000000001101110001100101;
assign LUT_2[55171] = 32'b00000000000000001010101001111110;
assign LUT_2[55172] = 32'b00000000000000000011010110010001;
assign LUT_2[55173] = 32'b00000000000000000000001110101010;
assign LUT_2[55174] = 32'b00000000000000001010001111001101;
assign LUT_2[55175] = 32'b00000000000000000111000111100110;
assign LUT_2[55176] = 32'b00000000000000000001101010000110;
assign LUT_2[55177] = 32'b11111111111111111110100010011111;
assign LUT_2[55178] = 32'b00000000000000001000100011000010;
assign LUT_2[55179] = 32'b00000000000000000101011011011011;
assign LUT_2[55180] = 32'b11111111111111111110000111101110;
assign LUT_2[55181] = 32'b11111111111111111011000000000111;
assign LUT_2[55182] = 32'b00000000000000000101000000101010;
assign LUT_2[55183] = 32'b00000000000000000001111001000011;
assign LUT_2[55184] = 32'b00000000000000000001011100110011;
assign LUT_2[55185] = 32'b11111111111111111110010101001100;
assign LUT_2[55186] = 32'b00000000000000001000010101101111;
assign LUT_2[55187] = 32'b00000000000000000101001110001000;
assign LUT_2[55188] = 32'b11111111111111111101111010011011;
assign LUT_2[55189] = 32'b11111111111111111010110010110100;
assign LUT_2[55190] = 32'b00000000000000000100110011010111;
assign LUT_2[55191] = 32'b00000000000000000001101011110000;
assign LUT_2[55192] = 32'b11111111111111111100001110010000;
assign LUT_2[55193] = 32'b11111111111111111001000110101001;
assign LUT_2[55194] = 32'b00000000000000000011000111001100;
assign LUT_2[55195] = 32'b11111111111111111111111111100101;
assign LUT_2[55196] = 32'b11111111111111111000101011111000;
assign LUT_2[55197] = 32'b11111111111111110101100100010001;
assign LUT_2[55198] = 32'b11111111111111111111100100110100;
assign LUT_2[55199] = 32'b11111111111111111100011101001101;
assign LUT_2[55200] = 32'b00000000000000000111010100010010;
assign LUT_2[55201] = 32'b00000000000000000100001100101011;
assign LUT_2[55202] = 32'b00000000000000001110001101001110;
assign LUT_2[55203] = 32'b00000000000000001011000101100111;
assign LUT_2[55204] = 32'b00000000000000000011110001111010;
assign LUT_2[55205] = 32'b00000000000000000000101010010011;
assign LUT_2[55206] = 32'b00000000000000001010101010110110;
assign LUT_2[55207] = 32'b00000000000000000111100011001111;
assign LUT_2[55208] = 32'b00000000000000000010000101101111;
assign LUT_2[55209] = 32'b11111111111111111110111110001000;
assign LUT_2[55210] = 32'b00000000000000001000111110101011;
assign LUT_2[55211] = 32'b00000000000000000101110111000100;
assign LUT_2[55212] = 32'b11111111111111111110100011010111;
assign LUT_2[55213] = 32'b11111111111111111011011011110000;
assign LUT_2[55214] = 32'b00000000000000000101011100010011;
assign LUT_2[55215] = 32'b00000000000000000010010100101100;
assign LUT_2[55216] = 32'b00000000000000000001111000011100;
assign LUT_2[55217] = 32'b11111111111111111110110000110101;
assign LUT_2[55218] = 32'b00000000000000001000110001011000;
assign LUT_2[55219] = 32'b00000000000000000101101001110001;
assign LUT_2[55220] = 32'b11111111111111111110010110000100;
assign LUT_2[55221] = 32'b11111111111111111011001110011101;
assign LUT_2[55222] = 32'b00000000000000000101001111000000;
assign LUT_2[55223] = 32'b00000000000000000010000111011001;
assign LUT_2[55224] = 32'b11111111111111111100101001111001;
assign LUT_2[55225] = 32'b11111111111111111001100010010010;
assign LUT_2[55226] = 32'b00000000000000000011100010110101;
assign LUT_2[55227] = 32'b00000000000000000000011011001110;
assign LUT_2[55228] = 32'b11111111111111111001000111100001;
assign LUT_2[55229] = 32'b11111111111111110101111111111010;
assign LUT_2[55230] = 32'b00000000000000000000000000011101;
assign LUT_2[55231] = 32'b11111111111111111100111000110110;
assign LUT_2[55232] = 32'b11111111111111111111000001001100;
assign LUT_2[55233] = 32'b11111111111111111011111001100101;
assign LUT_2[55234] = 32'b00000000000000000101111010001000;
assign LUT_2[55235] = 32'b00000000000000000010110010100001;
assign LUT_2[55236] = 32'b11111111111111111011011110110100;
assign LUT_2[55237] = 32'b11111111111111111000010111001101;
assign LUT_2[55238] = 32'b00000000000000000010010111110000;
assign LUT_2[55239] = 32'b11111111111111111111010000001001;
assign LUT_2[55240] = 32'b11111111111111111001110010101001;
assign LUT_2[55241] = 32'b11111111111111110110101011000010;
assign LUT_2[55242] = 32'b00000000000000000000101011100101;
assign LUT_2[55243] = 32'b11111111111111111101100011111110;
assign LUT_2[55244] = 32'b11111111111111110110010000010001;
assign LUT_2[55245] = 32'b11111111111111110011001000101010;
assign LUT_2[55246] = 32'b11111111111111111101001001001101;
assign LUT_2[55247] = 32'b11111111111111111010000001100110;
assign LUT_2[55248] = 32'b11111111111111111001100101010110;
assign LUT_2[55249] = 32'b11111111111111110110011101101111;
assign LUT_2[55250] = 32'b00000000000000000000011110010010;
assign LUT_2[55251] = 32'b11111111111111111101010110101011;
assign LUT_2[55252] = 32'b11111111111111110110000010111110;
assign LUT_2[55253] = 32'b11111111111111110010111011010111;
assign LUT_2[55254] = 32'b11111111111111111100111011111010;
assign LUT_2[55255] = 32'b11111111111111111001110100010011;
assign LUT_2[55256] = 32'b11111111111111110100010110110011;
assign LUT_2[55257] = 32'b11111111111111110001001111001100;
assign LUT_2[55258] = 32'b11111111111111111011001111101111;
assign LUT_2[55259] = 32'b11111111111111111000001000001000;
assign LUT_2[55260] = 32'b11111111111111110000110100011011;
assign LUT_2[55261] = 32'b11111111111111101101101100110100;
assign LUT_2[55262] = 32'b11111111111111110111101101010111;
assign LUT_2[55263] = 32'b11111111111111110100100101110000;
assign LUT_2[55264] = 32'b11111111111111111111011100110101;
assign LUT_2[55265] = 32'b11111111111111111100010101001110;
assign LUT_2[55266] = 32'b00000000000000000110010101110001;
assign LUT_2[55267] = 32'b00000000000000000011001110001010;
assign LUT_2[55268] = 32'b11111111111111111011111010011101;
assign LUT_2[55269] = 32'b11111111111111111000110010110110;
assign LUT_2[55270] = 32'b00000000000000000010110011011001;
assign LUT_2[55271] = 32'b11111111111111111111101011110010;
assign LUT_2[55272] = 32'b11111111111111111010001110010010;
assign LUT_2[55273] = 32'b11111111111111110111000110101011;
assign LUT_2[55274] = 32'b00000000000000000001000111001110;
assign LUT_2[55275] = 32'b11111111111111111101111111100111;
assign LUT_2[55276] = 32'b11111111111111110110101011111010;
assign LUT_2[55277] = 32'b11111111111111110011100100010011;
assign LUT_2[55278] = 32'b11111111111111111101100100110110;
assign LUT_2[55279] = 32'b11111111111111111010011101001111;
assign LUT_2[55280] = 32'b11111111111111111010000000111111;
assign LUT_2[55281] = 32'b11111111111111110110111001011000;
assign LUT_2[55282] = 32'b00000000000000000000111001111011;
assign LUT_2[55283] = 32'b11111111111111111101110010010100;
assign LUT_2[55284] = 32'b11111111111111110110011110100111;
assign LUT_2[55285] = 32'b11111111111111110011010111000000;
assign LUT_2[55286] = 32'b11111111111111111101010111100011;
assign LUT_2[55287] = 32'b11111111111111111010001111111100;
assign LUT_2[55288] = 32'b11111111111111110100110010011100;
assign LUT_2[55289] = 32'b11111111111111110001101010110101;
assign LUT_2[55290] = 32'b11111111111111111011101011011000;
assign LUT_2[55291] = 32'b11111111111111111000100011110001;
assign LUT_2[55292] = 32'b11111111111111110001010000000100;
assign LUT_2[55293] = 32'b11111111111111101110001000011101;
assign LUT_2[55294] = 32'b11111111111111111000001001000000;
assign LUT_2[55295] = 32'b11111111111111110101000001011001;
assign LUT_2[55296] = 32'b11111111111111101110111101111001;
assign LUT_2[55297] = 32'b11111111111111101011110110010010;
assign LUT_2[55298] = 32'b11111111111111110101110110110101;
assign LUT_2[55299] = 32'b11111111111111110010101111001110;
assign LUT_2[55300] = 32'b11111111111111101011011011100001;
assign LUT_2[55301] = 32'b11111111111111101000010011111010;
assign LUT_2[55302] = 32'b11111111111111110010010100011101;
assign LUT_2[55303] = 32'b11111111111111101111001100110110;
assign LUT_2[55304] = 32'b11111111111111101001101111010110;
assign LUT_2[55305] = 32'b11111111111111100110100111101111;
assign LUT_2[55306] = 32'b11111111111111110000101000010010;
assign LUT_2[55307] = 32'b11111111111111101101100000101011;
assign LUT_2[55308] = 32'b11111111111111100110001100111110;
assign LUT_2[55309] = 32'b11111111111111100011000101010111;
assign LUT_2[55310] = 32'b11111111111111101101000101111010;
assign LUT_2[55311] = 32'b11111111111111101001111110010011;
assign LUT_2[55312] = 32'b11111111111111101001100010000011;
assign LUT_2[55313] = 32'b11111111111111100110011010011100;
assign LUT_2[55314] = 32'b11111111111111110000011010111111;
assign LUT_2[55315] = 32'b11111111111111101101010011011000;
assign LUT_2[55316] = 32'b11111111111111100101111111101011;
assign LUT_2[55317] = 32'b11111111111111100010111000000100;
assign LUT_2[55318] = 32'b11111111111111101100111000100111;
assign LUT_2[55319] = 32'b11111111111111101001110001000000;
assign LUT_2[55320] = 32'b11111111111111100100010011100000;
assign LUT_2[55321] = 32'b11111111111111100001001011111001;
assign LUT_2[55322] = 32'b11111111111111101011001100011100;
assign LUT_2[55323] = 32'b11111111111111101000000100110101;
assign LUT_2[55324] = 32'b11111111111111100000110001001000;
assign LUT_2[55325] = 32'b11111111111111011101101001100001;
assign LUT_2[55326] = 32'b11111111111111100111101010000100;
assign LUT_2[55327] = 32'b11111111111111100100100010011101;
assign LUT_2[55328] = 32'b11111111111111101111011001100010;
assign LUT_2[55329] = 32'b11111111111111101100010001111011;
assign LUT_2[55330] = 32'b11111111111111110110010010011110;
assign LUT_2[55331] = 32'b11111111111111110011001010110111;
assign LUT_2[55332] = 32'b11111111111111101011110111001010;
assign LUT_2[55333] = 32'b11111111111111101000101111100011;
assign LUT_2[55334] = 32'b11111111111111110010110000000110;
assign LUT_2[55335] = 32'b11111111111111101111101000011111;
assign LUT_2[55336] = 32'b11111111111111101010001010111111;
assign LUT_2[55337] = 32'b11111111111111100111000011011000;
assign LUT_2[55338] = 32'b11111111111111110001000011111011;
assign LUT_2[55339] = 32'b11111111111111101101111100010100;
assign LUT_2[55340] = 32'b11111111111111100110101000100111;
assign LUT_2[55341] = 32'b11111111111111100011100001000000;
assign LUT_2[55342] = 32'b11111111111111101101100001100011;
assign LUT_2[55343] = 32'b11111111111111101010011001111100;
assign LUT_2[55344] = 32'b11111111111111101001111101101100;
assign LUT_2[55345] = 32'b11111111111111100110110110000101;
assign LUT_2[55346] = 32'b11111111111111110000110110101000;
assign LUT_2[55347] = 32'b11111111111111101101101111000001;
assign LUT_2[55348] = 32'b11111111111111100110011011010100;
assign LUT_2[55349] = 32'b11111111111111100011010011101101;
assign LUT_2[55350] = 32'b11111111111111101101010100010000;
assign LUT_2[55351] = 32'b11111111111111101010001100101001;
assign LUT_2[55352] = 32'b11111111111111100100101111001001;
assign LUT_2[55353] = 32'b11111111111111100001100111100010;
assign LUT_2[55354] = 32'b11111111111111101011101000000101;
assign LUT_2[55355] = 32'b11111111111111101000100000011110;
assign LUT_2[55356] = 32'b11111111111111100001001100110001;
assign LUT_2[55357] = 32'b11111111111111011110000101001010;
assign LUT_2[55358] = 32'b11111111111111101000000101101101;
assign LUT_2[55359] = 32'b11111111111111100100111110000110;
assign LUT_2[55360] = 32'b11111111111111100111000110011100;
assign LUT_2[55361] = 32'b11111111111111100011111110110101;
assign LUT_2[55362] = 32'b11111111111111101101111111011000;
assign LUT_2[55363] = 32'b11111111111111101010110111110001;
assign LUT_2[55364] = 32'b11111111111111100011100100000100;
assign LUT_2[55365] = 32'b11111111111111100000011100011101;
assign LUT_2[55366] = 32'b11111111111111101010011101000000;
assign LUT_2[55367] = 32'b11111111111111100111010101011001;
assign LUT_2[55368] = 32'b11111111111111100001110111111001;
assign LUT_2[55369] = 32'b11111111111111011110110000010010;
assign LUT_2[55370] = 32'b11111111111111101000110000110101;
assign LUT_2[55371] = 32'b11111111111111100101101001001110;
assign LUT_2[55372] = 32'b11111111111111011110010101100001;
assign LUT_2[55373] = 32'b11111111111111011011001101111010;
assign LUT_2[55374] = 32'b11111111111111100101001110011101;
assign LUT_2[55375] = 32'b11111111111111100010000110110110;
assign LUT_2[55376] = 32'b11111111111111100001101010100110;
assign LUT_2[55377] = 32'b11111111111111011110100010111111;
assign LUT_2[55378] = 32'b11111111111111101000100011100010;
assign LUT_2[55379] = 32'b11111111111111100101011011111011;
assign LUT_2[55380] = 32'b11111111111111011110001000001110;
assign LUT_2[55381] = 32'b11111111111111011011000000100111;
assign LUT_2[55382] = 32'b11111111111111100101000001001010;
assign LUT_2[55383] = 32'b11111111111111100001111001100011;
assign LUT_2[55384] = 32'b11111111111111011100011100000011;
assign LUT_2[55385] = 32'b11111111111111011001010100011100;
assign LUT_2[55386] = 32'b11111111111111100011010100111111;
assign LUT_2[55387] = 32'b11111111111111100000001101011000;
assign LUT_2[55388] = 32'b11111111111111011000111001101011;
assign LUT_2[55389] = 32'b11111111111111010101110010000100;
assign LUT_2[55390] = 32'b11111111111111011111110010100111;
assign LUT_2[55391] = 32'b11111111111111011100101011000000;
assign LUT_2[55392] = 32'b11111111111111100111100010000101;
assign LUT_2[55393] = 32'b11111111111111100100011010011110;
assign LUT_2[55394] = 32'b11111111111111101110011011000001;
assign LUT_2[55395] = 32'b11111111111111101011010011011010;
assign LUT_2[55396] = 32'b11111111111111100011111111101101;
assign LUT_2[55397] = 32'b11111111111111100000111000000110;
assign LUT_2[55398] = 32'b11111111111111101010111000101001;
assign LUT_2[55399] = 32'b11111111111111100111110001000010;
assign LUT_2[55400] = 32'b11111111111111100010010011100010;
assign LUT_2[55401] = 32'b11111111111111011111001011111011;
assign LUT_2[55402] = 32'b11111111111111101001001100011110;
assign LUT_2[55403] = 32'b11111111111111100110000100110111;
assign LUT_2[55404] = 32'b11111111111111011110110001001010;
assign LUT_2[55405] = 32'b11111111111111011011101001100011;
assign LUT_2[55406] = 32'b11111111111111100101101010000110;
assign LUT_2[55407] = 32'b11111111111111100010100010011111;
assign LUT_2[55408] = 32'b11111111111111100010000110001111;
assign LUT_2[55409] = 32'b11111111111111011110111110101000;
assign LUT_2[55410] = 32'b11111111111111101000111111001011;
assign LUT_2[55411] = 32'b11111111111111100101110111100100;
assign LUT_2[55412] = 32'b11111111111111011110100011110111;
assign LUT_2[55413] = 32'b11111111111111011011011100010000;
assign LUT_2[55414] = 32'b11111111111111100101011100110011;
assign LUT_2[55415] = 32'b11111111111111100010010101001100;
assign LUT_2[55416] = 32'b11111111111111011100110111101100;
assign LUT_2[55417] = 32'b11111111111111011001110000000101;
assign LUT_2[55418] = 32'b11111111111111100011110000101000;
assign LUT_2[55419] = 32'b11111111111111100000101001000001;
assign LUT_2[55420] = 32'b11111111111111011001010101010100;
assign LUT_2[55421] = 32'b11111111111111010110001101101101;
assign LUT_2[55422] = 32'b11111111111111100000001110010000;
assign LUT_2[55423] = 32'b11111111111111011101000110101001;
assign LUT_2[55424] = 32'b11111111111111110011010010001000;
assign LUT_2[55425] = 32'b11111111111111110000001010100001;
assign LUT_2[55426] = 32'b11111111111111111010001011000100;
assign LUT_2[55427] = 32'b11111111111111110111000011011101;
assign LUT_2[55428] = 32'b11111111111111101111101111110000;
assign LUT_2[55429] = 32'b11111111111111101100101000001001;
assign LUT_2[55430] = 32'b11111111111111110110101000101100;
assign LUT_2[55431] = 32'b11111111111111110011100001000101;
assign LUT_2[55432] = 32'b11111111111111101110000011100101;
assign LUT_2[55433] = 32'b11111111111111101010111011111110;
assign LUT_2[55434] = 32'b11111111111111110100111100100001;
assign LUT_2[55435] = 32'b11111111111111110001110100111010;
assign LUT_2[55436] = 32'b11111111111111101010100001001101;
assign LUT_2[55437] = 32'b11111111111111100111011001100110;
assign LUT_2[55438] = 32'b11111111111111110001011010001001;
assign LUT_2[55439] = 32'b11111111111111101110010010100010;
assign LUT_2[55440] = 32'b11111111111111101101110110010010;
assign LUT_2[55441] = 32'b11111111111111101010101110101011;
assign LUT_2[55442] = 32'b11111111111111110100101111001110;
assign LUT_2[55443] = 32'b11111111111111110001100111100111;
assign LUT_2[55444] = 32'b11111111111111101010010011111010;
assign LUT_2[55445] = 32'b11111111111111100111001100010011;
assign LUT_2[55446] = 32'b11111111111111110001001100110110;
assign LUT_2[55447] = 32'b11111111111111101110000101001111;
assign LUT_2[55448] = 32'b11111111111111101000100111101111;
assign LUT_2[55449] = 32'b11111111111111100101100000001000;
assign LUT_2[55450] = 32'b11111111111111101111100000101011;
assign LUT_2[55451] = 32'b11111111111111101100011001000100;
assign LUT_2[55452] = 32'b11111111111111100101000101010111;
assign LUT_2[55453] = 32'b11111111111111100001111101110000;
assign LUT_2[55454] = 32'b11111111111111101011111110010011;
assign LUT_2[55455] = 32'b11111111111111101000110110101100;
assign LUT_2[55456] = 32'b11111111111111110011101101110001;
assign LUT_2[55457] = 32'b11111111111111110000100110001010;
assign LUT_2[55458] = 32'b11111111111111111010100110101101;
assign LUT_2[55459] = 32'b11111111111111110111011111000110;
assign LUT_2[55460] = 32'b11111111111111110000001011011001;
assign LUT_2[55461] = 32'b11111111111111101101000011110010;
assign LUT_2[55462] = 32'b11111111111111110111000100010101;
assign LUT_2[55463] = 32'b11111111111111110011111100101110;
assign LUT_2[55464] = 32'b11111111111111101110011111001110;
assign LUT_2[55465] = 32'b11111111111111101011010111100111;
assign LUT_2[55466] = 32'b11111111111111110101011000001010;
assign LUT_2[55467] = 32'b11111111111111110010010000100011;
assign LUT_2[55468] = 32'b11111111111111101010111100110110;
assign LUT_2[55469] = 32'b11111111111111100111110101001111;
assign LUT_2[55470] = 32'b11111111111111110001110101110010;
assign LUT_2[55471] = 32'b11111111111111101110101110001011;
assign LUT_2[55472] = 32'b11111111111111101110010001111011;
assign LUT_2[55473] = 32'b11111111111111101011001010010100;
assign LUT_2[55474] = 32'b11111111111111110101001010110111;
assign LUT_2[55475] = 32'b11111111111111110010000011010000;
assign LUT_2[55476] = 32'b11111111111111101010101111100011;
assign LUT_2[55477] = 32'b11111111111111100111100111111100;
assign LUT_2[55478] = 32'b11111111111111110001101000011111;
assign LUT_2[55479] = 32'b11111111111111101110100000111000;
assign LUT_2[55480] = 32'b11111111111111101001000011011000;
assign LUT_2[55481] = 32'b11111111111111100101111011110001;
assign LUT_2[55482] = 32'b11111111111111101111111100010100;
assign LUT_2[55483] = 32'b11111111111111101100110100101101;
assign LUT_2[55484] = 32'b11111111111111100101100001000000;
assign LUT_2[55485] = 32'b11111111111111100010011001011001;
assign LUT_2[55486] = 32'b11111111111111101100011001111100;
assign LUT_2[55487] = 32'b11111111111111101001010010010101;
assign LUT_2[55488] = 32'b11111111111111101011011010101011;
assign LUT_2[55489] = 32'b11111111111111101000010011000100;
assign LUT_2[55490] = 32'b11111111111111110010010011100111;
assign LUT_2[55491] = 32'b11111111111111101111001100000000;
assign LUT_2[55492] = 32'b11111111111111100111111000010011;
assign LUT_2[55493] = 32'b11111111111111100100110000101100;
assign LUT_2[55494] = 32'b11111111111111101110110001001111;
assign LUT_2[55495] = 32'b11111111111111101011101001101000;
assign LUT_2[55496] = 32'b11111111111111100110001100001000;
assign LUT_2[55497] = 32'b11111111111111100011000100100001;
assign LUT_2[55498] = 32'b11111111111111101101000101000100;
assign LUT_2[55499] = 32'b11111111111111101001111101011101;
assign LUT_2[55500] = 32'b11111111111111100010101001110000;
assign LUT_2[55501] = 32'b11111111111111011111100010001001;
assign LUT_2[55502] = 32'b11111111111111101001100010101100;
assign LUT_2[55503] = 32'b11111111111111100110011011000101;
assign LUT_2[55504] = 32'b11111111111111100101111110110101;
assign LUT_2[55505] = 32'b11111111111111100010110111001110;
assign LUT_2[55506] = 32'b11111111111111101100110111110001;
assign LUT_2[55507] = 32'b11111111111111101001110000001010;
assign LUT_2[55508] = 32'b11111111111111100010011100011101;
assign LUT_2[55509] = 32'b11111111111111011111010100110110;
assign LUT_2[55510] = 32'b11111111111111101001010101011001;
assign LUT_2[55511] = 32'b11111111111111100110001101110010;
assign LUT_2[55512] = 32'b11111111111111100000110000010010;
assign LUT_2[55513] = 32'b11111111111111011101101000101011;
assign LUT_2[55514] = 32'b11111111111111100111101001001110;
assign LUT_2[55515] = 32'b11111111111111100100100001100111;
assign LUT_2[55516] = 32'b11111111111111011101001101111010;
assign LUT_2[55517] = 32'b11111111111111011010000110010011;
assign LUT_2[55518] = 32'b11111111111111100100000110110110;
assign LUT_2[55519] = 32'b11111111111111100000111111001111;
assign LUT_2[55520] = 32'b11111111111111101011110110010100;
assign LUT_2[55521] = 32'b11111111111111101000101110101101;
assign LUT_2[55522] = 32'b11111111111111110010101111010000;
assign LUT_2[55523] = 32'b11111111111111101111100111101001;
assign LUT_2[55524] = 32'b11111111111111101000010011111100;
assign LUT_2[55525] = 32'b11111111111111100101001100010101;
assign LUT_2[55526] = 32'b11111111111111101111001100111000;
assign LUT_2[55527] = 32'b11111111111111101100000101010001;
assign LUT_2[55528] = 32'b11111111111111100110100111110001;
assign LUT_2[55529] = 32'b11111111111111100011100000001010;
assign LUT_2[55530] = 32'b11111111111111101101100000101101;
assign LUT_2[55531] = 32'b11111111111111101010011001000110;
assign LUT_2[55532] = 32'b11111111111111100011000101011001;
assign LUT_2[55533] = 32'b11111111111111011111111101110010;
assign LUT_2[55534] = 32'b11111111111111101001111110010101;
assign LUT_2[55535] = 32'b11111111111111100110110110101110;
assign LUT_2[55536] = 32'b11111111111111100110011010011110;
assign LUT_2[55537] = 32'b11111111111111100011010010110111;
assign LUT_2[55538] = 32'b11111111111111101101010011011010;
assign LUT_2[55539] = 32'b11111111111111101010001011110011;
assign LUT_2[55540] = 32'b11111111111111100010111000000110;
assign LUT_2[55541] = 32'b11111111111111011111110000011111;
assign LUT_2[55542] = 32'b11111111111111101001110001000010;
assign LUT_2[55543] = 32'b11111111111111100110101001011011;
assign LUT_2[55544] = 32'b11111111111111100001001011111011;
assign LUT_2[55545] = 32'b11111111111111011110000100010100;
assign LUT_2[55546] = 32'b11111111111111101000000100110111;
assign LUT_2[55547] = 32'b11111111111111100100111101010000;
assign LUT_2[55548] = 32'b11111111111111011101101001100011;
assign LUT_2[55549] = 32'b11111111111111011010100001111100;
assign LUT_2[55550] = 32'b11111111111111100100100010011111;
assign LUT_2[55551] = 32'b11111111111111100001011010111000;
assign LUT_2[55552] = 32'b11111111111111110010111100011111;
assign LUT_2[55553] = 32'b11111111111111101111110100111000;
assign LUT_2[55554] = 32'b11111111111111111001110101011011;
assign LUT_2[55555] = 32'b11111111111111110110101101110100;
assign LUT_2[55556] = 32'b11111111111111101111011010000111;
assign LUT_2[55557] = 32'b11111111111111101100010010100000;
assign LUT_2[55558] = 32'b11111111111111110110010011000011;
assign LUT_2[55559] = 32'b11111111111111110011001011011100;
assign LUT_2[55560] = 32'b11111111111111101101101101111100;
assign LUT_2[55561] = 32'b11111111111111101010100110010101;
assign LUT_2[55562] = 32'b11111111111111110100100110111000;
assign LUT_2[55563] = 32'b11111111111111110001011111010001;
assign LUT_2[55564] = 32'b11111111111111101010001011100100;
assign LUT_2[55565] = 32'b11111111111111100111000011111101;
assign LUT_2[55566] = 32'b11111111111111110001000100100000;
assign LUT_2[55567] = 32'b11111111111111101101111100111001;
assign LUT_2[55568] = 32'b11111111111111101101100000101001;
assign LUT_2[55569] = 32'b11111111111111101010011001000010;
assign LUT_2[55570] = 32'b11111111111111110100011001100101;
assign LUT_2[55571] = 32'b11111111111111110001010001111110;
assign LUT_2[55572] = 32'b11111111111111101001111110010001;
assign LUT_2[55573] = 32'b11111111111111100110110110101010;
assign LUT_2[55574] = 32'b11111111111111110000110111001101;
assign LUT_2[55575] = 32'b11111111111111101101101111100110;
assign LUT_2[55576] = 32'b11111111111111101000010010000110;
assign LUT_2[55577] = 32'b11111111111111100101001010011111;
assign LUT_2[55578] = 32'b11111111111111101111001011000010;
assign LUT_2[55579] = 32'b11111111111111101100000011011011;
assign LUT_2[55580] = 32'b11111111111111100100101111101110;
assign LUT_2[55581] = 32'b11111111111111100001101000000111;
assign LUT_2[55582] = 32'b11111111111111101011101000101010;
assign LUT_2[55583] = 32'b11111111111111101000100001000011;
assign LUT_2[55584] = 32'b11111111111111110011011000001000;
assign LUT_2[55585] = 32'b11111111111111110000010000100001;
assign LUT_2[55586] = 32'b11111111111111111010010001000100;
assign LUT_2[55587] = 32'b11111111111111110111001001011101;
assign LUT_2[55588] = 32'b11111111111111101111110101110000;
assign LUT_2[55589] = 32'b11111111111111101100101110001001;
assign LUT_2[55590] = 32'b11111111111111110110101110101100;
assign LUT_2[55591] = 32'b11111111111111110011100111000101;
assign LUT_2[55592] = 32'b11111111111111101110001001100101;
assign LUT_2[55593] = 32'b11111111111111101011000001111110;
assign LUT_2[55594] = 32'b11111111111111110101000010100001;
assign LUT_2[55595] = 32'b11111111111111110001111010111010;
assign LUT_2[55596] = 32'b11111111111111101010100111001101;
assign LUT_2[55597] = 32'b11111111111111100111011111100110;
assign LUT_2[55598] = 32'b11111111111111110001100000001001;
assign LUT_2[55599] = 32'b11111111111111101110011000100010;
assign LUT_2[55600] = 32'b11111111111111101101111100010010;
assign LUT_2[55601] = 32'b11111111111111101010110100101011;
assign LUT_2[55602] = 32'b11111111111111110100110101001110;
assign LUT_2[55603] = 32'b11111111111111110001101101100111;
assign LUT_2[55604] = 32'b11111111111111101010011001111010;
assign LUT_2[55605] = 32'b11111111111111100111010010010011;
assign LUT_2[55606] = 32'b11111111111111110001010010110110;
assign LUT_2[55607] = 32'b11111111111111101110001011001111;
assign LUT_2[55608] = 32'b11111111111111101000101101101111;
assign LUT_2[55609] = 32'b11111111111111100101100110001000;
assign LUT_2[55610] = 32'b11111111111111101111100110101011;
assign LUT_2[55611] = 32'b11111111111111101100011111000100;
assign LUT_2[55612] = 32'b11111111111111100101001011010111;
assign LUT_2[55613] = 32'b11111111111111100010000011110000;
assign LUT_2[55614] = 32'b11111111111111101100000100010011;
assign LUT_2[55615] = 32'b11111111111111101000111100101100;
assign LUT_2[55616] = 32'b11111111111111101011000101000010;
assign LUT_2[55617] = 32'b11111111111111100111111101011011;
assign LUT_2[55618] = 32'b11111111111111110001111101111110;
assign LUT_2[55619] = 32'b11111111111111101110110110010111;
assign LUT_2[55620] = 32'b11111111111111100111100010101010;
assign LUT_2[55621] = 32'b11111111111111100100011011000011;
assign LUT_2[55622] = 32'b11111111111111101110011011100110;
assign LUT_2[55623] = 32'b11111111111111101011010011111111;
assign LUT_2[55624] = 32'b11111111111111100101110110011111;
assign LUT_2[55625] = 32'b11111111111111100010101110111000;
assign LUT_2[55626] = 32'b11111111111111101100101111011011;
assign LUT_2[55627] = 32'b11111111111111101001100111110100;
assign LUT_2[55628] = 32'b11111111111111100010010100000111;
assign LUT_2[55629] = 32'b11111111111111011111001100100000;
assign LUT_2[55630] = 32'b11111111111111101001001101000011;
assign LUT_2[55631] = 32'b11111111111111100110000101011100;
assign LUT_2[55632] = 32'b11111111111111100101101001001100;
assign LUT_2[55633] = 32'b11111111111111100010100001100101;
assign LUT_2[55634] = 32'b11111111111111101100100010001000;
assign LUT_2[55635] = 32'b11111111111111101001011010100001;
assign LUT_2[55636] = 32'b11111111111111100010000110110100;
assign LUT_2[55637] = 32'b11111111111111011110111111001101;
assign LUT_2[55638] = 32'b11111111111111101000111111110000;
assign LUT_2[55639] = 32'b11111111111111100101111000001001;
assign LUT_2[55640] = 32'b11111111111111100000011010101001;
assign LUT_2[55641] = 32'b11111111111111011101010011000010;
assign LUT_2[55642] = 32'b11111111111111100111010011100101;
assign LUT_2[55643] = 32'b11111111111111100100001011111110;
assign LUT_2[55644] = 32'b11111111111111011100111000010001;
assign LUT_2[55645] = 32'b11111111111111011001110000101010;
assign LUT_2[55646] = 32'b11111111111111100011110001001101;
assign LUT_2[55647] = 32'b11111111111111100000101001100110;
assign LUT_2[55648] = 32'b11111111111111101011100000101011;
assign LUT_2[55649] = 32'b11111111111111101000011001000100;
assign LUT_2[55650] = 32'b11111111111111110010011001100111;
assign LUT_2[55651] = 32'b11111111111111101111010010000000;
assign LUT_2[55652] = 32'b11111111111111100111111110010011;
assign LUT_2[55653] = 32'b11111111111111100100110110101100;
assign LUT_2[55654] = 32'b11111111111111101110110111001111;
assign LUT_2[55655] = 32'b11111111111111101011101111101000;
assign LUT_2[55656] = 32'b11111111111111100110010010001000;
assign LUT_2[55657] = 32'b11111111111111100011001010100001;
assign LUT_2[55658] = 32'b11111111111111101101001011000100;
assign LUT_2[55659] = 32'b11111111111111101010000011011101;
assign LUT_2[55660] = 32'b11111111111111100010101111110000;
assign LUT_2[55661] = 32'b11111111111111011111101000001001;
assign LUT_2[55662] = 32'b11111111111111101001101000101100;
assign LUT_2[55663] = 32'b11111111111111100110100001000101;
assign LUT_2[55664] = 32'b11111111111111100110000100110101;
assign LUT_2[55665] = 32'b11111111111111100010111101001110;
assign LUT_2[55666] = 32'b11111111111111101100111101110001;
assign LUT_2[55667] = 32'b11111111111111101001110110001010;
assign LUT_2[55668] = 32'b11111111111111100010100010011101;
assign LUT_2[55669] = 32'b11111111111111011111011010110110;
assign LUT_2[55670] = 32'b11111111111111101001011011011001;
assign LUT_2[55671] = 32'b11111111111111100110010011110010;
assign LUT_2[55672] = 32'b11111111111111100000110110010010;
assign LUT_2[55673] = 32'b11111111111111011101101110101011;
assign LUT_2[55674] = 32'b11111111111111100111101111001110;
assign LUT_2[55675] = 32'b11111111111111100100100111100111;
assign LUT_2[55676] = 32'b11111111111111011101010011111010;
assign LUT_2[55677] = 32'b11111111111111011010001100010011;
assign LUT_2[55678] = 32'b11111111111111100100001100110110;
assign LUT_2[55679] = 32'b11111111111111100001000101001111;
assign LUT_2[55680] = 32'b11111111111111110111010000101110;
assign LUT_2[55681] = 32'b11111111111111110100001001000111;
assign LUT_2[55682] = 32'b11111111111111111110001001101010;
assign LUT_2[55683] = 32'b11111111111111111011000010000011;
assign LUT_2[55684] = 32'b11111111111111110011101110010110;
assign LUT_2[55685] = 32'b11111111111111110000100110101111;
assign LUT_2[55686] = 32'b11111111111111111010100111010010;
assign LUT_2[55687] = 32'b11111111111111110111011111101011;
assign LUT_2[55688] = 32'b11111111111111110010000010001011;
assign LUT_2[55689] = 32'b11111111111111101110111010100100;
assign LUT_2[55690] = 32'b11111111111111111000111011000111;
assign LUT_2[55691] = 32'b11111111111111110101110011100000;
assign LUT_2[55692] = 32'b11111111111111101110011111110011;
assign LUT_2[55693] = 32'b11111111111111101011011000001100;
assign LUT_2[55694] = 32'b11111111111111110101011000101111;
assign LUT_2[55695] = 32'b11111111111111110010010001001000;
assign LUT_2[55696] = 32'b11111111111111110001110100111000;
assign LUT_2[55697] = 32'b11111111111111101110101101010001;
assign LUT_2[55698] = 32'b11111111111111111000101101110100;
assign LUT_2[55699] = 32'b11111111111111110101100110001101;
assign LUT_2[55700] = 32'b11111111111111101110010010100000;
assign LUT_2[55701] = 32'b11111111111111101011001010111001;
assign LUT_2[55702] = 32'b11111111111111110101001011011100;
assign LUT_2[55703] = 32'b11111111111111110010000011110101;
assign LUT_2[55704] = 32'b11111111111111101100100110010101;
assign LUT_2[55705] = 32'b11111111111111101001011110101110;
assign LUT_2[55706] = 32'b11111111111111110011011111010001;
assign LUT_2[55707] = 32'b11111111111111110000010111101010;
assign LUT_2[55708] = 32'b11111111111111101001000011111101;
assign LUT_2[55709] = 32'b11111111111111100101111100010110;
assign LUT_2[55710] = 32'b11111111111111101111111100111001;
assign LUT_2[55711] = 32'b11111111111111101100110101010010;
assign LUT_2[55712] = 32'b11111111111111110111101100010111;
assign LUT_2[55713] = 32'b11111111111111110100100100110000;
assign LUT_2[55714] = 32'b11111111111111111110100101010011;
assign LUT_2[55715] = 32'b11111111111111111011011101101100;
assign LUT_2[55716] = 32'b11111111111111110100001001111111;
assign LUT_2[55717] = 32'b11111111111111110001000010011000;
assign LUT_2[55718] = 32'b11111111111111111011000010111011;
assign LUT_2[55719] = 32'b11111111111111110111111011010100;
assign LUT_2[55720] = 32'b11111111111111110010011101110100;
assign LUT_2[55721] = 32'b11111111111111101111010110001101;
assign LUT_2[55722] = 32'b11111111111111111001010110110000;
assign LUT_2[55723] = 32'b11111111111111110110001111001001;
assign LUT_2[55724] = 32'b11111111111111101110111011011100;
assign LUT_2[55725] = 32'b11111111111111101011110011110101;
assign LUT_2[55726] = 32'b11111111111111110101110100011000;
assign LUT_2[55727] = 32'b11111111111111110010101100110001;
assign LUT_2[55728] = 32'b11111111111111110010010000100001;
assign LUT_2[55729] = 32'b11111111111111101111001000111010;
assign LUT_2[55730] = 32'b11111111111111111001001001011101;
assign LUT_2[55731] = 32'b11111111111111110110000001110110;
assign LUT_2[55732] = 32'b11111111111111101110101110001001;
assign LUT_2[55733] = 32'b11111111111111101011100110100010;
assign LUT_2[55734] = 32'b11111111111111110101100111000101;
assign LUT_2[55735] = 32'b11111111111111110010011111011110;
assign LUT_2[55736] = 32'b11111111111111101101000001111110;
assign LUT_2[55737] = 32'b11111111111111101001111010010111;
assign LUT_2[55738] = 32'b11111111111111110011111010111010;
assign LUT_2[55739] = 32'b11111111111111110000110011010011;
assign LUT_2[55740] = 32'b11111111111111101001011111100110;
assign LUT_2[55741] = 32'b11111111111111100110010111111111;
assign LUT_2[55742] = 32'b11111111111111110000011000100010;
assign LUT_2[55743] = 32'b11111111111111101101010000111011;
assign LUT_2[55744] = 32'b11111111111111101111011001010001;
assign LUT_2[55745] = 32'b11111111111111101100010001101010;
assign LUT_2[55746] = 32'b11111111111111110110010010001101;
assign LUT_2[55747] = 32'b11111111111111110011001010100110;
assign LUT_2[55748] = 32'b11111111111111101011110110111001;
assign LUT_2[55749] = 32'b11111111111111101000101111010010;
assign LUT_2[55750] = 32'b11111111111111110010101111110101;
assign LUT_2[55751] = 32'b11111111111111101111101000001110;
assign LUT_2[55752] = 32'b11111111111111101010001010101110;
assign LUT_2[55753] = 32'b11111111111111100111000011000111;
assign LUT_2[55754] = 32'b11111111111111110001000011101010;
assign LUT_2[55755] = 32'b11111111111111101101111100000011;
assign LUT_2[55756] = 32'b11111111111111100110101000010110;
assign LUT_2[55757] = 32'b11111111111111100011100000101111;
assign LUT_2[55758] = 32'b11111111111111101101100001010010;
assign LUT_2[55759] = 32'b11111111111111101010011001101011;
assign LUT_2[55760] = 32'b11111111111111101001111101011011;
assign LUT_2[55761] = 32'b11111111111111100110110101110100;
assign LUT_2[55762] = 32'b11111111111111110000110110010111;
assign LUT_2[55763] = 32'b11111111111111101101101110110000;
assign LUT_2[55764] = 32'b11111111111111100110011011000011;
assign LUT_2[55765] = 32'b11111111111111100011010011011100;
assign LUT_2[55766] = 32'b11111111111111101101010011111111;
assign LUT_2[55767] = 32'b11111111111111101010001100011000;
assign LUT_2[55768] = 32'b11111111111111100100101110111000;
assign LUT_2[55769] = 32'b11111111111111100001100111010001;
assign LUT_2[55770] = 32'b11111111111111101011100111110100;
assign LUT_2[55771] = 32'b11111111111111101000100000001101;
assign LUT_2[55772] = 32'b11111111111111100001001100100000;
assign LUT_2[55773] = 32'b11111111111111011110000100111001;
assign LUT_2[55774] = 32'b11111111111111101000000101011100;
assign LUT_2[55775] = 32'b11111111111111100100111101110101;
assign LUT_2[55776] = 32'b11111111111111101111110100111010;
assign LUT_2[55777] = 32'b11111111111111101100101101010011;
assign LUT_2[55778] = 32'b11111111111111110110101101110110;
assign LUT_2[55779] = 32'b11111111111111110011100110001111;
assign LUT_2[55780] = 32'b11111111111111101100010010100010;
assign LUT_2[55781] = 32'b11111111111111101001001010111011;
assign LUT_2[55782] = 32'b11111111111111110011001011011110;
assign LUT_2[55783] = 32'b11111111111111110000000011110111;
assign LUT_2[55784] = 32'b11111111111111101010100110010111;
assign LUT_2[55785] = 32'b11111111111111100111011110110000;
assign LUT_2[55786] = 32'b11111111111111110001011111010011;
assign LUT_2[55787] = 32'b11111111111111101110010111101100;
assign LUT_2[55788] = 32'b11111111111111100111000011111111;
assign LUT_2[55789] = 32'b11111111111111100011111100011000;
assign LUT_2[55790] = 32'b11111111111111101101111100111011;
assign LUT_2[55791] = 32'b11111111111111101010110101010100;
assign LUT_2[55792] = 32'b11111111111111101010011001000100;
assign LUT_2[55793] = 32'b11111111111111100111010001011101;
assign LUT_2[55794] = 32'b11111111111111110001010010000000;
assign LUT_2[55795] = 32'b11111111111111101110001010011001;
assign LUT_2[55796] = 32'b11111111111111100110110110101100;
assign LUT_2[55797] = 32'b11111111111111100011101111000101;
assign LUT_2[55798] = 32'b11111111111111101101101111101000;
assign LUT_2[55799] = 32'b11111111111111101010101000000001;
assign LUT_2[55800] = 32'b11111111111111100101001010100001;
assign LUT_2[55801] = 32'b11111111111111100010000010111010;
assign LUT_2[55802] = 32'b11111111111111101100000011011101;
assign LUT_2[55803] = 32'b11111111111111101000111011110110;
assign LUT_2[55804] = 32'b11111111111111100001101000001001;
assign LUT_2[55805] = 32'b11111111111111011110100000100010;
assign LUT_2[55806] = 32'b11111111111111101000100001000101;
assign LUT_2[55807] = 32'b11111111111111100101011001011110;
assign LUT_2[55808] = 32'b11111111111111110011101111101011;
assign LUT_2[55809] = 32'b11111111111111110000101000000100;
assign LUT_2[55810] = 32'b11111111111111111010101000100111;
assign LUT_2[55811] = 32'b11111111111111110111100001000000;
assign LUT_2[55812] = 32'b11111111111111110000001101010011;
assign LUT_2[55813] = 32'b11111111111111101101000101101100;
assign LUT_2[55814] = 32'b11111111111111110111000110001111;
assign LUT_2[55815] = 32'b11111111111111110011111110101000;
assign LUT_2[55816] = 32'b11111111111111101110100001001000;
assign LUT_2[55817] = 32'b11111111111111101011011001100001;
assign LUT_2[55818] = 32'b11111111111111110101011010000100;
assign LUT_2[55819] = 32'b11111111111111110010010010011101;
assign LUT_2[55820] = 32'b11111111111111101010111110110000;
assign LUT_2[55821] = 32'b11111111111111100111110111001001;
assign LUT_2[55822] = 32'b11111111111111110001110111101100;
assign LUT_2[55823] = 32'b11111111111111101110110000000101;
assign LUT_2[55824] = 32'b11111111111111101110010011110101;
assign LUT_2[55825] = 32'b11111111111111101011001100001110;
assign LUT_2[55826] = 32'b11111111111111110101001100110001;
assign LUT_2[55827] = 32'b11111111111111110010000101001010;
assign LUT_2[55828] = 32'b11111111111111101010110001011101;
assign LUT_2[55829] = 32'b11111111111111100111101001110110;
assign LUT_2[55830] = 32'b11111111111111110001101010011001;
assign LUT_2[55831] = 32'b11111111111111101110100010110010;
assign LUT_2[55832] = 32'b11111111111111101001000101010010;
assign LUT_2[55833] = 32'b11111111111111100101111101101011;
assign LUT_2[55834] = 32'b11111111111111101111111110001110;
assign LUT_2[55835] = 32'b11111111111111101100110110100111;
assign LUT_2[55836] = 32'b11111111111111100101100010111010;
assign LUT_2[55837] = 32'b11111111111111100010011011010011;
assign LUT_2[55838] = 32'b11111111111111101100011011110110;
assign LUT_2[55839] = 32'b11111111111111101001010100001111;
assign LUT_2[55840] = 32'b11111111111111110100001011010100;
assign LUT_2[55841] = 32'b11111111111111110001000011101101;
assign LUT_2[55842] = 32'b11111111111111111011000100010000;
assign LUT_2[55843] = 32'b11111111111111110111111100101001;
assign LUT_2[55844] = 32'b11111111111111110000101000111100;
assign LUT_2[55845] = 32'b11111111111111101101100001010101;
assign LUT_2[55846] = 32'b11111111111111110111100001111000;
assign LUT_2[55847] = 32'b11111111111111110100011010010001;
assign LUT_2[55848] = 32'b11111111111111101110111100110001;
assign LUT_2[55849] = 32'b11111111111111101011110101001010;
assign LUT_2[55850] = 32'b11111111111111110101110101101101;
assign LUT_2[55851] = 32'b11111111111111110010101110000110;
assign LUT_2[55852] = 32'b11111111111111101011011010011001;
assign LUT_2[55853] = 32'b11111111111111101000010010110010;
assign LUT_2[55854] = 32'b11111111111111110010010011010101;
assign LUT_2[55855] = 32'b11111111111111101111001011101110;
assign LUT_2[55856] = 32'b11111111111111101110101111011110;
assign LUT_2[55857] = 32'b11111111111111101011100111110111;
assign LUT_2[55858] = 32'b11111111111111110101101000011010;
assign LUT_2[55859] = 32'b11111111111111110010100000110011;
assign LUT_2[55860] = 32'b11111111111111101011001101000110;
assign LUT_2[55861] = 32'b11111111111111101000000101011111;
assign LUT_2[55862] = 32'b11111111111111110010000110000010;
assign LUT_2[55863] = 32'b11111111111111101110111110011011;
assign LUT_2[55864] = 32'b11111111111111101001100000111011;
assign LUT_2[55865] = 32'b11111111111111100110011001010100;
assign LUT_2[55866] = 32'b11111111111111110000011001110111;
assign LUT_2[55867] = 32'b11111111111111101101010010010000;
assign LUT_2[55868] = 32'b11111111111111100101111110100011;
assign LUT_2[55869] = 32'b11111111111111100010110110111100;
assign LUT_2[55870] = 32'b11111111111111101100110111011111;
assign LUT_2[55871] = 32'b11111111111111101001101111111000;
assign LUT_2[55872] = 32'b11111111111111101011111000001110;
assign LUT_2[55873] = 32'b11111111111111101000110000100111;
assign LUT_2[55874] = 32'b11111111111111110010110001001010;
assign LUT_2[55875] = 32'b11111111111111101111101001100011;
assign LUT_2[55876] = 32'b11111111111111101000010101110110;
assign LUT_2[55877] = 32'b11111111111111100101001110001111;
assign LUT_2[55878] = 32'b11111111111111101111001110110010;
assign LUT_2[55879] = 32'b11111111111111101100000111001011;
assign LUT_2[55880] = 32'b11111111111111100110101001101011;
assign LUT_2[55881] = 32'b11111111111111100011100010000100;
assign LUT_2[55882] = 32'b11111111111111101101100010100111;
assign LUT_2[55883] = 32'b11111111111111101010011011000000;
assign LUT_2[55884] = 32'b11111111111111100011000111010011;
assign LUT_2[55885] = 32'b11111111111111011111111111101100;
assign LUT_2[55886] = 32'b11111111111111101010000000001111;
assign LUT_2[55887] = 32'b11111111111111100110111000101000;
assign LUT_2[55888] = 32'b11111111111111100110011100011000;
assign LUT_2[55889] = 32'b11111111111111100011010100110001;
assign LUT_2[55890] = 32'b11111111111111101101010101010100;
assign LUT_2[55891] = 32'b11111111111111101010001101101101;
assign LUT_2[55892] = 32'b11111111111111100010111010000000;
assign LUT_2[55893] = 32'b11111111111111011111110010011001;
assign LUT_2[55894] = 32'b11111111111111101001110010111100;
assign LUT_2[55895] = 32'b11111111111111100110101011010101;
assign LUT_2[55896] = 32'b11111111111111100001001101110101;
assign LUT_2[55897] = 32'b11111111111111011110000110001110;
assign LUT_2[55898] = 32'b11111111111111101000000110110001;
assign LUT_2[55899] = 32'b11111111111111100100111111001010;
assign LUT_2[55900] = 32'b11111111111111011101101011011101;
assign LUT_2[55901] = 32'b11111111111111011010100011110110;
assign LUT_2[55902] = 32'b11111111111111100100100100011001;
assign LUT_2[55903] = 32'b11111111111111100001011100110010;
assign LUT_2[55904] = 32'b11111111111111101100010011110111;
assign LUT_2[55905] = 32'b11111111111111101001001100010000;
assign LUT_2[55906] = 32'b11111111111111110011001100110011;
assign LUT_2[55907] = 32'b11111111111111110000000101001100;
assign LUT_2[55908] = 32'b11111111111111101000110001011111;
assign LUT_2[55909] = 32'b11111111111111100101101001111000;
assign LUT_2[55910] = 32'b11111111111111101111101010011011;
assign LUT_2[55911] = 32'b11111111111111101100100010110100;
assign LUT_2[55912] = 32'b11111111111111100111000101010100;
assign LUT_2[55913] = 32'b11111111111111100011111101101101;
assign LUT_2[55914] = 32'b11111111111111101101111110010000;
assign LUT_2[55915] = 32'b11111111111111101010110110101001;
assign LUT_2[55916] = 32'b11111111111111100011100010111100;
assign LUT_2[55917] = 32'b11111111111111100000011011010101;
assign LUT_2[55918] = 32'b11111111111111101010011011111000;
assign LUT_2[55919] = 32'b11111111111111100111010100010001;
assign LUT_2[55920] = 32'b11111111111111100110111000000001;
assign LUT_2[55921] = 32'b11111111111111100011110000011010;
assign LUT_2[55922] = 32'b11111111111111101101110000111101;
assign LUT_2[55923] = 32'b11111111111111101010101001010110;
assign LUT_2[55924] = 32'b11111111111111100011010101101001;
assign LUT_2[55925] = 32'b11111111111111100000001110000010;
assign LUT_2[55926] = 32'b11111111111111101010001110100101;
assign LUT_2[55927] = 32'b11111111111111100111000110111110;
assign LUT_2[55928] = 32'b11111111111111100001101001011110;
assign LUT_2[55929] = 32'b11111111111111011110100001110111;
assign LUT_2[55930] = 32'b11111111111111101000100010011010;
assign LUT_2[55931] = 32'b11111111111111100101011010110011;
assign LUT_2[55932] = 32'b11111111111111011110000111000110;
assign LUT_2[55933] = 32'b11111111111111011010111111011111;
assign LUT_2[55934] = 32'b11111111111111100101000000000010;
assign LUT_2[55935] = 32'b11111111111111100001111000011011;
assign LUT_2[55936] = 32'b11111111111111111000000011111010;
assign LUT_2[55937] = 32'b11111111111111110100111100010011;
assign LUT_2[55938] = 32'b11111111111111111110111100110110;
assign LUT_2[55939] = 32'b11111111111111111011110101001111;
assign LUT_2[55940] = 32'b11111111111111110100100001100010;
assign LUT_2[55941] = 32'b11111111111111110001011001111011;
assign LUT_2[55942] = 32'b11111111111111111011011010011110;
assign LUT_2[55943] = 32'b11111111111111111000010010110111;
assign LUT_2[55944] = 32'b11111111111111110010110101010111;
assign LUT_2[55945] = 32'b11111111111111101111101101110000;
assign LUT_2[55946] = 32'b11111111111111111001101110010011;
assign LUT_2[55947] = 32'b11111111111111110110100110101100;
assign LUT_2[55948] = 32'b11111111111111101111010010111111;
assign LUT_2[55949] = 32'b11111111111111101100001011011000;
assign LUT_2[55950] = 32'b11111111111111110110001011111011;
assign LUT_2[55951] = 32'b11111111111111110011000100010100;
assign LUT_2[55952] = 32'b11111111111111110010101000000100;
assign LUT_2[55953] = 32'b11111111111111101111100000011101;
assign LUT_2[55954] = 32'b11111111111111111001100001000000;
assign LUT_2[55955] = 32'b11111111111111110110011001011001;
assign LUT_2[55956] = 32'b11111111111111101111000101101100;
assign LUT_2[55957] = 32'b11111111111111101011111110000101;
assign LUT_2[55958] = 32'b11111111111111110101111110101000;
assign LUT_2[55959] = 32'b11111111111111110010110111000001;
assign LUT_2[55960] = 32'b11111111111111101101011001100001;
assign LUT_2[55961] = 32'b11111111111111101010010001111010;
assign LUT_2[55962] = 32'b11111111111111110100010010011101;
assign LUT_2[55963] = 32'b11111111111111110001001010110110;
assign LUT_2[55964] = 32'b11111111111111101001110111001001;
assign LUT_2[55965] = 32'b11111111111111100110101111100010;
assign LUT_2[55966] = 32'b11111111111111110000110000000101;
assign LUT_2[55967] = 32'b11111111111111101101101000011110;
assign LUT_2[55968] = 32'b11111111111111111000011111100011;
assign LUT_2[55969] = 32'b11111111111111110101010111111100;
assign LUT_2[55970] = 32'b11111111111111111111011000011111;
assign LUT_2[55971] = 32'b11111111111111111100010000111000;
assign LUT_2[55972] = 32'b11111111111111110100111101001011;
assign LUT_2[55973] = 32'b11111111111111110001110101100100;
assign LUT_2[55974] = 32'b11111111111111111011110110000111;
assign LUT_2[55975] = 32'b11111111111111111000101110100000;
assign LUT_2[55976] = 32'b11111111111111110011010001000000;
assign LUT_2[55977] = 32'b11111111111111110000001001011001;
assign LUT_2[55978] = 32'b11111111111111111010001001111100;
assign LUT_2[55979] = 32'b11111111111111110111000010010101;
assign LUT_2[55980] = 32'b11111111111111101111101110101000;
assign LUT_2[55981] = 32'b11111111111111101100100111000001;
assign LUT_2[55982] = 32'b11111111111111110110100111100100;
assign LUT_2[55983] = 32'b11111111111111110011011111111101;
assign LUT_2[55984] = 32'b11111111111111110011000011101101;
assign LUT_2[55985] = 32'b11111111111111101111111100000110;
assign LUT_2[55986] = 32'b11111111111111111001111100101001;
assign LUT_2[55987] = 32'b11111111111111110110110101000010;
assign LUT_2[55988] = 32'b11111111111111101111100001010101;
assign LUT_2[55989] = 32'b11111111111111101100011001101110;
assign LUT_2[55990] = 32'b11111111111111110110011010010001;
assign LUT_2[55991] = 32'b11111111111111110011010010101010;
assign LUT_2[55992] = 32'b11111111111111101101110101001010;
assign LUT_2[55993] = 32'b11111111111111101010101101100011;
assign LUT_2[55994] = 32'b11111111111111110100101110000110;
assign LUT_2[55995] = 32'b11111111111111110001100110011111;
assign LUT_2[55996] = 32'b11111111111111101010010010110010;
assign LUT_2[55997] = 32'b11111111111111100111001011001011;
assign LUT_2[55998] = 32'b11111111111111110001001011101110;
assign LUT_2[55999] = 32'b11111111111111101110000100000111;
assign LUT_2[56000] = 32'b11111111111111110000001100011101;
assign LUT_2[56001] = 32'b11111111111111101101000100110110;
assign LUT_2[56002] = 32'b11111111111111110111000101011001;
assign LUT_2[56003] = 32'b11111111111111110011111101110010;
assign LUT_2[56004] = 32'b11111111111111101100101010000101;
assign LUT_2[56005] = 32'b11111111111111101001100010011110;
assign LUT_2[56006] = 32'b11111111111111110011100011000001;
assign LUT_2[56007] = 32'b11111111111111110000011011011010;
assign LUT_2[56008] = 32'b11111111111111101010111101111010;
assign LUT_2[56009] = 32'b11111111111111100111110110010011;
assign LUT_2[56010] = 32'b11111111111111110001110110110110;
assign LUT_2[56011] = 32'b11111111111111101110101111001111;
assign LUT_2[56012] = 32'b11111111111111100111011011100010;
assign LUT_2[56013] = 32'b11111111111111100100010011111011;
assign LUT_2[56014] = 32'b11111111111111101110010100011110;
assign LUT_2[56015] = 32'b11111111111111101011001100110111;
assign LUT_2[56016] = 32'b11111111111111101010110000100111;
assign LUT_2[56017] = 32'b11111111111111100111101001000000;
assign LUT_2[56018] = 32'b11111111111111110001101001100011;
assign LUT_2[56019] = 32'b11111111111111101110100001111100;
assign LUT_2[56020] = 32'b11111111111111100111001110001111;
assign LUT_2[56021] = 32'b11111111111111100100000110101000;
assign LUT_2[56022] = 32'b11111111111111101110000111001011;
assign LUT_2[56023] = 32'b11111111111111101010111111100100;
assign LUT_2[56024] = 32'b11111111111111100101100010000100;
assign LUT_2[56025] = 32'b11111111111111100010011010011101;
assign LUT_2[56026] = 32'b11111111111111101100011011000000;
assign LUT_2[56027] = 32'b11111111111111101001010011011001;
assign LUT_2[56028] = 32'b11111111111111100001111111101100;
assign LUT_2[56029] = 32'b11111111111111011110111000000101;
assign LUT_2[56030] = 32'b11111111111111101000111000101000;
assign LUT_2[56031] = 32'b11111111111111100101110001000001;
assign LUT_2[56032] = 32'b11111111111111110000101000000110;
assign LUT_2[56033] = 32'b11111111111111101101100000011111;
assign LUT_2[56034] = 32'b11111111111111110111100001000010;
assign LUT_2[56035] = 32'b11111111111111110100011001011011;
assign LUT_2[56036] = 32'b11111111111111101101000101101110;
assign LUT_2[56037] = 32'b11111111111111101001111110000111;
assign LUT_2[56038] = 32'b11111111111111110011111110101010;
assign LUT_2[56039] = 32'b11111111111111110000110111000011;
assign LUT_2[56040] = 32'b11111111111111101011011001100011;
assign LUT_2[56041] = 32'b11111111111111101000010001111100;
assign LUT_2[56042] = 32'b11111111111111110010010010011111;
assign LUT_2[56043] = 32'b11111111111111101111001010111000;
assign LUT_2[56044] = 32'b11111111111111100111110111001011;
assign LUT_2[56045] = 32'b11111111111111100100101111100100;
assign LUT_2[56046] = 32'b11111111111111101110110000000111;
assign LUT_2[56047] = 32'b11111111111111101011101000100000;
assign LUT_2[56048] = 32'b11111111111111101011001100010000;
assign LUT_2[56049] = 32'b11111111111111101000000100101001;
assign LUT_2[56050] = 32'b11111111111111110010000101001100;
assign LUT_2[56051] = 32'b11111111111111101110111101100101;
assign LUT_2[56052] = 32'b11111111111111100111101001111000;
assign LUT_2[56053] = 32'b11111111111111100100100010010001;
assign LUT_2[56054] = 32'b11111111111111101110100010110100;
assign LUT_2[56055] = 32'b11111111111111101011011011001101;
assign LUT_2[56056] = 32'b11111111111111100101111101101101;
assign LUT_2[56057] = 32'b11111111111111100010110110000110;
assign LUT_2[56058] = 32'b11111111111111101100110110101001;
assign LUT_2[56059] = 32'b11111111111111101001101111000010;
assign LUT_2[56060] = 32'b11111111111111100010011011010101;
assign LUT_2[56061] = 32'b11111111111111011111010011101110;
assign LUT_2[56062] = 32'b11111111111111101001010100010001;
assign LUT_2[56063] = 32'b11111111111111100110001100101010;
assign LUT_2[56064] = 32'b11111111111111110111101110010001;
assign LUT_2[56065] = 32'b11111111111111110100100110101010;
assign LUT_2[56066] = 32'b11111111111111111110100111001101;
assign LUT_2[56067] = 32'b11111111111111111011011111100110;
assign LUT_2[56068] = 32'b11111111111111110100001011111001;
assign LUT_2[56069] = 32'b11111111111111110001000100010010;
assign LUT_2[56070] = 32'b11111111111111111011000100110101;
assign LUT_2[56071] = 32'b11111111111111110111111101001110;
assign LUT_2[56072] = 32'b11111111111111110010011111101110;
assign LUT_2[56073] = 32'b11111111111111101111011000000111;
assign LUT_2[56074] = 32'b11111111111111111001011000101010;
assign LUT_2[56075] = 32'b11111111111111110110010001000011;
assign LUT_2[56076] = 32'b11111111111111101110111101010110;
assign LUT_2[56077] = 32'b11111111111111101011110101101111;
assign LUT_2[56078] = 32'b11111111111111110101110110010010;
assign LUT_2[56079] = 32'b11111111111111110010101110101011;
assign LUT_2[56080] = 32'b11111111111111110010010010011011;
assign LUT_2[56081] = 32'b11111111111111101111001010110100;
assign LUT_2[56082] = 32'b11111111111111111001001011010111;
assign LUT_2[56083] = 32'b11111111111111110110000011110000;
assign LUT_2[56084] = 32'b11111111111111101110110000000011;
assign LUT_2[56085] = 32'b11111111111111101011101000011100;
assign LUT_2[56086] = 32'b11111111111111110101101000111111;
assign LUT_2[56087] = 32'b11111111111111110010100001011000;
assign LUT_2[56088] = 32'b11111111111111101101000011111000;
assign LUT_2[56089] = 32'b11111111111111101001111100010001;
assign LUT_2[56090] = 32'b11111111111111110011111100110100;
assign LUT_2[56091] = 32'b11111111111111110000110101001101;
assign LUT_2[56092] = 32'b11111111111111101001100001100000;
assign LUT_2[56093] = 32'b11111111111111100110011001111001;
assign LUT_2[56094] = 32'b11111111111111110000011010011100;
assign LUT_2[56095] = 32'b11111111111111101101010010110101;
assign LUT_2[56096] = 32'b11111111111111111000001001111010;
assign LUT_2[56097] = 32'b11111111111111110101000010010011;
assign LUT_2[56098] = 32'b11111111111111111111000010110110;
assign LUT_2[56099] = 32'b11111111111111111011111011001111;
assign LUT_2[56100] = 32'b11111111111111110100100111100010;
assign LUT_2[56101] = 32'b11111111111111110001011111111011;
assign LUT_2[56102] = 32'b11111111111111111011100000011110;
assign LUT_2[56103] = 32'b11111111111111111000011000110111;
assign LUT_2[56104] = 32'b11111111111111110010111011010111;
assign LUT_2[56105] = 32'b11111111111111101111110011110000;
assign LUT_2[56106] = 32'b11111111111111111001110100010011;
assign LUT_2[56107] = 32'b11111111111111110110101100101100;
assign LUT_2[56108] = 32'b11111111111111101111011000111111;
assign LUT_2[56109] = 32'b11111111111111101100010001011000;
assign LUT_2[56110] = 32'b11111111111111110110010001111011;
assign LUT_2[56111] = 32'b11111111111111110011001010010100;
assign LUT_2[56112] = 32'b11111111111111110010101110000100;
assign LUT_2[56113] = 32'b11111111111111101111100110011101;
assign LUT_2[56114] = 32'b11111111111111111001100111000000;
assign LUT_2[56115] = 32'b11111111111111110110011111011001;
assign LUT_2[56116] = 32'b11111111111111101111001011101100;
assign LUT_2[56117] = 32'b11111111111111101100000100000101;
assign LUT_2[56118] = 32'b11111111111111110110000100101000;
assign LUT_2[56119] = 32'b11111111111111110010111101000001;
assign LUT_2[56120] = 32'b11111111111111101101011111100001;
assign LUT_2[56121] = 32'b11111111111111101010010111111010;
assign LUT_2[56122] = 32'b11111111111111110100011000011101;
assign LUT_2[56123] = 32'b11111111111111110001010000110110;
assign LUT_2[56124] = 32'b11111111111111101001111101001001;
assign LUT_2[56125] = 32'b11111111111111100110110101100010;
assign LUT_2[56126] = 32'b11111111111111110000110110000101;
assign LUT_2[56127] = 32'b11111111111111101101101110011110;
assign LUT_2[56128] = 32'b11111111111111101111110110110100;
assign LUT_2[56129] = 32'b11111111111111101100101111001101;
assign LUT_2[56130] = 32'b11111111111111110110101111110000;
assign LUT_2[56131] = 32'b11111111111111110011101000001001;
assign LUT_2[56132] = 32'b11111111111111101100010100011100;
assign LUT_2[56133] = 32'b11111111111111101001001100110101;
assign LUT_2[56134] = 32'b11111111111111110011001101011000;
assign LUT_2[56135] = 32'b11111111111111110000000101110001;
assign LUT_2[56136] = 32'b11111111111111101010101000010001;
assign LUT_2[56137] = 32'b11111111111111100111100000101010;
assign LUT_2[56138] = 32'b11111111111111110001100001001101;
assign LUT_2[56139] = 32'b11111111111111101110011001100110;
assign LUT_2[56140] = 32'b11111111111111100111000101111001;
assign LUT_2[56141] = 32'b11111111111111100011111110010010;
assign LUT_2[56142] = 32'b11111111111111101101111110110101;
assign LUT_2[56143] = 32'b11111111111111101010110111001110;
assign LUT_2[56144] = 32'b11111111111111101010011010111110;
assign LUT_2[56145] = 32'b11111111111111100111010011010111;
assign LUT_2[56146] = 32'b11111111111111110001010011111010;
assign LUT_2[56147] = 32'b11111111111111101110001100010011;
assign LUT_2[56148] = 32'b11111111111111100110111000100110;
assign LUT_2[56149] = 32'b11111111111111100011110000111111;
assign LUT_2[56150] = 32'b11111111111111101101110001100010;
assign LUT_2[56151] = 32'b11111111111111101010101001111011;
assign LUT_2[56152] = 32'b11111111111111100101001100011011;
assign LUT_2[56153] = 32'b11111111111111100010000100110100;
assign LUT_2[56154] = 32'b11111111111111101100000101010111;
assign LUT_2[56155] = 32'b11111111111111101000111101110000;
assign LUT_2[56156] = 32'b11111111111111100001101010000011;
assign LUT_2[56157] = 32'b11111111111111011110100010011100;
assign LUT_2[56158] = 32'b11111111111111101000100010111111;
assign LUT_2[56159] = 32'b11111111111111100101011011011000;
assign LUT_2[56160] = 32'b11111111111111110000010010011101;
assign LUT_2[56161] = 32'b11111111111111101101001010110110;
assign LUT_2[56162] = 32'b11111111111111110111001011011001;
assign LUT_2[56163] = 32'b11111111111111110100000011110010;
assign LUT_2[56164] = 32'b11111111111111101100110000000101;
assign LUT_2[56165] = 32'b11111111111111101001101000011110;
assign LUT_2[56166] = 32'b11111111111111110011101001000001;
assign LUT_2[56167] = 32'b11111111111111110000100001011010;
assign LUT_2[56168] = 32'b11111111111111101011000011111010;
assign LUT_2[56169] = 32'b11111111111111100111111100010011;
assign LUT_2[56170] = 32'b11111111111111110001111100110110;
assign LUT_2[56171] = 32'b11111111111111101110110101001111;
assign LUT_2[56172] = 32'b11111111111111100111100001100010;
assign LUT_2[56173] = 32'b11111111111111100100011001111011;
assign LUT_2[56174] = 32'b11111111111111101110011010011110;
assign LUT_2[56175] = 32'b11111111111111101011010010110111;
assign LUT_2[56176] = 32'b11111111111111101010110110100111;
assign LUT_2[56177] = 32'b11111111111111100111101111000000;
assign LUT_2[56178] = 32'b11111111111111110001101111100011;
assign LUT_2[56179] = 32'b11111111111111101110100111111100;
assign LUT_2[56180] = 32'b11111111111111100111010100001111;
assign LUT_2[56181] = 32'b11111111111111100100001100101000;
assign LUT_2[56182] = 32'b11111111111111101110001101001011;
assign LUT_2[56183] = 32'b11111111111111101011000101100100;
assign LUT_2[56184] = 32'b11111111111111100101101000000100;
assign LUT_2[56185] = 32'b11111111111111100010100000011101;
assign LUT_2[56186] = 32'b11111111111111101100100001000000;
assign LUT_2[56187] = 32'b11111111111111101001011001011001;
assign LUT_2[56188] = 32'b11111111111111100010000101101100;
assign LUT_2[56189] = 32'b11111111111111011110111110000101;
assign LUT_2[56190] = 32'b11111111111111101000111110101000;
assign LUT_2[56191] = 32'b11111111111111100101110111000001;
assign LUT_2[56192] = 32'b11111111111111111100000010100000;
assign LUT_2[56193] = 32'b11111111111111111000111010111001;
assign LUT_2[56194] = 32'b00000000000000000010111011011100;
assign LUT_2[56195] = 32'b11111111111111111111110011110101;
assign LUT_2[56196] = 32'b11111111111111111000100000001000;
assign LUT_2[56197] = 32'b11111111111111110101011000100001;
assign LUT_2[56198] = 32'b11111111111111111111011001000100;
assign LUT_2[56199] = 32'b11111111111111111100010001011101;
assign LUT_2[56200] = 32'b11111111111111110110110011111101;
assign LUT_2[56201] = 32'b11111111111111110011101100010110;
assign LUT_2[56202] = 32'b11111111111111111101101100111001;
assign LUT_2[56203] = 32'b11111111111111111010100101010010;
assign LUT_2[56204] = 32'b11111111111111110011010001100101;
assign LUT_2[56205] = 32'b11111111111111110000001001111110;
assign LUT_2[56206] = 32'b11111111111111111010001010100001;
assign LUT_2[56207] = 32'b11111111111111110111000010111010;
assign LUT_2[56208] = 32'b11111111111111110110100110101010;
assign LUT_2[56209] = 32'b11111111111111110011011111000011;
assign LUT_2[56210] = 32'b11111111111111111101011111100110;
assign LUT_2[56211] = 32'b11111111111111111010010111111111;
assign LUT_2[56212] = 32'b11111111111111110011000100010010;
assign LUT_2[56213] = 32'b11111111111111101111111100101011;
assign LUT_2[56214] = 32'b11111111111111111001111101001110;
assign LUT_2[56215] = 32'b11111111111111110110110101100111;
assign LUT_2[56216] = 32'b11111111111111110001011000000111;
assign LUT_2[56217] = 32'b11111111111111101110010000100000;
assign LUT_2[56218] = 32'b11111111111111111000010001000011;
assign LUT_2[56219] = 32'b11111111111111110101001001011100;
assign LUT_2[56220] = 32'b11111111111111101101110101101111;
assign LUT_2[56221] = 32'b11111111111111101010101110001000;
assign LUT_2[56222] = 32'b11111111111111110100101110101011;
assign LUT_2[56223] = 32'b11111111111111110001100111000100;
assign LUT_2[56224] = 32'b11111111111111111100011110001001;
assign LUT_2[56225] = 32'b11111111111111111001010110100010;
assign LUT_2[56226] = 32'b00000000000000000011010111000101;
assign LUT_2[56227] = 32'b00000000000000000000001111011110;
assign LUT_2[56228] = 32'b11111111111111111000111011110001;
assign LUT_2[56229] = 32'b11111111111111110101110100001010;
assign LUT_2[56230] = 32'b11111111111111111111110100101101;
assign LUT_2[56231] = 32'b11111111111111111100101101000110;
assign LUT_2[56232] = 32'b11111111111111110111001111100110;
assign LUT_2[56233] = 32'b11111111111111110100000111111111;
assign LUT_2[56234] = 32'b11111111111111111110001000100010;
assign LUT_2[56235] = 32'b11111111111111111011000000111011;
assign LUT_2[56236] = 32'b11111111111111110011101101001110;
assign LUT_2[56237] = 32'b11111111111111110000100101100111;
assign LUT_2[56238] = 32'b11111111111111111010100110001010;
assign LUT_2[56239] = 32'b11111111111111110111011110100011;
assign LUT_2[56240] = 32'b11111111111111110111000010010011;
assign LUT_2[56241] = 32'b11111111111111110011111010101100;
assign LUT_2[56242] = 32'b11111111111111111101111011001111;
assign LUT_2[56243] = 32'b11111111111111111010110011101000;
assign LUT_2[56244] = 32'b11111111111111110011011111111011;
assign LUT_2[56245] = 32'b11111111111111110000011000010100;
assign LUT_2[56246] = 32'b11111111111111111010011000110111;
assign LUT_2[56247] = 32'b11111111111111110111010001010000;
assign LUT_2[56248] = 32'b11111111111111110001110011110000;
assign LUT_2[56249] = 32'b11111111111111101110101100001001;
assign LUT_2[56250] = 32'b11111111111111111000101100101100;
assign LUT_2[56251] = 32'b11111111111111110101100101000101;
assign LUT_2[56252] = 32'b11111111111111101110010001011000;
assign LUT_2[56253] = 32'b11111111111111101011001001110001;
assign LUT_2[56254] = 32'b11111111111111110101001010010100;
assign LUT_2[56255] = 32'b11111111111111110010000010101101;
assign LUT_2[56256] = 32'b11111111111111110100001011000011;
assign LUT_2[56257] = 32'b11111111111111110001000011011100;
assign LUT_2[56258] = 32'b11111111111111111011000011111111;
assign LUT_2[56259] = 32'b11111111111111110111111100011000;
assign LUT_2[56260] = 32'b11111111111111110000101000101011;
assign LUT_2[56261] = 32'b11111111111111101101100001000100;
assign LUT_2[56262] = 32'b11111111111111110111100001100111;
assign LUT_2[56263] = 32'b11111111111111110100011010000000;
assign LUT_2[56264] = 32'b11111111111111101110111100100000;
assign LUT_2[56265] = 32'b11111111111111101011110100111001;
assign LUT_2[56266] = 32'b11111111111111110101110101011100;
assign LUT_2[56267] = 32'b11111111111111110010101101110101;
assign LUT_2[56268] = 32'b11111111111111101011011010001000;
assign LUT_2[56269] = 32'b11111111111111101000010010100001;
assign LUT_2[56270] = 32'b11111111111111110010010011000100;
assign LUT_2[56271] = 32'b11111111111111101111001011011101;
assign LUT_2[56272] = 32'b11111111111111101110101111001101;
assign LUT_2[56273] = 32'b11111111111111101011100111100110;
assign LUT_2[56274] = 32'b11111111111111110101101000001001;
assign LUT_2[56275] = 32'b11111111111111110010100000100010;
assign LUT_2[56276] = 32'b11111111111111101011001100110101;
assign LUT_2[56277] = 32'b11111111111111101000000101001110;
assign LUT_2[56278] = 32'b11111111111111110010000101110001;
assign LUT_2[56279] = 32'b11111111111111101110111110001010;
assign LUT_2[56280] = 32'b11111111111111101001100000101010;
assign LUT_2[56281] = 32'b11111111111111100110011001000011;
assign LUT_2[56282] = 32'b11111111111111110000011001100110;
assign LUT_2[56283] = 32'b11111111111111101101010001111111;
assign LUT_2[56284] = 32'b11111111111111100101111110010010;
assign LUT_2[56285] = 32'b11111111111111100010110110101011;
assign LUT_2[56286] = 32'b11111111111111101100110111001110;
assign LUT_2[56287] = 32'b11111111111111101001101111100111;
assign LUT_2[56288] = 32'b11111111111111110100100110101100;
assign LUT_2[56289] = 32'b11111111111111110001011111000101;
assign LUT_2[56290] = 32'b11111111111111111011011111101000;
assign LUT_2[56291] = 32'b11111111111111111000011000000001;
assign LUT_2[56292] = 32'b11111111111111110001000100010100;
assign LUT_2[56293] = 32'b11111111111111101101111100101101;
assign LUT_2[56294] = 32'b11111111111111110111111101010000;
assign LUT_2[56295] = 32'b11111111111111110100110101101001;
assign LUT_2[56296] = 32'b11111111111111101111011000001001;
assign LUT_2[56297] = 32'b11111111111111101100010000100010;
assign LUT_2[56298] = 32'b11111111111111110110010001000101;
assign LUT_2[56299] = 32'b11111111111111110011001001011110;
assign LUT_2[56300] = 32'b11111111111111101011110101110001;
assign LUT_2[56301] = 32'b11111111111111101000101110001010;
assign LUT_2[56302] = 32'b11111111111111110010101110101101;
assign LUT_2[56303] = 32'b11111111111111101111100111000110;
assign LUT_2[56304] = 32'b11111111111111101111001010110110;
assign LUT_2[56305] = 32'b11111111111111101100000011001111;
assign LUT_2[56306] = 32'b11111111111111110110000011110010;
assign LUT_2[56307] = 32'b11111111111111110010111100001011;
assign LUT_2[56308] = 32'b11111111111111101011101000011110;
assign LUT_2[56309] = 32'b11111111111111101000100000110111;
assign LUT_2[56310] = 32'b11111111111111110010100001011010;
assign LUT_2[56311] = 32'b11111111111111101111011001110011;
assign LUT_2[56312] = 32'b11111111111111101001111100010011;
assign LUT_2[56313] = 32'b11111111111111100110110100101100;
assign LUT_2[56314] = 32'b11111111111111110000110101001111;
assign LUT_2[56315] = 32'b11111111111111101101101101101000;
assign LUT_2[56316] = 32'b11111111111111100110011001111011;
assign LUT_2[56317] = 32'b11111111111111100011010010010100;
assign LUT_2[56318] = 32'b11111111111111101101010010110111;
assign LUT_2[56319] = 32'b11111111111111101010001011010000;
assign LUT_2[56320] = 32'b11111111111111110101101001111110;
assign LUT_2[56321] = 32'b11111111111111110010100010010111;
assign LUT_2[56322] = 32'b11111111111111111100100010111010;
assign LUT_2[56323] = 32'b11111111111111111001011011010011;
assign LUT_2[56324] = 32'b11111111111111110010000111100110;
assign LUT_2[56325] = 32'b11111111111111101110111111111111;
assign LUT_2[56326] = 32'b11111111111111111001000000100010;
assign LUT_2[56327] = 32'b11111111111111110101111000111011;
assign LUT_2[56328] = 32'b11111111111111110000011011011011;
assign LUT_2[56329] = 32'b11111111111111101101010011110100;
assign LUT_2[56330] = 32'b11111111111111110111010100010111;
assign LUT_2[56331] = 32'b11111111111111110100001100110000;
assign LUT_2[56332] = 32'b11111111111111101100111001000011;
assign LUT_2[56333] = 32'b11111111111111101001110001011100;
assign LUT_2[56334] = 32'b11111111111111110011110001111111;
assign LUT_2[56335] = 32'b11111111111111110000101010011000;
assign LUT_2[56336] = 32'b11111111111111110000001110001000;
assign LUT_2[56337] = 32'b11111111111111101101000110100001;
assign LUT_2[56338] = 32'b11111111111111110111000111000100;
assign LUT_2[56339] = 32'b11111111111111110011111111011101;
assign LUT_2[56340] = 32'b11111111111111101100101011110000;
assign LUT_2[56341] = 32'b11111111111111101001100100001001;
assign LUT_2[56342] = 32'b11111111111111110011100100101100;
assign LUT_2[56343] = 32'b11111111111111110000011101000101;
assign LUT_2[56344] = 32'b11111111111111101010111111100101;
assign LUT_2[56345] = 32'b11111111111111100111110111111110;
assign LUT_2[56346] = 32'b11111111111111110001111000100001;
assign LUT_2[56347] = 32'b11111111111111101110110000111010;
assign LUT_2[56348] = 32'b11111111111111100111011101001101;
assign LUT_2[56349] = 32'b11111111111111100100010101100110;
assign LUT_2[56350] = 32'b11111111111111101110010110001001;
assign LUT_2[56351] = 32'b11111111111111101011001110100010;
assign LUT_2[56352] = 32'b11111111111111110110000101100111;
assign LUT_2[56353] = 32'b11111111111111110010111110000000;
assign LUT_2[56354] = 32'b11111111111111111100111110100011;
assign LUT_2[56355] = 32'b11111111111111111001110110111100;
assign LUT_2[56356] = 32'b11111111111111110010100011001111;
assign LUT_2[56357] = 32'b11111111111111101111011011101000;
assign LUT_2[56358] = 32'b11111111111111111001011100001011;
assign LUT_2[56359] = 32'b11111111111111110110010100100100;
assign LUT_2[56360] = 32'b11111111111111110000110111000100;
assign LUT_2[56361] = 32'b11111111111111101101101111011101;
assign LUT_2[56362] = 32'b11111111111111110111110000000000;
assign LUT_2[56363] = 32'b11111111111111110100101000011001;
assign LUT_2[56364] = 32'b11111111111111101101010100101100;
assign LUT_2[56365] = 32'b11111111111111101010001101000101;
assign LUT_2[56366] = 32'b11111111111111110100001101101000;
assign LUT_2[56367] = 32'b11111111111111110001000110000001;
assign LUT_2[56368] = 32'b11111111111111110000101001110001;
assign LUT_2[56369] = 32'b11111111111111101101100010001010;
assign LUT_2[56370] = 32'b11111111111111110111100010101101;
assign LUT_2[56371] = 32'b11111111111111110100011011000110;
assign LUT_2[56372] = 32'b11111111111111101101000111011001;
assign LUT_2[56373] = 32'b11111111111111101001111111110010;
assign LUT_2[56374] = 32'b11111111111111110100000000010101;
assign LUT_2[56375] = 32'b11111111111111110000111000101110;
assign LUT_2[56376] = 32'b11111111111111101011011011001110;
assign LUT_2[56377] = 32'b11111111111111101000010011100111;
assign LUT_2[56378] = 32'b11111111111111110010010100001010;
assign LUT_2[56379] = 32'b11111111111111101111001100100011;
assign LUT_2[56380] = 32'b11111111111111100111111000110110;
assign LUT_2[56381] = 32'b11111111111111100100110001001111;
assign LUT_2[56382] = 32'b11111111111111101110110001110010;
assign LUT_2[56383] = 32'b11111111111111101011101010001011;
assign LUT_2[56384] = 32'b11111111111111101101110010100001;
assign LUT_2[56385] = 32'b11111111111111101010101010111010;
assign LUT_2[56386] = 32'b11111111111111110100101011011101;
assign LUT_2[56387] = 32'b11111111111111110001100011110110;
assign LUT_2[56388] = 32'b11111111111111101010010000001001;
assign LUT_2[56389] = 32'b11111111111111100111001000100010;
assign LUT_2[56390] = 32'b11111111111111110001001001000101;
assign LUT_2[56391] = 32'b11111111111111101110000001011110;
assign LUT_2[56392] = 32'b11111111111111101000100011111110;
assign LUT_2[56393] = 32'b11111111111111100101011100010111;
assign LUT_2[56394] = 32'b11111111111111101111011100111010;
assign LUT_2[56395] = 32'b11111111111111101100010101010011;
assign LUT_2[56396] = 32'b11111111111111100101000001100110;
assign LUT_2[56397] = 32'b11111111111111100001111001111111;
assign LUT_2[56398] = 32'b11111111111111101011111010100010;
assign LUT_2[56399] = 32'b11111111111111101000110010111011;
assign LUT_2[56400] = 32'b11111111111111101000010110101011;
assign LUT_2[56401] = 32'b11111111111111100101001111000100;
assign LUT_2[56402] = 32'b11111111111111101111001111100111;
assign LUT_2[56403] = 32'b11111111111111101100001000000000;
assign LUT_2[56404] = 32'b11111111111111100100110100010011;
assign LUT_2[56405] = 32'b11111111111111100001101100101100;
assign LUT_2[56406] = 32'b11111111111111101011101101001111;
assign LUT_2[56407] = 32'b11111111111111101000100101101000;
assign LUT_2[56408] = 32'b11111111111111100011001000001000;
assign LUT_2[56409] = 32'b11111111111111100000000000100001;
assign LUT_2[56410] = 32'b11111111111111101010000001000100;
assign LUT_2[56411] = 32'b11111111111111100110111001011101;
assign LUT_2[56412] = 32'b11111111111111011111100101110000;
assign LUT_2[56413] = 32'b11111111111111011100011110001001;
assign LUT_2[56414] = 32'b11111111111111100110011110101100;
assign LUT_2[56415] = 32'b11111111111111100011010111000101;
assign LUT_2[56416] = 32'b11111111111111101110001110001010;
assign LUT_2[56417] = 32'b11111111111111101011000110100011;
assign LUT_2[56418] = 32'b11111111111111110101000111000110;
assign LUT_2[56419] = 32'b11111111111111110001111111011111;
assign LUT_2[56420] = 32'b11111111111111101010101011110010;
assign LUT_2[56421] = 32'b11111111111111100111100100001011;
assign LUT_2[56422] = 32'b11111111111111110001100100101110;
assign LUT_2[56423] = 32'b11111111111111101110011101000111;
assign LUT_2[56424] = 32'b11111111111111101000111111100111;
assign LUT_2[56425] = 32'b11111111111111100101111000000000;
assign LUT_2[56426] = 32'b11111111111111101111111000100011;
assign LUT_2[56427] = 32'b11111111111111101100110000111100;
assign LUT_2[56428] = 32'b11111111111111100101011101001111;
assign LUT_2[56429] = 32'b11111111111111100010010101101000;
assign LUT_2[56430] = 32'b11111111111111101100010110001011;
assign LUT_2[56431] = 32'b11111111111111101001001110100100;
assign LUT_2[56432] = 32'b11111111111111101000110010010100;
assign LUT_2[56433] = 32'b11111111111111100101101010101101;
assign LUT_2[56434] = 32'b11111111111111101111101011010000;
assign LUT_2[56435] = 32'b11111111111111101100100011101001;
assign LUT_2[56436] = 32'b11111111111111100101001111111100;
assign LUT_2[56437] = 32'b11111111111111100010001000010101;
assign LUT_2[56438] = 32'b11111111111111101100001000111000;
assign LUT_2[56439] = 32'b11111111111111101001000001010001;
assign LUT_2[56440] = 32'b11111111111111100011100011110001;
assign LUT_2[56441] = 32'b11111111111111100000011100001010;
assign LUT_2[56442] = 32'b11111111111111101010011100101101;
assign LUT_2[56443] = 32'b11111111111111100111010101000110;
assign LUT_2[56444] = 32'b11111111111111100000000001011001;
assign LUT_2[56445] = 32'b11111111111111011100111001110010;
assign LUT_2[56446] = 32'b11111111111111100110111010010101;
assign LUT_2[56447] = 32'b11111111111111100011110010101110;
assign LUT_2[56448] = 32'b11111111111111111001111110001101;
assign LUT_2[56449] = 32'b11111111111111110110110110100110;
assign LUT_2[56450] = 32'b00000000000000000000110111001001;
assign LUT_2[56451] = 32'b11111111111111111101101111100010;
assign LUT_2[56452] = 32'b11111111111111110110011011110101;
assign LUT_2[56453] = 32'b11111111111111110011010100001110;
assign LUT_2[56454] = 32'b11111111111111111101010100110001;
assign LUT_2[56455] = 32'b11111111111111111010001101001010;
assign LUT_2[56456] = 32'b11111111111111110100101111101010;
assign LUT_2[56457] = 32'b11111111111111110001101000000011;
assign LUT_2[56458] = 32'b11111111111111111011101000100110;
assign LUT_2[56459] = 32'b11111111111111111000100000111111;
assign LUT_2[56460] = 32'b11111111111111110001001101010010;
assign LUT_2[56461] = 32'b11111111111111101110000101101011;
assign LUT_2[56462] = 32'b11111111111111111000000110001110;
assign LUT_2[56463] = 32'b11111111111111110100111110100111;
assign LUT_2[56464] = 32'b11111111111111110100100010010111;
assign LUT_2[56465] = 32'b11111111111111110001011010110000;
assign LUT_2[56466] = 32'b11111111111111111011011011010011;
assign LUT_2[56467] = 32'b11111111111111111000010011101100;
assign LUT_2[56468] = 32'b11111111111111110000111111111111;
assign LUT_2[56469] = 32'b11111111111111101101111000011000;
assign LUT_2[56470] = 32'b11111111111111110111111000111011;
assign LUT_2[56471] = 32'b11111111111111110100110001010100;
assign LUT_2[56472] = 32'b11111111111111101111010011110100;
assign LUT_2[56473] = 32'b11111111111111101100001100001101;
assign LUT_2[56474] = 32'b11111111111111110110001100110000;
assign LUT_2[56475] = 32'b11111111111111110011000101001001;
assign LUT_2[56476] = 32'b11111111111111101011110001011100;
assign LUT_2[56477] = 32'b11111111111111101000101001110101;
assign LUT_2[56478] = 32'b11111111111111110010101010011000;
assign LUT_2[56479] = 32'b11111111111111101111100010110001;
assign LUT_2[56480] = 32'b11111111111111111010011001110110;
assign LUT_2[56481] = 32'b11111111111111110111010010001111;
assign LUT_2[56482] = 32'b00000000000000000001010010110010;
assign LUT_2[56483] = 32'b11111111111111111110001011001011;
assign LUT_2[56484] = 32'b11111111111111110110110111011110;
assign LUT_2[56485] = 32'b11111111111111110011101111110111;
assign LUT_2[56486] = 32'b11111111111111111101110000011010;
assign LUT_2[56487] = 32'b11111111111111111010101000110011;
assign LUT_2[56488] = 32'b11111111111111110101001011010011;
assign LUT_2[56489] = 32'b11111111111111110010000011101100;
assign LUT_2[56490] = 32'b11111111111111111100000100001111;
assign LUT_2[56491] = 32'b11111111111111111000111100101000;
assign LUT_2[56492] = 32'b11111111111111110001101000111011;
assign LUT_2[56493] = 32'b11111111111111101110100001010100;
assign LUT_2[56494] = 32'b11111111111111111000100001110111;
assign LUT_2[56495] = 32'b11111111111111110101011010010000;
assign LUT_2[56496] = 32'b11111111111111110100111110000000;
assign LUT_2[56497] = 32'b11111111111111110001110110011001;
assign LUT_2[56498] = 32'b11111111111111111011110110111100;
assign LUT_2[56499] = 32'b11111111111111111000101111010101;
assign LUT_2[56500] = 32'b11111111111111110001011011101000;
assign LUT_2[56501] = 32'b11111111111111101110010100000001;
assign LUT_2[56502] = 32'b11111111111111111000010100100100;
assign LUT_2[56503] = 32'b11111111111111110101001100111101;
assign LUT_2[56504] = 32'b11111111111111101111101111011101;
assign LUT_2[56505] = 32'b11111111111111101100100111110110;
assign LUT_2[56506] = 32'b11111111111111110110101000011001;
assign LUT_2[56507] = 32'b11111111111111110011100000110010;
assign LUT_2[56508] = 32'b11111111111111101100001101000101;
assign LUT_2[56509] = 32'b11111111111111101001000101011110;
assign LUT_2[56510] = 32'b11111111111111110011000110000001;
assign LUT_2[56511] = 32'b11111111111111101111111110011010;
assign LUT_2[56512] = 32'b11111111111111110010000110110000;
assign LUT_2[56513] = 32'b11111111111111101110111111001001;
assign LUT_2[56514] = 32'b11111111111111111000111111101100;
assign LUT_2[56515] = 32'b11111111111111110101111000000101;
assign LUT_2[56516] = 32'b11111111111111101110100100011000;
assign LUT_2[56517] = 32'b11111111111111101011011100110001;
assign LUT_2[56518] = 32'b11111111111111110101011101010100;
assign LUT_2[56519] = 32'b11111111111111110010010101101101;
assign LUT_2[56520] = 32'b11111111111111101100111000001101;
assign LUT_2[56521] = 32'b11111111111111101001110000100110;
assign LUT_2[56522] = 32'b11111111111111110011110001001001;
assign LUT_2[56523] = 32'b11111111111111110000101001100010;
assign LUT_2[56524] = 32'b11111111111111101001010101110101;
assign LUT_2[56525] = 32'b11111111111111100110001110001110;
assign LUT_2[56526] = 32'b11111111111111110000001110110001;
assign LUT_2[56527] = 32'b11111111111111101101000111001010;
assign LUT_2[56528] = 32'b11111111111111101100101010111010;
assign LUT_2[56529] = 32'b11111111111111101001100011010011;
assign LUT_2[56530] = 32'b11111111111111110011100011110110;
assign LUT_2[56531] = 32'b11111111111111110000011100001111;
assign LUT_2[56532] = 32'b11111111111111101001001000100010;
assign LUT_2[56533] = 32'b11111111111111100110000000111011;
assign LUT_2[56534] = 32'b11111111111111110000000001011110;
assign LUT_2[56535] = 32'b11111111111111101100111001110111;
assign LUT_2[56536] = 32'b11111111111111100111011100010111;
assign LUT_2[56537] = 32'b11111111111111100100010100110000;
assign LUT_2[56538] = 32'b11111111111111101110010101010011;
assign LUT_2[56539] = 32'b11111111111111101011001101101100;
assign LUT_2[56540] = 32'b11111111111111100011111001111111;
assign LUT_2[56541] = 32'b11111111111111100000110010011000;
assign LUT_2[56542] = 32'b11111111111111101010110010111011;
assign LUT_2[56543] = 32'b11111111111111100111101011010100;
assign LUT_2[56544] = 32'b11111111111111110010100010011001;
assign LUT_2[56545] = 32'b11111111111111101111011010110010;
assign LUT_2[56546] = 32'b11111111111111111001011011010101;
assign LUT_2[56547] = 32'b11111111111111110110010011101110;
assign LUT_2[56548] = 32'b11111111111111101111000000000001;
assign LUT_2[56549] = 32'b11111111111111101011111000011010;
assign LUT_2[56550] = 32'b11111111111111110101111000111101;
assign LUT_2[56551] = 32'b11111111111111110010110001010110;
assign LUT_2[56552] = 32'b11111111111111101101010011110110;
assign LUT_2[56553] = 32'b11111111111111101010001100001111;
assign LUT_2[56554] = 32'b11111111111111110100001100110010;
assign LUT_2[56555] = 32'b11111111111111110001000101001011;
assign LUT_2[56556] = 32'b11111111111111101001110001011110;
assign LUT_2[56557] = 32'b11111111111111100110101001110111;
assign LUT_2[56558] = 32'b11111111111111110000101010011010;
assign LUT_2[56559] = 32'b11111111111111101101100010110011;
assign LUT_2[56560] = 32'b11111111111111101101000110100011;
assign LUT_2[56561] = 32'b11111111111111101001111110111100;
assign LUT_2[56562] = 32'b11111111111111110011111111011111;
assign LUT_2[56563] = 32'b11111111111111110000110111111000;
assign LUT_2[56564] = 32'b11111111111111101001100100001011;
assign LUT_2[56565] = 32'b11111111111111100110011100100100;
assign LUT_2[56566] = 32'b11111111111111110000011101000111;
assign LUT_2[56567] = 32'b11111111111111101101010101100000;
assign LUT_2[56568] = 32'b11111111111111100111111000000000;
assign LUT_2[56569] = 32'b11111111111111100100110000011001;
assign LUT_2[56570] = 32'b11111111111111101110110000111100;
assign LUT_2[56571] = 32'b11111111111111101011101001010101;
assign LUT_2[56572] = 32'b11111111111111100100010101101000;
assign LUT_2[56573] = 32'b11111111111111100001001110000001;
assign LUT_2[56574] = 32'b11111111111111101011001110100100;
assign LUT_2[56575] = 32'b11111111111111101000000110111101;
assign LUT_2[56576] = 32'b11111111111111111001101000100100;
assign LUT_2[56577] = 32'b11111111111111110110100000111101;
assign LUT_2[56578] = 32'b00000000000000000000100001100000;
assign LUT_2[56579] = 32'b11111111111111111101011001111001;
assign LUT_2[56580] = 32'b11111111111111110110000110001100;
assign LUT_2[56581] = 32'b11111111111111110010111110100101;
assign LUT_2[56582] = 32'b11111111111111111100111111001000;
assign LUT_2[56583] = 32'b11111111111111111001110111100001;
assign LUT_2[56584] = 32'b11111111111111110100011010000001;
assign LUT_2[56585] = 32'b11111111111111110001010010011010;
assign LUT_2[56586] = 32'b11111111111111111011010010111101;
assign LUT_2[56587] = 32'b11111111111111111000001011010110;
assign LUT_2[56588] = 32'b11111111111111110000110111101001;
assign LUT_2[56589] = 32'b11111111111111101101110000000010;
assign LUT_2[56590] = 32'b11111111111111110111110000100101;
assign LUT_2[56591] = 32'b11111111111111110100101000111110;
assign LUT_2[56592] = 32'b11111111111111110100001100101110;
assign LUT_2[56593] = 32'b11111111111111110001000101000111;
assign LUT_2[56594] = 32'b11111111111111111011000101101010;
assign LUT_2[56595] = 32'b11111111111111110111111110000011;
assign LUT_2[56596] = 32'b11111111111111110000101010010110;
assign LUT_2[56597] = 32'b11111111111111101101100010101111;
assign LUT_2[56598] = 32'b11111111111111110111100011010010;
assign LUT_2[56599] = 32'b11111111111111110100011011101011;
assign LUT_2[56600] = 32'b11111111111111101110111110001011;
assign LUT_2[56601] = 32'b11111111111111101011110110100100;
assign LUT_2[56602] = 32'b11111111111111110101110111000111;
assign LUT_2[56603] = 32'b11111111111111110010101111100000;
assign LUT_2[56604] = 32'b11111111111111101011011011110011;
assign LUT_2[56605] = 32'b11111111111111101000010100001100;
assign LUT_2[56606] = 32'b11111111111111110010010100101111;
assign LUT_2[56607] = 32'b11111111111111101111001101001000;
assign LUT_2[56608] = 32'b11111111111111111010000100001101;
assign LUT_2[56609] = 32'b11111111111111110110111100100110;
assign LUT_2[56610] = 32'b00000000000000000000111101001001;
assign LUT_2[56611] = 32'b11111111111111111101110101100010;
assign LUT_2[56612] = 32'b11111111111111110110100001110101;
assign LUT_2[56613] = 32'b11111111111111110011011010001110;
assign LUT_2[56614] = 32'b11111111111111111101011010110001;
assign LUT_2[56615] = 32'b11111111111111111010010011001010;
assign LUT_2[56616] = 32'b11111111111111110100110101101010;
assign LUT_2[56617] = 32'b11111111111111110001101110000011;
assign LUT_2[56618] = 32'b11111111111111111011101110100110;
assign LUT_2[56619] = 32'b11111111111111111000100110111111;
assign LUT_2[56620] = 32'b11111111111111110001010011010010;
assign LUT_2[56621] = 32'b11111111111111101110001011101011;
assign LUT_2[56622] = 32'b11111111111111111000001100001110;
assign LUT_2[56623] = 32'b11111111111111110101000100100111;
assign LUT_2[56624] = 32'b11111111111111110100101000010111;
assign LUT_2[56625] = 32'b11111111111111110001100000110000;
assign LUT_2[56626] = 32'b11111111111111111011100001010011;
assign LUT_2[56627] = 32'b11111111111111111000011001101100;
assign LUT_2[56628] = 32'b11111111111111110001000101111111;
assign LUT_2[56629] = 32'b11111111111111101101111110011000;
assign LUT_2[56630] = 32'b11111111111111110111111110111011;
assign LUT_2[56631] = 32'b11111111111111110100110111010100;
assign LUT_2[56632] = 32'b11111111111111101111011001110100;
assign LUT_2[56633] = 32'b11111111111111101100010010001101;
assign LUT_2[56634] = 32'b11111111111111110110010010110000;
assign LUT_2[56635] = 32'b11111111111111110011001011001001;
assign LUT_2[56636] = 32'b11111111111111101011110111011100;
assign LUT_2[56637] = 32'b11111111111111101000101111110101;
assign LUT_2[56638] = 32'b11111111111111110010110000011000;
assign LUT_2[56639] = 32'b11111111111111101111101000110001;
assign LUT_2[56640] = 32'b11111111111111110001110001000111;
assign LUT_2[56641] = 32'b11111111111111101110101001100000;
assign LUT_2[56642] = 32'b11111111111111111000101010000011;
assign LUT_2[56643] = 32'b11111111111111110101100010011100;
assign LUT_2[56644] = 32'b11111111111111101110001110101111;
assign LUT_2[56645] = 32'b11111111111111101011000111001000;
assign LUT_2[56646] = 32'b11111111111111110101000111101011;
assign LUT_2[56647] = 32'b11111111111111110010000000000100;
assign LUT_2[56648] = 32'b11111111111111101100100010100100;
assign LUT_2[56649] = 32'b11111111111111101001011010111101;
assign LUT_2[56650] = 32'b11111111111111110011011011100000;
assign LUT_2[56651] = 32'b11111111111111110000010011111001;
assign LUT_2[56652] = 32'b11111111111111101001000000001100;
assign LUT_2[56653] = 32'b11111111111111100101111000100101;
assign LUT_2[56654] = 32'b11111111111111101111111001001000;
assign LUT_2[56655] = 32'b11111111111111101100110001100001;
assign LUT_2[56656] = 32'b11111111111111101100010101010001;
assign LUT_2[56657] = 32'b11111111111111101001001101101010;
assign LUT_2[56658] = 32'b11111111111111110011001110001101;
assign LUT_2[56659] = 32'b11111111111111110000000110100110;
assign LUT_2[56660] = 32'b11111111111111101000110010111001;
assign LUT_2[56661] = 32'b11111111111111100101101011010010;
assign LUT_2[56662] = 32'b11111111111111101111101011110101;
assign LUT_2[56663] = 32'b11111111111111101100100100001110;
assign LUT_2[56664] = 32'b11111111111111100111000110101110;
assign LUT_2[56665] = 32'b11111111111111100011111111000111;
assign LUT_2[56666] = 32'b11111111111111101101111111101010;
assign LUT_2[56667] = 32'b11111111111111101010111000000011;
assign LUT_2[56668] = 32'b11111111111111100011100100010110;
assign LUT_2[56669] = 32'b11111111111111100000011100101111;
assign LUT_2[56670] = 32'b11111111111111101010011101010010;
assign LUT_2[56671] = 32'b11111111111111100111010101101011;
assign LUT_2[56672] = 32'b11111111111111110010001100110000;
assign LUT_2[56673] = 32'b11111111111111101111000101001001;
assign LUT_2[56674] = 32'b11111111111111111001000101101100;
assign LUT_2[56675] = 32'b11111111111111110101111110000101;
assign LUT_2[56676] = 32'b11111111111111101110101010011000;
assign LUT_2[56677] = 32'b11111111111111101011100010110001;
assign LUT_2[56678] = 32'b11111111111111110101100011010100;
assign LUT_2[56679] = 32'b11111111111111110010011011101101;
assign LUT_2[56680] = 32'b11111111111111101100111110001101;
assign LUT_2[56681] = 32'b11111111111111101001110110100110;
assign LUT_2[56682] = 32'b11111111111111110011110111001001;
assign LUT_2[56683] = 32'b11111111111111110000101111100010;
assign LUT_2[56684] = 32'b11111111111111101001011011110101;
assign LUT_2[56685] = 32'b11111111111111100110010100001110;
assign LUT_2[56686] = 32'b11111111111111110000010100110001;
assign LUT_2[56687] = 32'b11111111111111101101001101001010;
assign LUT_2[56688] = 32'b11111111111111101100110000111010;
assign LUT_2[56689] = 32'b11111111111111101001101001010011;
assign LUT_2[56690] = 32'b11111111111111110011101001110110;
assign LUT_2[56691] = 32'b11111111111111110000100010001111;
assign LUT_2[56692] = 32'b11111111111111101001001110100010;
assign LUT_2[56693] = 32'b11111111111111100110000110111011;
assign LUT_2[56694] = 32'b11111111111111110000000111011110;
assign LUT_2[56695] = 32'b11111111111111101100111111110111;
assign LUT_2[56696] = 32'b11111111111111100111100010010111;
assign LUT_2[56697] = 32'b11111111111111100100011010110000;
assign LUT_2[56698] = 32'b11111111111111101110011011010011;
assign LUT_2[56699] = 32'b11111111111111101011010011101100;
assign LUT_2[56700] = 32'b11111111111111100011111111111111;
assign LUT_2[56701] = 32'b11111111111111100000111000011000;
assign LUT_2[56702] = 32'b11111111111111101010111000111011;
assign LUT_2[56703] = 32'b11111111111111100111110001010100;
assign LUT_2[56704] = 32'b11111111111111111101111100110011;
assign LUT_2[56705] = 32'b11111111111111111010110101001100;
assign LUT_2[56706] = 32'b00000000000000000100110101101111;
assign LUT_2[56707] = 32'b00000000000000000001101110001000;
assign LUT_2[56708] = 32'b11111111111111111010011010011011;
assign LUT_2[56709] = 32'b11111111111111110111010010110100;
assign LUT_2[56710] = 32'b00000000000000000001010011010111;
assign LUT_2[56711] = 32'b11111111111111111110001011110000;
assign LUT_2[56712] = 32'b11111111111111111000101110010000;
assign LUT_2[56713] = 32'b11111111111111110101100110101001;
assign LUT_2[56714] = 32'b11111111111111111111100111001100;
assign LUT_2[56715] = 32'b11111111111111111100011111100101;
assign LUT_2[56716] = 32'b11111111111111110101001011111000;
assign LUT_2[56717] = 32'b11111111111111110010000100010001;
assign LUT_2[56718] = 32'b11111111111111111100000100110100;
assign LUT_2[56719] = 32'b11111111111111111000111101001101;
assign LUT_2[56720] = 32'b11111111111111111000100000111101;
assign LUT_2[56721] = 32'b11111111111111110101011001010110;
assign LUT_2[56722] = 32'b11111111111111111111011001111001;
assign LUT_2[56723] = 32'b11111111111111111100010010010010;
assign LUT_2[56724] = 32'b11111111111111110100111110100101;
assign LUT_2[56725] = 32'b11111111111111110001110110111110;
assign LUT_2[56726] = 32'b11111111111111111011110111100001;
assign LUT_2[56727] = 32'b11111111111111111000101111111010;
assign LUT_2[56728] = 32'b11111111111111110011010010011010;
assign LUT_2[56729] = 32'b11111111111111110000001010110011;
assign LUT_2[56730] = 32'b11111111111111111010001011010110;
assign LUT_2[56731] = 32'b11111111111111110111000011101111;
assign LUT_2[56732] = 32'b11111111111111101111110000000010;
assign LUT_2[56733] = 32'b11111111111111101100101000011011;
assign LUT_2[56734] = 32'b11111111111111110110101000111110;
assign LUT_2[56735] = 32'b11111111111111110011100001010111;
assign LUT_2[56736] = 32'b11111111111111111110011000011100;
assign LUT_2[56737] = 32'b11111111111111111011010000110101;
assign LUT_2[56738] = 32'b00000000000000000101010001011000;
assign LUT_2[56739] = 32'b00000000000000000010001001110001;
assign LUT_2[56740] = 32'b11111111111111111010110110000100;
assign LUT_2[56741] = 32'b11111111111111110111101110011101;
assign LUT_2[56742] = 32'b00000000000000000001101111000000;
assign LUT_2[56743] = 32'b11111111111111111110100111011001;
assign LUT_2[56744] = 32'b11111111111111111001001001111001;
assign LUT_2[56745] = 32'b11111111111111110110000010010010;
assign LUT_2[56746] = 32'b00000000000000000000000010110101;
assign LUT_2[56747] = 32'b11111111111111111100111011001110;
assign LUT_2[56748] = 32'b11111111111111110101100111100001;
assign LUT_2[56749] = 32'b11111111111111110010011111111010;
assign LUT_2[56750] = 32'b11111111111111111100100000011101;
assign LUT_2[56751] = 32'b11111111111111111001011000110110;
assign LUT_2[56752] = 32'b11111111111111111000111100100110;
assign LUT_2[56753] = 32'b11111111111111110101110100111111;
assign LUT_2[56754] = 32'b11111111111111111111110101100010;
assign LUT_2[56755] = 32'b11111111111111111100101101111011;
assign LUT_2[56756] = 32'b11111111111111110101011010001110;
assign LUT_2[56757] = 32'b11111111111111110010010010100111;
assign LUT_2[56758] = 32'b11111111111111111100010011001010;
assign LUT_2[56759] = 32'b11111111111111111001001011100011;
assign LUT_2[56760] = 32'b11111111111111110011101110000011;
assign LUT_2[56761] = 32'b11111111111111110000100110011100;
assign LUT_2[56762] = 32'b11111111111111111010100110111111;
assign LUT_2[56763] = 32'b11111111111111110111011111011000;
assign LUT_2[56764] = 32'b11111111111111110000001011101011;
assign LUT_2[56765] = 32'b11111111111111101101000100000100;
assign LUT_2[56766] = 32'b11111111111111110111000100100111;
assign LUT_2[56767] = 32'b11111111111111110011111101000000;
assign LUT_2[56768] = 32'b11111111111111110110000101010110;
assign LUT_2[56769] = 32'b11111111111111110010111101101111;
assign LUT_2[56770] = 32'b11111111111111111100111110010010;
assign LUT_2[56771] = 32'b11111111111111111001110110101011;
assign LUT_2[56772] = 32'b11111111111111110010100010111110;
assign LUT_2[56773] = 32'b11111111111111101111011011010111;
assign LUT_2[56774] = 32'b11111111111111111001011011111010;
assign LUT_2[56775] = 32'b11111111111111110110010100010011;
assign LUT_2[56776] = 32'b11111111111111110000110110110011;
assign LUT_2[56777] = 32'b11111111111111101101101111001100;
assign LUT_2[56778] = 32'b11111111111111110111101111101111;
assign LUT_2[56779] = 32'b11111111111111110100101000001000;
assign LUT_2[56780] = 32'b11111111111111101101010100011011;
assign LUT_2[56781] = 32'b11111111111111101010001100110100;
assign LUT_2[56782] = 32'b11111111111111110100001101010111;
assign LUT_2[56783] = 32'b11111111111111110001000101110000;
assign LUT_2[56784] = 32'b11111111111111110000101001100000;
assign LUT_2[56785] = 32'b11111111111111101101100001111001;
assign LUT_2[56786] = 32'b11111111111111110111100010011100;
assign LUT_2[56787] = 32'b11111111111111110100011010110101;
assign LUT_2[56788] = 32'b11111111111111101101000111001000;
assign LUT_2[56789] = 32'b11111111111111101001111111100001;
assign LUT_2[56790] = 32'b11111111111111110100000000000100;
assign LUT_2[56791] = 32'b11111111111111110000111000011101;
assign LUT_2[56792] = 32'b11111111111111101011011010111101;
assign LUT_2[56793] = 32'b11111111111111101000010011010110;
assign LUT_2[56794] = 32'b11111111111111110010010011111001;
assign LUT_2[56795] = 32'b11111111111111101111001100010010;
assign LUT_2[56796] = 32'b11111111111111100111111000100101;
assign LUT_2[56797] = 32'b11111111111111100100110000111110;
assign LUT_2[56798] = 32'b11111111111111101110110001100001;
assign LUT_2[56799] = 32'b11111111111111101011101001111010;
assign LUT_2[56800] = 32'b11111111111111110110100000111111;
assign LUT_2[56801] = 32'b11111111111111110011011001011000;
assign LUT_2[56802] = 32'b11111111111111111101011001111011;
assign LUT_2[56803] = 32'b11111111111111111010010010010100;
assign LUT_2[56804] = 32'b11111111111111110010111110100111;
assign LUT_2[56805] = 32'b11111111111111101111110111000000;
assign LUT_2[56806] = 32'b11111111111111111001110111100011;
assign LUT_2[56807] = 32'b11111111111111110110101111111100;
assign LUT_2[56808] = 32'b11111111111111110001010010011100;
assign LUT_2[56809] = 32'b11111111111111101110001010110101;
assign LUT_2[56810] = 32'b11111111111111111000001011011000;
assign LUT_2[56811] = 32'b11111111111111110101000011110001;
assign LUT_2[56812] = 32'b11111111111111101101110000000100;
assign LUT_2[56813] = 32'b11111111111111101010101000011101;
assign LUT_2[56814] = 32'b11111111111111110100101001000000;
assign LUT_2[56815] = 32'b11111111111111110001100001011001;
assign LUT_2[56816] = 32'b11111111111111110001000101001001;
assign LUT_2[56817] = 32'b11111111111111101101111101100010;
assign LUT_2[56818] = 32'b11111111111111110111111110000101;
assign LUT_2[56819] = 32'b11111111111111110100110110011110;
assign LUT_2[56820] = 32'b11111111111111101101100010110001;
assign LUT_2[56821] = 32'b11111111111111101010011011001010;
assign LUT_2[56822] = 32'b11111111111111110100011011101101;
assign LUT_2[56823] = 32'b11111111111111110001010100000110;
assign LUT_2[56824] = 32'b11111111111111101011110110100110;
assign LUT_2[56825] = 32'b11111111111111101000101110111111;
assign LUT_2[56826] = 32'b11111111111111110010101111100010;
assign LUT_2[56827] = 32'b11111111111111101111100111111011;
assign LUT_2[56828] = 32'b11111111111111101000010100001110;
assign LUT_2[56829] = 32'b11111111111111100101001100100111;
assign LUT_2[56830] = 32'b11111111111111101111001101001010;
assign LUT_2[56831] = 32'b11111111111111101100000101100011;
assign LUT_2[56832] = 32'b11111111111111111010011011110000;
assign LUT_2[56833] = 32'b11111111111111110111010100001001;
assign LUT_2[56834] = 32'b00000000000000000001010100101100;
assign LUT_2[56835] = 32'b11111111111111111110001101000101;
assign LUT_2[56836] = 32'b11111111111111110110111001011000;
assign LUT_2[56837] = 32'b11111111111111110011110001110001;
assign LUT_2[56838] = 32'b11111111111111111101110010010100;
assign LUT_2[56839] = 32'b11111111111111111010101010101101;
assign LUT_2[56840] = 32'b11111111111111110101001101001101;
assign LUT_2[56841] = 32'b11111111111111110010000101100110;
assign LUT_2[56842] = 32'b11111111111111111100000110001001;
assign LUT_2[56843] = 32'b11111111111111111000111110100010;
assign LUT_2[56844] = 32'b11111111111111110001101010110101;
assign LUT_2[56845] = 32'b11111111111111101110100011001110;
assign LUT_2[56846] = 32'b11111111111111111000100011110001;
assign LUT_2[56847] = 32'b11111111111111110101011100001010;
assign LUT_2[56848] = 32'b11111111111111110100111111111010;
assign LUT_2[56849] = 32'b11111111111111110001111000010011;
assign LUT_2[56850] = 32'b11111111111111111011111000110110;
assign LUT_2[56851] = 32'b11111111111111111000110001001111;
assign LUT_2[56852] = 32'b11111111111111110001011101100010;
assign LUT_2[56853] = 32'b11111111111111101110010101111011;
assign LUT_2[56854] = 32'b11111111111111111000010110011110;
assign LUT_2[56855] = 32'b11111111111111110101001110110111;
assign LUT_2[56856] = 32'b11111111111111101111110001010111;
assign LUT_2[56857] = 32'b11111111111111101100101001110000;
assign LUT_2[56858] = 32'b11111111111111110110101010010011;
assign LUT_2[56859] = 32'b11111111111111110011100010101100;
assign LUT_2[56860] = 32'b11111111111111101100001110111111;
assign LUT_2[56861] = 32'b11111111111111101001000111011000;
assign LUT_2[56862] = 32'b11111111111111110011000111111011;
assign LUT_2[56863] = 32'b11111111111111110000000000010100;
assign LUT_2[56864] = 32'b11111111111111111010110111011001;
assign LUT_2[56865] = 32'b11111111111111110111101111110010;
assign LUT_2[56866] = 32'b00000000000000000001110000010101;
assign LUT_2[56867] = 32'b11111111111111111110101000101110;
assign LUT_2[56868] = 32'b11111111111111110111010101000001;
assign LUT_2[56869] = 32'b11111111111111110100001101011010;
assign LUT_2[56870] = 32'b11111111111111111110001101111101;
assign LUT_2[56871] = 32'b11111111111111111011000110010110;
assign LUT_2[56872] = 32'b11111111111111110101101000110110;
assign LUT_2[56873] = 32'b11111111111111110010100001001111;
assign LUT_2[56874] = 32'b11111111111111111100100001110010;
assign LUT_2[56875] = 32'b11111111111111111001011010001011;
assign LUT_2[56876] = 32'b11111111111111110010000110011110;
assign LUT_2[56877] = 32'b11111111111111101110111110110111;
assign LUT_2[56878] = 32'b11111111111111111000111111011010;
assign LUT_2[56879] = 32'b11111111111111110101110111110011;
assign LUT_2[56880] = 32'b11111111111111110101011011100011;
assign LUT_2[56881] = 32'b11111111111111110010010011111100;
assign LUT_2[56882] = 32'b11111111111111111100010100011111;
assign LUT_2[56883] = 32'b11111111111111111001001100111000;
assign LUT_2[56884] = 32'b11111111111111110001111001001011;
assign LUT_2[56885] = 32'b11111111111111101110110001100100;
assign LUT_2[56886] = 32'b11111111111111111000110010000111;
assign LUT_2[56887] = 32'b11111111111111110101101010100000;
assign LUT_2[56888] = 32'b11111111111111110000001101000000;
assign LUT_2[56889] = 32'b11111111111111101101000101011001;
assign LUT_2[56890] = 32'b11111111111111110111000101111100;
assign LUT_2[56891] = 32'b11111111111111110011111110010101;
assign LUT_2[56892] = 32'b11111111111111101100101010101000;
assign LUT_2[56893] = 32'b11111111111111101001100011000001;
assign LUT_2[56894] = 32'b11111111111111110011100011100100;
assign LUT_2[56895] = 32'b11111111111111110000011011111101;
assign LUT_2[56896] = 32'b11111111111111110010100100010011;
assign LUT_2[56897] = 32'b11111111111111101111011100101100;
assign LUT_2[56898] = 32'b11111111111111111001011101001111;
assign LUT_2[56899] = 32'b11111111111111110110010101101000;
assign LUT_2[56900] = 32'b11111111111111101111000001111011;
assign LUT_2[56901] = 32'b11111111111111101011111010010100;
assign LUT_2[56902] = 32'b11111111111111110101111010110111;
assign LUT_2[56903] = 32'b11111111111111110010110011010000;
assign LUT_2[56904] = 32'b11111111111111101101010101110000;
assign LUT_2[56905] = 32'b11111111111111101010001110001001;
assign LUT_2[56906] = 32'b11111111111111110100001110101100;
assign LUT_2[56907] = 32'b11111111111111110001000111000101;
assign LUT_2[56908] = 32'b11111111111111101001110011011000;
assign LUT_2[56909] = 32'b11111111111111100110101011110001;
assign LUT_2[56910] = 32'b11111111111111110000101100010100;
assign LUT_2[56911] = 32'b11111111111111101101100100101101;
assign LUT_2[56912] = 32'b11111111111111101101001000011101;
assign LUT_2[56913] = 32'b11111111111111101010000000110110;
assign LUT_2[56914] = 32'b11111111111111110100000001011001;
assign LUT_2[56915] = 32'b11111111111111110000111001110010;
assign LUT_2[56916] = 32'b11111111111111101001100110000101;
assign LUT_2[56917] = 32'b11111111111111100110011110011110;
assign LUT_2[56918] = 32'b11111111111111110000011111000001;
assign LUT_2[56919] = 32'b11111111111111101101010111011010;
assign LUT_2[56920] = 32'b11111111111111100111111001111010;
assign LUT_2[56921] = 32'b11111111111111100100110010010011;
assign LUT_2[56922] = 32'b11111111111111101110110010110110;
assign LUT_2[56923] = 32'b11111111111111101011101011001111;
assign LUT_2[56924] = 32'b11111111111111100100010111100010;
assign LUT_2[56925] = 32'b11111111111111100001001111111011;
assign LUT_2[56926] = 32'b11111111111111101011010000011110;
assign LUT_2[56927] = 32'b11111111111111101000001000110111;
assign LUT_2[56928] = 32'b11111111111111110010111111111100;
assign LUT_2[56929] = 32'b11111111111111101111111000010101;
assign LUT_2[56930] = 32'b11111111111111111001111000111000;
assign LUT_2[56931] = 32'b11111111111111110110110001010001;
assign LUT_2[56932] = 32'b11111111111111101111011101100100;
assign LUT_2[56933] = 32'b11111111111111101100010101111101;
assign LUT_2[56934] = 32'b11111111111111110110010110100000;
assign LUT_2[56935] = 32'b11111111111111110011001110111001;
assign LUT_2[56936] = 32'b11111111111111101101110001011001;
assign LUT_2[56937] = 32'b11111111111111101010101001110010;
assign LUT_2[56938] = 32'b11111111111111110100101010010101;
assign LUT_2[56939] = 32'b11111111111111110001100010101110;
assign LUT_2[56940] = 32'b11111111111111101010001111000001;
assign LUT_2[56941] = 32'b11111111111111100111000111011010;
assign LUT_2[56942] = 32'b11111111111111110001000111111101;
assign LUT_2[56943] = 32'b11111111111111101110000000010110;
assign LUT_2[56944] = 32'b11111111111111101101100100000110;
assign LUT_2[56945] = 32'b11111111111111101010011100011111;
assign LUT_2[56946] = 32'b11111111111111110100011101000010;
assign LUT_2[56947] = 32'b11111111111111110001010101011011;
assign LUT_2[56948] = 32'b11111111111111101010000001101110;
assign LUT_2[56949] = 32'b11111111111111100110111010000111;
assign LUT_2[56950] = 32'b11111111111111110000111010101010;
assign LUT_2[56951] = 32'b11111111111111101101110011000011;
assign LUT_2[56952] = 32'b11111111111111101000010101100011;
assign LUT_2[56953] = 32'b11111111111111100101001101111100;
assign LUT_2[56954] = 32'b11111111111111101111001110011111;
assign LUT_2[56955] = 32'b11111111111111101100000110111000;
assign LUT_2[56956] = 32'b11111111111111100100110011001011;
assign LUT_2[56957] = 32'b11111111111111100001101011100100;
assign LUT_2[56958] = 32'b11111111111111101011101100000111;
assign LUT_2[56959] = 32'b11111111111111101000100100100000;
assign LUT_2[56960] = 32'b11111111111111111110101111111111;
assign LUT_2[56961] = 32'b11111111111111111011101000011000;
assign LUT_2[56962] = 32'b00000000000000000101101000111011;
assign LUT_2[56963] = 32'b00000000000000000010100001010100;
assign LUT_2[56964] = 32'b11111111111111111011001101100111;
assign LUT_2[56965] = 32'b11111111111111111000000110000000;
assign LUT_2[56966] = 32'b00000000000000000010000110100011;
assign LUT_2[56967] = 32'b11111111111111111110111110111100;
assign LUT_2[56968] = 32'b11111111111111111001100001011100;
assign LUT_2[56969] = 32'b11111111111111110110011001110101;
assign LUT_2[56970] = 32'b00000000000000000000011010011000;
assign LUT_2[56971] = 32'b11111111111111111101010010110001;
assign LUT_2[56972] = 32'b11111111111111110101111111000100;
assign LUT_2[56973] = 32'b11111111111111110010110111011101;
assign LUT_2[56974] = 32'b11111111111111111100111000000000;
assign LUT_2[56975] = 32'b11111111111111111001110000011001;
assign LUT_2[56976] = 32'b11111111111111111001010100001001;
assign LUT_2[56977] = 32'b11111111111111110110001100100010;
assign LUT_2[56978] = 32'b00000000000000000000001101000101;
assign LUT_2[56979] = 32'b11111111111111111101000101011110;
assign LUT_2[56980] = 32'b11111111111111110101110001110001;
assign LUT_2[56981] = 32'b11111111111111110010101010001010;
assign LUT_2[56982] = 32'b11111111111111111100101010101101;
assign LUT_2[56983] = 32'b11111111111111111001100011000110;
assign LUT_2[56984] = 32'b11111111111111110100000101100110;
assign LUT_2[56985] = 32'b11111111111111110000111101111111;
assign LUT_2[56986] = 32'b11111111111111111010111110100010;
assign LUT_2[56987] = 32'b11111111111111110111110110111011;
assign LUT_2[56988] = 32'b11111111111111110000100011001110;
assign LUT_2[56989] = 32'b11111111111111101101011011100111;
assign LUT_2[56990] = 32'b11111111111111110111011100001010;
assign LUT_2[56991] = 32'b11111111111111110100010100100011;
assign LUT_2[56992] = 32'b11111111111111111111001011101000;
assign LUT_2[56993] = 32'b11111111111111111100000100000001;
assign LUT_2[56994] = 32'b00000000000000000110000100100100;
assign LUT_2[56995] = 32'b00000000000000000010111100111101;
assign LUT_2[56996] = 32'b11111111111111111011101001010000;
assign LUT_2[56997] = 32'b11111111111111111000100001101001;
assign LUT_2[56998] = 32'b00000000000000000010100010001100;
assign LUT_2[56999] = 32'b11111111111111111111011010100101;
assign LUT_2[57000] = 32'b11111111111111111001111101000101;
assign LUT_2[57001] = 32'b11111111111111110110110101011110;
assign LUT_2[57002] = 32'b00000000000000000000110110000001;
assign LUT_2[57003] = 32'b11111111111111111101101110011010;
assign LUT_2[57004] = 32'b11111111111111110110011010101101;
assign LUT_2[57005] = 32'b11111111111111110011010011000110;
assign LUT_2[57006] = 32'b11111111111111111101010011101001;
assign LUT_2[57007] = 32'b11111111111111111010001100000010;
assign LUT_2[57008] = 32'b11111111111111111001101111110010;
assign LUT_2[57009] = 32'b11111111111111110110101000001011;
assign LUT_2[57010] = 32'b00000000000000000000101000101110;
assign LUT_2[57011] = 32'b11111111111111111101100001000111;
assign LUT_2[57012] = 32'b11111111111111110110001101011010;
assign LUT_2[57013] = 32'b11111111111111110011000101110011;
assign LUT_2[57014] = 32'b11111111111111111101000110010110;
assign LUT_2[57015] = 32'b11111111111111111001111110101111;
assign LUT_2[57016] = 32'b11111111111111110100100001001111;
assign LUT_2[57017] = 32'b11111111111111110001011001101000;
assign LUT_2[57018] = 32'b11111111111111111011011010001011;
assign LUT_2[57019] = 32'b11111111111111111000010010100100;
assign LUT_2[57020] = 32'b11111111111111110000111110110111;
assign LUT_2[57021] = 32'b11111111111111101101110111010000;
assign LUT_2[57022] = 32'b11111111111111110111110111110011;
assign LUT_2[57023] = 32'b11111111111111110100110000001100;
assign LUT_2[57024] = 32'b11111111111111110110111000100010;
assign LUT_2[57025] = 32'b11111111111111110011110000111011;
assign LUT_2[57026] = 32'b11111111111111111101110001011110;
assign LUT_2[57027] = 32'b11111111111111111010101001110111;
assign LUT_2[57028] = 32'b11111111111111110011010110001010;
assign LUT_2[57029] = 32'b11111111111111110000001110100011;
assign LUT_2[57030] = 32'b11111111111111111010001111000110;
assign LUT_2[57031] = 32'b11111111111111110111000111011111;
assign LUT_2[57032] = 32'b11111111111111110001101001111111;
assign LUT_2[57033] = 32'b11111111111111101110100010011000;
assign LUT_2[57034] = 32'b11111111111111111000100010111011;
assign LUT_2[57035] = 32'b11111111111111110101011011010100;
assign LUT_2[57036] = 32'b11111111111111101110000111100111;
assign LUT_2[57037] = 32'b11111111111111101011000000000000;
assign LUT_2[57038] = 32'b11111111111111110101000000100011;
assign LUT_2[57039] = 32'b11111111111111110001111000111100;
assign LUT_2[57040] = 32'b11111111111111110001011100101100;
assign LUT_2[57041] = 32'b11111111111111101110010101000101;
assign LUT_2[57042] = 32'b11111111111111111000010101101000;
assign LUT_2[57043] = 32'b11111111111111110101001110000001;
assign LUT_2[57044] = 32'b11111111111111101101111010010100;
assign LUT_2[57045] = 32'b11111111111111101010110010101101;
assign LUT_2[57046] = 32'b11111111111111110100110011010000;
assign LUT_2[57047] = 32'b11111111111111110001101011101001;
assign LUT_2[57048] = 32'b11111111111111101100001110001001;
assign LUT_2[57049] = 32'b11111111111111101001000110100010;
assign LUT_2[57050] = 32'b11111111111111110011000111000101;
assign LUT_2[57051] = 32'b11111111111111101111111111011110;
assign LUT_2[57052] = 32'b11111111111111101000101011110001;
assign LUT_2[57053] = 32'b11111111111111100101100100001010;
assign LUT_2[57054] = 32'b11111111111111101111100100101101;
assign LUT_2[57055] = 32'b11111111111111101100011101000110;
assign LUT_2[57056] = 32'b11111111111111110111010100001011;
assign LUT_2[57057] = 32'b11111111111111110100001100100100;
assign LUT_2[57058] = 32'b11111111111111111110001101000111;
assign LUT_2[57059] = 32'b11111111111111111011000101100000;
assign LUT_2[57060] = 32'b11111111111111110011110001110011;
assign LUT_2[57061] = 32'b11111111111111110000101010001100;
assign LUT_2[57062] = 32'b11111111111111111010101010101111;
assign LUT_2[57063] = 32'b11111111111111110111100011001000;
assign LUT_2[57064] = 32'b11111111111111110010000101101000;
assign LUT_2[57065] = 32'b11111111111111101110111110000001;
assign LUT_2[57066] = 32'b11111111111111111000111110100100;
assign LUT_2[57067] = 32'b11111111111111110101110110111101;
assign LUT_2[57068] = 32'b11111111111111101110100011010000;
assign LUT_2[57069] = 32'b11111111111111101011011011101001;
assign LUT_2[57070] = 32'b11111111111111110101011100001100;
assign LUT_2[57071] = 32'b11111111111111110010010100100101;
assign LUT_2[57072] = 32'b11111111111111110001111000010101;
assign LUT_2[57073] = 32'b11111111111111101110110000101110;
assign LUT_2[57074] = 32'b11111111111111111000110001010001;
assign LUT_2[57075] = 32'b11111111111111110101101001101010;
assign LUT_2[57076] = 32'b11111111111111101110010101111101;
assign LUT_2[57077] = 32'b11111111111111101011001110010110;
assign LUT_2[57078] = 32'b11111111111111110101001110111001;
assign LUT_2[57079] = 32'b11111111111111110010000111010010;
assign LUT_2[57080] = 32'b11111111111111101100101001110010;
assign LUT_2[57081] = 32'b11111111111111101001100010001011;
assign LUT_2[57082] = 32'b11111111111111110011100010101110;
assign LUT_2[57083] = 32'b11111111111111110000011011000111;
assign LUT_2[57084] = 32'b11111111111111101001000111011010;
assign LUT_2[57085] = 32'b11111111111111100101111111110011;
assign LUT_2[57086] = 32'b11111111111111110000000000010110;
assign LUT_2[57087] = 32'b11111111111111101100111000101111;
assign LUT_2[57088] = 32'b11111111111111111110011010010110;
assign LUT_2[57089] = 32'b11111111111111111011010010101111;
assign LUT_2[57090] = 32'b00000000000000000101010011010010;
assign LUT_2[57091] = 32'b00000000000000000010001011101011;
assign LUT_2[57092] = 32'b11111111111111111010110111111110;
assign LUT_2[57093] = 32'b11111111111111110111110000010111;
assign LUT_2[57094] = 32'b00000000000000000001110000111010;
assign LUT_2[57095] = 32'b11111111111111111110101001010011;
assign LUT_2[57096] = 32'b11111111111111111001001011110011;
assign LUT_2[57097] = 32'b11111111111111110110000100001100;
assign LUT_2[57098] = 32'b00000000000000000000000100101111;
assign LUT_2[57099] = 32'b11111111111111111100111101001000;
assign LUT_2[57100] = 32'b11111111111111110101101001011011;
assign LUT_2[57101] = 32'b11111111111111110010100001110100;
assign LUT_2[57102] = 32'b11111111111111111100100010010111;
assign LUT_2[57103] = 32'b11111111111111111001011010110000;
assign LUT_2[57104] = 32'b11111111111111111000111110100000;
assign LUT_2[57105] = 32'b11111111111111110101110110111001;
assign LUT_2[57106] = 32'b11111111111111111111110111011100;
assign LUT_2[57107] = 32'b11111111111111111100101111110101;
assign LUT_2[57108] = 32'b11111111111111110101011100001000;
assign LUT_2[57109] = 32'b11111111111111110010010100100001;
assign LUT_2[57110] = 32'b11111111111111111100010101000100;
assign LUT_2[57111] = 32'b11111111111111111001001101011101;
assign LUT_2[57112] = 32'b11111111111111110011101111111101;
assign LUT_2[57113] = 32'b11111111111111110000101000010110;
assign LUT_2[57114] = 32'b11111111111111111010101000111001;
assign LUT_2[57115] = 32'b11111111111111110111100001010010;
assign LUT_2[57116] = 32'b11111111111111110000001101100101;
assign LUT_2[57117] = 32'b11111111111111101101000101111110;
assign LUT_2[57118] = 32'b11111111111111110111000110100001;
assign LUT_2[57119] = 32'b11111111111111110011111110111010;
assign LUT_2[57120] = 32'b11111111111111111110110101111111;
assign LUT_2[57121] = 32'b11111111111111111011101110011000;
assign LUT_2[57122] = 32'b00000000000000000101101110111011;
assign LUT_2[57123] = 32'b00000000000000000010100111010100;
assign LUT_2[57124] = 32'b11111111111111111011010011100111;
assign LUT_2[57125] = 32'b11111111111111111000001100000000;
assign LUT_2[57126] = 32'b00000000000000000010001100100011;
assign LUT_2[57127] = 32'b11111111111111111111000100111100;
assign LUT_2[57128] = 32'b11111111111111111001100111011100;
assign LUT_2[57129] = 32'b11111111111111110110011111110101;
assign LUT_2[57130] = 32'b00000000000000000000100000011000;
assign LUT_2[57131] = 32'b11111111111111111101011000110001;
assign LUT_2[57132] = 32'b11111111111111110110000101000100;
assign LUT_2[57133] = 32'b11111111111111110010111101011101;
assign LUT_2[57134] = 32'b11111111111111111100111110000000;
assign LUT_2[57135] = 32'b11111111111111111001110110011001;
assign LUT_2[57136] = 32'b11111111111111111001011010001001;
assign LUT_2[57137] = 32'b11111111111111110110010010100010;
assign LUT_2[57138] = 32'b00000000000000000000010011000101;
assign LUT_2[57139] = 32'b11111111111111111101001011011110;
assign LUT_2[57140] = 32'b11111111111111110101110111110001;
assign LUT_2[57141] = 32'b11111111111111110010110000001010;
assign LUT_2[57142] = 32'b11111111111111111100110000101101;
assign LUT_2[57143] = 32'b11111111111111111001101001000110;
assign LUT_2[57144] = 32'b11111111111111110100001011100110;
assign LUT_2[57145] = 32'b11111111111111110001000011111111;
assign LUT_2[57146] = 32'b11111111111111111011000100100010;
assign LUT_2[57147] = 32'b11111111111111110111111100111011;
assign LUT_2[57148] = 32'b11111111111111110000101001001110;
assign LUT_2[57149] = 32'b11111111111111101101100001100111;
assign LUT_2[57150] = 32'b11111111111111110111100010001010;
assign LUT_2[57151] = 32'b11111111111111110100011010100011;
assign LUT_2[57152] = 32'b11111111111111110110100010111001;
assign LUT_2[57153] = 32'b11111111111111110011011011010010;
assign LUT_2[57154] = 32'b11111111111111111101011011110101;
assign LUT_2[57155] = 32'b11111111111111111010010100001110;
assign LUT_2[57156] = 32'b11111111111111110011000000100001;
assign LUT_2[57157] = 32'b11111111111111101111111000111010;
assign LUT_2[57158] = 32'b11111111111111111001111001011101;
assign LUT_2[57159] = 32'b11111111111111110110110001110110;
assign LUT_2[57160] = 32'b11111111111111110001010100010110;
assign LUT_2[57161] = 32'b11111111111111101110001100101111;
assign LUT_2[57162] = 32'b11111111111111111000001101010010;
assign LUT_2[57163] = 32'b11111111111111110101000101101011;
assign LUT_2[57164] = 32'b11111111111111101101110001111110;
assign LUT_2[57165] = 32'b11111111111111101010101010010111;
assign LUT_2[57166] = 32'b11111111111111110100101010111010;
assign LUT_2[57167] = 32'b11111111111111110001100011010011;
assign LUT_2[57168] = 32'b11111111111111110001000111000011;
assign LUT_2[57169] = 32'b11111111111111101101111111011100;
assign LUT_2[57170] = 32'b11111111111111110111111111111111;
assign LUT_2[57171] = 32'b11111111111111110100111000011000;
assign LUT_2[57172] = 32'b11111111111111101101100100101011;
assign LUT_2[57173] = 32'b11111111111111101010011101000100;
assign LUT_2[57174] = 32'b11111111111111110100011101100111;
assign LUT_2[57175] = 32'b11111111111111110001010110000000;
assign LUT_2[57176] = 32'b11111111111111101011111000100000;
assign LUT_2[57177] = 32'b11111111111111101000110000111001;
assign LUT_2[57178] = 32'b11111111111111110010110001011100;
assign LUT_2[57179] = 32'b11111111111111101111101001110101;
assign LUT_2[57180] = 32'b11111111111111101000010110001000;
assign LUT_2[57181] = 32'b11111111111111100101001110100001;
assign LUT_2[57182] = 32'b11111111111111101111001111000100;
assign LUT_2[57183] = 32'b11111111111111101100000111011101;
assign LUT_2[57184] = 32'b11111111111111110110111110100010;
assign LUT_2[57185] = 32'b11111111111111110011110110111011;
assign LUT_2[57186] = 32'b11111111111111111101110111011110;
assign LUT_2[57187] = 32'b11111111111111111010101111110111;
assign LUT_2[57188] = 32'b11111111111111110011011100001010;
assign LUT_2[57189] = 32'b11111111111111110000010100100011;
assign LUT_2[57190] = 32'b11111111111111111010010101000110;
assign LUT_2[57191] = 32'b11111111111111110111001101011111;
assign LUT_2[57192] = 32'b11111111111111110001101111111111;
assign LUT_2[57193] = 32'b11111111111111101110101000011000;
assign LUT_2[57194] = 32'b11111111111111111000101000111011;
assign LUT_2[57195] = 32'b11111111111111110101100001010100;
assign LUT_2[57196] = 32'b11111111111111101110001101100111;
assign LUT_2[57197] = 32'b11111111111111101011000110000000;
assign LUT_2[57198] = 32'b11111111111111110101000110100011;
assign LUT_2[57199] = 32'b11111111111111110001111110111100;
assign LUT_2[57200] = 32'b11111111111111110001100010101100;
assign LUT_2[57201] = 32'b11111111111111101110011011000101;
assign LUT_2[57202] = 32'b11111111111111111000011011101000;
assign LUT_2[57203] = 32'b11111111111111110101010100000001;
assign LUT_2[57204] = 32'b11111111111111101110000000010100;
assign LUT_2[57205] = 32'b11111111111111101010111000101101;
assign LUT_2[57206] = 32'b11111111111111110100111001010000;
assign LUT_2[57207] = 32'b11111111111111110001110001101001;
assign LUT_2[57208] = 32'b11111111111111101100010100001001;
assign LUT_2[57209] = 32'b11111111111111101001001100100010;
assign LUT_2[57210] = 32'b11111111111111110011001101000101;
assign LUT_2[57211] = 32'b11111111111111110000000101011110;
assign LUT_2[57212] = 32'b11111111111111101000110001110001;
assign LUT_2[57213] = 32'b11111111111111100101101010001010;
assign LUT_2[57214] = 32'b11111111111111101111101010101101;
assign LUT_2[57215] = 32'b11111111111111101100100011000110;
assign LUT_2[57216] = 32'b00000000000000000010101110100101;
assign LUT_2[57217] = 32'b11111111111111111111100110111110;
assign LUT_2[57218] = 32'b00000000000000001001100111100001;
assign LUT_2[57219] = 32'b00000000000000000110011111111010;
assign LUT_2[57220] = 32'b11111111111111111111001100001101;
assign LUT_2[57221] = 32'b11111111111111111100000100100110;
assign LUT_2[57222] = 32'b00000000000000000110000101001001;
assign LUT_2[57223] = 32'b00000000000000000010111101100010;
assign LUT_2[57224] = 32'b11111111111111111101100000000010;
assign LUT_2[57225] = 32'b11111111111111111010011000011011;
assign LUT_2[57226] = 32'b00000000000000000100011000111110;
assign LUT_2[57227] = 32'b00000000000000000001010001010111;
assign LUT_2[57228] = 32'b11111111111111111001111101101010;
assign LUT_2[57229] = 32'b11111111111111110110110110000011;
assign LUT_2[57230] = 32'b00000000000000000000110110100110;
assign LUT_2[57231] = 32'b11111111111111111101101110111111;
assign LUT_2[57232] = 32'b11111111111111111101010010101111;
assign LUT_2[57233] = 32'b11111111111111111010001011001000;
assign LUT_2[57234] = 32'b00000000000000000100001011101011;
assign LUT_2[57235] = 32'b00000000000000000001000100000100;
assign LUT_2[57236] = 32'b11111111111111111001110000010111;
assign LUT_2[57237] = 32'b11111111111111110110101000110000;
assign LUT_2[57238] = 32'b00000000000000000000101001010011;
assign LUT_2[57239] = 32'b11111111111111111101100001101100;
assign LUT_2[57240] = 32'b11111111111111111000000100001100;
assign LUT_2[57241] = 32'b11111111111111110100111100100101;
assign LUT_2[57242] = 32'b11111111111111111110111101001000;
assign LUT_2[57243] = 32'b11111111111111111011110101100001;
assign LUT_2[57244] = 32'b11111111111111110100100001110100;
assign LUT_2[57245] = 32'b11111111111111110001011010001101;
assign LUT_2[57246] = 32'b11111111111111111011011010110000;
assign LUT_2[57247] = 32'b11111111111111111000010011001001;
assign LUT_2[57248] = 32'b00000000000000000011001010001110;
assign LUT_2[57249] = 32'b00000000000000000000000010100111;
assign LUT_2[57250] = 32'b00000000000000001010000011001010;
assign LUT_2[57251] = 32'b00000000000000000110111011100011;
assign LUT_2[57252] = 32'b11111111111111111111100111110110;
assign LUT_2[57253] = 32'b11111111111111111100100000001111;
assign LUT_2[57254] = 32'b00000000000000000110100000110010;
assign LUT_2[57255] = 32'b00000000000000000011011001001011;
assign LUT_2[57256] = 32'b11111111111111111101111011101011;
assign LUT_2[57257] = 32'b11111111111111111010110100000100;
assign LUT_2[57258] = 32'b00000000000000000100110100100111;
assign LUT_2[57259] = 32'b00000000000000000001101101000000;
assign LUT_2[57260] = 32'b11111111111111111010011001010011;
assign LUT_2[57261] = 32'b11111111111111110111010001101100;
assign LUT_2[57262] = 32'b00000000000000000001010010001111;
assign LUT_2[57263] = 32'b11111111111111111110001010101000;
assign LUT_2[57264] = 32'b11111111111111111101101110011000;
assign LUT_2[57265] = 32'b11111111111111111010100110110001;
assign LUT_2[57266] = 32'b00000000000000000100100111010100;
assign LUT_2[57267] = 32'b00000000000000000001011111101101;
assign LUT_2[57268] = 32'b11111111111111111010001100000000;
assign LUT_2[57269] = 32'b11111111111111110111000100011001;
assign LUT_2[57270] = 32'b00000000000000000001000100111100;
assign LUT_2[57271] = 32'b11111111111111111101111101010101;
assign LUT_2[57272] = 32'b11111111111111111000011111110101;
assign LUT_2[57273] = 32'b11111111111111110101011000001110;
assign LUT_2[57274] = 32'b11111111111111111111011000110001;
assign LUT_2[57275] = 32'b11111111111111111100010001001010;
assign LUT_2[57276] = 32'b11111111111111110100111101011101;
assign LUT_2[57277] = 32'b11111111111111110001110101110110;
assign LUT_2[57278] = 32'b11111111111111111011110110011001;
assign LUT_2[57279] = 32'b11111111111111111000101110110010;
assign LUT_2[57280] = 32'b11111111111111111010110111001000;
assign LUT_2[57281] = 32'b11111111111111110111101111100001;
assign LUT_2[57282] = 32'b00000000000000000001110000000100;
assign LUT_2[57283] = 32'b11111111111111111110101000011101;
assign LUT_2[57284] = 32'b11111111111111110111010100110000;
assign LUT_2[57285] = 32'b11111111111111110100001101001001;
assign LUT_2[57286] = 32'b11111111111111111110001101101100;
assign LUT_2[57287] = 32'b11111111111111111011000110000101;
assign LUT_2[57288] = 32'b11111111111111110101101000100101;
assign LUT_2[57289] = 32'b11111111111111110010100000111110;
assign LUT_2[57290] = 32'b11111111111111111100100001100001;
assign LUT_2[57291] = 32'b11111111111111111001011001111010;
assign LUT_2[57292] = 32'b11111111111111110010000110001101;
assign LUT_2[57293] = 32'b11111111111111101110111110100110;
assign LUT_2[57294] = 32'b11111111111111111000111111001001;
assign LUT_2[57295] = 32'b11111111111111110101110111100010;
assign LUT_2[57296] = 32'b11111111111111110101011011010010;
assign LUT_2[57297] = 32'b11111111111111110010010011101011;
assign LUT_2[57298] = 32'b11111111111111111100010100001110;
assign LUT_2[57299] = 32'b11111111111111111001001100100111;
assign LUT_2[57300] = 32'b11111111111111110001111000111010;
assign LUT_2[57301] = 32'b11111111111111101110110001010011;
assign LUT_2[57302] = 32'b11111111111111111000110001110110;
assign LUT_2[57303] = 32'b11111111111111110101101010001111;
assign LUT_2[57304] = 32'b11111111111111110000001100101111;
assign LUT_2[57305] = 32'b11111111111111101101000101001000;
assign LUT_2[57306] = 32'b11111111111111110111000101101011;
assign LUT_2[57307] = 32'b11111111111111110011111110000100;
assign LUT_2[57308] = 32'b11111111111111101100101010010111;
assign LUT_2[57309] = 32'b11111111111111101001100010110000;
assign LUT_2[57310] = 32'b11111111111111110011100011010011;
assign LUT_2[57311] = 32'b11111111111111110000011011101100;
assign LUT_2[57312] = 32'b11111111111111111011010010110001;
assign LUT_2[57313] = 32'b11111111111111111000001011001010;
assign LUT_2[57314] = 32'b00000000000000000010001011101101;
assign LUT_2[57315] = 32'b11111111111111111111000100000110;
assign LUT_2[57316] = 32'b11111111111111110111110000011001;
assign LUT_2[57317] = 32'b11111111111111110100101000110010;
assign LUT_2[57318] = 32'b11111111111111111110101001010101;
assign LUT_2[57319] = 32'b11111111111111111011100001101110;
assign LUT_2[57320] = 32'b11111111111111110110000100001110;
assign LUT_2[57321] = 32'b11111111111111110010111100100111;
assign LUT_2[57322] = 32'b11111111111111111100111101001010;
assign LUT_2[57323] = 32'b11111111111111111001110101100011;
assign LUT_2[57324] = 32'b11111111111111110010100001110110;
assign LUT_2[57325] = 32'b11111111111111101111011010001111;
assign LUT_2[57326] = 32'b11111111111111111001011010110010;
assign LUT_2[57327] = 32'b11111111111111110110010011001011;
assign LUT_2[57328] = 32'b11111111111111110101110110111011;
assign LUT_2[57329] = 32'b11111111111111110010101111010100;
assign LUT_2[57330] = 32'b11111111111111111100101111110111;
assign LUT_2[57331] = 32'b11111111111111111001101000010000;
assign LUT_2[57332] = 32'b11111111111111110010010100100011;
assign LUT_2[57333] = 32'b11111111111111101111001100111100;
assign LUT_2[57334] = 32'b11111111111111111001001101011111;
assign LUT_2[57335] = 32'b11111111111111110110000101111000;
assign LUT_2[57336] = 32'b11111111111111110000101000011000;
assign LUT_2[57337] = 32'b11111111111111101101100000110001;
assign LUT_2[57338] = 32'b11111111111111110111100001010100;
assign LUT_2[57339] = 32'b11111111111111110100011001101101;
assign LUT_2[57340] = 32'b11111111111111101101000110000000;
assign LUT_2[57341] = 32'b11111111111111101001111110011001;
assign LUT_2[57342] = 32'b11111111111111110011111110111100;
assign LUT_2[57343] = 32'b11111111111111110000110111010101;
assign LUT_2[57344] = 32'b11111111111111101101011001110000;
assign LUT_2[57345] = 32'b11111111111111101010010010001001;
assign LUT_2[57346] = 32'b11111111111111110100010010101100;
assign LUT_2[57347] = 32'b11111111111111110001001011000101;
assign LUT_2[57348] = 32'b11111111111111101001110111011000;
assign LUT_2[57349] = 32'b11111111111111100110101111110001;
assign LUT_2[57350] = 32'b11111111111111110000110000010100;
assign LUT_2[57351] = 32'b11111111111111101101101000101101;
assign LUT_2[57352] = 32'b11111111111111101000001011001101;
assign LUT_2[57353] = 32'b11111111111111100101000011100110;
assign LUT_2[57354] = 32'b11111111111111101111000100001001;
assign LUT_2[57355] = 32'b11111111111111101011111100100010;
assign LUT_2[57356] = 32'b11111111111111100100101000110101;
assign LUT_2[57357] = 32'b11111111111111100001100001001110;
assign LUT_2[57358] = 32'b11111111111111101011100001110001;
assign LUT_2[57359] = 32'b11111111111111101000011010001010;
assign LUT_2[57360] = 32'b11111111111111100111111101111010;
assign LUT_2[57361] = 32'b11111111111111100100110110010011;
assign LUT_2[57362] = 32'b11111111111111101110110110110110;
assign LUT_2[57363] = 32'b11111111111111101011101111001111;
assign LUT_2[57364] = 32'b11111111111111100100011011100010;
assign LUT_2[57365] = 32'b11111111111111100001010011111011;
assign LUT_2[57366] = 32'b11111111111111101011010100011110;
assign LUT_2[57367] = 32'b11111111111111101000001100110111;
assign LUT_2[57368] = 32'b11111111111111100010101111010111;
assign LUT_2[57369] = 32'b11111111111111011111100111110000;
assign LUT_2[57370] = 32'b11111111111111101001101000010011;
assign LUT_2[57371] = 32'b11111111111111100110100000101100;
assign LUT_2[57372] = 32'b11111111111111011111001100111111;
assign LUT_2[57373] = 32'b11111111111111011100000101011000;
assign LUT_2[57374] = 32'b11111111111111100110000101111011;
assign LUT_2[57375] = 32'b11111111111111100010111110010100;
assign LUT_2[57376] = 32'b11111111111111101101110101011001;
assign LUT_2[57377] = 32'b11111111111111101010101101110010;
assign LUT_2[57378] = 32'b11111111111111110100101110010101;
assign LUT_2[57379] = 32'b11111111111111110001100110101110;
assign LUT_2[57380] = 32'b11111111111111101010010011000001;
assign LUT_2[57381] = 32'b11111111111111100111001011011010;
assign LUT_2[57382] = 32'b11111111111111110001001011111101;
assign LUT_2[57383] = 32'b11111111111111101110000100010110;
assign LUT_2[57384] = 32'b11111111111111101000100110110110;
assign LUT_2[57385] = 32'b11111111111111100101011111001111;
assign LUT_2[57386] = 32'b11111111111111101111011111110010;
assign LUT_2[57387] = 32'b11111111111111101100011000001011;
assign LUT_2[57388] = 32'b11111111111111100101000100011110;
assign LUT_2[57389] = 32'b11111111111111100001111100110111;
assign LUT_2[57390] = 32'b11111111111111101011111101011010;
assign LUT_2[57391] = 32'b11111111111111101000110101110011;
assign LUT_2[57392] = 32'b11111111111111101000011001100011;
assign LUT_2[57393] = 32'b11111111111111100101010001111100;
assign LUT_2[57394] = 32'b11111111111111101111010010011111;
assign LUT_2[57395] = 32'b11111111111111101100001010111000;
assign LUT_2[57396] = 32'b11111111111111100100110111001011;
assign LUT_2[57397] = 32'b11111111111111100001101111100100;
assign LUT_2[57398] = 32'b11111111111111101011110000000111;
assign LUT_2[57399] = 32'b11111111111111101000101000100000;
assign LUT_2[57400] = 32'b11111111111111100011001011000000;
assign LUT_2[57401] = 32'b11111111111111100000000011011001;
assign LUT_2[57402] = 32'b11111111111111101010000011111100;
assign LUT_2[57403] = 32'b11111111111111100110111100010101;
assign LUT_2[57404] = 32'b11111111111111011111101000101000;
assign LUT_2[57405] = 32'b11111111111111011100100001000001;
assign LUT_2[57406] = 32'b11111111111111100110100001100100;
assign LUT_2[57407] = 32'b11111111111111100011011001111101;
assign LUT_2[57408] = 32'b11111111111111100101100010010011;
assign LUT_2[57409] = 32'b11111111111111100010011010101100;
assign LUT_2[57410] = 32'b11111111111111101100011011001111;
assign LUT_2[57411] = 32'b11111111111111101001010011101000;
assign LUT_2[57412] = 32'b11111111111111100001111111111011;
assign LUT_2[57413] = 32'b11111111111111011110111000010100;
assign LUT_2[57414] = 32'b11111111111111101000111000110111;
assign LUT_2[57415] = 32'b11111111111111100101110001010000;
assign LUT_2[57416] = 32'b11111111111111100000010011110000;
assign LUT_2[57417] = 32'b11111111111111011101001100001001;
assign LUT_2[57418] = 32'b11111111111111100111001100101100;
assign LUT_2[57419] = 32'b11111111111111100100000101000101;
assign LUT_2[57420] = 32'b11111111111111011100110001011000;
assign LUT_2[57421] = 32'b11111111111111011001101001110001;
assign LUT_2[57422] = 32'b11111111111111100011101010010100;
assign LUT_2[57423] = 32'b11111111111111100000100010101101;
assign LUT_2[57424] = 32'b11111111111111100000000110011101;
assign LUT_2[57425] = 32'b11111111111111011100111110110110;
assign LUT_2[57426] = 32'b11111111111111100110111111011001;
assign LUT_2[57427] = 32'b11111111111111100011110111110010;
assign LUT_2[57428] = 32'b11111111111111011100100100000101;
assign LUT_2[57429] = 32'b11111111111111011001011100011110;
assign LUT_2[57430] = 32'b11111111111111100011011101000001;
assign LUT_2[57431] = 32'b11111111111111100000010101011010;
assign LUT_2[57432] = 32'b11111111111111011010110111111010;
assign LUT_2[57433] = 32'b11111111111111010111110000010011;
assign LUT_2[57434] = 32'b11111111111111100001110000110110;
assign LUT_2[57435] = 32'b11111111111111011110101001001111;
assign LUT_2[57436] = 32'b11111111111111010111010101100010;
assign LUT_2[57437] = 32'b11111111111111010100001101111011;
assign LUT_2[57438] = 32'b11111111111111011110001110011110;
assign LUT_2[57439] = 32'b11111111111111011011000110110111;
assign LUT_2[57440] = 32'b11111111111111100101111101111100;
assign LUT_2[57441] = 32'b11111111111111100010110110010101;
assign LUT_2[57442] = 32'b11111111111111101100110110111000;
assign LUT_2[57443] = 32'b11111111111111101001101111010001;
assign LUT_2[57444] = 32'b11111111111111100010011011100100;
assign LUT_2[57445] = 32'b11111111111111011111010011111101;
assign LUT_2[57446] = 32'b11111111111111101001010100100000;
assign LUT_2[57447] = 32'b11111111111111100110001100111001;
assign LUT_2[57448] = 32'b11111111111111100000101111011001;
assign LUT_2[57449] = 32'b11111111111111011101100111110010;
assign LUT_2[57450] = 32'b11111111111111100111101000010101;
assign LUT_2[57451] = 32'b11111111111111100100100000101110;
assign LUT_2[57452] = 32'b11111111111111011101001101000001;
assign LUT_2[57453] = 32'b11111111111111011010000101011010;
assign LUT_2[57454] = 32'b11111111111111100100000101111101;
assign LUT_2[57455] = 32'b11111111111111100000111110010110;
assign LUT_2[57456] = 32'b11111111111111100000100010000110;
assign LUT_2[57457] = 32'b11111111111111011101011010011111;
assign LUT_2[57458] = 32'b11111111111111100111011011000010;
assign LUT_2[57459] = 32'b11111111111111100100010011011011;
assign LUT_2[57460] = 32'b11111111111111011100111111101110;
assign LUT_2[57461] = 32'b11111111111111011001111000000111;
assign LUT_2[57462] = 32'b11111111111111100011111000101010;
assign LUT_2[57463] = 32'b11111111111111100000110001000011;
assign LUT_2[57464] = 32'b11111111111111011011010011100011;
assign LUT_2[57465] = 32'b11111111111111011000001011111100;
assign LUT_2[57466] = 32'b11111111111111100010001100011111;
assign LUT_2[57467] = 32'b11111111111111011111000100111000;
assign LUT_2[57468] = 32'b11111111111111010111110001001011;
assign LUT_2[57469] = 32'b11111111111111010100101001100100;
assign LUT_2[57470] = 32'b11111111111111011110101010000111;
assign LUT_2[57471] = 32'b11111111111111011011100010100000;
assign LUT_2[57472] = 32'b11111111111111110001101101111111;
assign LUT_2[57473] = 32'b11111111111111101110100110011000;
assign LUT_2[57474] = 32'b11111111111111111000100110111011;
assign LUT_2[57475] = 32'b11111111111111110101011111010100;
assign LUT_2[57476] = 32'b11111111111111101110001011100111;
assign LUT_2[57477] = 32'b11111111111111101011000100000000;
assign LUT_2[57478] = 32'b11111111111111110101000100100011;
assign LUT_2[57479] = 32'b11111111111111110001111100111100;
assign LUT_2[57480] = 32'b11111111111111101100011111011100;
assign LUT_2[57481] = 32'b11111111111111101001010111110101;
assign LUT_2[57482] = 32'b11111111111111110011011000011000;
assign LUT_2[57483] = 32'b11111111111111110000010000110001;
assign LUT_2[57484] = 32'b11111111111111101000111101000100;
assign LUT_2[57485] = 32'b11111111111111100101110101011101;
assign LUT_2[57486] = 32'b11111111111111101111110110000000;
assign LUT_2[57487] = 32'b11111111111111101100101110011001;
assign LUT_2[57488] = 32'b11111111111111101100010010001001;
assign LUT_2[57489] = 32'b11111111111111101001001010100010;
assign LUT_2[57490] = 32'b11111111111111110011001011000101;
assign LUT_2[57491] = 32'b11111111111111110000000011011110;
assign LUT_2[57492] = 32'b11111111111111101000101111110001;
assign LUT_2[57493] = 32'b11111111111111100101101000001010;
assign LUT_2[57494] = 32'b11111111111111101111101000101101;
assign LUT_2[57495] = 32'b11111111111111101100100001000110;
assign LUT_2[57496] = 32'b11111111111111100111000011100110;
assign LUT_2[57497] = 32'b11111111111111100011111011111111;
assign LUT_2[57498] = 32'b11111111111111101101111100100010;
assign LUT_2[57499] = 32'b11111111111111101010110100111011;
assign LUT_2[57500] = 32'b11111111111111100011100001001110;
assign LUT_2[57501] = 32'b11111111111111100000011001100111;
assign LUT_2[57502] = 32'b11111111111111101010011010001010;
assign LUT_2[57503] = 32'b11111111111111100111010010100011;
assign LUT_2[57504] = 32'b11111111111111110010001001101000;
assign LUT_2[57505] = 32'b11111111111111101111000010000001;
assign LUT_2[57506] = 32'b11111111111111111001000010100100;
assign LUT_2[57507] = 32'b11111111111111110101111010111101;
assign LUT_2[57508] = 32'b11111111111111101110100111010000;
assign LUT_2[57509] = 32'b11111111111111101011011111101001;
assign LUT_2[57510] = 32'b11111111111111110101100000001100;
assign LUT_2[57511] = 32'b11111111111111110010011000100101;
assign LUT_2[57512] = 32'b11111111111111101100111011000101;
assign LUT_2[57513] = 32'b11111111111111101001110011011110;
assign LUT_2[57514] = 32'b11111111111111110011110100000001;
assign LUT_2[57515] = 32'b11111111111111110000101100011010;
assign LUT_2[57516] = 32'b11111111111111101001011000101101;
assign LUT_2[57517] = 32'b11111111111111100110010001000110;
assign LUT_2[57518] = 32'b11111111111111110000010001101001;
assign LUT_2[57519] = 32'b11111111111111101101001010000010;
assign LUT_2[57520] = 32'b11111111111111101100101101110010;
assign LUT_2[57521] = 32'b11111111111111101001100110001011;
assign LUT_2[57522] = 32'b11111111111111110011100110101110;
assign LUT_2[57523] = 32'b11111111111111110000011111000111;
assign LUT_2[57524] = 32'b11111111111111101001001011011010;
assign LUT_2[57525] = 32'b11111111111111100110000011110011;
assign LUT_2[57526] = 32'b11111111111111110000000100010110;
assign LUT_2[57527] = 32'b11111111111111101100111100101111;
assign LUT_2[57528] = 32'b11111111111111100111011111001111;
assign LUT_2[57529] = 32'b11111111111111100100010111101000;
assign LUT_2[57530] = 32'b11111111111111101110011000001011;
assign LUT_2[57531] = 32'b11111111111111101011010000100100;
assign LUT_2[57532] = 32'b11111111111111100011111100110111;
assign LUT_2[57533] = 32'b11111111111111100000110101010000;
assign LUT_2[57534] = 32'b11111111111111101010110101110011;
assign LUT_2[57535] = 32'b11111111111111100111101110001100;
assign LUT_2[57536] = 32'b11111111111111101001110110100010;
assign LUT_2[57537] = 32'b11111111111111100110101110111011;
assign LUT_2[57538] = 32'b11111111111111110000101111011110;
assign LUT_2[57539] = 32'b11111111111111101101100111110111;
assign LUT_2[57540] = 32'b11111111111111100110010100001010;
assign LUT_2[57541] = 32'b11111111111111100011001100100011;
assign LUT_2[57542] = 32'b11111111111111101101001101000110;
assign LUT_2[57543] = 32'b11111111111111101010000101011111;
assign LUT_2[57544] = 32'b11111111111111100100100111111111;
assign LUT_2[57545] = 32'b11111111111111100001100000011000;
assign LUT_2[57546] = 32'b11111111111111101011100000111011;
assign LUT_2[57547] = 32'b11111111111111101000011001010100;
assign LUT_2[57548] = 32'b11111111111111100001000101100111;
assign LUT_2[57549] = 32'b11111111111111011101111110000000;
assign LUT_2[57550] = 32'b11111111111111100111111110100011;
assign LUT_2[57551] = 32'b11111111111111100100110110111100;
assign LUT_2[57552] = 32'b11111111111111100100011010101100;
assign LUT_2[57553] = 32'b11111111111111100001010011000101;
assign LUT_2[57554] = 32'b11111111111111101011010011101000;
assign LUT_2[57555] = 32'b11111111111111101000001100000001;
assign LUT_2[57556] = 32'b11111111111111100000111000010100;
assign LUT_2[57557] = 32'b11111111111111011101110000101101;
assign LUT_2[57558] = 32'b11111111111111100111110001010000;
assign LUT_2[57559] = 32'b11111111111111100100101001101001;
assign LUT_2[57560] = 32'b11111111111111011111001100001001;
assign LUT_2[57561] = 32'b11111111111111011100000100100010;
assign LUT_2[57562] = 32'b11111111111111100110000101000101;
assign LUT_2[57563] = 32'b11111111111111100010111101011110;
assign LUT_2[57564] = 32'b11111111111111011011101001110001;
assign LUT_2[57565] = 32'b11111111111111011000100010001010;
assign LUT_2[57566] = 32'b11111111111111100010100010101101;
assign LUT_2[57567] = 32'b11111111111111011111011011000110;
assign LUT_2[57568] = 32'b11111111111111101010010010001011;
assign LUT_2[57569] = 32'b11111111111111100111001010100100;
assign LUT_2[57570] = 32'b11111111111111110001001011000111;
assign LUT_2[57571] = 32'b11111111111111101110000011100000;
assign LUT_2[57572] = 32'b11111111111111100110101111110011;
assign LUT_2[57573] = 32'b11111111111111100011101000001100;
assign LUT_2[57574] = 32'b11111111111111101101101000101111;
assign LUT_2[57575] = 32'b11111111111111101010100001001000;
assign LUT_2[57576] = 32'b11111111111111100101000011101000;
assign LUT_2[57577] = 32'b11111111111111100001111100000001;
assign LUT_2[57578] = 32'b11111111111111101011111100100100;
assign LUT_2[57579] = 32'b11111111111111101000110100111101;
assign LUT_2[57580] = 32'b11111111111111100001100001010000;
assign LUT_2[57581] = 32'b11111111111111011110011001101001;
assign LUT_2[57582] = 32'b11111111111111101000011010001100;
assign LUT_2[57583] = 32'b11111111111111100101010010100101;
assign LUT_2[57584] = 32'b11111111111111100100110110010101;
assign LUT_2[57585] = 32'b11111111111111100001101110101110;
assign LUT_2[57586] = 32'b11111111111111101011101111010001;
assign LUT_2[57587] = 32'b11111111111111101000100111101010;
assign LUT_2[57588] = 32'b11111111111111100001010011111101;
assign LUT_2[57589] = 32'b11111111111111011110001100010110;
assign LUT_2[57590] = 32'b11111111111111101000001100111001;
assign LUT_2[57591] = 32'b11111111111111100101000101010010;
assign LUT_2[57592] = 32'b11111111111111011111100111110010;
assign LUT_2[57593] = 32'b11111111111111011100100000001011;
assign LUT_2[57594] = 32'b11111111111111100110100000101110;
assign LUT_2[57595] = 32'b11111111111111100011011001000111;
assign LUT_2[57596] = 32'b11111111111111011100000101011010;
assign LUT_2[57597] = 32'b11111111111111011000111101110011;
assign LUT_2[57598] = 32'b11111111111111100010111110010110;
assign LUT_2[57599] = 32'b11111111111111011111110110101111;
assign LUT_2[57600] = 32'b11111111111111110001011000010110;
assign LUT_2[57601] = 32'b11111111111111101110010000101111;
assign LUT_2[57602] = 32'b11111111111111111000010001010010;
assign LUT_2[57603] = 32'b11111111111111110101001001101011;
assign LUT_2[57604] = 32'b11111111111111101101110101111110;
assign LUT_2[57605] = 32'b11111111111111101010101110010111;
assign LUT_2[57606] = 32'b11111111111111110100101110111010;
assign LUT_2[57607] = 32'b11111111111111110001100111010011;
assign LUT_2[57608] = 32'b11111111111111101100001001110011;
assign LUT_2[57609] = 32'b11111111111111101001000010001100;
assign LUT_2[57610] = 32'b11111111111111110011000010101111;
assign LUT_2[57611] = 32'b11111111111111101111111011001000;
assign LUT_2[57612] = 32'b11111111111111101000100111011011;
assign LUT_2[57613] = 32'b11111111111111100101011111110100;
assign LUT_2[57614] = 32'b11111111111111101111100000010111;
assign LUT_2[57615] = 32'b11111111111111101100011000110000;
assign LUT_2[57616] = 32'b11111111111111101011111100100000;
assign LUT_2[57617] = 32'b11111111111111101000110100111001;
assign LUT_2[57618] = 32'b11111111111111110010110101011100;
assign LUT_2[57619] = 32'b11111111111111101111101101110101;
assign LUT_2[57620] = 32'b11111111111111101000011010001000;
assign LUT_2[57621] = 32'b11111111111111100101010010100001;
assign LUT_2[57622] = 32'b11111111111111101111010011000100;
assign LUT_2[57623] = 32'b11111111111111101100001011011101;
assign LUT_2[57624] = 32'b11111111111111100110101101111101;
assign LUT_2[57625] = 32'b11111111111111100011100110010110;
assign LUT_2[57626] = 32'b11111111111111101101100110111001;
assign LUT_2[57627] = 32'b11111111111111101010011111010010;
assign LUT_2[57628] = 32'b11111111111111100011001011100101;
assign LUT_2[57629] = 32'b11111111111111100000000011111110;
assign LUT_2[57630] = 32'b11111111111111101010000100100001;
assign LUT_2[57631] = 32'b11111111111111100110111100111010;
assign LUT_2[57632] = 32'b11111111111111110001110011111111;
assign LUT_2[57633] = 32'b11111111111111101110101100011000;
assign LUT_2[57634] = 32'b11111111111111111000101100111011;
assign LUT_2[57635] = 32'b11111111111111110101100101010100;
assign LUT_2[57636] = 32'b11111111111111101110010001100111;
assign LUT_2[57637] = 32'b11111111111111101011001010000000;
assign LUT_2[57638] = 32'b11111111111111110101001010100011;
assign LUT_2[57639] = 32'b11111111111111110010000010111100;
assign LUT_2[57640] = 32'b11111111111111101100100101011100;
assign LUT_2[57641] = 32'b11111111111111101001011101110101;
assign LUT_2[57642] = 32'b11111111111111110011011110011000;
assign LUT_2[57643] = 32'b11111111111111110000010110110001;
assign LUT_2[57644] = 32'b11111111111111101001000011000100;
assign LUT_2[57645] = 32'b11111111111111100101111011011101;
assign LUT_2[57646] = 32'b11111111111111101111111100000000;
assign LUT_2[57647] = 32'b11111111111111101100110100011001;
assign LUT_2[57648] = 32'b11111111111111101100011000001001;
assign LUT_2[57649] = 32'b11111111111111101001010000100010;
assign LUT_2[57650] = 32'b11111111111111110011010001000101;
assign LUT_2[57651] = 32'b11111111111111110000001001011110;
assign LUT_2[57652] = 32'b11111111111111101000110101110001;
assign LUT_2[57653] = 32'b11111111111111100101101110001010;
assign LUT_2[57654] = 32'b11111111111111101111101110101101;
assign LUT_2[57655] = 32'b11111111111111101100100111000110;
assign LUT_2[57656] = 32'b11111111111111100111001001100110;
assign LUT_2[57657] = 32'b11111111111111100100000001111111;
assign LUT_2[57658] = 32'b11111111111111101110000010100010;
assign LUT_2[57659] = 32'b11111111111111101010111010111011;
assign LUT_2[57660] = 32'b11111111111111100011100111001110;
assign LUT_2[57661] = 32'b11111111111111100000011111100111;
assign LUT_2[57662] = 32'b11111111111111101010100000001010;
assign LUT_2[57663] = 32'b11111111111111100111011000100011;
assign LUT_2[57664] = 32'b11111111111111101001100000111001;
assign LUT_2[57665] = 32'b11111111111111100110011001010010;
assign LUT_2[57666] = 32'b11111111111111110000011001110101;
assign LUT_2[57667] = 32'b11111111111111101101010010001110;
assign LUT_2[57668] = 32'b11111111111111100101111110100001;
assign LUT_2[57669] = 32'b11111111111111100010110110111010;
assign LUT_2[57670] = 32'b11111111111111101100110111011101;
assign LUT_2[57671] = 32'b11111111111111101001101111110110;
assign LUT_2[57672] = 32'b11111111111111100100010010010110;
assign LUT_2[57673] = 32'b11111111111111100001001010101111;
assign LUT_2[57674] = 32'b11111111111111101011001011010010;
assign LUT_2[57675] = 32'b11111111111111101000000011101011;
assign LUT_2[57676] = 32'b11111111111111100000101111111110;
assign LUT_2[57677] = 32'b11111111111111011101101000010111;
assign LUT_2[57678] = 32'b11111111111111100111101000111010;
assign LUT_2[57679] = 32'b11111111111111100100100001010011;
assign LUT_2[57680] = 32'b11111111111111100100000101000011;
assign LUT_2[57681] = 32'b11111111111111100000111101011100;
assign LUT_2[57682] = 32'b11111111111111101010111101111111;
assign LUT_2[57683] = 32'b11111111111111100111110110011000;
assign LUT_2[57684] = 32'b11111111111111100000100010101011;
assign LUT_2[57685] = 32'b11111111111111011101011011000100;
assign LUT_2[57686] = 32'b11111111111111100111011011100111;
assign LUT_2[57687] = 32'b11111111111111100100010100000000;
assign LUT_2[57688] = 32'b11111111111111011110110110100000;
assign LUT_2[57689] = 32'b11111111111111011011101110111001;
assign LUT_2[57690] = 32'b11111111111111100101101111011100;
assign LUT_2[57691] = 32'b11111111111111100010100111110101;
assign LUT_2[57692] = 32'b11111111111111011011010100001000;
assign LUT_2[57693] = 32'b11111111111111011000001100100001;
assign LUT_2[57694] = 32'b11111111111111100010001101000100;
assign LUT_2[57695] = 32'b11111111111111011111000101011101;
assign LUT_2[57696] = 32'b11111111111111101001111100100010;
assign LUT_2[57697] = 32'b11111111111111100110110100111011;
assign LUT_2[57698] = 32'b11111111111111110000110101011110;
assign LUT_2[57699] = 32'b11111111111111101101101101110111;
assign LUT_2[57700] = 32'b11111111111111100110011010001010;
assign LUT_2[57701] = 32'b11111111111111100011010010100011;
assign LUT_2[57702] = 32'b11111111111111101101010011000110;
assign LUT_2[57703] = 32'b11111111111111101010001011011111;
assign LUT_2[57704] = 32'b11111111111111100100101101111111;
assign LUT_2[57705] = 32'b11111111111111100001100110011000;
assign LUT_2[57706] = 32'b11111111111111101011100110111011;
assign LUT_2[57707] = 32'b11111111111111101000011111010100;
assign LUT_2[57708] = 32'b11111111111111100001001011100111;
assign LUT_2[57709] = 32'b11111111111111011110000100000000;
assign LUT_2[57710] = 32'b11111111111111101000000100100011;
assign LUT_2[57711] = 32'b11111111111111100100111100111100;
assign LUT_2[57712] = 32'b11111111111111100100100000101100;
assign LUT_2[57713] = 32'b11111111111111100001011001000101;
assign LUT_2[57714] = 32'b11111111111111101011011001101000;
assign LUT_2[57715] = 32'b11111111111111101000010010000001;
assign LUT_2[57716] = 32'b11111111111111100000111110010100;
assign LUT_2[57717] = 32'b11111111111111011101110110101101;
assign LUT_2[57718] = 32'b11111111111111100111110111010000;
assign LUT_2[57719] = 32'b11111111111111100100101111101001;
assign LUT_2[57720] = 32'b11111111111111011111010010001001;
assign LUT_2[57721] = 32'b11111111111111011100001010100010;
assign LUT_2[57722] = 32'b11111111111111100110001011000101;
assign LUT_2[57723] = 32'b11111111111111100011000011011110;
assign LUT_2[57724] = 32'b11111111111111011011101111110001;
assign LUT_2[57725] = 32'b11111111111111011000101000001010;
assign LUT_2[57726] = 32'b11111111111111100010101000101101;
assign LUT_2[57727] = 32'b11111111111111011111100001000110;
assign LUT_2[57728] = 32'b11111111111111110101101100100101;
assign LUT_2[57729] = 32'b11111111111111110010100100111110;
assign LUT_2[57730] = 32'b11111111111111111100100101100001;
assign LUT_2[57731] = 32'b11111111111111111001011101111010;
assign LUT_2[57732] = 32'b11111111111111110010001010001101;
assign LUT_2[57733] = 32'b11111111111111101111000010100110;
assign LUT_2[57734] = 32'b11111111111111111001000011001001;
assign LUT_2[57735] = 32'b11111111111111110101111011100010;
assign LUT_2[57736] = 32'b11111111111111110000011110000010;
assign LUT_2[57737] = 32'b11111111111111101101010110011011;
assign LUT_2[57738] = 32'b11111111111111110111010110111110;
assign LUT_2[57739] = 32'b11111111111111110100001111010111;
assign LUT_2[57740] = 32'b11111111111111101100111011101010;
assign LUT_2[57741] = 32'b11111111111111101001110100000011;
assign LUT_2[57742] = 32'b11111111111111110011110100100110;
assign LUT_2[57743] = 32'b11111111111111110000101100111111;
assign LUT_2[57744] = 32'b11111111111111110000010000101111;
assign LUT_2[57745] = 32'b11111111111111101101001001001000;
assign LUT_2[57746] = 32'b11111111111111110111001001101011;
assign LUT_2[57747] = 32'b11111111111111110100000010000100;
assign LUT_2[57748] = 32'b11111111111111101100101110010111;
assign LUT_2[57749] = 32'b11111111111111101001100110110000;
assign LUT_2[57750] = 32'b11111111111111110011100111010011;
assign LUT_2[57751] = 32'b11111111111111110000011111101100;
assign LUT_2[57752] = 32'b11111111111111101011000010001100;
assign LUT_2[57753] = 32'b11111111111111100111111010100101;
assign LUT_2[57754] = 32'b11111111111111110001111011001000;
assign LUT_2[57755] = 32'b11111111111111101110110011100001;
assign LUT_2[57756] = 32'b11111111111111100111011111110100;
assign LUT_2[57757] = 32'b11111111111111100100011000001101;
assign LUT_2[57758] = 32'b11111111111111101110011000110000;
assign LUT_2[57759] = 32'b11111111111111101011010001001001;
assign LUT_2[57760] = 32'b11111111111111110110001000001110;
assign LUT_2[57761] = 32'b11111111111111110011000000100111;
assign LUT_2[57762] = 32'b11111111111111111101000001001010;
assign LUT_2[57763] = 32'b11111111111111111001111001100011;
assign LUT_2[57764] = 32'b11111111111111110010100101110110;
assign LUT_2[57765] = 32'b11111111111111101111011110001111;
assign LUT_2[57766] = 32'b11111111111111111001011110110010;
assign LUT_2[57767] = 32'b11111111111111110110010111001011;
assign LUT_2[57768] = 32'b11111111111111110000111001101011;
assign LUT_2[57769] = 32'b11111111111111101101110010000100;
assign LUT_2[57770] = 32'b11111111111111110111110010100111;
assign LUT_2[57771] = 32'b11111111111111110100101011000000;
assign LUT_2[57772] = 32'b11111111111111101101010111010011;
assign LUT_2[57773] = 32'b11111111111111101010001111101100;
assign LUT_2[57774] = 32'b11111111111111110100010000001111;
assign LUT_2[57775] = 32'b11111111111111110001001000101000;
assign LUT_2[57776] = 32'b11111111111111110000101100011000;
assign LUT_2[57777] = 32'b11111111111111101101100100110001;
assign LUT_2[57778] = 32'b11111111111111110111100101010100;
assign LUT_2[57779] = 32'b11111111111111110100011101101101;
assign LUT_2[57780] = 32'b11111111111111101101001010000000;
assign LUT_2[57781] = 32'b11111111111111101010000010011001;
assign LUT_2[57782] = 32'b11111111111111110100000010111100;
assign LUT_2[57783] = 32'b11111111111111110000111011010101;
assign LUT_2[57784] = 32'b11111111111111101011011101110101;
assign LUT_2[57785] = 32'b11111111111111101000010110001110;
assign LUT_2[57786] = 32'b11111111111111110010010110110001;
assign LUT_2[57787] = 32'b11111111111111101111001111001010;
assign LUT_2[57788] = 32'b11111111111111100111111011011101;
assign LUT_2[57789] = 32'b11111111111111100100110011110110;
assign LUT_2[57790] = 32'b11111111111111101110110100011001;
assign LUT_2[57791] = 32'b11111111111111101011101100110010;
assign LUT_2[57792] = 32'b11111111111111101101110101001000;
assign LUT_2[57793] = 32'b11111111111111101010101101100001;
assign LUT_2[57794] = 32'b11111111111111110100101110000100;
assign LUT_2[57795] = 32'b11111111111111110001100110011101;
assign LUT_2[57796] = 32'b11111111111111101010010010110000;
assign LUT_2[57797] = 32'b11111111111111100111001011001001;
assign LUT_2[57798] = 32'b11111111111111110001001011101100;
assign LUT_2[57799] = 32'b11111111111111101110000100000101;
assign LUT_2[57800] = 32'b11111111111111101000100110100101;
assign LUT_2[57801] = 32'b11111111111111100101011110111110;
assign LUT_2[57802] = 32'b11111111111111101111011111100001;
assign LUT_2[57803] = 32'b11111111111111101100010111111010;
assign LUT_2[57804] = 32'b11111111111111100101000100001101;
assign LUT_2[57805] = 32'b11111111111111100001111100100110;
assign LUT_2[57806] = 32'b11111111111111101011111101001001;
assign LUT_2[57807] = 32'b11111111111111101000110101100010;
assign LUT_2[57808] = 32'b11111111111111101000011001010010;
assign LUT_2[57809] = 32'b11111111111111100101010001101011;
assign LUT_2[57810] = 32'b11111111111111101111010010001110;
assign LUT_2[57811] = 32'b11111111111111101100001010100111;
assign LUT_2[57812] = 32'b11111111111111100100110110111010;
assign LUT_2[57813] = 32'b11111111111111100001101111010011;
assign LUT_2[57814] = 32'b11111111111111101011101111110110;
assign LUT_2[57815] = 32'b11111111111111101000101000001111;
assign LUT_2[57816] = 32'b11111111111111100011001010101111;
assign LUT_2[57817] = 32'b11111111111111100000000011001000;
assign LUT_2[57818] = 32'b11111111111111101010000011101011;
assign LUT_2[57819] = 32'b11111111111111100110111100000100;
assign LUT_2[57820] = 32'b11111111111111011111101000010111;
assign LUT_2[57821] = 32'b11111111111111011100100000110000;
assign LUT_2[57822] = 32'b11111111111111100110100001010011;
assign LUT_2[57823] = 32'b11111111111111100011011001101100;
assign LUT_2[57824] = 32'b11111111111111101110010000110001;
assign LUT_2[57825] = 32'b11111111111111101011001001001010;
assign LUT_2[57826] = 32'b11111111111111110101001001101101;
assign LUT_2[57827] = 32'b11111111111111110010000010000110;
assign LUT_2[57828] = 32'b11111111111111101010101110011001;
assign LUT_2[57829] = 32'b11111111111111100111100110110010;
assign LUT_2[57830] = 32'b11111111111111110001100111010101;
assign LUT_2[57831] = 32'b11111111111111101110011111101110;
assign LUT_2[57832] = 32'b11111111111111101001000010001110;
assign LUT_2[57833] = 32'b11111111111111100101111010100111;
assign LUT_2[57834] = 32'b11111111111111101111111011001010;
assign LUT_2[57835] = 32'b11111111111111101100110011100011;
assign LUT_2[57836] = 32'b11111111111111100101011111110110;
assign LUT_2[57837] = 32'b11111111111111100010011000001111;
assign LUT_2[57838] = 32'b11111111111111101100011000110010;
assign LUT_2[57839] = 32'b11111111111111101001010001001011;
assign LUT_2[57840] = 32'b11111111111111101000110100111011;
assign LUT_2[57841] = 32'b11111111111111100101101101010100;
assign LUT_2[57842] = 32'b11111111111111101111101101110111;
assign LUT_2[57843] = 32'b11111111111111101100100110010000;
assign LUT_2[57844] = 32'b11111111111111100101010010100011;
assign LUT_2[57845] = 32'b11111111111111100010001010111100;
assign LUT_2[57846] = 32'b11111111111111101100001011011111;
assign LUT_2[57847] = 32'b11111111111111101001000011111000;
assign LUT_2[57848] = 32'b11111111111111100011100110011000;
assign LUT_2[57849] = 32'b11111111111111100000011110110001;
assign LUT_2[57850] = 32'b11111111111111101010011111010100;
assign LUT_2[57851] = 32'b11111111111111100111010111101101;
assign LUT_2[57852] = 32'b11111111111111100000000100000000;
assign LUT_2[57853] = 32'b11111111111111011100111100011001;
assign LUT_2[57854] = 32'b11111111111111100110111100111100;
assign LUT_2[57855] = 32'b11111111111111100011110101010101;
assign LUT_2[57856] = 32'b11111111111111110010001011100010;
assign LUT_2[57857] = 32'b11111111111111101111000011111011;
assign LUT_2[57858] = 32'b11111111111111111001000100011110;
assign LUT_2[57859] = 32'b11111111111111110101111100110111;
assign LUT_2[57860] = 32'b11111111111111101110101001001010;
assign LUT_2[57861] = 32'b11111111111111101011100001100011;
assign LUT_2[57862] = 32'b11111111111111110101100010000110;
assign LUT_2[57863] = 32'b11111111111111110010011010011111;
assign LUT_2[57864] = 32'b11111111111111101100111100111111;
assign LUT_2[57865] = 32'b11111111111111101001110101011000;
assign LUT_2[57866] = 32'b11111111111111110011110101111011;
assign LUT_2[57867] = 32'b11111111111111110000101110010100;
assign LUT_2[57868] = 32'b11111111111111101001011010100111;
assign LUT_2[57869] = 32'b11111111111111100110010011000000;
assign LUT_2[57870] = 32'b11111111111111110000010011100011;
assign LUT_2[57871] = 32'b11111111111111101101001011111100;
assign LUT_2[57872] = 32'b11111111111111101100101111101100;
assign LUT_2[57873] = 32'b11111111111111101001101000000101;
assign LUT_2[57874] = 32'b11111111111111110011101000101000;
assign LUT_2[57875] = 32'b11111111111111110000100001000001;
assign LUT_2[57876] = 32'b11111111111111101001001101010100;
assign LUT_2[57877] = 32'b11111111111111100110000101101101;
assign LUT_2[57878] = 32'b11111111111111110000000110010000;
assign LUT_2[57879] = 32'b11111111111111101100111110101001;
assign LUT_2[57880] = 32'b11111111111111100111100001001001;
assign LUT_2[57881] = 32'b11111111111111100100011001100010;
assign LUT_2[57882] = 32'b11111111111111101110011010000101;
assign LUT_2[57883] = 32'b11111111111111101011010010011110;
assign LUT_2[57884] = 32'b11111111111111100011111110110001;
assign LUT_2[57885] = 32'b11111111111111100000110111001010;
assign LUT_2[57886] = 32'b11111111111111101010110111101101;
assign LUT_2[57887] = 32'b11111111111111100111110000000110;
assign LUT_2[57888] = 32'b11111111111111110010100111001011;
assign LUT_2[57889] = 32'b11111111111111101111011111100100;
assign LUT_2[57890] = 32'b11111111111111111001100000000111;
assign LUT_2[57891] = 32'b11111111111111110110011000100000;
assign LUT_2[57892] = 32'b11111111111111101111000100110011;
assign LUT_2[57893] = 32'b11111111111111101011111101001100;
assign LUT_2[57894] = 32'b11111111111111110101111101101111;
assign LUT_2[57895] = 32'b11111111111111110010110110001000;
assign LUT_2[57896] = 32'b11111111111111101101011000101000;
assign LUT_2[57897] = 32'b11111111111111101010010001000001;
assign LUT_2[57898] = 32'b11111111111111110100010001100100;
assign LUT_2[57899] = 32'b11111111111111110001001001111101;
assign LUT_2[57900] = 32'b11111111111111101001110110010000;
assign LUT_2[57901] = 32'b11111111111111100110101110101001;
assign LUT_2[57902] = 32'b11111111111111110000101111001100;
assign LUT_2[57903] = 32'b11111111111111101101100111100101;
assign LUT_2[57904] = 32'b11111111111111101101001011010101;
assign LUT_2[57905] = 32'b11111111111111101010000011101110;
assign LUT_2[57906] = 32'b11111111111111110100000100010001;
assign LUT_2[57907] = 32'b11111111111111110000111100101010;
assign LUT_2[57908] = 32'b11111111111111101001101000111101;
assign LUT_2[57909] = 32'b11111111111111100110100001010110;
assign LUT_2[57910] = 32'b11111111111111110000100001111001;
assign LUT_2[57911] = 32'b11111111111111101101011010010010;
assign LUT_2[57912] = 32'b11111111111111100111111100110010;
assign LUT_2[57913] = 32'b11111111111111100100110101001011;
assign LUT_2[57914] = 32'b11111111111111101110110101101110;
assign LUT_2[57915] = 32'b11111111111111101011101110000111;
assign LUT_2[57916] = 32'b11111111111111100100011010011010;
assign LUT_2[57917] = 32'b11111111111111100001010010110011;
assign LUT_2[57918] = 32'b11111111111111101011010011010110;
assign LUT_2[57919] = 32'b11111111111111101000001011101111;
assign LUT_2[57920] = 32'b11111111111111101010010100000101;
assign LUT_2[57921] = 32'b11111111111111100111001100011110;
assign LUT_2[57922] = 32'b11111111111111110001001101000001;
assign LUT_2[57923] = 32'b11111111111111101110000101011010;
assign LUT_2[57924] = 32'b11111111111111100110110001101101;
assign LUT_2[57925] = 32'b11111111111111100011101010000110;
assign LUT_2[57926] = 32'b11111111111111101101101010101001;
assign LUT_2[57927] = 32'b11111111111111101010100011000010;
assign LUT_2[57928] = 32'b11111111111111100101000101100010;
assign LUT_2[57929] = 32'b11111111111111100001111101111011;
assign LUT_2[57930] = 32'b11111111111111101011111110011110;
assign LUT_2[57931] = 32'b11111111111111101000110110110111;
assign LUT_2[57932] = 32'b11111111111111100001100011001010;
assign LUT_2[57933] = 32'b11111111111111011110011011100011;
assign LUT_2[57934] = 32'b11111111111111101000011100000110;
assign LUT_2[57935] = 32'b11111111111111100101010100011111;
assign LUT_2[57936] = 32'b11111111111111100100111000001111;
assign LUT_2[57937] = 32'b11111111111111100001110000101000;
assign LUT_2[57938] = 32'b11111111111111101011110001001011;
assign LUT_2[57939] = 32'b11111111111111101000101001100100;
assign LUT_2[57940] = 32'b11111111111111100001010101110111;
assign LUT_2[57941] = 32'b11111111111111011110001110010000;
assign LUT_2[57942] = 32'b11111111111111101000001110110011;
assign LUT_2[57943] = 32'b11111111111111100101000111001100;
assign LUT_2[57944] = 32'b11111111111111011111101001101100;
assign LUT_2[57945] = 32'b11111111111111011100100010000101;
assign LUT_2[57946] = 32'b11111111111111100110100010101000;
assign LUT_2[57947] = 32'b11111111111111100011011011000001;
assign LUT_2[57948] = 32'b11111111111111011100000111010100;
assign LUT_2[57949] = 32'b11111111111111011000111111101101;
assign LUT_2[57950] = 32'b11111111111111100011000000010000;
assign LUT_2[57951] = 32'b11111111111111011111111000101001;
assign LUT_2[57952] = 32'b11111111111111101010101111101110;
assign LUT_2[57953] = 32'b11111111111111100111101000000111;
assign LUT_2[57954] = 32'b11111111111111110001101000101010;
assign LUT_2[57955] = 32'b11111111111111101110100001000011;
assign LUT_2[57956] = 32'b11111111111111100111001101010110;
assign LUT_2[57957] = 32'b11111111111111100100000101101111;
assign LUT_2[57958] = 32'b11111111111111101110000110010010;
assign LUT_2[57959] = 32'b11111111111111101010111110101011;
assign LUT_2[57960] = 32'b11111111111111100101100001001011;
assign LUT_2[57961] = 32'b11111111111111100010011001100100;
assign LUT_2[57962] = 32'b11111111111111101100011010000111;
assign LUT_2[57963] = 32'b11111111111111101001010010100000;
assign LUT_2[57964] = 32'b11111111111111100001111110110011;
assign LUT_2[57965] = 32'b11111111111111011110110111001100;
assign LUT_2[57966] = 32'b11111111111111101000110111101111;
assign LUT_2[57967] = 32'b11111111111111100101110000001000;
assign LUT_2[57968] = 32'b11111111111111100101010011111000;
assign LUT_2[57969] = 32'b11111111111111100010001100010001;
assign LUT_2[57970] = 32'b11111111111111101100001100110100;
assign LUT_2[57971] = 32'b11111111111111101001000101001101;
assign LUT_2[57972] = 32'b11111111111111100001110001100000;
assign LUT_2[57973] = 32'b11111111111111011110101001111001;
assign LUT_2[57974] = 32'b11111111111111101000101010011100;
assign LUT_2[57975] = 32'b11111111111111100101100010110101;
assign LUT_2[57976] = 32'b11111111111111100000000101010101;
assign LUT_2[57977] = 32'b11111111111111011100111101101110;
assign LUT_2[57978] = 32'b11111111111111100110111110010001;
assign LUT_2[57979] = 32'b11111111111111100011110110101010;
assign LUT_2[57980] = 32'b11111111111111011100100010111101;
assign LUT_2[57981] = 32'b11111111111111011001011011010110;
assign LUT_2[57982] = 32'b11111111111111100011011011111001;
assign LUT_2[57983] = 32'b11111111111111100000010100010010;
assign LUT_2[57984] = 32'b11111111111111110110011111110001;
assign LUT_2[57985] = 32'b11111111111111110011011000001010;
assign LUT_2[57986] = 32'b11111111111111111101011000101101;
assign LUT_2[57987] = 32'b11111111111111111010010001000110;
assign LUT_2[57988] = 32'b11111111111111110010111101011001;
assign LUT_2[57989] = 32'b11111111111111101111110101110010;
assign LUT_2[57990] = 32'b11111111111111111001110110010101;
assign LUT_2[57991] = 32'b11111111111111110110101110101110;
assign LUT_2[57992] = 32'b11111111111111110001010001001110;
assign LUT_2[57993] = 32'b11111111111111101110001001100111;
assign LUT_2[57994] = 32'b11111111111111111000001010001010;
assign LUT_2[57995] = 32'b11111111111111110101000010100011;
assign LUT_2[57996] = 32'b11111111111111101101101110110110;
assign LUT_2[57997] = 32'b11111111111111101010100111001111;
assign LUT_2[57998] = 32'b11111111111111110100100111110010;
assign LUT_2[57999] = 32'b11111111111111110001100000001011;
assign LUT_2[58000] = 32'b11111111111111110001000011111011;
assign LUT_2[58001] = 32'b11111111111111101101111100010100;
assign LUT_2[58002] = 32'b11111111111111110111111100110111;
assign LUT_2[58003] = 32'b11111111111111110100110101010000;
assign LUT_2[58004] = 32'b11111111111111101101100001100011;
assign LUT_2[58005] = 32'b11111111111111101010011001111100;
assign LUT_2[58006] = 32'b11111111111111110100011010011111;
assign LUT_2[58007] = 32'b11111111111111110001010010111000;
assign LUT_2[58008] = 32'b11111111111111101011110101011000;
assign LUT_2[58009] = 32'b11111111111111101000101101110001;
assign LUT_2[58010] = 32'b11111111111111110010101110010100;
assign LUT_2[58011] = 32'b11111111111111101111100110101101;
assign LUT_2[58012] = 32'b11111111111111101000010011000000;
assign LUT_2[58013] = 32'b11111111111111100101001011011001;
assign LUT_2[58014] = 32'b11111111111111101111001011111100;
assign LUT_2[58015] = 32'b11111111111111101100000100010101;
assign LUT_2[58016] = 32'b11111111111111110110111011011010;
assign LUT_2[58017] = 32'b11111111111111110011110011110011;
assign LUT_2[58018] = 32'b11111111111111111101110100010110;
assign LUT_2[58019] = 32'b11111111111111111010101100101111;
assign LUT_2[58020] = 32'b11111111111111110011011001000010;
assign LUT_2[58021] = 32'b11111111111111110000010001011011;
assign LUT_2[58022] = 32'b11111111111111111010010001111110;
assign LUT_2[58023] = 32'b11111111111111110111001010010111;
assign LUT_2[58024] = 32'b11111111111111110001101100110111;
assign LUT_2[58025] = 32'b11111111111111101110100101010000;
assign LUT_2[58026] = 32'b11111111111111111000100101110011;
assign LUT_2[58027] = 32'b11111111111111110101011110001100;
assign LUT_2[58028] = 32'b11111111111111101110001010011111;
assign LUT_2[58029] = 32'b11111111111111101011000010111000;
assign LUT_2[58030] = 32'b11111111111111110101000011011011;
assign LUT_2[58031] = 32'b11111111111111110001111011110100;
assign LUT_2[58032] = 32'b11111111111111110001011111100100;
assign LUT_2[58033] = 32'b11111111111111101110010111111101;
assign LUT_2[58034] = 32'b11111111111111111000011000100000;
assign LUT_2[58035] = 32'b11111111111111110101010000111001;
assign LUT_2[58036] = 32'b11111111111111101101111101001100;
assign LUT_2[58037] = 32'b11111111111111101010110101100101;
assign LUT_2[58038] = 32'b11111111111111110100110110001000;
assign LUT_2[58039] = 32'b11111111111111110001101110100001;
assign LUT_2[58040] = 32'b11111111111111101100010001000001;
assign LUT_2[58041] = 32'b11111111111111101001001001011010;
assign LUT_2[58042] = 32'b11111111111111110011001001111101;
assign LUT_2[58043] = 32'b11111111111111110000000010010110;
assign LUT_2[58044] = 32'b11111111111111101000101110101001;
assign LUT_2[58045] = 32'b11111111111111100101100111000010;
assign LUT_2[58046] = 32'b11111111111111101111100111100101;
assign LUT_2[58047] = 32'b11111111111111101100011111111110;
assign LUT_2[58048] = 32'b11111111111111101110101000010100;
assign LUT_2[58049] = 32'b11111111111111101011100000101101;
assign LUT_2[58050] = 32'b11111111111111110101100001010000;
assign LUT_2[58051] = 32'b11111111111111110010011001101001;
assign LUT_2[58052] = 32'b11111111111111101011000101111100;
assign LUT_2[58053] = 32'b11111111111111100111111110010101;
assign LUT_2[58054] = 32'b11111111111111110001111110111000;
assign LUT_2[58055] = 32'b11111111111111101110110111010001;
assign LUT_2[58056] = 32'b11111111111111101001011001110001;
assign LUT_2[58057] = 32'b11111111111111100110010010001010;
assign LUT_2[58058] = 32'b11111111111111110000010010101101;
assign LUT_2[58059] = 32'b11111111111111101101001011000110;
assign LUT_2[58060] = 32'b11111111111111100101110111011001;
assign LUT_2[58061] = 32'b11111111111111100010101111110010;
assign LUT_2[58062] = 32'b11111111111111101100110000010101;
assign LUT_2[58063] = 32'b11111111111111101001101000101110;
assign LUT_2[58064] = 32'b11111111111111101001001100011110;
assign LUT_2[58065] = 32'b11111111111111100110000100110111;
assign LUT_2[58066] = 32'b11111111111111110000000101011010;
assign LUT_2[58067] = 32'b11111111111111101100111101110011;
assign LUT_2[58068] = 32'b11111111111111100101101010000110;
assign LUT_2[58069] = 32'b11111111111111100010100010011111;
assign LUT_2[58070] = 32'b11111111111111101100100011000010;
assign LUT_2[58071] = 32'b11111111111111101001011011011011;
assign LUT_2[58072] = 32'b11111111111111100011111101111011;
assign LUT_2[58073] = 32'b11111111111111100000110110010100;
assign LUT_2[58074] = 32'b11111111111111101010110110110111;
assign LUT_2[58075] = 32'b11111111111111100111101111010000;
assign LUT_2[58076] = 32'b11111111111111100000011011100011;
assign LUT_2[58077] = 32'b11111111111111011101010011111100;
assign LUT_2[58078] = 32'b11111111111111100111010100011111;
assign LUT_2[58079] = 32'b11111111111111100100001100111000;
assign LUT_2[58080] = 32'b11111111111111101111000011111101;
assign LUT_2[58081] = 32'b11111111111111101011111100010110;
assign LUT_2[58082] = 32'b11111111111111110101111100111001;
assign LUT_2[58083] = 32'b11111111111111110010110101010010;
assign LUT_2[58084] = 32'b11111111111111101011100001100101;
assign LUT_2[58085] = 32'b11111111111111101000011001111110;
assign LUT_2[58086] = 32'b11111111111111110010011010100001;
assign LUT_2[58087] = 32'b11111111111111101111010010111010;
assign LUT_2[58088] = 32'b11111111111111101001110101011010;
assign LUT_2[58089] = 32'b11111111111111100110101101110011;
assign LUT_2[58090] = 32'b11111111111111110000101110010110;
assign LUT_2[58091] = 32'b11111111111111101101100110101111;
assign LUT_2[58092] = 32'b11111111111111100110010011000010;
assign LUT_2[58093] = 32'b11111111111111100011001011011011;
assign LUT_2[58094] = 32'b11111111111111101101001011111110;
assign LUT_2[58095] = 32'b11111111111111101010000100010111;
assign LUT_2[58096] = 32'b11111111111111101001101000000111;
assign LUT_2[58097] = 32'b11111111111111100110100000100000;
assign LUT_2[58098] = 32'b11111111111111110000100001000011;
assign LUT_2[58099] = 32'b11111111111111101101011001011100;
assign LUT_2[58100] = 32'b11111111111111100110000101101111;
assign LUT_2[58101] = 32'b11111111111111100010111110001000;
assign LUT_2[58102] = 32'b11111111111111101100111110101011;
assign LUT_2[58103] = 32'b11111111111111101001110111000100;
assign LUT_2[58104] = 32'b11111111111111100100011001100100;
assign LUT_2[58105] = 32'b11111111111111100001010001111101;
assign LUT_2[58106] = 32'b11111111111111101011010010100000;
assign LUT_2[58107] = 32'b11111111111111101000001010111001;
assign LUT_2[58108] = 32'b11111111111111100000110111001100;
assign LUT_2[58109] = 32'b11111111111111011101101111100101;
assign LUT_2[58110] = 32'b11111111111111100111110000001000;
assign LUT_2[58111] = 32'b11111111111111100100101000100001;
assign LUT_2[58112] = 32'b11111111111111110110001010001000;
assign LUT_2[58113] = 32'b11111111111111110011000010100001;
assign LUT_2[58114] = 32'b11111111111111111101000011000100;
assign LUT_2[58115] = 32'b11111111111111111001111011011101;
assign LUT_2[58116] = 32'b11111111111111110010100111110000;
assign LUT_2[58117] = 32'b11111111111111101111100000001001;
assign LUT_2[58118] = 32'b11111111111111111001100000101100;
assign LUT_2[58119] = 32'b11111111111111110110011001000101;
assign LUT_2[58120] = 32'b11111111111111110000111011100101;
assign LUT_2[58121] = 32'b11111111111111101101110011111110;
assign LUT_2[58122] = 32'b11111111111111110111110100100001;
assign LUT_2[58123] = 32'b11111111111111110100101100111010;
assign LUT_2[58124] = 32'b11111111111111101101011001001101;
assign LUT_2[58125] = 32'b11111111111111101010010001100110;
assign LUT_2[58126] = 32'b11111111111111110100010010001001;
assign LUT_2[58127] = 32'b11111111111111110001001010100010;
assign LUT_2[58128] = 32'b11111111111111110000101110010010;
assign LUT_2[58129] = 32'b11111111111111101101100110101011;
assign LUT_2[58130] = 32'b11111111111111110111100111001110;
assign LUT_2[58131] = 32'b11111111111111110100011111100111;
assign LUT_2[58132] = 32'b11111111111111101101001011111010;
assign LUT_2[58133] = 32'b11111111111111101010000100010011;
assign LUT_2[58134] = 32'b11111111111111110100000100110110;
assign LUT_2[58135] = 32'b11111111111111110000111101001111;
assign LUT_2[58136] = 32'b11111111111111101011011111101111;
assign LUT_2[58137] = 32'b11111111111111101000011000001000;
assign LUT_2[58138] = 32'b11111111111111110010011000101011;
assign LUT_2[58139] = 32'b11111111111111101111010001000100;
assign LUT_2[58140] = 32'b11111111111111100111111101010111;
assign LUT_2[58141] = 32'b11111111111111100100110101110000;
assign LUT_2[58142] = 32'b11111111111111101110110110010011;
assign LUT_2[58143] = 32'b11111111111111101011101110101100;
assign LUT_2[58144] = 32'b11111111111111110110100101110001;
assign LUT_2[58145] = 32'b11111111111111110011011110001010;
assign LUT_2[58146] = 32'b11111111111111111101011110101101;
assign LUT_2[58147] = 32'b11111111111111111010010111000110;
assign LUT_2[58148] = 32'b11111111111111110011000011011001;
assign LUT_2[58149] = 32'b11111111111111101111111011110010;
assign LUT_2[58150] = 32'b11111111111111111001111100010101;
assign LUT_2[58151] = 32'b11111111111111110110110100101110;
assign LUT_2[58152] = 32'b11111111111111110001010111001110;
assign LUT_2[58153] = 32'b11111111111111101110001111100111;
assign LUT_2[58154] = 32'b11111111111111111000010000001010;
assign LUT_2[58155] = 32'b11111111111111110101001000100011;
assign LUT_2[58156] = 32'b11111111111111101101110100110110;
assign LUT_2[58157] = 32'b11111111111111101010101101001111;
assign LUT_2[58158] = 32'b11111111111111110100101101110010;
assign LUT_2[58159] = 32'b11111111111111110001100110001011;
assign LUT_2[58160] = 32'b11111111111111110001001001111011;
assign LUT_2[58161] = 32'b11111111111111101110000010010100;
assign LUT_2[58162] = 32'b11111111111111111000000010110111;
assign LUT_2[58163] = 32'b11111111111111110100111011010000;
assign LUT_2[58164] = 32'b11111111111111101101100111100011;
assign LUT_2[58165] = 32'b11111111111111101010011111111100;
assign LUT_2[58166] = 32'b11111111111111110100100000011111;
assign LUT_2[58167] = 32'b11111111111111110001011000111000;
assign LUT_2[58168] = 32'b11111111111111101011111011011000;
assign LUT_2[58169] = 32'b11111111111111101000110011110001;
assign LUT_2[58170] = 32'b11111111111111110010110100010100;
assign LUT_2[58171] = 32'b11111111111111101111101100101101;
assign LUT_2[58172] = 32'b11111111111111101000011001000000;
assign LUT_2[58173] = 32'b11111111111111100101010001011001;
assign LUT_2[58174] = 32'b11111111111111101111010001111100;
assign LUT_2[58175] = 32'b11111111111111101100001010010101;
assign LUT_2[58176] = 32'b11111111111111101110010010101011;
assign LUT_2[58177] = 32'b11111111111111101011001011000100;
assign LUT_2[58178] = 32'b11111111111111110101001011100111;
assign LUT_2[58179] = 32'b11111111111111110010000100000000;
assign LUT_2[58180] = 32'b11111111111111101010110000010011;
assign LUT_2[58181] = 32'b11111111111111100111101000101100;
assign LUT_2[58182] = 32'b11111111111111110001101001001111;
assign LUT_2[58183] = 32'b11111111111111101110100001101000;
assign LUT_2[58184] = 32'b11111111111111101001000100001000;
assign LUT_2[58185] = 32'b11111111111111100101111100100001;
assign LUT_2[58186] = 32'b11111111111111101111111101000100;
assign LUT_2[58187] = 32'b11111111111111101100110101011101;
assign LUT_2[58188] = 32'b11111111111111100101100001110000;
assign LUT_2[58189] = 32'b11111111111111100010011010001001;
assign LUT_2[58190] = 32'b11111111111111101100011010101100;
assign LUT_2[58191] = 32'b11111111111111101001010011000101;
assign LUT_2[58192] = 32'b11111111111111101000110110110101;
assign LUT_2[58193] = 32'b11111111111111100101101111001110;
assign LUT_2[58194] = 32'b11111111111111101111101111110001;
assign LUT_2[58195] = 32'b11111111111111101100101000001010;
assign LUT_2[58196] = 32'b11111111111111100101010100011101;
assign LUT_2[58197] = 32'b11111111111111100010001100110110;
assign LUT_2[58198] = 32'b11111111111111101100001101011001;
assign LUT_2[58199] = 32'b11111111111111101001000101110010;
assign LUT_2[58200] = 32'b11111111111111100011101000010010;
assign LUT_2[58201] = 32'b11111111111111100000100000101011;
assign LUT_2[58202] = 32'b11111111111111101010100001001110;
assign LUT_2[58203] = 32'b11111111111111100111011001100111;
assign LUT_2[58204] = 32'b11111111111111100000000101111010;
assign LUT_2[58205] = 32'b11111111111111011100111110010011;
assign LUT_2[58206] = 32'b11111111111111100110111110110110;
assign LUT_2[58207] = 32'b11111111111111100011110111001111;
assign LUT_2[58208] = 32'b11111111111111101110101110010100;
assign LUT_2[58209] = 32'b11111111111111101011100110101101;
assign LUT_2[58210] = 32'b11111111111111110101100111010000;
assign LUT_2[58211] = 32'b11111111111111110010011111101001;
assign LUT_2[58212] = 32'b11111111111111101011001011111100;
assign LUT_2[58213] = 32'b11111111111111101000000100010101;
assign LUT_2[58214] = 32'b11111111111111110010000100111000;
assign LUT_2[58215] = 32'b11111111111111101110111101010001;
assign LUT_2[58216] = 32'b11111111111111101001011111110001;
assign LUT_2[58217] = 32'b11111111111111100110011000001010;
assign LUT_2[58218] = 32'b11111111111111110000011000101101;
assign LUT_2[58219] = 32'b11111111111111101101010001000110;
assign LUT_2[58220] = 32'b11111111111111100101111101011001;
assign LUT_2[58221] = 32'b11111111111111100010110101110010;
assign LUT_2[58222] = 32'b11111111111111101100110110010101;
assign LUT_2[58223] = 32'b11111111111111101001101110101110;
assign LUT_2[58224] = 32'b11111111111111101001010010011110;
assign LUT_2[58225] = 32'b11111111111111100110001010110111;
assign LUT_2[58226] = 32'b11111111111111110000001011011010;
assign LUT_2[58227] = 32'b11111111111111101101000011110011;
assign LUT_2[58228] = 32'b11111111111111100101110000000110;
assign LUT_2[58229] = 32'b11111111111111100010101000011111;
assign LUT_2[58230] = 32'b11111111111111101100101001000010;
assign LUT_2[58231] = 32'b11111111111111101001100001011011;
assign LUT_2[58232] = 32'b11111111111111100100000011111011;
assign LUT_2[58233] = 32'b11111111111111100000111100010100;
assign LUT_2[58234] = 32'b11111111111111101010111100110111;
assign LUT_2[58235] = 32'b11111111111111100111110101010000;
assign LUT_2[58236] = 32'b11111111111111100000100001100011;
assign LUT_2[58237] = 32'b11111111111111011101011001111100;
assign LUT_2[58238] = 32'b11111111111111100111011010011111;
assign LUT_2[58239] = 32'b11111111111111100100010010111000;
assign LUT_2[58240] = 32'b11111111111111111010011110010111;
assign LUT_2[58241] = 32'b11111111111111110111010110110000;
assign LUT_2[58242] = 32'b00000000000000000001010111010011;
assign LUT_2[58243] = 32'b11111111111111111110001111101100;
assign LUT_2[58244] = 32'b11111111111111110110111011111111;
assign LUT_2[58245] = 32'b11111111111111110011110100011000;
assign LUT_2[58246] = 32'b11111111111111111101110100111011;
assign LUT_2[58247] = 32'b11111111111111111010101101010100;
assign LUT_2[58248] = 32'b11111111111111110101001111110100;
assign LUT_2[58249] = 32'b11111111111111110010001000001101;
assign LUT_2[58250] = 32'b11111111111111111100001000110000;
assign LUT_2[58251] = 32'b11111111111111111001000001001001;
assign LUT_2[58252] = 32'b11111111111111110001101101011100;
assign LUT_2[58253] = 32'b11111111111111101110100101110101;
assign LUT_2[58254] = 32'b11111111111111111000100110011000;
assign LUT_2[58255] = 32'b11111111111111110101011110110001;
assign LUT_2[58256] = 32'b11111111111111110101000010100001;
assign LUT_2[58257] = 32'b11111111111111110001111010111010;
assign LUT_2[58258] = 32'b11111111111111111011111011011101;
assign LUT_2[58259] = 32'b11111111111111111000110011110110;
assign LUT_2[58260] = 32'b11111111111111110001100000001001;
assign LUT_2[58261] = 32'b11111111111111101110011000100010;
assign LUT_2[58262] = 32'b11111111111111111000011001000101;
assign LUT_2[58263] = 32'b11111111111111110101010001011110;
assign LUT_2[58264] = 32'b11111111111111101111110011111110;
assign LUT_2[58265] = 32'b11111111111111101100101100010111;
assign LUT_2[58266] = 32'b11111111111111110110101100111010;
assign LUT_2[58267] = 32'b11111111111111110011100101010011;
assign LUT_2[58268] = 32'b11111111111111101100010001100110;
assign LUT_2[58269] = 32'b11111111111111101001001001111111;
assign LUT_2[58270] = 32'b11111111111111110011001010100010;
assign LUT_2[58271] = 32'b11111111111111110000000010111011;
assign LUT_2[58272] = 32'b11111111111111111010111010000000;
assign LUT_2[58273] = 32'b11111111111111110111110010011001;
assign LUT_2[58274] = 32'b00000000000000000001110010111100;
assign LUT_2[58275] = 32'b11111111111111111110101011010101;
assign LUT_2[58276] = 32'b11111111111111110111010111101000;
assign LUT_2[58277] = 32'b11111111111111110100010000000001;
assign LUT_2[58278] = 32'b11111111111111111110010000100100;
assign LUT_2[58279] = 32'b11111111111111111011001000111101;
assign LUT_2[58280] = 32'b11111111111111110101101011011101;
assign LUT_2[58281] = 32'b11111111111111110010100011110110;
assign LUT_2[58282] = 32'b11111111111111111100100100011001;
assign LUT_2[58283] = 32'b11111111111111111001011100110010;
assign LUT_2[58284] = 32'b11111111111111110010001001000101;
assign LUT_2[58285] = 32'b11111111111111101111000001011110;
assign LUT_2[58286] = 32'b11111111111111111001000010000001;
assign LUT_2[58287] = 32'b11111111111111110101111010011010;
assign LUT_2[58288] = 32'b11111111111111110101011110001010;
assign LUT_2[58289] = 32'b11111111111111110010010110100011;
assign LUT_2[58290] = 32'b11111111111111111100010111000110;
assign LUT_2[58291] = 32'b11111111111111111001001111011111;
assign LUT_2[58292] = 32'b11111111111111110001111011110010;
assign LUT_2[58293] = 32'b11111111111111101110110100001011;
assign LUT_2[58294] = 32'b11111111111111111000110100101110;
assign LUT_2[58295] = 32'b11111111111111110101101101000111;
assign LUT_2[58296] = 32'b11111111111111110000001111100111;
assign LUT_2[58297] = 32'b11111111111111101101001000000000;
assign LUT_2[58298] = 32'b11111111111111110111001000100011;
assign LUT_2[58299] = 32'b11111111111111110100000000111100;
assign LUT_2[58300] = 32'b11111111111111101100101101001111;
assign LUT_2[58301] = 32'b11111111111111101001100101101000;
assign LUT_2[58302] = 32'b11111111111111110011100110001011;
assign LUT_2[58303] = 32'b11111111111111110000011110100100;
assign LUT_2[58304] = 32'b11111111111111110010100110111010;
assign LUT_2[58305] = 32'b11111111111111101111011111010011;
assign LUT_2[58306] = 32'b11111111111111111001011111110110;
assign LUT_2[58307] = 32'b11111111111111110110011000001111;
assign LUT_2[58308] = 32'b11111111111111101111000100100010;
assign LUT_2[58309] = 32'b11111111111111101011111100111011;
assign LUT_2[58310] = 32'b11111111111111110101111101011110;
assign LUT_2[58311] = 32'b11111111111111110010110101110111;
assign LUT_2[58312] = 32'b11111111111111101101011000010111;
assign LUT_2[58313] = 32'b11111111111111101010010000110000;
assign LUT_2[58314] = 32'b11111111111111110100010001010011;
assign LUT_2[58315] = 32'b11111111111111110001001001101100;
assign LUT_2[58316] = 32'b11111111111111101001110101111111;
assign LUT_2[58317] = 32'b11111111111111100110101110011000;
assign LUT_2[58318] = 32'b11111111111111110000101110111011;
assign LUT_2[58319] = 32'b11111111111111101101100111010100;
assign LUT_2[58320] = 32'b11111111111111101101001011000100;
assign LUT_2[58321] = 32'b11111111111111101010000011011101;
assign LUT_2[58322] = 32'b11111111111111110100000100000000;
assign LUT_2[58323] = 32'b11111111111111110000111100011001;
assign LUT_2[58324] = 32'b11111111111111101001101000101100;
assign LUT_2[58325] = 32'b11111111111111100110100001000101;
assign LUT_2[58326] = 32'b11111111111111110000100001101000;
assign LUT_2[58327] = 32'b11111111111111101101011010000001;
assign LUT_2[58328] = 32'b11111111111111100111111100100001;
assign LUT_2[58329] = 32'b11111111111111100100110100111010;
assign LUT_2[58330] = 32'b11111111111111101110110101011101;
assign LUT_2[58331] = 32'b11111111111111101011101101110110;
assign LUT_2[58332] = 32'b11111111111111100100011010001001;
assign LUT_2[58333] = 32'b11111111111111100001010010100010;
assign LUT_2[58334] = 32'b11111111111111101011010011000101;
assign LUT_2[58335] = 32'b11111111111111101000001011011110;
assign LUT_2[58336] = 32'b11111111111111110011000010100011;
assign LUT_2[58337] = 32'b11111111111111101111111010111100;
assign LUT_2[58338] = 32'b11111111111111111001111011011111;
assign LUT_2[58339] = 32'b11111111111111110110110011111000;
assign LUT_2[58340] = 32'b11111111111111101111100000001011;
assign LUT_2[58341] = 32'b11111111111111101100011000100100;
assign LUT_2[58342] = 32'b11111111111111110110011001000111;
assign LUT_2[58343] = 32'b11111111111111110011010001100000;
assign LUT_2[58344] = 32'b11111111111111101101110100000000;
assign LUT_2[58345] = 32'b11111111111111101010101100011001;
assign LUT_2[58346] = 32'b11111111111111110100101100111100;
assign LUT_2[58347] = 32'b11111111111111110001100101010101;
assign LUT_2[58348] = 32'b11111111111111101010010001101000;
assign LUT_2[58349] = 32'b11111111111111100111001010000001;
assign LUT_2[58350] = 32'b11111111111111110001001010100100;
assign LUT_2[58351] = 32'b11111111111111101110000010111101;
assign LUT_2[58352] = 32'b11111111111111101101100110101101;
assign LUT_2[58353] = 32'b11111111111111101010011111000110;
assign LUT_2[58354] = 32'b11111111111111110100011111101001;
assign LUT_2[58355] = 32'b11111111111111110001011000000010;
assign LUT_2[58356] = 32'b11111111111111101010000100010101;
assign LUT_2[58357] = 32'b11111111111111100110111100101110;
assign LUT_2[58358] = 32'b11111111111111110000111101010001;
assign LUT_2[58359] = 32'b11111111111111101101110101101010;
assign LUT_2[58360] = 32'b11111111111111101000011000001010;
assign LUT_2[58361] = 32'b11111111111111100101010000100011;
assign LUT_2[58362] = 32'b11111111111111101111010001000110;
assign LUT_2[58363] = 32'b11111111111111101100001001011111;
assign LUT_2[58364] = 32'b11111111111111100100110101110010;
assign LUT_2[58365] = 32'b11111111111111100001101110001011;
assign LUT_2[58366] = 32'b11111111111111101011101110101110;
assign LUT_2[58367] = 32'b11111111111111101000100111000111;
assign LUT_2[58368] = 32'b11111111111111110100000101110101;
assign LUT_2[58369] = 32'b11111111111111110000111110001110;
assign LUT_2[58370] = 32'b11111111111111111010111110110001;
assign LUT_2[58371] = 32'b11111111111111110111110111001010;
assign LUT_2[58372] = 32'b11111111111111110000100011011101;
assign LUT_2[58373] = 32'b11111111111111101101011011110110;
assign LUT_2[58374] = 32'b11111111111111110111011100011001;
assign LUT_2[58375] = 32'b11111111111111110100010100110010;
assign LUT_2[58376] = 32'b11111111111111101110110111010010;
assign LUT_2[58377] = 32'b11111111111111101011101111101011;
assign LUT_2[58378] = 32'b11111111111111110101110000001110;
assign LUT_2[58379] = 32'b11111111111111110010101000100111;
assign LUT_2[58380] = 32'b11111111111111101011010100111010;
assign LUT_2[58381] = 32'b11111111111111101000001101010011;
assign LUT_2[58382] = 32'b11111111111111110010001101110110;
assign LUT_2[58383] = 32'b11111111111111101111000110001111;
assign LUT_2[58384] = 32'b11111111111111101110101001111111;
assign LUT_2[58385] = 32'b11111111111111101011100010011000;
assign LUT_2[58386] = 32'b11111111111111110101100010111011;
assign LUT_2[58387] = 32'b11111111111111110010011011010100;
assign LUT_2[58388] = 32'b11111111111111101011000111100111;
assign LUT_2[58389] = 32'b11111111111111101000000000000000;
assign LUT_2[58390] = 32'b11111111111111110010000000100011;
assign LUT_2[58391] = 32'b11111111111111101110111000111100;
assign LUT_2[58392] = 32'b11111111111111101001011011011100;
assign LUT_2[58393] = 32'b11111111111111100110010011110101;
assign LUT_2[58394] = 32'b11111111111111110000010100011000;
assign LUT_2[58395] = 32'b11111111111111101101001100110001;
assign LUT_2[58396] = 32'b11111111111111100101111001000100;
assign LUT_2[58397] = 32'b11111111111111100010110001011101;
assign LUT_2[58398] = 32'b11111111111111101100110010000000;
assign LUT_2[58399] = 32'b11111111111111101001101010011001;
assign LUT_2[58400] = 32'b11111111111111110100100001011110;
assign LUT_2[58401] = 32'b11111111111111110001011001110111;
assign LUT_2[58402] = 32'b11111111111111111011011010011010;
assign LUT_2[58403] = 32'b11111111111111111000010010110011;
assign LUT_2[58404] = 32'b11111111111111110000111111000110;
assign LUT_2[58405] = 32'b11111111111111101101110111011111;
assign LUT_2[58406] = 32'b11111111111111110111111000000010;
assign LUT_2[58407] = 32'b11111111111111110100110000011011;
assign LUT_2[58408] = 32'b11111111111111101111010010111011;
assign LUT_2[58409] = 32'b11111111111111101100001011010100;
assign LUT_2[58410] = 32'b11111111111111110110001011110111;
assign LUT_2[58411] = 32'b11111111111111110011000100010000;
assign LUT_2[58412] = 32'b11111111111111101011110000100011;
assign LUT_2[58413] = 32'b11111111111111101000101000111100;
assign LUT_2[58414] = 32'b11111111111111110010101001011111;
assign LUT_2[58415] = 32'b11111111111111101111100001111000;
assign LUT_2[58416] = 32'b11111111111111101111000101101000;
assign LUT_2[58417] = 32'b11111111111111101011111110000001;
assign LUT_2[58418] = 32'b11111111111111110101111110100100;
assign LUT_2[58419] = 32'b11111111111111110010110110111101;
assign LUT_2[58420] = 32'b11111111111111101011100011010000;
assign LUT_2[58421] = 32'b11111111111111101000011011101001;
assign LUT_2[58422] = 32'b11111111111111110010011100001100;
assign LUT_2[58423] = 32'b11111111111111101111010100100101;
assign LUT_2[58424] = 32'b11111111111111101001110111000101;
assign LUT_2[58425] = 32'b11111111111111100110101111011110;
assign LUT_2[58426] = 32'b11111111111111110000110000000001;
assign LUT_2[58427] = 32'b11111111111111101101101000011010;
assign LUT_2[58428] = 32'b11111111111111100110010100101101;
assign LUT_2[58429] = 32'b11111111111111100011001101000110;
assign LUT_2[58430] = 32'b11111111111111101101001101101001;
assign LUT_2[58431] = 32'b11111111111111101010000110000010;
assign LUT_2[58432] = 32'b11111111111111101100001110011000;
assign LUT_2[58433] = 32'b11111111111111101001000110110001;
assign LUT_2[58434] = 32'b11111111111111110011000111010100;
assign LUT_2[58435] = 32'b11111111111111101111111111101101;
assign LUT_2[58436] = 32'b11111111111111101000101100000000;
assign LUT_2[58437] = 32'b11111111111111100101100100011001;
assign LUT_2[58438] = 32'b11111111111111101111100100111100;
assign LUT_2[58439] = 32'b11111111111111101100011101010101;
assign LUT_2[58440] = 32'b11111111111111100110111111110101;
assign LUT_2[58441] = 32'b11111111111111100011111000001110;
assign LUT_2[58442] = 32'b11111111111111101101111000110001;
assign LUT_2[58443] = 32'b11111111111111101010110001001010;
assign LUT_2[58444] = 32'b11111111111111100011011101011101;
assign LUT_2[58445] = 32'b11111111111111100000010101110110;
assign LUT_2[58446] = 32'b11111111111111101010010110011001;
assign LUT_2[58447] = 32'b11111111111111100111001110110010;
assign LUT_2[58448] = 32'b11111111111111100110110010100010;
assign LUT_2[58449] = 32'b11111111111111100011101010111011;
assign LUT_2[58450] = 32'b11111111111111101101101011011110;
assign LUT_2[58451] = 32'b11111111111111101010100011110111;
assign LUT_2[58452] = 32'b11111111111111100011010000001010;
assign LUT_2[58453] = 32'b11111111111111100000001000100011;
assign LUT_2[58454] = 32'b11111111111111101010001001000110;
assign LUT_2[58455] = 32'b11111111111111100111000001011111;
assign LUT_2[58456] = 32'b11111111111111100001100011111111;
assign LUT_2[58457] = 32'b11111111111111011110011100011000;
assign LUT_2[58458] = 32'b11111111111111101000011100111011;
assign LUT_2[58459] = 32'b11111111111111100101010101010100;
assign LUT_2[58460] = 32'b11111111111111011110000001100111;
assign LUT_2[58461] = 32'b11111111111111011010111010000000;
assign LUT_2[58462] = 32'b11111111111111100100111010100011;
assign LUT_2[58463] = 32'b11111111111111100001110010111100;
assign LUT_2[58464] = 32'b11111111111111101100101010000001;
assign LUT_2[58465] = 32'b11111111111111101001100010011010;
assign LUT_2[58466] = 32'b11111111111111110011100010111101;
assign LUT_2[58467] = 32'b11111111111111110000011011010110;
assign LUT_2[58468] = 32'b11111111111111101001000111101001;
assign LUT_2[58469] = 32'b11111111111111100110000000000010;
assign LUT_2[58470] = 32'b11111111111111110000000000100101;
assign LUT_2[58471] = 32'b11111111111111101100111000111110;
assign LUT_2[58472] = 32'b11111111111111100111011011011110;
assign LUT_2[58473] = 32'b11111111111111100100010011110111;
assign LUT_2[58474] = 32'b11111111111111101110010100011010;
assign LUT_2[58475] = 32'b11111111111111101011001100110011;
assign LUT_2[58476] = 32'b11111111111111100011111001000110;
assign LUT_2[58477] = 32'b11111111111111100000110001011111;
assign LUT_2[58478] = 32'b11111111111111101010110010000010;
assign LUT_2[58479] = 32'b11111111111111100111101010011011;
assign LUT_2[58480] = 32'b11111111111111100111001110001011;
assign LUT_2[58481] = 32'b11111111111111100100000110100100;
assign LUT_2[58482] = 32'b11111111111111101110000111000111;
assign LUT_2[58483] = 32'b11111111111111101010111111100000;
assign LUT_2[58484] = 32'b11111111111111100011101011110011;
assign LUT_2[58485] = 32'b11111111111111100000100100001100;
assign LUT_2[58486] = 32'b11111111111111101010100100101111;
assign LUT_2[58487] = 32'b11111111111111100111011101001000;
assign LUT_2[58488] = 32'b11111111111111100001111111101000;
assign LUT_2[58489] = 32'b11111111111111011110111000000001;
assign LUT_2[58490] = 32'b11111111111111101000111000100100;
assign LUT_2[58491] = 32'b11111111111111100101110000111101;
assign LUT_2[58492] = 32'b11111111111111011110011101010000;
assign LUT_2[58493] = 32'b11111111111111011011010101101001;
assign LUT_2[58494] = 32'b11111111111111100101010110001100;
assign LUT_2[58495] = 32'b11111111111111100010001110100101;
assign LUT_2[58496] = 32'b11111111111111111000011010000100;
assign LUT_2[58497] = 32'b11111111111111110101010010011101;
assign LUT_2[58498] = 32'b11111111111111111111010011000000;
assign LUT_2[58499] = 32'b11111111111111111100001011011001;
assign LUT_2[58500] = 32'b11111111111111110100110111101100;
assign LUT_2[58501] = 32'b11111111111111110001110000000101;
assign LUT_2[58502] = 32'b11111111111111111011110000101000;
assign LUT_2[58503] = 32'b11111111111111111000101001000001;
assign LUT_2[58504] = 32'b11111111111111110011001011100001;
assign LUT_2[58505] = 32'b11111111111111110000000011111010;
assign LUT_2[58506] = 32'b11111111111111111010000100011101;
assign LUT_2[58507] = 32'b11111111111111110110111100110110;
assign LUT_2[58508] = 32'b11111111111111101111101001001001;
assign LUT_2[58509] = 32'b11111111111111101100100001100010;
assign LUT_2[58510] = 32'b11111111111111110110100010000101;
assign LUT_2[58511] = 32'b11111111111111110011011010011110;
assign LUT_2[58512] = 32'b11111111111111110010111110001110;
assign LUT_2[58513] = 32'b11111111111111101111110110100111;
assign LUT_2[58514] = 32'b11111111111111111001110111001010;
assign LUT_2[58515] = 32'b11111111111111110110101111100011;
assign LUT_2[58516] = 32'b11111111111111101111011011110110;
assign LUT_2[58517] = 32'b11111111111111101100010100001111;
assign LUT_2[58518] = 32'b11111111111111110110010100110010;
assign LUT_2[58519] = 32'b11111111111111110011001101001011;
assign LUT_2[58520] = 32'b11111111111111101101101111101011;
assign LUT_2[58521] = 32'b11111111111111101010101000000100;
assign LUT_2[58522] = 32'b11111111111111110100101000100111;
assign LUT_2[58523] = 32'b11111111111111110001100001000000;
assign LUT_2[58524] = 32'b11111111111111101010001101010011;
assign LUT_2[58525] = 32'b11111111111111100111000101101100;
assign LUT_2[58526] = 32'b11111111111111110001000110001111;
assign LUT_2[58527] = 32'b11111111111111101101111110101000;
assign LUT_2[58528] = 32'b11111111111111111000110101101101;
assign LUT_2[58529] = 32'b11111111111111110101101110000110;
assign LUT_2[58530] = 32'b11111111111111111111101110101001;
assign LUT_2[58531] = 32'b11111111111111111100100111000010;
assign LUT_2[58532] = 32'b11111111111111110101010011010101;
assign LUT_2[58533] = 32'b11111111111111110010001011101110;
assign LUT_2[58534] = 32'b11111111111111111100001100010001;
assign LUT_2[58535] = 32'b11111111111111111001000100101010;
assign LUT_2[58536] = 32'b11111111111111110011100111001010;
assign LUT_2[58537] = 32'b11111111111111110000011111100011;
assign LUT_2[58538] = 32'b11111111111111111010100000000110;
assign LUT_2[58539] = 32'b11111111111111110111011000011111;
assign LUT_2[58540] = 32'b11111111111111110000000100110010;
assign LUT_2[58541] = 32'b11111111111111101100111101001011;
assign LUT_2[58542] = 32'b11111111111111110110111101101110;
assign LUT_2[58543] = 32'b11111111111111110011110110000111;
assign LUT_2[58544] = 32'b11111111111111110011011001110111;
assign LUT_2[58545] = 32'b11111111111111110000010010010000;
assign LUT_2[58546] = 32'b11111111111111111010010010110011;
assign LUT_2[58547] = 32'b11111111111111110111001011001100;
assign LUT_2[58548] = 32'b11111111111111101111110111011111;
assign LUT_2[58549] = 32'b11111111111111101100101111111000;
assign LUT_2[58550] = 32'b11111111111111110110110000011011;
assign LUT_2[58551] = 32'b11111111111111110011101000110100;
assign LUT_2[58552] = 32'b11111111111111101110001011010100;
assign LUT_2[58553] = 32'b11111111111111101011000011101101;
assign LUT_2[58554] = 32'b11111111111111110101000100010000;
assign LUT_2[58555] = 32'b11111111111111110001111100101001;
assign LUT_2[58556] = 32'b11111111111111101010101000111100;
assign LUT_2[58557] = 32'b11111111111111100111100001010101;
assign LUT_2[58558] = 32'b11111111111111110001100001111000;
assign LUT_2[58559] = 32'b11111111111111101110011010010001;
assign LUT_2[58560] = 32'b11111111111111110000100010100111;
assign LUT_2[58561] = 32'b11111111111111101101011011000000;
assign LUT_2[58562] = 32'b11111111111111110111011011100011;
assign LUT_2[58563] = 32'b11111111111111110100010011111100;
assign LUT_2[58564] = 32'b11111111111111101101000000001111;
assign LUT_2[58565] = 32'b11111111111111101001111000101000;
assign LUT_2[58566] = 32'b11111111111111110011111001001011;
assign LUT_2[58567] = 32'b11111111111111110000110001100100;
assign LUT_2[58568] = 32'b11111111111111101011010100000100;
assign LUT_2[58569] = 32'b11111111111111101000001100011101;
assign LUT_2[58570] = 32'b11111111111111110010001101000000;
assign LUT_2[58571] = 32'b11111111111111101111000101011001;
assign LUT_2[58572] = 32'b11111111111111100111110001101100;
assign LUT_2[58573] = 32'b11111111111111100100101010000101;
assign LUT_2[58574] = 32'b11111111111111101110101010101000;
assign LUT_2[58575] = 32'b11111111111111101011100011000001;
assign LUT_2[58576] = 32'b11111111111111101011000110110001;
assign LUT_2[58577] = 32'b11111111111111100111111111001010;
assign LUT_2[58578] = 32'b11111111111111110001111111101101;
assign LUT_2[58579] = 32'b11111111111111101110111000000110;
assign LUT_2[58580] = 32'b11111111111111100111100100011001;
assign LUT_2[58581] = 32'b11111111111111100100011100110010;
assign LUT_2[58582] = 32'b11111111111111101110011101010101;
assign LUT_2[58583] = 32'b11111111111111101011010101101110;
assign LUT_2[58584] = 32'b11111111111111100101111000001110;
assign LUT_2[58585] = 32'b11111111111111100010110000100111;
assign LUT_2[58586] = 32'b11111111111111101100110001001010;
assign LUT_2[58587] = 32'b11111111111111101001101001100011;
assign LUT_2[58588] = 32'b11111111111111100010010101110110;
assign LUT_2[58589] = 32'b11111111111111011111001110001111;
assign LUT_2[58590] = 32'b11111111111111101001001110110010;
assign LUT_2[58591] = 32'b11111111111111100110000111001011;
assign LUT_2[58592] = 32'b11111111111111110000111110010000;
assign LUT_2[58593] = 32'b11111111111111101101110110101001;
assign LUT_2[58594] = 32'b11111111111111110111110111001100;
assign LUT_2[58595] = 32'b11111111111111110100101111100101;
assign LUT_2[58596] = 32'b11111111111111101101011011111000;
assign LUT_2[58597] = 32'b11111111111111101010010100010001;
assign LUT_2[58598] = 32'b11111111111111110100010100110100;
assign LUT_2[58599] = 32'b11111111111111110001001101001101;
assign LUT_2[58600] = 32'b11111111111111101011101111101101;
assign LUT_2[58601] = 32'b11111111111111101000101000000110;
assign LUT_2[58602] = 32'b11111111111111110010101000101001;
assign LUT_2[58603] = 32'b11111111111111101111100001000010;
assign LUT_2[58604] = 32'b11111111111111101000001101010101;
assign LUT_2[58605] = 32'b11111111111111100101000101101110;
assign LUT_2[58606] = 32'b11111111111111101111000110010001;
assign LUT_2[58607] = 32'b11111111111111101011111110101010;
assign LUT_2[58608] = 32'b11111111111111101011100010011010;
assign LUT_2[58609] = 32'b11111111111111101000011010110011;
assign LUT_2[58610] = 32'b11111111111111110010011011010110;
assign LUT_2[58611] = 32'b11111111111111101111010011101111;
assign LUT_2[58612] = 32'b11111111111111101000000000000010;
assign LUT_2[58613] = 32'b11111111111111100100111000011011;
assign LUT_2[58614] = 32'b11111111111111101110111000111110;
assign LUT_2[58615] = 32'b11111111111111101011110001010111;
assign LUT_2[58616] = 32'b11111111111111100110010011110111;
assign LUT_2[58617] = 32'b11111111111111100011001100010000;
assign LUT_2[58618] = 32'b11111111111111101101001100110011;
assign LUT_2[58619] = 32'b11111111111111101010000101001100;
assign LUT_2[58620] = 32'b11111111111111100010110001011111;
assign LUT_2[58621] = 32'b11111111111111011111101001111000;
assign LUT_2[58622] = 32'b11111111111111101001101010011011;
assign LUT_2[58623] = 32'b11111111111111100110100010110100;
assign LUT_2[58624] = 32'b11111111111111111000000100011011;
assign LUT_2[58625] = 32'b11111111111111110100111100110100;
assign LUT_2[58626] = 32'b11111111111111111110111101010111;
assign LUT_2[58627] = 32'b11111111111111111011110101110000;
assign LUT_2[58628] = 32'b11111111111111110100100010000011;
assign LUT_2[58629] = 32'b11111111111111110001011010011100;
assign LUT_2[58630] = 32'b11111111111111111011011010111111;
assign LUT_2[58631] = 32'b11111111111111111000010011011000;
assign LUT_2[58632] = 32'b11111111111111110010110101111000;
assign LUT_2[58633] = 32'b11111111111111101111101110010001;
assign LUT_2[58634] = 32'b11111111111111111001101110110100;
assign LUT_2[58635] = 32'b11111111111111110110100111001101;
assign LUT_2[58636] = 32'b11111111111111101111010011100000;
assign LUT_2[58637] = 32'b11111111111111101100001011111001;
assign LUT_2[58638] = 32'b11111111111111110110001100011100;
assign LUT_2[58639] = 32'b11111111111111110011000100110101;
assign LUT_2[58640] = 32'b11111111111111110010101000100101;
assign LUT_2[58641] = 32'b11111111111111101111100000111110;
assign LUT_2[58642] = 32'b11111111111111111001100001100001;
assign LUT_2[58643] = 32'b11111111111111110110011001111010;
assign LUT_2[58644] = 32'b11111111111111101111000110001101;
assign LUT_2[58645] = 32'b11111111111111101011111110100110;
assign LUT_2[58646] = 32'b11111111111111110101111111001001;
assign LUT_2[58647] = 32'b11111111111111110010110111100010;
assign LUT_2[58648] = 32'b11111111111111101101011010000010;
assign LUT_2[58649] = 32'b11111111111111101010010010011011;
assign LUT_2[58650] = 32'b11111111111111110100010010111110;
assign LUT_2[58651] = 32'b11111111111111110001001011010111;
assign LUT_2[58652] = 32'b11111111111111101001110111101010;
assign LUT_2[58653] = 32'b11111111111111100110110000000011;
assign LUT_2[58654] = 32'b11111111111111110000110000100110;
assign LUT_2[58655] = 32'b11111111111111101101101000111111;
assign LUT_2[58656] = 32'b11111111111111111000100000000100;
assign LUT_2[58657] = 32'b11111111111111110101011000011101;
assign LUT_2[58658] = 32'b11111111111111111111011001000000;
assign LUT_2[58659] = 32'b11111111111111111100010001011001;
assign LUT_2[58660] = 32'b11111111111111110100111101101100;
assign LUT_2[58661] = 32'b11111111111111110001110110000101;
assign LUT_2[58662] = 32'b11111111111111111011110110101000;
assign LUT_2[58663] = 32'b11111111111111111000101111000001;
assign LUT_2[58664] = 32'b11111111111111110011010001100001;
assign LUT_2[58665] = 32'b11111111111111110000001001111010;
assign LUT_2[58666] = 32'b11111111111111111010001010011101;
assign LUT_2[58667] = 32'b11111111111111110111000010110110;
assign LUT_2[58668] = 32'b11111111111111101111101111001001;
assign LUT_2[58669] = 32'b11111111111111101100100111100010;
assign LUT_2[58670] = 32'b11111111111111110110101000000101;
assign LUT_2[58671] = 32'b11111111111111110011100000011110;
assign LUT_2[58672] = 32'b11111111111111110011000100001110;
assign LUT_2[58673] = 32'b11111111111111101111111100100111;
assign LUT_2[58674] = 32'b11111111111111111001111101001010;
assign LUT_2[58675] = 32'b11111111111111110110110101100011;
assign LUT_2[58676] = 32'b11111111111111101111100001110110;
assign LUT_2[58677] = 32'b11111111111111101100011010001111;
assign LUT_2[58678] = 32'b11111111111111110110011010110010;
assign LUT_2[58679] = 32'b11111111111111110011010011001011;
assign LUT_2[58680] = 32'b11111111111111101101110101101011;
assign LUT_2[58681] = 32'b11111111111111101010101110000100;
assign LUT_2[58682] = 32'b11111111111111110100101110100111;
assign LUT_2[58683] = 32'b11111111111111110001100111000000;
assign LUT_2[58684] = 32'b11111111111111101010010011010011;
assign LUT_2[58685] = 32'b11111111111111100111001011101100;
assign LUT_2[58686] = 32'b11111111111111110001001100001111;
assign LUT_2[58687] = 32'b11111111111111101110000100101000;
assign LUT_2[58688] = 32'b11111111111111110000001100111110;
assign LUT_2[58689] = 32'b11111111111111101101000101010111;
assign LUT_2[58690] = 32'b11111111111111110111000101111010;
assign LUT_2[58691] = 32'b11111111111111110011111110010011;
assign LUT_2[58692] = 32'b11111111111111101100101010100110;
assign LUT_2[58693] = 32'b11111111111111101001100010111111;
assign LUT_2[58694] = 32'b11111111111111110011100011100010;
assign LUT_2[58695] = 32'b11111111111111110000011011111011;
assign LUT_2[58696] = 32'b11111111111111101010111110011011;
assign LUT_2[58697] = 32'b11111111111111100111110110110100;
assign LUT_2[58698] = 32'b11111111111111110001110111010111;
assign LUT_2[58699] = 32'b11111111111111101110101111110000;
assign LUT_2[58700] = 32'b11111111111111100111011100000011;
assign LUT_2[58701] = 32'b11111111111111100100010100011100;
assign LUT_2[58702] = 32'b11111111111111101110010100111111;
assign LUT_2[58703] = 32'b11111111111111101011001101011000;
assign LUT_2[58704] = 32'b11111111111111101010110001001000;
assign LUT_2[58705] = 32'b11111111111111100111101001100001;
assign LUT_2[58706] = 32'b11111111111111110001101010000100;
assign LUT_2[58707] = 32'b11111111111111101110100010011101;
assign LUT_2[58708] = 32'b11111111111111100111001110110000;
assign LUT_2[58709] = 32'b11111111111111100100000111001001;
assign LUT_2[58710] = 32'b11111111111111101110000111101100;
assign LUT_2[58711] = 32'b11111111111111101011000000000101;
assign LUT_2[58712] = 32'b11111111111111100101100010100101;
assign LUT_2[58713] = 32'b11111111111111100010011010111110;
assign LUT_2[58714] = 32'b11111111111111101100011011100001;
assign LUT_2[58715] = 32'b11111111111111101001010011111010;
assign LUT_2[58716] = 32'b11111111111111100010000000001101;
assign LUT_2[58717] = 32'b11111111111111011110111000100110;
assign LUT_2[58718] = 32'b11111111111111101000111001001001;
assign LUT_2[58719] = 32'b11111111111111100101110001100010;
assign LUT_2[58720] = 32'b11111111111111110000101000100111;
assign LUT_2[58721] = 32'b11111111111111101101100001000000;
assign LUT_2[58722] = 32'b11111111111111110111100001100011;
assign LUT_2[58723] = 32'b11111111111111110100011001111100;
assign LUT_2[58724] = 32'b11111111111111101101000110001111;
assign LUT_2[58725] = 32'b11111111111111101001111110101000;
assign LUT_2[58726] = 32'b11111111111111110011111111001011;
assign LUT_2[58727] = 32'b11111111111111110000110111100100;
assign LUT_2[58728] = 32'b11111111111111101011011010000100;
assign LUT_2[58729] = 32'b11111111111111101000010010011101;
assign LUT_2[58730] = 32'b11111111111111110010010011000000;
assign LUT_2[58731] = 32'b11111111111111101111001011011001;
assign LUT_2[58732] = 32'b11111111111111100111110111101100;
assign LUT_2[58733] = 32'b11111111111111100100110000000101;
assign LUT_2[58734] = 32'b11111111111111101110110000101000;
assign LUT_2[58735] = 32'b11111111111111101011101001000001;
assign LUT_2[58736] = 32'b11111111111111101011001100110001;
assign LUT_2[58737] = 32'b11111111111111101000000101001010;
assign LUT_2[58738] = 32'b11111111111111110010000101101101;
assign LUT_2[58739] = 32'b11111111111111101110111110000110;
assign LUT_2[58740] = 32'b11111111111111100111101010011001;
assign LUT_2[58741] = 32'b11111111111111100100100010110010;
assign LUT_2[58742] = 32'b11111111111111101110100011010101;
assign LUT_2[58743] = 32'b11111111111111101011011011101110;
assign LUT_2[58744] = 32'b11111111111111100101111110001110;
assign LUT_2[58745] = 32'b11111111111111100010110110100111;
assign LUT_2[58746] = 32'b11111111111111101100110111001010;
assign LUT_2[58747] = 32'b11111111111111101001101111100011;
assign LUT_2[58748] = 32'b11111111111111100010011011110110;
assign LUT_2[58749] = 32'b11111111111111011111010100001111;
assign LUT_2[58750] = 32'b11111111111111101001010100110010;
assign LUT_2[58751] = 32'b11111111111111100110001101001011;
assign LUT_2[58752] = 32'b11111111111111111100011000101010;
assign LUT_2[58753] = 32'b11111111111111111001010001000011;
assign LUT_2[58754] = 32'b00000000000000000011010001100110;
assign LUT_2[58755] = 32'b00000000000000000000001001111111;
assign LUT_2[58756] = 32'b11111111111111111000110110010010;
assign LUT_2[58757] = 32'b11111111111111110101101110101011;
assign LUT_2[58758] = 32'b11111111111111111111101111001110;
assign LUT_2[58759] = 32'b11111111111111111100100111100111;
assign LUT_2[58760] = 32'b11111111111111110111001010000111;
assign LUT_2[58761] = 32'b11111111111111110100000010100000;
assign LUT_2[58762] = 32'b11111111111111111110000011000011;
assign LUT_2[58763] = 32'b11111111111111111010111011011100;
assign LUT_2[58764] = 32'b11111111111111110011100111101111;
assign LUT_2[58765] = 32'b11111111111111110000100000001000;
assign LUT_2[58766] = 32'b11111111111111111010100000101011;
assign LUT_2[58767] = 32'b11111111111111110111011001000100;
assign LUT_2[58768] = 32'b11111111111111110110111100110100;
assign LUT_2[58769] = 32'b11111111111111110011110101001101;
assign LUT_2[58770] = 32'b11111111111111111101110101110000;
assign LUT_2[58771] = 32'b11111111111111111010101110001001;
assign LUT_2[58772] = 32'b11111111111111110011011010011100;
assign LUT_2[58773] = 32'b11111111111111110000010010110101;
assign LUT_2[58774] = 32'b11111111111111111010010011011000;
assign LUT_2[58775] = 32'b11111111111111110111001011110001;
assign LUT_2[58776] = 32'b11111111111111110001101110010001;
assign LUT_2[58777] = 32'b11111111111111101110100110101010;
assign LUT_2[58778] = 32'b11111111111111111000100111001101;
assign LUT_2[58779] = 32'b11111111111111110101011111100110;
assign LUT_2[58780] = 32'b11111111111111101110001011111001;
assign LUT_2[58781] = 32'b11111111111111101011000100010010;
assign LUT_2[58782] = 32'b11111111111111110101000100110101;
assign LUT_2[58783] = 32'b11111111111111110001111101001110;
assign LUT_2[58784] = 32'b11111111111111111100110100010011;
assign LUT_2[58785] = 32'b11111111111111111001101100101100;
assign LUT_2[58786] = 32'b00000000000000000011101101001111;
assign LUT_2[58787] = 32'b00000000000000000000100101101000;
assign LUT_2[58788] = 32'b11111111111111111001010001111011;
assign LUT_2[58789] = 32'b11111111111111110110001010010100;
assign LUT_2[58790] = 32'b00000000000000000000001010110111;
assign LUT_2[58791] = 32'b11111111111111111101000011010000;
assign LUT_2[58792] = 32'b11111111111111110111100101110000;
assign LUT_2[58793] = 32'b11111111111111110100011110001001;
assign LUT_2[58794] = 32'b11111111111111111110011110101100;
assign LUT_2[58795] = 32'b11111111111111111011010111000101;
assign LUT_2[58796] = 32'b11111111111111110100000011011000;
assign LUT_2[58797] = 32'b11111111111111110000111011110001;
assign LUT_2[58798] = 32'b11111111111111111010111100010100;
assign LUT_2[58799] = 32'b11111111111111110111110100101101;
assign LUT_2[58800] = 32'b11111111111111110111011000011101;
assign LUT_2[58801] = 32'b11111111111111110100010000110110;
assign LUT_2[58802] = 32'b11111111111111111110010001011001;
assign LUT_2[58803] = 32'b11111111111111111011001001110010;
assign LUT_2[58804] = 32'b11111111111111110011110110000101;
assign LUT_2[58805] = 32'b11111111111111110000101110011110;
assign LUT_2[58806] = 32'b11111111111111111010101111000001;
assign LUT_2[58807] = 32'b11111111111111110111100111011010;
assign LUT_2[58808] = 32'b11111111111111110010001001111010;
assign LUT_2[58809] = 32'b11111111111111101111000010010011;
assign LUT_2[58810] = 32'b11111111111111111001000010110110;
assign LUT_2[58811] = 32'b11111111111111110101111011001111;
assign LUT_2[58812] = 32'b11111111111111101110100111100010;
assign LUT_2[58813] = 32'b11111111111111101011011111111011;
assign LUT_2[58814] = 32'b11111111111111110101100000011110;
assign LUT_2[58815] = 32'b11111111111111110010011000110111;
assign LUT_2[58816] = 32'b11111111111111110100100001001101;
assign LUT_2[58817] = 32'b11111111111111110001011001100110;
assign LUT_2[58818] = 32'b11111111111111111011011010001001;
assign LUT_2[58819] = 32'b11111111111111111000010010100010;
assign LUT_2[58820] = 32'b11111111111111110000111110110101;
assign LUT_2[58821] = 32'b11111111111111101101110111001110;
assign LUT_2[58822] = 32'b11111111111111110111110111110001;
assign LUT_2[58823] = 32'b11111111111111110100110000001010;
assign LUT_2[58824] = 32'b11111111111111101111010010101010;
assign LUT_2[58825] = 32'b11111111111111101100001011000011;
assign LUT_2[58826] = 32'b11111111111111110110001011100110;
assign LUT_2[58827] = 32'b11111111111111110011000011111111;
assign LUT_2[58828] = 32'b11111111111111101011110000010010;
assign LUT_2[58829] = 32'b11111111111111101000101000101011;
assign LUT_2[58830] = 32'b11111111111111110010101001001110;
assign LUT_2[58831] = 32'b11111111111111101111100001100111;
assign LUT_2[58832] = 32'b11111111111111101111000101010111;
assign LUT_2[58833] = 32'b11111111111111101011111101110000;
assign LUT_2[58834] = 32'b11111111111111110101111110010011;
assign LUT_2[58835] = 32'b11111111111111110010110110101100;
assign LUT_2[58836] = 32'b11111111111111101011100010111111;
assign LUT_2[58837] = 32'b11111111111111101000011011011000;
assign LUT_2[58838] = 32'b11111111111111110010011011111011;
assign LUT_2[58839] = 32'b11111111111111101111010100010100;
assign LUT_2[58840] = 32'b11111111111111101001110110110100;
assign LUT_2[58841] = 32'b11111111111111100110101111001101;
assign LUT_2[58842] = 32'b11111111111111110000101111110000;
assign LUT_2[58843] = 32'b11111111111111101101101000001001;
assign LUT_2[58844] = 32'b11111111111111100110010100011100;
assign LUT_2[58845] = 32'b11111111111111100011001100110101;
assign LUT_2[58846] = 32'b11111111111111101101001101011000;
assign LUT_2[58847] = 32'b11111111111111101010000101110001;
assign LUT_2[58848] = 32'b11111111111111110100111100110110;
assign LUT_2[58849] = 32'b11111111111111110001110101001111;
assign LUT_2[58850] = 32'b11111111111111111011110101110010;
assign LUT_2[58851] = 32'b11111111111111111000101110001011;
assign LUT_2[58852] = 32'b11111111111111110001011010011110;
assign LUT_2[58853] = 32'b11111111111111101110010010110111;
assign LUT_2[58854] = 32'b11111111111111111000010011011010;
assign LUT_2[58855] = 32'b11111111111111110101001011110011;
assign LUT_2[58856] = 32'b11111111111111101111101110010011;
assign LUT_2[58857] = 32'b11111111111111101100100110101100;
assign LUT_2[58858] = 32'b11111111111111110110100111001111;
assign LUT_2[58859] = 32'b11111111111111110011011111101000;
assign LUT_2[58860] = 32'b11111111111111101100001011111011;
assign LUT_2[58861] = 32'b11111111111111101001000100010100;
assign LUT_2[58862] = 32'b11111111111111110011000100110111;
assign LUT_2[58863] = 32'b11111111111111101111111101010000;
assign LUT_2[58864] = 32'b11111111111111101111100001000000;
assign LUT_2[58865] = 32'b11111111111111101100011001011001;
assign LUT_2[58866] = 32'b11111111111111110110011001111100;
assign LUT_2[58867] = 32'b11111111111111110011010010010101;
assign LUT_2[58868] = 32'b11111111111111101011111110101000;
assign LUT_2[58869] = 32'b11111111111111101000110111000001;
assign LUT_2[58870] = 32'b11111111111111110010110111100100;
assign LUT_2[58871] = 32'b11111111111111101111101111111101;
assign LUT_2[58872] = 32'b11111111111111101010010010011101;
assign LUT_2[58873] = 32'b11111111111111100111001010110110;
assign LUT_2[58874] = 32'b11111111111111110001001011011001;
assign LUT_2[58875] = 32'b11111111111111101110000011110010;
assign LUT_2[58876] = 32'b11111111111111100110110000000101;
assign LUT_2[58877] = 32'b11111111111111100011101000011110;
assign LUT_2[58878] = 32'b11111111111111101101101001000001;
assign LUT_2[58879] = 32'b11111111111111101010100001011010;
assign LUT_2[58880] = 32'b11111111111111111000110111100111;
assign LUT_2[58881] = 32'b11111111111111110101110000000000;
assign LUT_2[58882] = 32'b11111111111111111111110000100011;
assign LUT_2[58883] = 32'b11111111111111111100101000111100;
assign LUT_2[58884] = 32'b11111111111111110101010101001111;
assign LUT_2[58885] = 32'b11111111111111110010001101101000;
assign LUT_2[58886] = 32'b11111111111111111100001110001011;
assign LUT_2[58887] = 32'b11111111111111111001000110100100;
assign LUT_2[58888] = 32'b11111111111111110011101001000100;
assign LUT_2[58889] = 32'b11111111111111110000100001011101;
assign LUT_2[58890] = 32'b11111111111111111010100010000000;
assign LUT_2[58891] = 32'b11111111111111110111011010011001;
assign LUT_2[58892] = 32'b11111111111111110000000110101100;
assign LUT_2[58893] = 32'b11111111111111101100111111000101;
assign LUT_2[58894] = 32'b11111111111111110110111111101000;
assign LUT_2[58895] = 32'b11111111111111110011111000000001;
assign LUT_2[58896] = 32'b11111111111111110011011011110001;
assign LUT_2[58897] = 32'b11111111111111110000010100001010;
assign LUT_2[58898] = 32'b11111111111111111010010100101101;
assign LUT_2[58899] = 32'b11111111111111110111001101000110;
assign LUT_2[58900] = 32'b11111111111111101111111001011001;
assign LUT_2[58901] = 32'b11111111111111101100110001110010;
assign LUT_2[58902] = 32'b11111111111111110110110010010101;
assign LUT_2[58903] = 32'b11111111111111110011101010101110;
assign LUT_2[58904] = 32'b11111111111111101110001101001110;
assign LUT_2[58905] = 32'b11111111111111101011000101100111;
assign LUT_2[58906] = 32'b11111111111111110101000110001010;
assign LUT_2[58907] = 32'b11111111111111110001111110100011;
assign LUT_2[58908] = 32'b11111111111111101010101010110110;
assign LUT_2[58909] = 32'b11111111111111100111100011001111;
assign LUT_2[58910] = 32'b11111111111111110001100011110010;
assign LUT_2[58911] = 32'b11111111111111101110011100001011;
assign LUT_2[58912] = 32'b11111111111111111001010011010000;
assign LUT_2[58913] = 32'b11111111111111110110001011101001;
assign LUT_2[58914] = 32'b00000000000000000000001100001100;
assign LUT_2[58915] = 32'b11111111111111111101000100100101;
assign LUT_2[58916] = 32'b11111111111111110101110000111000;
assign LUT_2[58917] = 32'b11111111111111110010101001010001;
assign LUT_2[58918] = 32'b11111111111111111100101001110100;
assign LUT_2[58919] = 32'b11111111111111111001100010001101;
assign LUT_2[58920] = 32'b11111111111111110100000100101101;
assign LUT_2[58921] = 32'b11111111111111110000111101000110;
assign LUT_2[58922] = 32'b11111111111111111010111101101001;
assign LUT_2[58923] = 32'b11111111111111110111110110000010;
assign LUT_2[58924] = 32'b11111111111111110000100010010101;
assign LUT_2[58925] = 32'b11111111111111101101011010101110;
assign LUT_2[58926] = 32'b11111111111111110111011011010001;
assign LUT_2[58927] = 32'b11111111111111110100010011101010;
assign LUT_2[58928] = 32'b11111111111111110011110111011010;
assign LUT_2[58929] = 32'b11111111111111110000101111110011;
assign LUT_2[58930] = 32'b11111111111111111010110000010110;
assign LUT_2[58931] = 32'b11111111111111110111101000101111;
assign LUT_2[58932] = 32'b11111111111111110000010101000010;
assign LUT_2[58933] = 32'b11111111111111101101001101011011;
assign LUT_2[58934] = 32'b11111111111111110111001101111110;
assign LUT_2[58935] = 32'b11111111111111110100000110010111;
assign LUT_2[58936] = 32'b11111111111111101110101000110111;
assign LUT_2[58937] = 32'b11111111111111101011100001010000;
assign LUT_2[58938] = 32'b11111111111111110101100001110011;
assign LUT_2[58939] = 32'b11111111111111110010011010001100;
assign LUT_2[58940] = 32'b11111111111111101011000110011111;
assign LUT_2[58941] = 32'b11111111111111100111111110111000;
assign LUT_2[58942] = 32'b11111111111111110001111111011011;
assign LUT_2[58943] = 32'b11111111111111101110110111110100;
assign LUT_2[58944] = 32'b11111111111111110001000000001010;
assign LUT_2[58945] = 32'b11111111111111101101111000100011;
assign LUT_2[58946] = 32'b11111111111111110111111001000110;
assign LUT_2[58947] = 32'b11111111111111110100110001011111;
assign LUT_2[58948] = 32'b11111111111111101101011101110010;
assign LUT_2[58949] = 32'b11111111111111101010010110001011;
assign LUT_2[58950] = 32'b11111111111111110100010110101110;
assign LUT_2[58951] = 32'b11111111111111110001001111000111;
assign LUT_2[58952] = 32'b11111111111111101011110001100111;
assign LUT_2[58953] = 32'b11111111111111101000101010000000;
assign LUT_2[58954] = 32'b11111111111111110010101010100011;
assign LUT_2[58955] = 32'b11111111111111101111100010111100;
assign LUT_2[58956] = 32'b11111111111111101000001111001111;
assign LUT_2[58957] = 32'b11111111111111100101000111101000;
assign LUT_2[58958] = 32'b11111111111111101111001000001011;
assign LUT_2[58959] = 32'b11111111111111101100000000100100;
assign LUT_2[58960] = 32'b11111111111111101011100100010100;
assign LUT_2[58961] = 32'b11111111111111101000011100101101;
assign LUT_2[58962] = 32'b11111111111111110010011101010000;
assign LUT_2[58963] = 32'b11111111111111101111010101101001;
assign LUT_2[58964] = 32'b11111111111111101000000001111100;
assign LUT_2[58965] = 32'b11111111111111100100111010010101;
assign LUT_2[58966] = 32'b11111111111111101110111010111000;
assign LUT_2[58967] = 32'b11111111111111101011110011010001;
assign LUT_2[58968] = 32'b11111111111111100110010101110001;
assign LUT_2[58969] = 32'b11111111111111100011001110001010;
assign LUT_2[58970] = 32'b11111111111111101101001110101101;
assign LUT_2[58971] = 32'b11111111111111101010000111000110;
assign LUT_2[58972] = 32'b11111111111111100010110011011001;
assign LUT_2[58973] = 32'b11111111111111011111101011110010;
assign LUT_2[58974] = 32'b11111111111111101001101100010101;
assign LUT_2[58975] = 32'b11111111111111100110100100101110;
assign LUT_2[58976] = 32'b11111111111111110001011011110011;
assign LUT_2[58977] = 32'b11111111111111101110010100001100;
assign LUT_2[58978] = 32'b11111111111111111000010100101111;
assign LUT_2[58979] = 32'b11111111111111110101001101001000;
assign LUT_2[58980] = 32'b11111111111111101101111001011011;
assign LUT_2[58981] = 32'b11111111111111101010110001110100;
assign LUT_2[58982] = 32'b11111111111111110100110010010111;
assign LUT_2[58983] = 32'b11111111111111110001101010110000;
assign LUT_2[58984] = 32'b11111111111111101100001101010000;
assign LUT_2[58985] = 32'b11111111111111101001000101101001;
assign LUT_2[58986] = 32'b11111111111111110011000110001100;
assign LUT_2[58987] = 32'b11111111111111101111111110100101;
assign LUT_2[58988] = 32'b11111111111111101000101010111000;
assign LUT_2[58989] = 32'b11111111111111100101100011010001;
assign LUT_2[58990] = 32'b11111111111111101111100011110100;
assign LUT_2[58991] = 32'b11111111111111101100011100001101;
assign LUT_2[58992] = 32'b11111111111111101011111111111101;
assign LUT_2[58993] = 32'b11111111111111101000111000010110;
assign LUT_2[58994] = 32'b11111111111111110010111000111001;
assign LUT_2[58995] = 32'b11111111111111101111110001010010;
assign LUT_2[58996] = 32'b11111111111111101000011101100101;
assign LUT_2[58997] = 32'b11111111111111100101010101111110;
assign LUT_2[58998] = 32'b11111111111111101111010110100001;
assign LUT_2[58999] = 32'b11111111111111101100001110111010;
assign LUT_2[59000] = 32'b11111111111111100110110001011010;
assign LUT_2[59001] = 32'b11111111111111100011101001110011;
assign LUT_2[59002] = 32'b11111111111111101101101010010110;
assign LUT_2[59003] = 32'b11111111111111101010100010101111;
assign LUT_2[59004] = 32'b11111111111111100011001111000010;
assign LUT_2[59005] = 32'b11111111111111100000000111011011;
assign LUT_2[59006] = 32'b11111111111111101010000111111110;
assign LUT_2[59007] = 32'b11111111111111100111000000010111;
assign LUT_2[59008] = 32'b11111111111111111101001011110110;
assign LUT_2[59009] = 32'b11111111111111111010000100001111;
assign LUT_2[59010] = 32'b00000000000000000100000100110010;
assign LUT_2[59011] = 32'b00000000000000000000111101001011;
assign LUT_2[59012] = 32'b11111111111111111001101001011110;
assign LUT_2[59013] = 32'b11111111111111110110100001110111;
assign LUT_2[59014] = 32'b00000000000000000000100010011010;
assign LUT_2[59015] = 32'b11111111111111111101011010110011;
assign LUT_2[59016] = 32'b11111111111111110111111101010011;
assign LUT_2[59017] = 32'b11111111111111110100110101101100;
assign LUT_2[59018] = 32'b11111111111111111110110110001111;
assign LUT_2[59019] = 32'b11111111111111111011101110101000;
assign LUT_2[59020] = 32'b11111111111111110100011010111011;
assign LUT_2[59021] = 32'b11111111111111110001010011010100;
assign LUT_2[59022] = 32'b11111111111111111011010011110111;
assign LUT_2[59023] = 32'b11111111111111111000001100010000;
assign LUT_2[59024] = 32'b11111111111111110111110000000000;
assign LUT_2[59025] = 32'b11111111111111110100101000011001;
assign LUT_2[59026] = 32'b11111111111111111110101000111100;
assign LUT_2[59027] = 32'b11111111111111111011100001010101;
assign LUT_2[59028] = 32'b11111111111111110100001101101000;
assign LUT_2[59029] = 32'b11111111111111110001000110000001;
assign LUT_2[59030] = 32'b11111111111111111011000110100100;
assign LUT_2[59031] = 32'b11111111111111110111111110111101;
assign LUT_2[59032] = 32'b11111111111111110010100001011101;
assign LUT_2[59033] = 32'b11111111111111101111011001110110;
assign LUT_2[59034] = 32'b11111111111111111001011010011001;
assign LUT_2[59035] = 32'b11111111111111110110010010110010;
assign LUT_2[59036] = 32'b11111111111111101110111111000101;
assign LUT_2[59037] = 32'b11111111111111101011110111011110;
assign LUT_2[59038] = 32'b11111111111111110101111000000001;
assign LUT_2[59039] = 32'b11111111111111110010110000011010;
assign LUT_2[59040] = 32'b11111111111111111101100111011111;
assign LUT_2[59041] = 32'b11111111111111111010011111111000;
assign LUT_2[59042] = 32'b00000000000000000100100000011011;
assign LUT_2[59043] = 32'b00000000000000000001011000110100;
assign LUT_2[59044] = 32'b11111111111111111010000101000111;
assign LUT_2[59045] = 32'b11111111111111110110111101100000;
assign LUT_2[59046] = 32'b00000000000000000000111110000011;
assign LUT_2[59047] = 32'b11111111111111111101110110011100;
assign LUT_2[59048] = 32'b11111111111111111000011000111100;
assign LUT_2[59049] = 32'b11111111111111110101010001010101;
assign LUT_2[59050] = 32'b11111111111111111111010001111000;
assign LUT_2[59051] = 32'b11111111111111111100001010010001;
assign LUT_2[59052] = 32'b11111111111111110100110110100100;
assign LUT_2[59053] = 32'b11111111111111110001101110111101;
assign LUT_2[59054] = 32'b11111111111111111011101111100000;
assign LUT_2[59055] = 32'b11111111111111111000100111111001;
assign LUT_2[59056] = 32'b11111111111111111000001011101001;
assign LUT_2[59057] = 32'b11111111111111110101000100000010;
assign LUT_2[59058] = 32'b11111111111111111111000100100101;
assign LUT_2[59059] = 32'b11111111111111111011111100111110;
assign LUT_2[59060] = 32'b11111111111111110100101001010001;
assign LUT_2[59061] = 32'b11111111111111110001100001101010;
assign LUT_2[59062] = 32'b11111111111111111011100010001101;
assign LUT_2[59063] = 32'b11111111111111111000011010100110;
assign LUT_2[59064] = 32'b11111111111111110010111101000110;
assign LUT_2[59065] = 32'b11111111111111101111110101011111;
assign LUT_2[59066] = 32'b11111111111111111001110110000010;
assign LUT_2[59067] = 32'b11111111111111110110101110011011;
assign LUT_2[59068] = 32'b11111111111111101111011010101110;
assign LUT_2[59069] = 32'b11111111111111101100010011000111;
assign LUT_2[59070] = 32'b11111111111111110110010011101010;
assign LUT_2[59071] = 32'b11111111111111110011001100000011;
assign LUT_2[59072] = 32'b11111111111111110101010100011001;
assign LUT_2[59073] = 32'b11111111111111110010001100110010;
assign LUT_2[59074] = 32'b11111111111111111100001101010101;
assign LUT_2[59075] = 32'b11111111111111111001000101101110;
assign LUT_2[59076] = 32'b11111111111111110001110010000001;
assign LUT_2[59077] = 32'b11111111111111101110101010011010;
assign LUT_2[59078] = 32'b11111111111111111000101010111101;
assign LUT_2[59079] = 32'b11111111111111110101100011010110;
assign LUT_2[59080] = 32'b11111111111111110000000101110110;
assign LUT_2[59081] = 32'b11111111111111101100111110001111;
assign LUT_2[59082] = 32'b11111111111111110110111110110010;
assign LUT_2[59083] = 32'b11111111111111110011110111001011;
assign LUT_2[59084] = 32'b11111111111111101100100011011110;
assign LUT_2[59085] = 32'b11111111111111101001011011110111;
assign LUT_2[59086] = 32'b11111111111111110011011100011010;
assign LUT_2[59087] = 32'b11111111111111110000010100110011;
assign LUT_2[59088] = 32'b11111111111111101111111000100011;
assign LUT_2[59089] = 32'b11111111111111101100110000111100;
assign LUT_2[59090] = 32'b11111111111111110110110001011111;
assign LUT_2[59091] = 32'b11111111111111110011101001111000;
assign LUT_2[59092] = 32'b11111111111111101100010110001011;
assign LUT_2[59093] = 32'b11111111111111101001001110100100;
assign LUT_2[59094] = 32'b11111111111111110011001111000111;
assign LUT_2[59095] = 32'b11111111111111110000000111100000;
assign LUT_2[59096] = 32'b11111111111111101010101010000000;
assign LUT_2[59097] = 32'b11111111111111100111100010011001;
assign LUT_2[59098] = 32'b11111111111111110001100010111100;
assign LUT_2[59099] = 32'b11111111111111101110011011010101;
assign LUT_2[59100] = 32'b11111111111111100111000111101000;
assign LUT_2[59101] = 32'b11111111111111100100000000000001;
assign LUT_2[59102] = 32'b11111111111111101110000000100100;
assign LUT_2[59103] = 32'b11111111111111101010111000111101;
assign LUT_2[59104] = 32'b11111111111111110101110000000010;
assign LUT_2[59105] = 32'b11111111111111110010101000011011;
assign LUT_2[59106] = 32'b11111111111111111100101000111110;
assign LUT_2[59107] = 32'b11111111111111111001100001010111;
assign LUT_2[59108] = 32'b11111111111111110010001101101010;
assign LUT_2[59109] = 32'b11111111111111101111000110000011;
assign LUT_2[59110] = 32'b11111111111111111001000110100110;
assign LUT_2[59111] = 32'b11111111111111110101111110111111;
assign LUT_2[59112] = 32'b11111111111111110000100001011111;
assign LUT_2[59113] = 32'b11111111111111101101011001111000;
assign LUT_2[59114] = 32'b11111111111111110111011010011011;
assign LUT_2[59115] = 32'b11111111111111110100010010110100;
assign LUT_2[59116] = 32'b11111111111111101100111111000111;
assign LUT_2[59117] = 32'b11111111111111101001110111100000;
assign LUT_2[59118] = 32'b11111111111111110011111000000011;
assign LUT_2[59119] = 32'b11111111111111110000110000011100;
assign LUT_2[59120] = 32'b11111111111111110000010100001100;
assign LUT_2[59121] = 32'b11111111111111101101001100100101;
assign LUT_2[59122] = 32'b11111111111111110111001101001000;
assign LUT_2[59123] = 32'b11111111111111110100000101100001;
assign LUT_2[59124] = 32'b11111111111111101100110001110100;
assign LUT_2[59125] = 32'b11111111111111101001101010001101;
assign LUT_2[59126] = 32'b11111111111111110011101010110000;
assign LUT_2[59127] = 32'b11111111111111110000100011001001;
assign LUT_2[59128] = 32'b11111111111111101011000101101001;
assign LUT_2[59129] = 32'b11111111111111100111111110000010;
assign LUT_2[59130] = 32'b11111111111111110001111110100101;
assign LUT_2[59131] = 32'b11111111111111101110110110111110;
assign LUT_2[59132] = 32'b11111111111111100111100011010001;
assign LUT_2[59133] = 32'b11111111111111100100011011101010;
assign LUT_2[59134] = 32'b11111111111111101110011100001101;
assign LUT_2[59135] = 32'b11111111111111101011010100100110;
assign LUT_2[59136] = 32'b11111111111111111100110110001101;
assign LUT_2[59137] = 32'b11111111111111111001101110100110;
assign LUT_2[59138] = 32'b00000000000000000011101111001001;
assign LUT_2[59139] = 32'b00000000000000000000100111100010;
assign LUT_2[59140] = 32'b11111111111111111001010011110101;
assign LUT_2[59141] = 32'b11111111111111110110001100001110;
assign LUT_2[59142] = 32'b00000000000000000000001100110001;
assign LUT_2[59143] = 32'b11111111111111111101000101001010;
assign LUT_2[59144] = 32'b11111111111111110111100111101010;
assign LUT_2[59145] = 32'b11111111111111110100100000000011;
assign LUT_2[59146] = 32'b11111111111111111110100000100110;
assign LUT_2[59147] = 32'b11111111111111111011011000111111;
assign LUT_2[59148] = 32'b11111111111111110100000101010010;
assign LUT_2[59149] = 32'b11111111111111110000111101101011;
assign LUT_2[59150] = 32'b11111111111111111010111110001110;
assign LUT_2[59151] = 32'b11111111111111110111110110100111;
assign LUT_2[59152] = 32'b11111111111111110111011010010111;
assign LUT_2[59153] = 32'b11111111111111110100010010110000;
assign LUT_2[59154] = 32'b11111111111111111110010011010011;
assign LUT_2[59155] = 32'b11111111111111111011001011101100;
assign LUT_2[59156] = 32'b11111111111111110011110111111111;
assign LUT_2[59157] = 32'b11111111111111110000110000011000;
assign LUT_2[59158] = 32'b11111111111111111010110000111011;
assign LUT_2[59159] = 32'b11111111111111110111101001010100;
assign LUT_2[59160] = 32'b11111111111111110010001011110100;
assign LUT_2[59161] = 32'b11111111111111101111000100001101;
assign LUT_2[59162] = 32'b11111111111111111001000100110000;
assign LUT_2[59163] = 32'b11111111111111110101111101001001;
assign LUT_2[59164] = 32'b11111111111111101110101001011100;
assign LUT_2[59165] = 32'b11111111111111101011100001110101;
assign LUT_2[59166] = 32'b11111111111111110101100010011000;
assign LUT_2[59167] = 32'b11111111111111110010011010110001;
assign LUT_2[59168] = 32'b11111111111111111101010001110110;
assign LUT_2[59169] = 32'b11111111111111111010001010001111;
assign LUT_2[59170] = 32'b00000000000000000100001010110010;
assign LUT_2[59171] = 32'b00000000000000000001000011001011;
assign LUT_2[59172] = 32'b11111111111111111001101111011110;
assign LUT_2[59173] = 32'b11111111111111110110100111110111;
assign LUT_2[59174] = 32'b00000000000000000000101000011010;
assign LUT_2[59175] = 32'b11111111111111111101100000110011;
assign LUT_2[59176] = 32'b11111111111111111000000011010011;
assign LUT_2[59177] = 32'b11111111111111110100111011101100;
assign LUT_2[59178] = 32'b11111111111111111110111100001111;
assign LUT_2[59179] = 32'b11111111111111111011110100101000;
assign LUT_2[59180] = 32'b11111111111111110100100000111011;
assign LUT_2[59181] = 32'b11111111111111110001011001010100;
assign LUT_2[59182] = 32'b11111111111111111011011001110111;
assign LUT_2[59183] = 32'b11111111111111111000010010010000;
assign LUT_2[59184] = 32'b11111111111111110111110110000000;
assign LUT_2[59185] = 32'b11111111111111110100101110011001;
assign LUT_2[59186] = 32'b11111111111111111110101110111100;
assign LUT_2[59187] = 32'b11111111111111111011100111010101;
assign LUT_2[59188] = 32'b11111111111111110100010011101000;
assign LUT_2[59189] = 32'b11111111111111110001001100000001;
assign LUT_2[59190] = 32'b11111111111111111011001100100100;
assign LUT_2[59191] = 32'b11111111111111111000000100111101;
assign LUT_2[59192] = 32'b11111111111111110010100111011101;
assign LUT_2[59193] = 32'b11111111111111101111011111110110;
assign LUT_2[59194] = 32'b11111111111111111001100000011001;
assign LUT_2[59195] = 32'b11111111111111110110011000110010;
assign LUT_2[59196] = 32'b11111111111111101111000101000101;
assign LUT_2[59197] = 32'b11111111111111101011111101011110;
assign LUT_2[59198] = 32'b11111111111111110101111110000001;
assign LUT_2[59199] = 32'b11111111111111110010110110011010;
assign LUT_2[59200] = 32'b11111111111111110100111110110000;
assign LUT_2[59201] = 32'b11111111111111110001110111001001;
assign LUT_2[59202] = 32'b11111111111111111011110111101100;
assign LUT_2[59203] = 32'b11111111111111111000110000000101;
assign LUT_2[59204] = 32'b11111111111111110001011100011000;
assign LUT_2[59205] = 32'b11111111111111101110010100110001;
assign LUT_2[59206] = 32'b11111111111111111000010101010100;
assign LUT_2[59207] = 32'b11111111111111110101001101101101;
assign LUT_2[59208] = 32'b11111111111111101111110000001101;
assign LUT_2[59209] = 32'b11111111111111101100101000100110;
assign LUT_2[59210] = 32'b11111111111111110110101001001001;
assign LUT_2[59211] = 32'b11111111111111110011100001100010;
assign LUT_2[59212] = 32'b11111111111111101100001101110101;
assign LUT_2[59213] = 32'b11111111111111101001000110001110;
assign LUT_2[59214] = 32'b11111111111111110011000110110001;
assign LUT_2[59215] = 32'b11111111111111101111111111001010;
assign LUT_2[59216] = 32'b11111111111111101111100010111010;
assign LUT_2[59217] = 32'b11111111111111101100011011010011;
assign LUT_2[59218] = 32'b11111111111111110110011011110110;
assign LUT_2[59219] = 32'b11111111111111110011010100001111;
assign LUT_2[59220] = 32'b11111111111111101100000000100010;
assign LUT_2[59221] = 32'b11111111111111101000111000111011;
assign LUT_2[59222] = 32'b11111111111111110010111001011110;
assign LUT_2[59223] = 32'b11111111111111101111110001110111;
assign LUT_2[59224] = 32'b11111111111111101010010100010111;
assign LUT_2[59225] = 32'b11111111111111100111001100110000;
assign LUT_2[59226] = 32'b11111111111111110001001101010011;
assign LUT_2[59227] = 32'b11111111111111101110000101101100;
assign LUT_2[59228] = 32'b11111111111111100110110001111111;
assign LUT_2[59229] = 32'b11111111111111100011101010011000;
assign LUT_2[59230] = 32'b11111111111111101101101010111011;
assign LUT_2[59231] = 32'b11111111111111101010100011010100;
assign LUT_2[59232] = 32'b11111111111111110101011010011001;
assign LUT_2[59233] = 32'b11111111111111110010010010110010;
assign LUT_2[59234] = 32'b11111111111111111100010011010101;
assign LUT_2[59235] = 32'b11111111111111111001001011101110;
assign LUT_2[59236] = 32'b11111111111111110001111000000001;
assign LUT_2[59237] = 32'b11111111111111101110110000011010;
assign LUT_2[59238] = 32'b11111111111111111000110000111101;
assign LUT_2[59239] = 32'b11111111111111110101101001010110;
assign LUT_2[59240] = 32'b11111111111111110000001011110110;
assign LUT_2[59241] = 32'b11111111111111101101000100001111;
assign LUT_2[59242] = 32'b11111111111111110111000100110010;
assign LUT_2[59243] = 32'b11111111111111110011111101001011;
assign LUT_2[59244] = 32'b11111111111111101100101001011110;
assign LUT_2[59245] = 32'b11111111111111101001100001110111;
assign LUT_2[59246] = 32'b11111111111111110011100010011010;
assign LUT_2[59247] = 32'b11111111111111110000011010110011;
assign LUT_2[59248] = 32'b11111111111111101111111110100011;
assign LUT_2[59249] = 32'b11111111111111101100110110111100;
assign LUT_2[59250] = 32'b11111111111111110110110111011111;
assign LUT_2[59251] = 32'b11111111111111110011101111111000;
assign LUT_2[59252] = 32'b11111111111111101100011100001011;
assign LUT_2[59253] = 32'b11111111111111101001010100100100;
assign LUT_2[59254] = 32'b11111111111111110011010101000111;
assign LUT_2[59255] = 32'b11111111111111110000001101100000;
assign LUT_2[59256] = 32'b11111111111111101010110000000000;
assign LUT_2[59257] = 32'b11111111111111100111101000011001;
assign LUT_2[59258] = 32'b11111111111111110001101000111100;
assign LUT_2[59259] = 32'b11111111111111101110100001010101;
assign LUT_2[59260] = 32'b11111111111111100111001101101000;
assign LUT_2[59261] = 32'b11111111111111100100000110000001;
assign LUT_2[59262] = 32'b11111111111111101110000110100100;
assign LUT_2[59263] = 32'b11111111111111101010111110111101;
assign LUT_2[59264] = 32'b00000000000000000001001010011100;
assign LUT_2[59265] = 32'b11111111111111111110000010110101;
assign LUT_2[59266] = 32'b00000000000000001000000011011000;
assign LUT_2[59267] = 32'b00000000000000000100111011110001;
assign LUT_2[59268] = 32'b11111111111111111101101000000100;
assign LUT_2[59269] = 32'b11111111111111111010100000011101;
assign LUT_2[59270] = 32'b00000000000000000100100001000000;
assign LUT_2[59271] = 32'b00000000000000000001011001011001;
assign LUT_2[59272] = 32'b11111111111111111011111011111001;
assign LUT_2[59273] = 32'b11111111111111111000110100010010;
assign LUT_2[59274] = 32'b00000000000000000010110100110101;
assign LUT_2[59275] = 32'b11111111111111111111101101001110;
assign LUT_2[59276] = 32'b11111111111111111000011001100001;
assign LUT_2[59277] = 32'b11111111111111110101010001111010;
assign LUT_2[59278] = 32'b11111111111111111111010010011101;
assign LUT_2[59279] = 32'b11111111111111111100001010110110;
assign LUT_2[59280] = 32'b11111111111111111011101110100110;
assign LUT_2[59281] = 32'b11111111111111111000100110111111;
assign LUT_2[59282] = 32'b00000000000000000010100111100010;
assign LUT_2[59283] = 32'b11111111111111111111011111111011;
assign LUT_2[59284] = 32'b11111111111111111000001100001110;
assign LUT_2[59285] = 32'b11111111111111110101000100100111;
assign LUT_2[59286] = 32'b11111111111111111111000101001010;
assign LUT_2[59287] = 32'b11111111111111111011111101100011;
assign LUT_2[59288] = 32'b11111111111111110110100000000011;
assign LUT_2[59289] = 32'b11111111111111110011011000011100;
assign LUT_2[59290] = 32'b11111111111111111101011000111111;
assign LUT_2[59291] = 32'b11111111111111111010010001011000;
assign LUT_2[59292] = 32'b11111111111111110010111101101011;
assign LUT_2[59293] = 32'b11111111111111101111110110000100;
assign LUT_2[59294] = 32'b11111111111111111001110110100111;
assign LUT_2[59295] = 32'b11111111111111110110101111000000;
assign LUT_2[59296] = 32'b00000000000000000001100110000101;
assign LUT_2[59297] = 32'b11111111111111111110011110011110;
assign LUT_2[59298] = 32'b00000000000000001000011111000001;
assign LUT_2[59299] = 32'b00000000000000000101010111011010;
assign LUT_2[59300] = 32'b11111111111111111110000011101101;
assign LUT_2[59301] = 32'b11111111111111111010111100000110;
assign LUT_2[59302] = 32'b00000000000000000100111100101001;
assign LUT_2[59303] = 32'b00000000000000000001110101000010;
assign LUT_2[59304] = 32'b11111111111111111100010111100010;
assign LUT_2[59305] = 32'b11111111111111111001001111111011;
assign LUT_2[59306] = 32'b00000000000000000011010000011110;
assign LUT_2[59307] = 32'b00000000000000000000001000110111;
assign LUT_2[59308] = 32'b11111111111111111000110101001010;
assign LUT_2[59309] = 32'b11111111111111110101101101100011;
assign LUT_2[59310] = 32'b11111111111111111111101110000110;
assign LUT_2[59311] = 32'b11111111111111111100100110011111;
assign LUT_2[59312] = 32'b11111111111111111100001010001111;
assign LUT_2[59313] = 32'b11111111111111111001000010101000;
assign LUT_2[59314] = 32'b00000000000000000011000011001011;
assign LUT_2[59315] = 32'b11111111111111111111111011100100;
assign LUT_2[59316] = 32'b11111111111111111000100111110111;
assign LUT_2[59317] = 32'b11111111111111110101100000010000;
assign LUT_2[59318] = 32'b11111111111111111111100000110011;
assign LUT_2[59319] = 32'b11111111111111111100011001001100;
assign LUT_2[59320] = 32'b11111111111111110110111011101100;
assign LUT_2[59321] = 32'b11111111111111110011110100000101;
assign LUT_2[59322] = 32'b11111111111111111101110100101000;
assign LUT_2[59323] = 32'b11111111111111111010101101000001;
assign LUT_2[59324] = 32'b11111111111111110011011001010100;
assign LUT_2[59325] = 32'b11111111111111110000010001101101;
assign LUT_2[59326] = 32'b11111111111111111010010010010000;
assign LUT_2[59327] = 32'b11111111111111110111001010101001;
assign LUT_2[59328] = 32'b11111111111111111001010010111111;
assign LUT_2[59329] = 32'b11111111111111110110001011011000;
assign LUT_2[59330] = 32'b00000000000000000000001011111011;
assign LUT_2[59331] = 32'b11111111111111111101000100010100;
assign LUT_2[59332] = 32'b11111111111111110101110000100111;
assign LUT_2[59333] = 32'b11111111111111110010101001000000;
assign LUT_2[59334] = 32'b11111111111111111100101001100011;
assign LUT_2[59335] = 32'b11111111111111111001100001111100;
assign LUT_2[59336] = 32'b11111111111111110100000100011100;
assign LUT_2[59337] = 32'b11111111111111110000111100110101;
assign LUT_2[59338] = 32'b11111111111111111010111101011000;
assign LUT_2[59339] = 32'b11111111111111110111110101110001;
assign LUT_2[59340] = 32'b11111111111111110000100010000100;
assign LUT_2[59341] = 32'b11111111111111101101011010011101;
assign LUT_2[59342] = 32'b11111111111111110111011011000000;
assign LUT_2[59343] = 32'b11111111111111110100010011011001;
assign LUT_2[59344] = 32'b11111111111111110011110111001001;
assign LUT_2[59345] = 32'b11111111111111110000101111100010;
assign LUT_2[59346] = 32'b11111111111111111010110000000101;
assign LUT_2[59347] = 32'b11111111111111110111101000011110;
assign LUT_2[59348] = 32'b11111111111111110000010100110001;
assign LUT_2[59349] = 32'b11111111111111101101001101001010;
assign LUT_2[59350] = 32'b11111111111111110111001101101101;
assign LUT_2[59351] = 32'b11111111111111110100000110000110;
assign LUT_2[59352] = 32'b11111111111111101110101000100110;
assign LUT_2[59353] = 32'b11111111111111101011100000111111;
assign LUT_2[59354] = 32'b11111111111111110101100001100010;
assign LUT_2[59355] = 32'b11111111111111110010011001111011;
assign LUT_2[59356] = 32'b11111111111111101011000110001110;
assign LUT_2[59357] = 32'b11111111111111100111111110100111;
assign LUT_2[59358] = 32'b11111111111111110001111111001010;
assign LUT_2[59359] = 32'b11111111111111101110110111100011;
assign LUT_2[59360] = 32'b11111111111111111001101110101000;
assign LUT_2[59361] = 32'b11111111111111110110100111000001;
assign LUT_2[59362] = 32'b00000000000000000000100111100100;
assign LUT_2[59363] = 32'b11111111111111111101011111111101;
assign LUT_2[59364] = 32'b11111111111111110110001100010000;
assign LUT_2[59365] = 32'b11111111111111110011000100101001;
assign LUT_2[59366] = 32'b11111111111111111101000101001100;
assign LUT_2[59367] = 32'b11111111111111111001111101100101;
assign LUT_2[59368] = 32'b11111111111111110100100000000101;
assign LUT_2[59369] = 32'b11111111111111110001011000011110;
assign LUT_2[59370] = 32'b11111111111111111011011001000001;
assign LUT_2[59371] = 32'b11111111111111111000010001011010;
assign LUT_2[59372] = 32'b11111111111111110000111101101101;
assign LUT_2[59373] = 32'b11111111111111101101110110000110;
assign LUT_2[59374] = 32'b11111111111111110111110110101001;
assign LUT_2[59375] = 32'b11111111111111110100101111000010;
assign LUT_2[59376] = 32'b11111111111111110100010010110010;
assign LUT_2[59377] = 32'b11111111111111110001001011001011;
assign LUT_2[59378] = 32'b11111111111111111011001011101110;
assign LUT_2[59379] = 32'b11111111111111111000000100000111;
assign LUT_2[59380] = 32'b11111111111111110000110000011010;
assign LUT_2[59381] = 32'b11111111111111101101101000110011;
assign LUT_2[59382] = 32'b11111111111111110111101001010110;
assign LUT_2[59383] = 32'b11111111111111110100100001101111;
assign LUT_2[59384] = 32'b11111111111111101111000100001111;
assign LUT_2[59385] = 32'b11111111111111101011111100101000;
assign LUT_2[59386] = 32'b11111111111111110101111101001011;
assign LUT_2[59387] = 32'b11111111111111110010110101100100;
assign LUT_2[59388] = 32'b11111111111111101011100001110111;
assign LUT_2[59389] = 32'b11111111111111101000011010010000;
assign LUT_2[59390] = 32'b11111111111111110010011010110011;
assign LUT_2[59391] = 32'b11111111111111101111010011001100;
assign LUT_2[59392] = 32'b11111111111111101001001111101100;
assign LUT_2[59393] = 32'b11111111111111100110001000000101;
assign LUT_2[59394] = 32'b11111111111111110000001000101000;
assign LUT_2[59395] = 32'b11111111111111101101000001000001;
assign LUT_2[59396] = 32'b11111111111111100101101101010100;
assign LUT_2[59397] = 32'b11111111111111100010100101101101;
assign LUT_2[59398] = 32'b11111111111111101100100110010000;
assign LUT_2[59399] = 32'b11111111111111101001011110101001;
assign LUT_2[59400] = 32'b11111111111111100100000001001001;
assign LUT_2[59401] = 32'b11111111111111100000111001100010;
assign LUT_2[59402] = 32'b11111111111111101010111010000101;
assign LUT_2[59403] = 32'b11111111111111100111110010011110;
assign LUT_2[59404] = 32'b11111111111111100000011110110001;
assign LUT_2[59405] = 32'b11111111111111011101010111001010;
assign LUT_2[59406] = 32'b11111111111111100111010111101101;
assign LUT_2[59407] = 32'b11111111111111100100010000000110;
assign LUT_2[59408] = 32'b11111111111111100011110011110110;
assign LUT_2[59409] = 32'b11111111111111100000101100001111;
assign LUT_2[59410] = 32'b11111111111111101010101100110010;
assign LUT_2[59411] = 32'b11111111111111100111100101001011;
assign LUT_2[59412] = 32'b11111111111111100000010001011110;
assign LUT_2[59413] = 32'b11111111111111011101001001110111;
assign LUT_2[59414] = 32'b11111111111111100111001010011010;
assign LUT_2[59415] = 32'b11111111111111100100000010110011;
assign LUT_2[59416] = 32'b11111111111111011110100101010011;
assign LUT_2[59417] = 32'b11111111111111011011011101101100;
assign LUT_2[59418] = 32'b11111111111111100101011110001111;
assign LUT_2[59419] = 32'b11111111111111100010010110101000;
assign LUT_2[59420] = 32'b11111111111111011011000010111011;
assign LUT_2[59421] = 32'b11111111111111010111111011010100;
assign LUT_2[59422] = 32'b11111111111111100001111011110111;
assign LUT_2[59423] = 32'b11111111111111011110110100010000;
assign LUT_2[59424] = 32'b11111111111111101001101011010101;
assign LUT_2[59425] = 32'b11111111111111100110100011101110;
assign LUT_2[59426] = 32'b11111111111111110000100100010001;
assign LUT_2[59427] = 32'b11111111111111101101011100101010;
assign LUT_2[59428] = 32'b11111111111111100110001000111101;
assign LUT_2[59429] = 32'b11111111111111100011000001010110;
assign LUT_2[59430] = 32'b11111111111111101101000001111001;
assign LUT_2[59431] = 32'b11111111111111101001111010010010;
assign LUT_2[59432] = 32'b11111111111111100100011100110010;
assign LUT_2[59433] = 32'b11111111111111100001010101001011;
assign LUT_2[59434] = 32'b11111111111111101011010101101110;
assign LUT_2[59435] = 32'b11111111111111101000001110000111;
assign LUT_2[59436] = 32'b11111111111111100000111010011010;
assign LUT_2[59437] = 32'b11111111111111011101110010110011;
assign LUT_2[59438] = 32'b11111111111111100111110011010110;
assign LUT_2[59439] = 32'b11111111111111100100101011101111;
assign LUT_2[59440] = 32'b11111111111111100100001111011111;
assign LUT_2[59441] = 32'b11111111111111100001000111111000;
assign LUT_2[59442] = 32'b11111111111111101011001000011011;
assign LUT_2[59443] = 32'b11111111111111101000000000110100;
assign LUT_2[59444] = 32'b11111111111111100000101101000111;
assign LUT_2[59445] = 32'b11111111111111011101100101100000;
assign LUT_2[59446] = 32'b11111111111111100111100110000011;
assign LUT_2[59447] = 32'b11111111111111100100011110011100;
assign LUT_2[59448] = 32'b11111111111111011111000000111100;
assign LUT_2[59449] = 32'b11111111111111011011111001010101;
assign LUT_2[59450] = 32'b11111111111111100101111001111000;
assign LUT_2[59451] = 32'b11111111111111100010110010010001;
assign LUT_2[59452] = 32'b11111111111111011011011110100100;
assign LUT_2[59453] = 32'b11111111111111011000010110111101;
assign LUT_2[59454] = 32'b11111111111111100010010111100000;
assign LUT_2[59455] = 32'b11111111111111011111001111111001;
assign LUT_2[59456] = 32'b11111111111111100001011000001111;
assign LUT_2[59457] = 32'b11111111111111011110010000101000;
assign LUT_2[59458] = 32'b11111111111111101000010001001011;
assign LUT_2[59459] = 32'b11111111111111100101001001100100;
assign LUT_2[59460] = 32'b11111111111111011101110101110111;
assign LUT_2[59461] = 32'b11111111111111011010101110010000;
assign LUT_2[59462] = 32'b11111111111111100100101110110011;
assign LUT_2[59463] = 32'b11111111111111100001100111001100;
assign LUT_2[59464] = 32'b11111111111111011100001001101100;
assign LUT_2[59465] = 32'b11111111111111011001000010000101;
assign LUT_2[59466] = 32'b11111111111111100011000010101000;
assign LUT_2[59467] = 32'b11111111111111011111111011000001;
assign LUT_2[59468] = 32'b11111111111111011000100111010100;
assign LUT_2[59469] = 32'b11111111111111010101011111101101;
assign LUT_2[59470] = 32'b11111111111111011111100000010000;
assign LUT_2[59471] = 32'b11111111111111011100011000101001;
assign LUT_2[59472] = 32'b11111111111111011011111100011001;
assign LUT_2[59473] = 32'b11111111111111011000110100110010;
assign LUT_2[59474] = 32'b11111111111111100010110101010101;
assign LUT_2[59475] = 32'b11111111111111011111101101101110;
assign LUT_2[59476] = 32'b11111111111111011000011010000001;
assign LUT_2[59477] = 32'b11111111111111010101010010011010;
assign LUT_2[59478] = 32'b11111111111111011111010010111101;
assign LUT_2[59479] = 32'b11111111111111011100001011010110;
assign LUT_2[59480] = 32'b11111111111111010110101101110110;
assign LUT_2[59481] = 32'b11111111111111010011100110001111;
assign LUT_2[59482] = 32'b11111111111111011101100110110010;
assign LUT_2[59483] = 32'b11111111111111011010011111001011;
assign LUT_2[59484] = 32'b11111111111111010011001011011110;
assign LUT_2[59485] = 32'b11111111111111010000000011110111;
assign LUT_2[59486] = 32'b11111111111111011010000100011010;
assign LUT_2[59487] = 32'b11111111111111010110111100110011;
assign LUT_2[59488] = 32'b11111111111111100001110011111000;
assign LUT_2[59489] = 32'b11111111111111011110101100010001;
assign LUT_2[59490] = 32'b11111111111111101000101100110100;
assign LUT_2[59491] = 32'b11111111111111100101100101001101;
assign LUT_2[59492] = 32'b11111111111111011110010001100000;
assign LUT_2[59493] = 32'b11111111111111011011001001111001;
assign LUT_2[59494] = 32'b11111111111111100101001010011100;
assign LUT_2[59495] = 32'b11111111111111100010000010110101;
assign LUT_2[59496] = 32'b11111111111111011100100101010101;
assign LUT_2[59497] = 32'b11111111111111011001011101101110;
assign LUT_2[59498] = 32'b11111111111111100011011110010001;
assign LUT_2[59499] = 32'b11111111111111100000010110101010;
assign LUT_2[59500] = 32'b11111111111111011001000010111101;
assign LUT_2[59501] = 32'b11111111111111010101111011010110;
assign LUT_2[59502] = 32'b11111111111111011111111011111001;
assign LUT_2[59503] = 32'b11111111111111011100110100010010;
assign LUT_2[59504] = 32'b11111111111111011100011000000010;
assign LUT_2[59505] = 32'b11111111111111011001010000011011;
assign LUT_2[59506] = 32'b11111111111111100011010000111110;
assign LUT_2[59507] = 32'b11111111111111100000001001010111;
assign LUT_2[59508] = 32'b11111111111111011000110101101010;
assign LUT_2[59509] = 32'b11111111111111010101101110000011;
assign LUT_2[59510] = 32'b11111111111111011111101110100110;
assign LUT_2[59511] = 32'b11111111111111011100100110111111;
assign LUT_2[59512] = 32'b11111111111111010111001001011111;
assign LUT_2[59513] = 32'b11111111111111010100000001111000;
assign LUT_2[59514] = 32'b11111111111111011110000010011011;
assign LUT_2[59515] = 32'b11111111111111011010111010110100;
assign LUT_2[59516] = 32'b11111111111111010011100111000111;
assign LUT_2[59517] = 32'b11111111111111010000011111100000;
assign LUT_2[59518] = 32'b11111111111111011010100000000011;
assign LUT_2[59519] = 32'b11111111111111010111011000011100;
assign LUT_2[59520] = 32'b11111111111111101101100011111011;
assign LUT_2[59521] = 32'b11111111111111101010011100010100;
assign LUT_2[59522] = 32'b11111111111111110100011100110111;
assign LUT_2[59523] = 32'b11111111111111110001010101010000;
assign LUT_2[59524] = 32'b11111111111111101010000001100011;
assign LUT_2[59525] = 32'b11111111111111100110111001111100;
assign LUT_2[59526] = 32'b11111111111111110000111010011111;
assign LUT_2[59527] = 32'b11111111111111101101110010111000;
assign LUT_2[59528] = 32'b11111111111111101000010101011000;
assign LUT_2[59529] = 32'b11111111111111100101001101110001;
assign LUT_2[59530] = 32'b11111111111111101111001110010100;
assign LUT_2[59531] = 32'b11111111111111101100000110101101;
assign LUT_2[59532] = 32'b11111111111111100100110011000000;
assign LUT_2[59533] = 32'b11111111111111100001101011011001;
assign LUT_2[59534] = 32'b11111111111111101011101011111100;
assign LUT_2[59535] = 32'b11111111111111101000100100010101;
assign LUT_2[59536] = 32'b11111111111111101000001000000101;
assign LUT_2[59537] = 32'b11111111111111100101000000011110;
assign LUT_2[59538] = 32'b11111111111111101111000001000001;
assign LUT_2[59539] = 32'b11111111111111101011111001011010;
assign LUT_2[59540] = 32'b11111111111111100100100101101101;
assign LUT_2[59541] = 32'b11111111111111100001011110000110;
assign LUT_2[59542] = 32'b11111111111111101011011110101001;
assign LUT_2[59543] = 32'b11111111111111101000010111000010;
assign LUT_2[59544] = 32'b11111111111111100010111001100010;
assign LUT_2[59545] = 32'b11111111111111011111110001111011;
assign LUT_2[59546] = 32'b11111111111111101001110010011110;
assign LUT_2[59547] = 32'b11111111111111100110101010110111;
assign LUT_2[59548] = 32'b11111111111111011111010111001010;
assign LUT_2[59549] = 32'b11111111111111011100001111100011;
assign LUT_2[59550] = 32'b11111111111111100110010000000110;
assign LUT_2[59551] = 32'b11111111111111100011001000011111;
assign LUT_2[59552] = 32'b11111111111111101101111111100100;
assign LUT_2[59553] = 32'b11111111111111101010110111111101;
assign LUT_2[59554] = 32'b11111111111111110100111000100000;
assign LUT_2[59555] = 32'b11111111111111110001110000111001;
assign LUT_2[59556] = 32'b11111111111111101010011101001100;
assign LUT_2[59557] = 32'b11111111111111100111010101100101;
assign LUT_2[59558] = 32'b11111111111111110001010110001000;
assign LUT_2[59559] = 32'b11111111111111101110001110100001;
assign LUT_2[59560] = 32'b11111111111111101000110001000001;
assign LUT_2[59561] = 32'b11111111111111100101101001011010;
assign LUT_2[59562] = 32'b11111111111111101111101001111101;
assign LUT_2[59563] = 32'b11111111111111101100100010010110;
assign LUT_2[59564] = 32'b11111111111111100101001110101001;
assign LUT_2[59565] = 32'b11111111111111100010000111000010;
assign LUT_2[59566] = 32'b11111111111111101100000111100101;
assign LUT_2[59567] = 32'b11111111111111101000111111111110;
assign LUT_2[59568] = 32'b11111111111111101000100011101110;
assign LUT_2[59569] = 32'b11111111111111100101011100000111;
assign LUT_2[59570] = 32'b11111111111111101111011100101010;
assign LUT_2[59571] = 32'b11111111111111101100010101000011;
assign LUT_2[59572] = 32'b11111111111111100101000001010110;
assign LUT_2[59573] = 32'b11111111111111100001111001101111;
assign LUT_2[59574] = 32'b11111111111111101011111010010010;
assign LUT_2[59575] = 32'b11111111111111101000110010101011;
assign LUT_2[59576] = 32'b11111111111111100011010101001011;
assign LUT_2[59577] = 32'b11111111111111100000001101100100;
assign LUT_2[59578] = 32'b11111111111111101010001110000111;
assign LUT_2[59579] = 32'b11111111111111100111000110100000;
assign LUT_2[59580] = 32'b11111111111111011111110010110011;
assign LUT_2[59581] = 32'b11111111111111011100101011001100;
assign LUT_2[59582] = 32'b11111111111111100110101011101111;
assign LUT_2[59583] = 32'b11111111111111100011100100001000;
assign LUT_2[59584] = 32'b11111111111111100101101100011110;
assign LUT_2[59585] = 32'b11111111111111100010100100110111;
assign LUT_2[59586] = 32'b11111111111111101100100101011010;
assign LUT_2[59587] = 32'b11111111111111101001011101110011;
assign LUT_2[59588] = 32'b11111111111111100010001010000110;
assign LUT_2[59589] = 32'b11111111111111011111000010011111;
assign LUT_2[59590] = 32'b11111111111111101001000011000010;
assign LUT_2[59591] = 32'b11111111111111100101111011011011;
assign LUT_2[59592] = 32'b11111111111111100000011101111011;
assign LUT_2[59593] = 32'b11111111111111011101010110010100;
assign LUT_2[59594] = 32'b11111111111111100111010110110111;
assign LUT_2[59595] = 32'b11111111111111100100001111010000;
assign LUT_2[59596] = 32'b11111111111111011100111011100011;
assign LUT_2[59597] = 32'b11111111111111011001110011111100;
assign LUT_2[59598] = 32'b11111111111111100011110100011111;
assign LUT_2[59599] = 32'b11111111111111100000101100111000;
assign LUT_2[59600] = 32'b11111111111111100000010000101000;
assign LUT_2[59601] = 32'b11111111111111011101001001000001;
assign LUT_2[59602] = 32'b11111111111111100111001001100100;
assign LUT_2[59603] = 32'b11111111111111100100000001111101;
assign LUT_2[59604] = 32'b11111111111111011100101110010000;
assign LUT_2[59605] = 32'b11111111111111011001100110101001;
assign LUT_2[59606] = 32'b11111111111111100011100111001100;
assign LUT_2[59607] = 32'b11111111111111100000011111100101;
assign LUT_2[59608] = 32'b11111111111111011011000010000101;
assign LUT_2[59609] = 32'b11111111111111010111111010011110;
assign LUT_2[59610] = 32'b11111111111111100001111011000001;
assign LUT_2[59611] = 32'b11111111111111011110110011011010;
assign LUT_2[59612] = 32'b11111111111111010111011111101101;
assign LUT_2[59613] = 32'b11111111111111010100011000000110;
assign LUT_2[59614] = 32'b11111111111111011110011000101001;
assign LUT_2[59615] = 32'b11111111111111011011010001000010;
assign LUT_2[59616] = 32'b11111111111111100110001000000111;
assign LUT_2[59617] = 32'b11111111111111100011000000100000;
assign LUT_2[59618] = 32'b11111111111111101101000001000011;
assign LUT_2[59619] = 32'b11111111111111101001111001011100;
assign LUT_2[59620] = 32'b11111111111111100010100101101111;
assign LUT_2[59621] = 32'b11111111111111011111011110001000;
assign LUT_2[59622] = 32'b11111111111111101001011110101011;
assign LUT_2[59623] = 32'b11111111111111100110010111000100;
assign LUT_2[59624] = 32'b11111111111111100000111001100100;
assign LUT_2[59625] = 32'b11111111111111011101110001111101;
assign LUT_2[59626] = 32'b11111111111111100111110010100000;
assign LUT_2[59627] = 32'b11111111111111100100101010111001;
assign LUT_2[59628] = 32'b11111111111111011101010111001100;
assign LUT_2[59629] = 32'b11111111111111011010001111100101;
assign LUT_2[59630] = 32'b11111111111111100100010000001000;
assign LUT_2[59631] = 32'b11111111111111100001001000100001;
assign LUT_2[59632] = 32'b11111111111111100000101100010001;
assign LUT_2[59633] = 32'b11111111111111011101100100101010;
assign LUT_2[59634] = 32'b11111111111111100111100101001101;
assign LUT_2[59635] = 32'b11111111111111100100011101100110;
assign LUT_2[59636] = 32'b11111111111111011101001001111001;
assign LUT_2[59637] = 32'b11111111111111011010000010010010;
assign LUT_2[59638] = 32'b11111111111111100100000010110101;
assign LUT_2[59639] = 32'b11111111111111100000111011001110;
assign LUT_2[59640] = 32'b11111111111111011011011101101110;
assign LUT_2[59641] = 32'b11111111111111011000010110000111;
assign LUT_2[59642] = 32'b11111111111111100010010110101010;
assign LUT_2[59643] = 32'b11111111111111011111001111000011;
assign LUT_2[59644] = 32'b11111111111111010111111011010110;
assign LUT_2[59645] = 32'b11111111111111010100110011101111;
assign LUT_2[59646] = 32'b11111111111111011110110100010010;
assign LUT_2[59647] = 32'b11111111111111011011101100101011;
assign LUT_2[59648] = 32'b11111111111111101101001110010010;
assign LUT_2[59649] = 32'b11111111111111101010000110101011;
assign LUT_2[59650] = 32'b11111111111111110100000111001110;
assign LUT_2[59651] = 32'b11111111111111110000111111100111;
assign LUT_2[59652] = 32'b11111111111111101001101011111010;
assign LUT_2[59653] = 32'b11111111111111100110100100010011;
assign LUT_2[59654] = 32'b11111111111111110000100100110110;
assign LUT_2[59655] = 32'b11111111111111101101011101001111;
assign LUT_2[59656] = 32'b11111111111111100111111111101111;
assign LUT_2[59657] = 32'b11111111111111100100111000001000;
assign LUT_2[59658] = 32'b11111111111111101110111000101011;
assign LUT_2[59659] = 32'b11111111111111101011110001000100;
assign LUT_2[59660] = 32'b11111111111111100100011101010111;
assign LUT_2[59661] = 32'b11111111111111100001010101110000;
assign LUT_2[59662] = 32'b11111111111111101011010110010011;
assign LUT_2[59663] = 32'b11111111111111101000001110101100;
assign LUT_2[59664] = 32'b11111111111111100111110010011100;
assign LUT_2[59665] = 32'b11111111111111100100101010110101;
assign LUT_2[59666] = 32'b11111111111111101110101011011000;
assign LUT_2[59667] = 32'b11111111111111101011100011110001;
assign LUT_2[59668] = 32'b11111111111111100100010000000100;
assign LUT_2[59669] = 32'b11111111111111100001001000011101;
assign LUT_2[59670] = 32'b11111111111111101011001001000000;
assign LUT_2[59671] = 32'b11111111111111101000000001011001;
assign LUT_2[59672] = 32'b11111111111111100010100011111001;
assign LUT_2[59673] = 32'b11111111111111011111011100010010;
assign LUT_2[59674] = 32'b11111111111111101001011100110101;
assign LUT_2[59675] = 32'b11111111111111100110010101001110;
assign LUT_2[59676] = 32'b11111111111111011111000001100001;
assign LUT_2[59677] = 32'b11111111111111011011111001111010;
assign LUT_2[59678] = 32'b11111111111111100101111010011101;
assign LUT_2[59679] = 32'b11111111111111100010110010110110;
assign LUT_2[59680] = 32'b11111111111111101101101001111011;
assign LUT_2[59681] = 32'b11111111111111101010100010010100;
assign LUT_2[59682] = 32'b11111111111111110100100010110111;
assign LUT_2[59683] = 32'b11111111111111110001011011010000;
assign LUT_2[59684] = 32'b11111111111111101010000111100011;
assign LUT_2[59685] = 32'b11111111111111100110111111111100;
assign LUT_2[59686] = 32'b11111111111111110001000000011111;
assign LUT_2[59687] = 32'b11111111111111101101111000111000;
assign LUT_2[59688] = 32'b11111111111111101000011011011000;
assign LUT_2[59689] = 32'b11111111111111100101010011110001;
assign LUT_2[59690] = 32'b11111111111111101111010100010100;
assign LUT_2[59691] = 32'b11111111111111101100001100101101;
assign LUT_2[59692] = 32'b11111111111111100100111001000000;
assign LUT_2[59693] = 32'b11111111111111100001110001011001;
assign LUT_2[59694] = 32'b11111111111111101011110001111100;
assign LUT_2[59695] = 32'b11111111111111101000101010010101;
assign LUT_2[59696] = 32'b11111111111111101000001110000101;
assign LUT_2[59697] = 32'b11111111111111100101000110011110;
assign LUT_2[59698] = 32'b11111111111111101111000111000001;
assign LUT_2[59699] = 32'b11111111111111101011111111011010;
assign LUT_2[59700] = 32'b11111111111111100100101011101101;
assign LUT_2[59701] = 32'b11111111111111100001100100000110;
assign LUT_2[59702] = 32'b11111111111111101011100100101001;
assign LUT_2[59703] = 32'b11111111111111101000011101000010;
assign LUT_2[59704] = 32'b11111111111111100010111111100010;
assign LUT_2[59705] = 32'b11111111111111011111110111111011;
assign LUT_2[59706] = 32'b11111111111111101001111000011110;
assign LUT_2[59707] = 32'b11111111111111100110110000110111;
assign LUT_2[59708] = 32'b11111111111111011111011101001010;
assign LUT_2[59709] = 32'b11111111111111011100010101100011;
assign LUT_2[59710] = 32'b11111111111111100110010110000110;
assign LUT_2[59711] = 32'b11111111111111100011001110011111;
assign LUT_2[59712] = 32'b11111111111111100101010110110101;
assign LUT_2[59713] = 32'b11111111111111100010001111001110;
assign LUT_2[59714] = 32'b11111111111111101100001111110001;
assign LUT_2[59715] = 32'b11111111111111101001001000001010;
assign LUT_2[59716] = 32'b11111111111111100001110100011101;
assign LUT_2[59717] = 32'b11111111111111011110101100110110;
assign LUT_2[59718] = 32'b11111111111111101000101101011001;
assign LUT_2[59719] = 32'b11111111111111100101100101110010;
assign LUT_2[59720] = 32'b11111111111111100000001000010010;
assign LUT_2[59721] = 32'b11111111111111011101000000101011;
assign LUT_2[59722] = 32'b11111111111111100111000001001110;
assign LUT_2[59723] = 32'b11111111111111100011111001100111;
assign LUT_2[59724] = 32'b11111111111111011100100101111010;
assign LUT_2[59725] = 32'b11111111111111011001011110010011;
assign LUT_2[59726] = 32'b11111111111111100011011110110110;
assign LUT_2[59727] = 32'b11111111111111100000010111001111;
assign LUT_2[59728] = 32'b11111111111111011111111010111111;
assign LUT_2[59729] = 32'b11111111111111011100110011011000;
assign LUT_2[59730] = 32'b11111111111111100110110011111011;
assign LUT_2[59731] = 32'b11111111111111100011101100010100;
assign LUT_2[59732] = 32'b11111111111111011100011000100111;
assign LUT_2[59733] = 32'b11111111111111011001010001000000;
assign LUT_2[59734] = 32'b11111111111111100011010001100011;
assign LUT_2[59735] = 32'b11111111111111100000001001111100;
assign LUT_2[59736] = 32'b11111111111111011010101100011100;
assign LUT_2[59737] = 32'b11111111111111010111100100110101;
assign LUT_2[59738] = 32'b11111111111111100001100101011000;
assign LUT_2[59739] = 32'b11111111111111011110011101110001;
assign LUT_2[59740] = 32'b11111111111111010111001010000100;
assign LUT_2[59741] = 32'b11111111111111010100000010011101;
assign LUT_2[59742] = 32'b11111111111111011110000011000000;
assign LUT_2[59743] = 32'b11111111111111011010111011011001;
assign LUT_2[59744] = 32'b11111111111111100101110010011110;
assign LUT_2[59745] = 32'b11111111111111100010101010110111;
assign LUT_2[59746] = 32'b11111111111111101100101011011010;
assign LUT_2[59747] = 32'b11111111111111101001100011110011;
assign LUT_2[59748] = 32'b11111111111111100010010000000110;
assign LUT_2[59749] = 32'b11111111111111011111001000011111;
assign LUT_2[59750] = 32'b11111111111111101001001001000010;
assign LUT_2[59751] = 32'b11111111111111100110000001011011;
assign LUT_2[59752] = 32'b11111111111111100000100011111011;
assign LUT_2[59753] = 32'b11111111111111011101011100010100;
assign LUT_2[59754] = 32'b11111111111111100111011100110111;
assign LUT_2[59755] = 32'b11111111111111100100010101010000;
assign LUT_2[59756] = 32'b11111111111111011101000001100011;
assign LUT_2[59757] = 32'b11111111111111011001111001111100;
assign LUT_2[59758] = 32'b11111111111111100011111010011111;
assign LUT_2[59759] = 32'b11111111111111100000110010111000;
assign LUT_2[59760] = 32'b11111111111111100000010110101000;
assign LUT_2[59761] = 32'b11111111111111011101001111000001;
assign LUT_2[59762] = 32'b11111111111111100111001111100100;
assign LUT_2[59763] = 32'b11111111111111100100000111111101;
assign LUT_2[59764] = 32'b11111111111111011100110100010000;
assign LUT_2[59765] = 32'b11111111111111011001101100101001;
assign LUT_2[59766] = 32'b11111111111111100011101101001100;
assign LUT_2[59767] = 32'b11111111111111100000100101100101;
assign LUT_2[59768] = 32'b11111111111111011011001000000101;
assign LUT_2[59769] = 32'b11111111111111011000000000011110;
assign LUT_2[59770] = 32'b11111111111111100010000001000001;
assign LUT_2[59771] = 32'b11111111111111011110111001011010;
assign LUT_2[59772] = 32'b11111111111111010111100101101101;
assign LUT_2[59773] = 32'b11111111111111010100011110000110;
assign LUT_2[59774] = 32'b11111111111111011110011110101001;
assign LUT_2[59775] = 32'b11111111111111011011010111000010;
assign LUT_2[59776] = 32'b11111111111111110001100010100001;
assign LUT_2[59777] = 32'b11111111111111101110011010111010;
assign LUT_2[59778] = 32'b11111111111111111000011011011101;
assign LUT_2[59779] = 32'b11111111111111110101010011110110;
assign LUT_2[59780] = 32'b11111111111111101110000000001001;
assign LUT_2[59781] = 32'b11111111111111101010111000100010;
assign LUT_2[59782] = 32'b11111111111111110100111001000101;
assign LUT_2[59783] = 32'b11111111111111110001110001011110;
assign LUT_2[59784] = 32'b11111111111111101100010011111110;
assign LUT_2[59785] = 32'b11111111111111101001001100010111;
assign LUT_2[59786] = 32'b11111111111111110011001100111010;
assign LUT_2[59787] = 32'b11111111111111110000000101010011;
assign LUT_2[59788] = 32'b11111111111111101000110001100110;
assign LUT_2[59789] = 32'b11111111111111100101101001111111;
assign LUT_2[59790] = 32'b11111111111111101111101010100010;
assign LUT_2[59791] = 32'b11111111111111101100100010111011;
assign LUT_2[59792] = 32'b11111111111111101100000110101011;
assign LUT_2[59793] = 32'b11111111111111101000111111000100;
assign LUT_2[59794] = 32'b11111111111111110010111111100111;
assign LUT_2[59795] = 32'b11111111111111101111111000000000;
assign LUT_2[59796] = 32'b11111111111111101000100100010011;
assign LUT_2[59797] = 32'b11111111111111100101011100101100;
assign LUT_2[59798] = 32'b11111111111111101111011101001111;
assign LUT_2[59799] = 32'b11111111111111101100010101101000;
assign LUT_2[59800] = 32'b11111111111111100110111000001000;
assign LUT_2[59801] = 32'b11111111111111100011110000100001;
assign LUT_2[59802] = 32'b11111111111111101101110001000100;
assign LUT_2[59803] = 32'b11111111111111101010101001011101;
assign LUT_2[59804] = 32'b11111111111111100011010101110000;
assign LUT_2[59805] = 32'b11111111111111100000001110001001;
assign LUT_2[59806] = 32'b11111111111111101010001110101100;
assign LUT_2[59807] = 32'b11111111111111100111000111000101;
assign LUT_2[59808] = 32'b11111111111111110001111110001010;
assign LUT_2[59809] = 32'b11111111111111101110110110100011;
assign LUT_2[59810] = 32'b11111111111111111000110111000110;
assign LUT_2[59811] = 32'b11111111111111110101101111011111;
assign LUT_2[59812] = 32'b11111111111111101110011011110010;
assign LUT_2[59813] = 32'b11111111111111101011010100001011;
assign LUT_2[59814] = 32'b11111111111111110101010100101110;
assign LUT_2[59815] = 32'b11111111111111110010001101000111;
assign LUT_2[59816] = 32'b11111111111111101100101111100111;
assign LUT_2[59817] = 32'b11111111111111101001101000000000;
assign LUT_2[59818] = 32'b11111111111111110011101000100011;
assign LUT_2[59819] = 32'b11111111111111110000100000111100;
assign LUT_2[59820] = 32'b11111111111111101001001101001111;
assign LUT_2[59821] = 32'b11111111111111100110000101101000;
assign LUT_2[59822] = 32'b11111111111111110000000110001011;
assign LUT_2[59823] = 32'b11111111111111101100111110100100;
assign LUT_2[59824] = 32'b11111111111111101100100010010100;
assign LUT_2[59825] = 32'b11111111111111101001011010101101;
assign LUT_2[59826] = 32'b11111111111111110011011011010000;
assign LUT_2[59827] = 32'b11111111111111110000010011101001;
assign LUT_2[59828] = 32'b11111111111111101000111111111100;
assign LUT_2[59829] = 32'b11111111111111100101111000010101;
assign LUT_2[59830] = 32'b11111111111111101111111000111000;
assign LUT_2[59831] = 32'b11111111111111101100110001010001;
assign LUT_2[59832] = 32'b11111111111111100111010011110001;
assign LUT_2[59833] = 32'b11111111111111100100001100001010;
assign LUT_2[59834] = 32'b11111111111111101110001100101101;
assign LUT_2[59835] = 32'b11111111111111101011000101000110;
assign LUT_2[59836] = 32'b11111111111111100011110001011001;
assign LUT_2[59837] = 32'b11111111111111100000101001110010;
assign LUT_2[59838] = 32'b11111111111111101010101010010101;
assign LUT_2[59839] = 32'b11111111111111100111100010101110;
assign LUT_2[59840] = 32'b11111111111111101001101011000100;
assign LUT_2[59841] = 32'b11111111111111100110100011011101;
assign LUT_2[59842] = 32'b11111111111111110000100100000000;
assign LUT_2[59843] = 32'b11111111111111101101011100011001;
assign LUT_2[59844] = 32'b11111111111111100110001000101100;
assign LUT_2[59845] = 32'b11111111111111100011000001000101;
assign LUT_2[59846] = 32'b11111111111111101101000001101000;
assign LUT_2[59847] = 32'b11111111111111101001111010000001;
assign LUT_2[59848] = 32'b11111111111111100100011100100001;
assign LUT_2[59849] = 32'b11111111111111100001010100111010;
assign LUT_2[59850] = 32'b11111111111111101011010101011101;
assign LUT_2[59851] = 32'b11111111111111101000001101110110;
assign LUT_2[59852] = 32'b11111111111111100000111010001001;
assign LUT_2[59853] = 32'b11111111111111011101110010100010;
assign LUT_2[59854] = 32'b11111111111111100111110011000101;
assign LUT_2[59855] = 32'b11111111111111100100101011011110;
assign LUT_2[59856] = 32'b11111111111111100100001111001110;
assign LUT_2[59857] = 32'b11111111111111100001000111100111;
assign LUT_2[59858] = 32'b11111111111111101011001000001010;
assign LUT_2[59859] = 32'b11111111111111101000000000100011;
assign LUT_2[59860] = 32'b11111111111111100000101100110110;
assign LUT_2[59861] = 32'b11111111111111011101100101001111;
assign LUT_2[59862] = 32'b11111111111111100111100101110010;
assign LUT_2[59863] = 32'b11111111111111100100011110001011;
assign LUT_2[59864] = 32'b11111111111111011111000000101011;
assign LUT_2[59865] = 32'b11111111111111011011111001000100;
assign LUT_2[59866] = 32'b11111111111111100101111001100111;
assign LUT_2[59867] = 32'b11111111111111100010110010000000;
assign LUT_2[59868] = 32'b11111111111111011011011110010011;
assign LUT_2[59869] = 32'b11111111111111011000010110101100;
assign LUT_2[59870] = 32'b11111111111111100010010111001111;
assign LUT_2[59871] = 32'b11111111111111011111001111101000;
assign LUT_2[59872] = 32'b11111111111111101010000110101101;
assign LUT_2[59873] = 32'b11111111111111100110111111000110;
assign LUT_2[59874] = 32'b11111111111111110000111111101001;
assign LUT_2[59875] = 32'b11111111111111101101111000000010;
assign LUT_2[59876] = 32'b11111111111111100110100100010101;
assign LUT_2[59877] = 32'b11111111111111100011011100101110;
assign LUT_2[59878] = 32'b11111111111111101101011101010001;
assign LUT_2[59879] = 32'b11111111111111101010010101101010;
assign LUT_2[59880] = 32'b11111111111111100100111000001010;
assign LUT_2[59881] = 32'b11111111111111100001110000100011;
assign LUT_2[59882] = 32'b11111111111111101011110001000110;
assign LUT_2[59883] = 32'b11111111111111101000101001011111;
assign LUT_2[59884] = 32'b11111111111111100001010101110010;
assign LUT_2[59885] = 32'b11111111111111011110001110001011;
assign LUT_2[59886] = 32'b11111111111111101000001110101110;
assign LUT_2[59887] = 32'b11111111111111100101000111000111;
assign LUT_2[59888] = 32'b11111111111111100100101010110111;
assign LUT_2[59889] = 32'b11111111111111100001100011010000;
assign LUT_2[59890] = 32'b11111111111111101011100011110011;
assign LUT_2[59891] = 32'b11111111111111101000011100001100;
assign LUT_2[59892] = 32'b11111111111111100001001000011111;
assign LUT_2[59893] = 32'b11111111111111011110000000111000;
assign LUT_2[59894] = 32'b11111111111111101000000001011011;
assign LUT_2[59895] = 32'b11111111111111100100111001110100;
assign LUT_2[59896] = 32'b11111111111111011111011100010100;
assign LUT_2[59897] = 32'b11111111111111011100010100101101;
assign LUT_2[59898] = 32'b11111111111111100110010101010000;
assign LUT_2[59899] = 32'b11111111111111100011001101101001;
assign LUT_2[59900] = 32'b11111111111111011011111001111100;
assign LUT_2[59901] = 32'b11111111111111011000110010010101;
assign LUT_2[59902] = 32'b11111111111111100010110010111000;
assign LUT_2[59903] = 32'b11111111111111011111101011010001;
assign LUT_2[59904] = 32'b11111111111111101110000001011110;
assign LUT_2[59905] = 32'b11111111111111101010111001110111;
assign LUT_2[59906] = 32'b11111111111111110100111010011010;
assign LUT_2[59907] = 32'b11111111111111110001110010110011;
assign LUT_2[59908] = 32'b11111111111111101010011111000110;
assign LUT_2[59909] = 32'b11111111111111100111010111011111;
assign LUT_2[59910] = 32'b11111111111111110001011000000010;
assign LUT_2[59911] = 32'b11111111111111101110010000011011;
assign LUT_2[59912] = 32'b11111111111111101000110010111011;
assign LUT_2[59913] = 32'b11111111111111100101101011010100;
assign LUT_2[59914] = 32'b11111111111111101111101011110111;
assign LUT_2[59915] = 32'b11111111111111101100100100010000;
assign LUT_2[59916] = 32'b11111111111111100101010000100011;
assign LUT_2[59917] = 32'b11111111111111100010001000111100;
assign LUT_2[59918] = 32'b11111111111111101100001001011111;
assign LUT_2[59919] = 32'b11111111111111101001000001111000;
assign LUT_2[59920] = 32'b11111111111111101000100101101000;
assign LUT_2[59921] = 32'b11111111111111100101011110000001;
assign LUT_2[59922] = 32'b11111111111111101111011110100100;
assign LUT_2[59923] = 32'b11111111111111101100010110111101;
assign LUT_2[59924] = 32'b11111111111111100101000011010000;
assign LUT_2[59925] = 32'b11111111111111100001111011101001;
assign LUT_2[59926] = 32'b11111111111111101011111100001100;
assign LUT_2[59927] = 32'b11111111111111101000110100100101;
assign LUT_2[59928] = 32'b11111111111111100011010111000101;
assign LUT_2[59929] = 32'b11111111111111100000001111011110;
assign LUT_2[59930] = 32'b11111111111111101010010000000001;
assign LUT_2[59931] = 32'b11111111111111100111001000011010;
assign LUT_2[59932] = 32'b11111111111111011111110100101101;
assign LUT_2[59933] = 32'b11111111111111011100101101000110;
assign LUT_2[59934] = 32'b11111111111111100110101101101001;
assign LUT_2[59935] = 32'b11111111111111100011100110000010;
assign LUT_2[59936] = 32'b11111111111111101110011101000111;
assign LUT_2[59937] = 32'b11111111111111101011010101100000;
assign LUT_2[59938] = 32'b11111111111111110101010110000011;
assign LUT_2[59939] = 32'b11111111111111110010001110011100;
assign LUT_2[59940] = 32'b11111111111111101010111010101111;
assign LUT_2[59941] = 32'b11111111111111100111110011001000;
assign LUT_2[59942] = 32'b11111111111111110001110011101011;
assign LUT_2[59943] = 32'b11111111111111101110101100000100;
assign LUT_2[59944] = 32'b11111111111111101001001110100100;
assign LUT_2[59945] = 32'b11111111111111100110000110111101;
assign LUT_2[59946] = 32'b11111111111111110000000111100000;
assign LUT_2[59947] = 32'b11111111111111101100111111111001;
assign LUT_2[59948] = 32'b11111111111111100101101100001100;
assign LUT_2[59949] = 32'b11111111111111100010100100100101;
assign LUT_2[59950] = 32'b11111111111111101100100101001000;
assign LUT_2[59951] = 32'b11111111111111101001011101100001;
assign LUT_2[59952] = 32'b11111111111111101001000001010001;
assign LUT_2[59953] = 32'b11111111111111100101111001101010;
assign LUT_2[59954] = 32'b11111111111111101111111010001101;
assign LUT_2[59955] = 32'b11111111111111101100110010100110;
assign LUT_2[59956] = 32'b11111111111111100101011110111001;
assign LUT_2[59957] = 32'b11111111111111100010010111010010;
assign LUT_2[59958] = 32'b11111111111111101100010111110101;
assign LUT_2[59959] = 32'b11111111111111101001010000001110;
assign LUT_2[59960] = 32'b11111111111111100011110010101110;
assign LUT_2[59961] = 32'b11111111111111100000101011000111;
assign LUT_2[59962] = 32'b11111111111111101010101011101010;
assign LUT_2[59963] = 32'b11111111111111100111100100000011;
assign LUT_2[59964] = 32'b11111111111111100000010000010110;
assign LUT_2[59965] = 32'b11111111111111011101001000101111;
assign LUT_2[59966] = 32'b11111111111111100111001001010010;
assign LUT_2[59967] = 32'b11111111111111100100000001101011;
assign LUT_2[59968] = 32'b11111111111111100110001010000001;
assign LUT_2[59969] = 32'b11111111111111100011000010011010;
assign LUT_2[59970] = 32'b11111111111111101101000010111101;
assign LUT_2[59971] = 32'b11111111111111101001111011010110;
assign LUT_2[59972] = 32'b11111111111111100010100111101001;
assign LUT_2[59973] = 32'b11111111111111011111100000000010;
assign LUT_2[59974] = 32'b11111111111111101001100000100101;
assign LUT_2[59975] = 32'b11111111111111100110011000111110;
assign LUT_2[59976] = 32'b11111111111111100000111011011110;
assign LUT_2[59977] = 32'b11111111111111011101110011110111;
assign LUT_2[59978] = 32'b11111111111111100111110100011010;
assign LUT_2[59979] = 32'b11111111111111100100101100110011;
assign LUT_2[59980] = 32'b11111111111111011101011001000110;
assign LUT_2[59981] = 32'b11111111111111011010010001011111;
assign LUT_2[59982] = 32'b11111111111111100100010010000010;
assign LUT_2[59983] = 32'b11111111111111100001001010011011;
assign LUT_2[59984] = 32'b11111111111111100000101110001011;
assign LUT_2[59985] = 32'b11111111111111011101100110100100;
assign LUT_2[59986] = 32'b11111111111111100111100111000111;
assign LUT_2[59987] = 32'b11111111111111100100011111100000;
assign LUT_2[59988] = 32'b11111111111111011101001011110011;
assign LUT_2[59989] = 32'b11111111111111011010000100001100;
assign LUT_2[59990] = 32'b11111111111111100100000100101111;
assign LUT_2[59991] = 32'b11111111111111100000111101001000;
assign LUT_2[59992] = 32'b11111111111111011011011111101000;
assign LUT_2[59993] = 32'b11111111111111011000011000000001;
assign LUT_2[59994] = 32'b11111111111111100010011000100100;
assign LUT_2[59995] = 32'b11111111111111011111010000111101;
assign LUT_2[59996] = 32'b11111111111111010111111101010000;
assign LUT_2[59997] = 32'b11111111111111010100110101101001;
assign LUT_2[59998] = 32'b11111111111111011110110110001100;
assign LUT_2[59999] = 32'b11111111111111011011101110100101;
assign LUT_2[60000] = 32'b11111111111111100110100101101010;
assign LUT_2[60001] = 32'b11111111111111100011011110000011;
assign LUT_2[60002] = 32'b11111111111111101101011110100110;
assign LUT_2[60003] = 32'b11111111111111101010010110111111;
assign LUT_2[60004] = 32'b11111111111111100011000011010010;
assign LUT_2[60005] = 32'b11111111111111011111111011101011;
assign LUT_2[60006] = 32'b11111111111111101001111100001110;
assign LUT_2[60007] = 32'b11111111111111100110110100100111;
assign LUT_2[60008] = 32'b11111111111111100001010111000111;
assign LUT_2[60009] = 32'b11111111111111011110001111100000;
assign LUT_2[60010] = 32'b11111111111111101000010000000011;
assign LUT_2[60011] = 32'b11111111111111100101001000011100;
assign LUT_2[60012] = 32'b11111111111111011101110100101111;
assign LUT_2[60013] = 32'b11111111111111011010101101001000;
assign LUT_2[60014] = 32'b11111111111111100100101101101011;
assign LUT_2[60015] = 32'b11111111111111100001100110000100;
assign LUT_2[60016] = 32'b11111111111111100001001001110100;
assign LUT_2[60017] = 32'b11111111111111011110000010001101;
assign LUT_2[60018] = 32'b11111111111111101000000010110000;
assign LUT_2[60019] = 32'b11111111111111100100111011001001;
assign LUT_2[60020] = 32'b11111111111111011101100111011100;
assign LUT_2[60021] = 32'b11111111111111011010011111110101;
assign LUT_2[60022] = 32'b11111111111111100100100000011000;
assign LUT_2[60023] = 32'b11111111111111100001011000110001;
assign LUT_2[60024] = 32'b11111111111111011011111011010001;
assign LUT_2[60025] = 32'b11111111111111011000110011101010;
assign LUT_2[60026] = 32'b11111111111111100010110100001101;
assign LUT_2[60027] = 32'b11111111111111011111101100100110;
assign LUT_2[60028] = 32'b11111111111111011000011000111001;
assign LUT_2[60029] = 32'b11111111111111010101010001010010;
assign LUT_2[60030] = 32'b11111111111111011111010001110101;
assign LUT_2[60031] = 32'b11111111111111011100001010001110;
assign LUT_2[60032] = 32'b11111111111111110010010101101101;
assign LUT_2[60033] = 32'b11111111111111101111001110000110;
assign LUT_2[60034] = 32'b11111111111111111001001110101001;
assign LUT_2[60035] = 32'b11111111111111110110000111000010;
assign LUT_2[60036] = 32'b11111111111111101110110011010101;
assign LUT_2[60037] = 32'b11111111111111101011101011101110;
assign LUT_2[60038] = 32'b11111111111111110101101100010001;
assign LUT_2[60039] = 32'b11111111111111110010100100101010;
assign LUT_2[60040] = 32'b11111111111111101101000111001010;
assign LUT_2[60041] = 32'b11111111111111101001111111100011;
assign LUT_2[60042] = 32'b11111111111111110100000000000110;
assign LUT_2[60043] = 32'b11111111111111110000111000011111;
assign LUT_2[60044] = 32'b11111111111111101001100100110010;
assign LUT_2[60045] = 32'b11111111111111100110011101001011;
assign LUT_2[60046] = 32'b11111111111111110000011101101110;
assign LUT_2[60047] = 32'b11111111111111101101010110000111;
assign LUT_2[60048] = 32'b11111111111111101100111001110111;
assign LUT_2[60049] = 32'b11111111111111101001110010010000;
assign LUT_2[60050] = 32'b11111111111111110011110010110011;
assign LUT_2[60051] = 32'b11111111111111110000101011001100;
assign LUT_2[60052] = 32'b11111111111111101001010111011111;
assign LUT_2[60053] = 32'b11111111111111100110001111111000;
assign LUT_2[60054] = 32'b11111111111111110000010000011011;
assign LUT_2[60055] = 32'b11111111111111101101001000110100;
assign LUT_2[60056] = 32'b11111111111111100111101011010100;
assign LUT_2[60057] = 32'b11111111111111100100100011101101;
assign LUT_2[60058] = 32'b11111111111111101110100100010000;
assign LUT_2[60059] = 32'b11111111111111101011011100101001;
assign LUT_2[60060] = 32'b11111111111111100100001000111100;
assign LUT_2[60061] = 32'b11111111111111100001000001010101;
assign LUT_2[60062] = 32'b11111111111111101011000001111000;
assign LUT_2[60063] = 32'b11111111111111100111111010010001;
assign LUT_2[60064] = 32'b11111111111111110010110001010110;
assign LUT_2[60065] = 32'b11111111111111101111101001101111;
assign LUT_2[60066] = 32'b11111111111111111001101010010010;
assign LUT_2[60067] = 32'b11111111111111110110100010101011;
assign LUT_2[60068] = 32'b11111111111111101111001110111110;
assign LUT_2[60069] = 32'b11111111111111101100000111010111;
assign LUT_2[60070] = 32'b11111111111111110110000111111010;
assign LUT_2[60071] = 32'b11111111111111110011000000010011;
assign LUT_2[60072] = 32'b11111111111111101101100010110011;
assign LUT_2[60073] = 32'b11111111111111101010011011001100;
assign LUT_2[60074] = 32'b11111111111111110100011011101111;
assign LUT_2[60075] = 32'b11111111111111110001010100001000;
assign LUT_2[60076] = 32'b11111111111111101010000000011011;
assign LUT_2[60077] = 32'b11111111111111100110111000110100;
assign LUT_2[60078] = 32'b11111111111111110000111001010111;
assign LUT_2[60079] = 32'b11111111111111101101110001110000;
assign LUT_2[60080] = 32'b11111111111111101101010101100000;
assign LUT_2[60081] = 32'b11111111111111101010001101111001;
assign LUT_2[60082] = 32'b11111111111111110100001110011100;
assign LUT_2[60083] = 32'b11111111111111110001000110110101;
assign LUT_2[60084] = 32'b11111111111111101001110011001000;
assign LUT_2[60085] = 32'b11111111111111100110101011100001;
assign LUT_2[60086] = 32'b11111111111111110000101100000100;
assign LUT_2[60087] = 32'b11111111111111101101100100011101;
assign LUT_2[60088] = 32'b11111111111111101000000110111101;
assign LUT_2[60089] = 32'b11111111111111100100111111010110;
assign LUT_2[60090] = 32'b11111111111111101110111111111001;
assign LUT_2[60091] = 32'b11111111111111101011111000010010;
assign LUT_2[60092] = 32'b11111111111111100100100100100101;
assign LUT_2[60093] = 32'b11111111111111100001011100111110;
assign LUT_2[60094] = 32'b11111111111111101011011101100001;
assign LUT_2[60095] = 32'b11111111111111101000010101111010;
assign LUT_2[60096] = 32'b11111111111111101010011110010000;
assign LUT_2[60097] = 32'b11111111111111100111010110101001;
assign LUT_2[60098] = 32'b11111111111111110001010111001100;
assign LUT_2[60099] = 32'b11111111111111101110001111100101;
assign LUT_2[60100] = 32'b11111111111111100110111011111000;
assign LUT_2[60101] = 32'b11111111111111100011110100010001;
assign LUT_2[60102] = 32'b11111111111111101101110100110100;
assign LUT_2[60103] = 32'b11111111111111101010101101001101;
assign LUT_2[60104] = 32'b11111111111111100101001111101101;
assign LUT_2[60105] = 32'b11111111111111100010001000000110;
assign LUT_2[60106] = 32'b11111111111111101100001000101001;
assign LUT_2[60107] = 32'b11111111111111101001000001000010;
assign LUT_2[60108] = 32'b11111111111111100001101101010101;
assign LUT_2[60109] = 32'b11111111111111011110100101101110;
assign LUT_2[60110] = 32'b11111111111111101000100110010001;
assign LUT_2[60111] = 32'b11111111111111100101011110101010;
assign LUT_2[60112] = 32'b11111111111111100101000010011010;
assign LUT_2[60113] = 32'b11111111111111100001111010110011;
assign LUT_2[60114] = 32'b11111111111111101011111011010110;
assign LUT_2[60115] = 32'b11111111111111101000110011101111;
assign LUT_2[60116] = 32'b11111111111111100001100000000010;
assign LUT_2[60117] = 32'b11111111111111011110011000011011;
assign LUT_2[60118] = 32'b11111111111111101000011000111110;
assign LUT_2[60119] = 32'b11111111111111100101010001010111;
assign LUT_2[60120] = 32'b11111111111111011111110011110111;
assign LUT_2[60121] = 32'b11111111111111011100101100010000;
assign LUT_2[60122] = 32'b11111111111111100110101100110011;
assign LUT_2[60123] = 32'b11111111111111100011100101001100;
assign LUT_2[60124] = 32'b11111111111111011100010001011111;
assign LUT_2[60125] = 32'b11111111111111011001001001111000;
assign LUT_2[60126] = 32'b11111111111111100011001010011011;
assign LUT_2[60127] = 32'b11111111111111100000000010110100;
assign LUT_2[60128] = 32'b11111111111111101010111001111001;
assign LUT_2[60129] = 32'b11111111111111100111110010010010;
assign LUT_2[60130] = 32'b11111111111111110001110010110101;
assign LUT_2[60131] = 32'b11111111111111101110101011001110;
assign LUT_2[60132] = 32'b11111111111111100111010111100001;
assign LUT_2[60133] = 32'b11111111111111100100001111111010;
assign LUT_2[60134] = 32'b11111111111111101110010000011101;
assign LUT_2[60135] = 32'b11111111111111101011001000110110;
assign LUT_2[60136] = 32'b11111111111111100101101011010110;
assign LUT_2[60137] = 32'b11111111111111100010100011101111;
assign LUT_2[60138] = 32'b11111111111111101100100100010010;
assign LUT_2[60139] = 32'b11111111111111101001011100101011;
assign LUT_2[60140] = 32'b11111111111111100010001000111110;
assign LUT_2[60141] = 32'b11111111111111011111000001010111;
assign LUT_2[60142] = 32'b11111111111111101001000001111010;
assign LUT_2[60143] = 32'b11111111111111100101111010010011;
assign LUT_2[60144] = 32'b11111111111111100101011110000011;
assign LUT_2[60145] = 32'b11111111111111100010010110011100;
assign LUT_2[60146] = 32'b11111111111111101100010110111111;
assign LUT_2[60147] = 32'b11111111111111101001001111011000;
assign LUT_2[60148] = 32'b11111111111111100001111011101011;
assign LUT_2[60149] = 32'b11111111111111011110110100000100;
assign LUT_2[60150] = 32'b11111111111111101000110100100111;
assign LUT_2[60151] = 32'b11111111111111100101101101000000;
assign LUT_2[60152] = 32'b11111111111111100000001111100000;
assign LUT_2[60153] = 32'b11111111111111011101000111111001;
assign LUT_2[60154] = 32'b11111111111111100111001000011100;
assign LUT_2[60155] = 32'b11111111111111100100000000110101;
assign LUT_2[60156] = 32'b11111111111111011100101101001000;
assign LUT_2[60157] = 32'b11111111111111011001100101100001;
assign LUT_2[60158] = 32'b11111111111111100011100110000100;
assign LUT_2[60159] = 32'b11111111111111100000011110011101;
assign LUT_2[60160] = 32'b11111111111111110010000000000100;
assign LUT_2[60161] = 32'b11111111111111101110111000011101;
assign LUT_2[60162] = 32'b11111111111111111000111001000000;
assign LUT_2[60163] = 32'b11111111111111110101110001011001;
assign LUT_2[60164] = 32'b11111111111111101110011101101100;
assign LUT_2[60165] = 32'b11111111111111101011010110000101;
assign LUT_2[60166] = 32'b11111111111111110101010110101000;
assign LUT_2[60167] = 32'b11111111111111110010001111000001;
assign LUT_2[60168] = 32'b11111111111111101100110001100001;
assign LUT_2[60169] = 32'b11111111111111101001101001111010;
assign LUT_2[60170] = 32'b11111111111111110011101010011101;
assign LUT_2[60171] = 32'b11111111111111110000100010110110;
assign LUT_2[60172] = 32'b11111111111111101001001111001001;
assign LUT_2[60173] = 32'b11111111111111100110000111100010;
assign LUT_2[60174] = 32'b11111111111111110000001000000101;
assign LUT_2[60175] = 32'b11111111111111101101000000011110;
assign LUT_2[60176] = 32'b11111111111111101100100100001110;
assign LUT_2[60177] = 32'b11111111111111101001011100100111;
assign LUT_2[60178] = 32'b11111111111111110011011101001010;
assign LUT_2[60179] = 32'b11111111111111110000010101100011;
assign LUT_2[60180] = 32'b11111111111111101001000001110110;
assign LUT_2[60181] = 32'b11111111111111100101111010001111;
assign LUT_2[60182] = 32'b11111111111111101111111010110010;
assign LUT_2[60183] = 32'b11111111111111101100110011001011;
assign LUT_2[60184] = 32'b11111111111111100111010101101011;
assign LUT_2[60185] = 32'b11111111111111100100001110000100;
assign LUT_2[60186] = 32'b11111111111111101110001110100111;
assign LUT_2[60187] = 32'b11111111111111101011000111000000;
assign LUT_2[60188] = 32'b11111111111111100011110011010011;
assign LUT_2[60189] = 32'b11111111111111100000101011101100;
assign LUT_2[60190] = 32'b11111111111111101010101100001111;
assign LUT_2[60191] = 32'b11111111111111100111100100101000;
assign LUT_2[60192] = 32'b11111111111111110010011011101101;
assign LUT_2[60193] = 32'b11111111111111101111010100000110;
assign LUT_2[60194] = 32'b11111111111111111001010100101001;
assign LUT_2[60195] = 32'b11111111111111110110001101000010;
assign LUT_2[60196] = 32'b11111111111111101110111001010101;
assign LUT_2[60197] = 32'b11111111111111101011110001101110;
assign LUT_2[60198] = 32'b11111111111111110101110010010001;
assign LUT_2[60199] = 32'b11111111111111110010101010101010;
assign LUT_2[60200] = 32'b11111111111111101101001101001010;
assign LUT_2[60201] = 32'b11111111111111101010000101100011;
assign LUT_2[60202] = 32'b11111111111111110100000110000110;
assign LUT_2[60203] = 32'b11111111111111110000111110011111;
assign LUT_2[60204] = 32'b11111111111111101001101010110010;
assign LUT_2[60205] = 32'b11111111111111100110100011001011;
assign LUT_2[60206] = 32'b11111111111111110000100011101110;
assign LUT_2[60207] = 32'b11111111111111101101011100000111;
assign LUT_2[60208] = 32'b11111111111111101100111111110111;
assign LUT_2[60209] = 32'b11111111111111101001111000010000;
assign LUT_2[60210] = 32'b11111111111111110011111000110011;
assign LUT_2[60211] = 32'b11111111111111110000110001001100;
assign LUT_2[60212] = 32'b11111111111111101001011101011111;
assign LUT_2[60213] = 32'b11111111111111100110010101111000;
assign LUT_2[60214] = 32'b11111111111111110000010110011011;
assign LUT_2[60215] = 32'b11111111111111101101001110110100;
assign LUT_2[60216] = 32'b11111111111111100111110001010100;
assign LUT_2[60217] = 32'b11111111111111100100101001101101;
assign LUT_2[60218] = 32'b11111111111111101110101010010000;
assign LUT_2[60219] = 32'b11111111111111101011100010101001;
assign LUT_2[60220] = 32'b11111111111111100100001110111100;
assign LUT_2[60221] = 32'b11111111111111100001000111010101;
assign LUT_2[60222] = 32'b11111111111111101011000111111000;
assign LUT_2[60223] = 32'b11111111111111101000000000010001;
assign LUT_2[60224] = 32'b11111111111111101010001000100111;
assign LUT_2[60225] = 32'b11111111111111100111000001000000;
assign LUT_2[60226] = 32'b11111111111111110001000001100011;
assign LUT_2[60227] = 32'b11111111111111101101111001111100;
assign LUT_2[60228] = 32'b11111111111111100110100110001111;
assign LUT_2[60229] = 32'b11111111111111100011011110101000;
assign LUT_2[60230] = 32'b11111111111111101101011111001011;
assign LUT_2[60231] = 32'b11111111111111101010010111100100;
assign LUT_2[60232] = 32'b11111111111111100100111010000100;
assign LUT_2[60233] = 32'b11111111111111100001110010011101;
assign LUT_2[60234] = 32'b11111111111111101011110011000000;
assign LUT_2[60235] = 32'b11111111111111101000101011011001;
assign LUT_2[60236] = 32'b11111111111111100001010111101100;
assign LUT_2[60237] = 32'b11111111111111011110010000000101;
assign LUT_2[60238] = 32'b11111111111111101000010000101000;
assign LUT_2[60239] = 32'b11111111111111100101001001000001;
assign LUT_2[60240] = 32'b11111111111111100100101100110001;
assign LUT_2[60241] = 32'b11111111111111100001100101001010;
assign LUT_2[60242] = 32'b11111111111111101011100101101101;
assign LUT_2[60243] = 32'b11111111111111101000011110000110;
assign LUT_2[60244] = 32'b11111111111111100001001010011001;
assign LUT_2[60245] = 32'b11111111111111011110000010110010;
assign LUT_2[60246] = 32'b11111111111111101000000011010101;
assign LUT_2[60247] = 32'b11111111111111100100111011101110;
assign LUT_2[60248] = 32'b11111111111111011111011110001110;
assign LUT_2[60249] = 32'b11111111111111011100010110100111;
assign LUT_2[60250] = 32'b11111111111111100110010111001010;
assign LUT_2[60251] = 32'b11111111111111100011001111100011;
assign LUT_2[60252] = 32'b11111111111111011011111011110110;
assign LUT_2[60253] = 32'b11111111111111011000110100001111;
assign LUT_2[60254] = 32'b11111111111111100010110100110010;
assign LUT_2[60255] = 32'b11111111111111011111101101001011;
assign LUT_2[60256] = 32'b11111111111111101010100100010000;
assign LUT_2[60257] = 32'b11111111111111100111011100101001;
assign LUT_2[60258] = 32'b11111111111111110001011101001100;
assign LUT_2[60259] = 32'b11111111111111101110010101100101;
assign LUT_2[60260] = 32'b11111111111111100111000001111000;
assign LUT_2[60261] = 32'b11111111111111100011111010010001;
assign LUT_2[60262] = 32'b11111111111111101101111010110100;
assign LUT_2[60263] = 32'b11111111111111101010110011001101;
assign LUT_2[60264] = 32'b11111111111111100101010101101101;
assign LUT_2[60265] = 32'b11111111111111100010001110000110;
assign LUT_2[60266] = 32'b11111111111111101100001110101001;
assign LUT_2[60267] = 32'b11111111111111101001000111000010;
assign LUT_2[60268] = 32'b11111111111111100001110011010101;
assign LUT_2[60269] = 32'b11111111111111011110101011101110;
assign LUT_2[60270] = 32'b11111111111111101000101100010001;
assign LUT_2[60271] = 32'b11111111111111100101100100101010;
assign LUT_2[60272] = 32'b11111111111111100101001000011010;
assign LUT_2[60273] = 32'b11111111111111100010000000110011;
assign LUT_2[60274] = 32'b11111111111111101100000001010110;
assign LUT_2[60275] = 32'b11111111111111101000111001101111;
assign LUT_2[60276] = 32'b11111111111111100001100110000010;
assign LUT_2[60277] = 32'b11111111111111011110011110011011;
assign LUT_2[60278] = 32'b11111111111111101000011110111110;
assign LUT_2[60279] = 32'b11111111111111100101010111010111;
assign LUT_2[60280] = 32'b11111111111111011111111001110111;
assign LUT_2[60281] = 32'b11111111111111011100110010010000;
assign LUT_2[60282] = 32'b11111111111111100110110010110011;
assign LUT_2[60283] = 32'b11111111111111100011101011001100;
assign LUT_2[60284] = 32'b11111111111111011100010111011111;
assign LUT_2[60285] = 32'b11111111111111011001001111111000;
assign LUT_2[60286] = 32'b11111111111111100011010000011011;
assign LUT_2[60287] = 32'b11111111111111100000001000110100;
assign LUT_2[60288] = 32'b11111111111111110110010100010011;
assign LUT_2[60289] = 32'b11111111111111110011001100101100;
assign LUT_2[60290] = 32'b11111111111111111101001101001111;
assign LUT_2[60291] = 32'b11111111111111111010000101101000;
assign LUT_2[60292] = 32'b11111111111111110010110001111011;
assign LUT_2[60293] = 32'b11111111111111101111101010010100;
assign LUT_2[60294] = 32'b11111111111111111001101010110111;
assign LUT_2[60295] = 32'b11111111111111110110100011010000;
assign LUT_2[60296] = 32'b11111111111111110001000101110000;
assign LUT_2[60297] = 32'b11111111111111101101111110001001;
assign LUT_2[60298] = 32'b11111111111111110111111110101100;
assign LUT_2[60299] = 32'b11111111111111110100110111000101;
assign LUT_2[60300] = 32'b11111111111111101101100011011000;
assign LUT_2[60301] = 32'b11111111111111101010011011110001;
assign LUT_2[60302] = 32'b11111111111111110100011100010100;
assign LUT_2[60303] = 32'b11111111111111110001010100101101;
assign LUT_2[60304] = 32'b11111111111111110000111000011101;
assign LUT_2[60305] = 32'b11111111111111101101110000110110;
assign LUT_2[60306] = 32'b11111111111111110111110001011001;
assign LUT_2[60307] = 32'b11111111111111110100101001110010;
assign LUT_2[60308] = 32'b11111111111111101101010110000101;
assign LUT_2[60309] = 32'b11111111111111101010001110011110;
assign LUT_2[60310] = 32'b11111111111111110100001111000001;
assign LUT_2[60311] = 32'b11111111111111110001000111011010;
assign LUT_2[60312] = 32'b11111111111111101011101001111010;
assign LUT_2[60313] = 32'b11111111111111101000100010010011;
assign LUT_2[60314] = 32'b11111111111111110010100010110110;
assign LUT_2[60315] = 32'b11111111111111101111011011001111;
assign LUT_2[60316] = 32'b11111111111111101000000111100010;
assign LUT_2[60317] = 32'b11111111111111100100111111111011;
assign LUT_2[60318] = 32'b11111111111111101111000000011110;
assign LUT_2[60319] = 32'b11111111111111101011111000110111;
assign LUT_2[60320] = 32'b11111111111111110110101111111100;
assign LUT_2[60321] = 32'b11111111111111110011101000010101;
assign LUT_2[60322] = 32'b11111111111111111101101000111000;
assign LUT_2[60323] = 32'b11111111111111111010100001010001;
assign LUT_2[60324] = 32'b11111111111111110011001101100100;
assign LUT_2[60325] = 32'b11111111111111110000000101111101;
assign LUT_2[60326] = 32'b11111111111111111010000110100000;
assign LUT_2[60327] = 32'b11111111111111110110111110111001;
assign LUT_2[60328] = 32'b11111111111111110001100001011001;
assign LUT_2[60329] = 32'b11111111111111101110011001110010;
assign LUT_2[60330] = 32'b11111111111111111000011010010101;
assign LUT_2[60331] = 32'b11111111111111110101010010101110;
assign LUT_2[60332] = 32'b11111111111111101101111111000001;
assign LUT_2[60333] = 32'b11111111111111101010110111011010;
assign LUT_2[60334] = 32'b11111111111111110100110111111101;
assign LUT_2[60335] = 32'b11111111111111110001110000010110;
assign LUT_2[60336] = 32'b11111111111111110001010100000110;
assign LUT_2[60337] = 32'b11111111111111101110001100011111;
assign LUT_2[60338] = 32'b11111111111111111000001101000010;
assign LUT_2[60339] = 32'b11111111111111110101000101011011;
assign LUT_2[60340] = 32'b11111111111111101101110001101110;
assign LUT_2[60341] = 32'b11111111111111101010101010000111;
assign LUT_2[60342] = 32'b11111111111111110100101010101010;
assign LUT_2[60343] = 32'b11111111111111110001100011000011;
assign LUT_2[60344] = 32'b11111111111111101100000101100011;
assign LUT_2[60345] = 32'b11111111111111101000111101111100;
assign LUT_2[60346] = 32'b11111111111111110010111110011111;
assign LUT_2[60347] = 32'b11111111111111101111110110111000;
assign LUT_2[60348] = 32'b11111111111111101000100011001011;
assign LUT_2[60349] = 32'b11111111111111100101011011100100;
assign LUT_2[60350] = 32'b11111111111111101111011100000111;
assign LUT_2[60351] = 32'b11111111111111101100010100100000;
assign LUT_2[60352] = 32'b11111111111111101110011100110110;
assign LUT_2[60353] = 32'b11111111111111101011010101001111;
assign LUT_2[60354] = 32'b11111111111111110101010101110010;
assign LUT_2[60355] = 32'b11111111111111110010001110001011;
assign LUT_2[60356] = 32'b11111111111111101010111010011110;
assign LUT_2[60357] = 32'b11111111111111100111110010110111;
assign LUT_2[60358] = 32'b11111111111111110001110011011010;
assign LUT_2[60359] = 32'b11111111111111101110101011110011;
assign LUT_2[60360] = 32'b11111111111111101001001110010011;
assign LUT_2[60361] = 32'b11111111111111100110000110101100;
assign LUT_2[60362] = 32'b11111111111111110000000111001111;
assign LUT_2[60363] = 32'b11111111111111101100111111101000;
assign LUT_2[60364] = 32'b11111111111111100101101011111011;
assign LUT_2[60365] = 32'b11111111111111100010100100010100;
assign LUT_2[60366] = 32'b11111111111111101100100100110111;
assign LUT_2[60367] = 32'b11111111111111101001011101010000;
assign LUT_2[60368] = 32'b11111111111111101001000001000000;
assign LUT_2[60369] = 32'b11111111111111100101111001011001;
assign LUT_2[60370] = 32'b11111111111111101111111001111100;
assign LUT_2[60371] = 32'b11111111111111101100110010010101;
assign LUT_2[60372] = 32'b11111111111111100101011110101000;
assign LUT_2[60373] = 32'b11111111111111100010010111000001;
assign LUT_2[60374] = 32'b11111111111111101100010111100100;
assign LUT_2[60375] = 32'b11111111111111101001001111111101;
assign LUT_2[60376] = 32'b11111111111111100011110010011101;
assign LUT_2[60377] = 32'b11111111111111100000101010110110;
assign LUT_2[60378] = 32'b11111111111111101010101011011001;
assign LUT_2[60379] = 32'b11111111111111100111100011110010;
assign LUT_2[60380] = 32'b11111111111111100000010000000101;
assign LUT_2[60381] = 32'b11111111111111011101001000011110;
assign LUT_2[60382] = 32'b11111111111111100111001001000001;
assign LUT_2[60383] = 32'b11111111111111100100000001011010;
assign LUT_2[60384] = 32'b11111111111111101110111000011111;
assign LUT_2[60385] = 32'b11111111111111101011110000111000;
assign LUT_2[60386] = 32'b11111111111111110101110001011011;
assign LUT_2[60387] = 32'b11111111111111110010101001110100;
assign LUT_2[60388] = 32'b11111111111111101011010110000111;
assign LUT_2[60389] = 32'b11111111111111101000001110100000;
assign LUT_2[60390] = 32'b11111111111111110010001111000011;
assign LUT_2[60391] = 32'b11111111111111101111000111011100;
assign LUT_2[60392] = 32'b11111111111111101001101001111100;
assign LUT_2[60393] = 32'b11111111111111100110100010010101;
assign LUT_2[60394] = 32'b11111111111111110000100010111000;
assign LUT_2[60395] = 32'b11111111111111101101011011010001;
assign LUT_2[60396] = 32'b11111111111111100110000111100100;
assign LUT_2[60397] = 32'b11111111111111100010111111111101;
assign LUT_2[60398] = 32'b11111111111111101101000000100000;
assign LUT_2[60399] = 32'b11111111111111101001111000111001;
assign LUT_2[60400] = 32'b11111111111111101001011100101001;
assign LUT_2[60401] = 32'b11111111111111100110010101000010;
assign LUT_2[60402] = 32'b11111111111111110000010101100101;
assign LUT_2[60403] = 32'b11111111111111101101001101111110;
assign LUT_2[60404] = 32'b11111111111111100101111010010001;
assign LUT_2[60405] = 32'b11111111111111100010110010101010;
assign LUT_2[60406] = 32'b11111111111111101100110011001101;
assign LUT_2[60407] = 32'b11111111111111101001101011100110;
assign LUT_2[60408] = 32'b11111111111111100100001110000110;
assign LUT_2[60409] = 32'b11111111111111100001000110011111;
assign LUT_2[60410] = 32'b11111111111111101011000111000010;
assign LUT_2[60411] = 32'b11111111111111100111111111011011;
assign LUT_2[60412] = 32'b11111111111111100000101011101110;
assign LUT_2[60413] = 32'b11111111111111011101100100000111;
assign LUT_2[60414] = 32'b11111111111111100111100100101010;
assign LUT_2[60415] = 32'b11111111111111100100011101000011;
assign LUT_2[60416] = 32'b11111111111111101111111011110001;
assign LUT_2[60417] = 32'b11111111111111101100110100001010;
assign LUT_2[60418] = 32'b11111111111111110110110100101101;
assign LUT_2[60419] = 32'b11111111111111110011101101000110;
assign LUT_2[60420] = 32'b11111111111111101100011001011001;
assign LUT_2[60421] = 32'b11111111111111101001010001110010;
assign LUT_2[60422] = 32'b11111111111111110011010010010101;
assign LUT_2[60423] = 32'b11111111111111110000001010101110;
assign LUT_2[60424] = 32'b11111111111111101010101101001110;
assign LUT_2[60425] = 32'b11111111111111100111100101100111;
assign LUT_2[60426] = 32'b11111111111111110001100110001010;
assign LUT_2[60427] = 32'b11111111111111101110011110100011;
assign LUT_2[60428] = 32'b11111111111111100111001010110110;
assign LUT_2[60429] = 32'b11111111111111100100000011001111;
assign LUT_2[60430] = 32'b11111111111111101110000011110010;
assign LUT_2[60431] = 32'b11111111111111101010111100001011;
assign LUT_2[60432] = 32'b11111111111111101010011111111011;
assign LUT_2[60433] = 32'b11111111111111100111011000010100;
assign LUT_2[60434] = 32'b11111111111111110001011000110111;
assign LUT_2[60435] = 32'b11111111111111101110010001010000;
assign LUT_2[60436] = 32'b11111111111111100110111101100011;
assign LUT_2[60437] = 32'b11111111111111100011110101111100;
assign LUT_2[60438] = 32'b11111111111111101101110110011111;
assign LUT_2[60439] = 32'b11111111111111101010101110111000;
assign LUT_2[60440] = 32'b11111111111111100101010001011000;
assign LUT_2[60441] = 32'b11111111111111100010001001110001;
assign LUT_2[60442] = 32'b11111111111111101100001010010100;
assign LUT_2[60443] = 32'b11111111111111101001000010101101;
assign LUT_2[60444] = 32'b11111111111111100001101111000000;
assign LUT_2[60445] = 32'b11111111111111011110100111011001;
assign LUT_2[60446] = 32'b11111111111111101000100111111100;
assign LUT_2[60447] = 32'b11111111111111100101100000010101;
assign LUT_2[60448] = 32'b11111111111111110000010111011010;
assign LUT_2[60449] = 32'b11111111111111101101001111110011;
assign LUT_2[60450] = 32'b11111111111111110111010000010110;
assign LUT_2[60451] = 32'b11111111111111110100001000101111;
assign LUT_2[60452] = 32'b11111111111111101100110101000010;
assign LUT_2[60453] = 32'b11111111111111101001101101011011;
assign LUT_2[60454] = 32'b11111111111111110011101101111110;
assign LUT_2[60455] = 32'b11111111111111110000100110010111;
assign LUT_2[60456] = 32'b11111111111111101011001000110111;
assign LUT_2[60457] = 32'b11111111111111101000000001010000;
assign LUT_2[60458] = 32'b11111111111111110010000001110011;
assign LUT_2[60459] = 32'b11111111111111101110111010001100;
assign LUT_2[60460] = 32'b11111111111111100111100110011111;
assign LUT_2[60461] = 32'b11111111111111100100011110111000;
assign LUT_2[60462] = 32'b11111111111111101110011111011011;
assign LUT_2[60463] = 32'b11111111111111101011010111110100;
assign LUT_2[60464] = 32'b11111111111111101010111011100100;
assign LUT_2[60465] = 32'b11111111111111100111110011111101;
assign LUT_2[60466] = 32'b11111111111111110001110100100000;
assign LUT_2[60467] = 32'b11111111111111101110101100111001;
assign LUT_2[60468] = 32'b11111111111111100111011001001100;
assign LUT_2[60469] = 32'b11111111111111100100010001100101;
assign LUT_2[60470] = 32'b11111111111111101110010010001000;
assign LUT_2[60471] = 32'b11111111111111101011001010100001;
assign LUT_2[60472] = 32'b11111111111111100101101101000001;
assign LUT_2[60473] = 32'b11111111111111100010100101011010;
assign LUT_2[60474] = 32'b11111111111111101100100101111101;
assign LUT_2[60475] = 32'b11111111111111101001011110010110;
assign LUT_2[60476] = 32'b11111111111111100010001010101001;
assign LUT_2[60477] = 32'b11111111111111011111000011000010;
assign LUT_2[60478] = 32'b11111111111111101001000011100101;
assign LUT_2[60479] = 32'b11111111111111100101111011111110;
assign LUT_2[60480] = 32'b11111111111111101000000100010100;
assign LUT_2[60481] = 32'b11111111111111100100111100101101;
assign LUT_2[60482] = 32'b11111111111111101110111101010000;
assign LUT_2[60483] = 32'b11111111111111101011110101101001;
assign LUT_2[60484] = 32'b11111111111111100100100001111100;
assign LUT_2[60485] = 32'b11111111111111100001011010010101;
assign LUT_2[60486] = 32'b11111111111111101011011010111000;
assign LUT_2[60487] = 32'b11111111111111101000010011010001;
assign LUT_2[60488] = 32'b11111111111111100010110101110001;
assign LUT_2[60489] = 32'b11111111111111011111101110001010;
assign LUT_2[60490] = 32'b11111111111111101001101110101101;
assign LUT_2[60491] = 32'b11111111111111100110100111000110;
assign LUT_2[60492] = 32'b11111111111111011111010011011001;
assign LUT_2[60493] = 32'b11111111111111011100001011110010;
assign LUT_2[60494] = 32'b11111111111111100110001100010101;
assign LUT_2[60495] = 32'b11111111111111100011000100101110;
assign LUT_2[60496] = 32'b11111111111111100010101000011110;
assign LUT_2[60497] = 32'b11111111111111011111100000110111;
assign LUT_2[60498] = 32'b11111111111111101001100001011010;
assign LUT_2[60499] = 32'b11111111111111100110011001110011;
assign LUT_2[60500] = 32'b11111111111111011111000110000110;
assign LUT_2[60501] = 32'b11111111111111011011111110011111;
assign LUT_2[60502] = 32'b11111111111111100101111111000010;
assign LUT_2[60503] = 32'b11111111111111100010110111011011;
assign LUT_2[60504] = 32'b11111111111111011101011001111011;
assign LUT_2[60505] = 32'b11111111111111011010010010010100;
assign LUT_2[60506] = 32'b11111111111111100100010010110111;
assign LUT_2[60507] = 32'b11111111111111100001001011010000;
assign LUT_2[60508] = 32'b11111111111111011001110111100011;
assign LUT_2[60509] = 32'b11111111111111010110101111111100;
assign LUT_2[60510] = 32'b11111111111111100000110000011111;
assign LUT_2[60511] = 32'b11111111111111011101101000111000;
assign LUT_2[60512] = 32'b11111111111111101000011111111101;
assign LUT_2[60513] = 32'b11111111111111100101011000010110;
assign LUT_2[60514] = 32'b11111111111111101111011000111001;
assign LUT_2[60515] = 32'b11111111111111101100010001010010;
assign LUT_2[60516] = 32'b11111111111111100100111101100101;
assign LUT_2[60517] = 32'b11111111111111100001110101111110;
assign LUT_2[60518] = 32'b11111111111111101011110110100001;
assign LUT_2[60519] = 32'b11111111111111101000101110111010;
assign LUT_2[60520] = 32'b11111111111111100011010001011010;
assign LUT_2[60521] = 32'b11111111111111100000001001110011;
assign LUT_2[60522] = 32'b11111111111111101010001010010110;
assign LUT_2[60523] = 32'b11111111111111100111000010101111;
assign LUT_2[60524] = 32'b11111111111111011111101111000010;
assign LUT_2[60525] = 32'b11111111111111011100100111011011;
assign LUT_2[60526] = 32'b11111111111111100110100111111110;
assign LUT_2[60527] = 32'b11111111111111100011100000010111;
assign LUT_2[60528] = 32'b11111111111111100011000100000111;
assign LUT_2[60529] = 32'b11111111111111011111111100100000;
assign LUT_2[60530] = 32'b11111111111111101001111101000011;
assign LUT_2[60531] = 32'b11111111111111100110110101011100;
assign LUT_2[60532] = 32'b11111111111111011111100001101111;
assign LUT_2[60533] = 32'b11111111111111011100011010001000;
assign LUT_2[60534] = 32'b11111111111111100110011010101011;
assign LUT_2[60535] = 32'b11111111111111100011010011000100;
assign LUT_2[60536] = 32'b11111111111111011101110101100100;
assign LUT_2[60537] = 32'b11111111111111011010101101111101;
assign LUT_2[60538] = 32'b11111111111111100100101110100000;
assign LUT_2[60539] = 32'b11111111111111100001100110111001;
assign LUT_2[60540] = 32'b11111111111111011010010011001100;
assign LUT_2[60541] = 32'b11111111111111010111001011100101;
assign LUT_2[60542] = 32'b11111111111111100001001100001000;
assign LUT_2[60543] = 32'b11111111111111011110000100100001;
assign LUT_2[60544] = 32'b11111111111111110100010000000000;
assign LUT_2[60545] = 32'b11111111111111110001001000011001;
assign LUT_2[60546] = 32'b11111111111111111011001000111100;
assign LUT_2[60547] = 32'b11111111111111111000000001010101;
assign LUT_2[60548] = 32'b11111111111111110000101101101000;
assign LUT_2[60549] = 32'b11111111111111101101100110000001;
assign LUT_2[60550] = 32'b11111111111111110111100110100100;
assign LUT_2[60551] = 32'b11111111111111110100011110111101;
assign LUT_2[60552] = 32'b11111111111111101111000001011101;
assign LUT_2[60553] = 32'b11111111111111101011111001110110;
assign LUT_2[60554] = 32'b11111111111111110101111010011001;
assign LUT_2[60555] = 32'b11111111111111110010110010110010;
assign LUT_2[60556] = 32'b11111111111111101011011111000101;
assign LUT_2[60557] = 32'b11111111111111101000010111011110;
assign LUT_2[60558] = 32'b11111111111111110010011000000001;
assign LUT_2[60559] = 32'b11111111111111101111010000011010;
assign LUT_2[60560] = 32'b11111111111111101110110100001010;
assign LUT_2[60561] = 32'b11111111111111101011101100100011;
assign LUT_2[60562] = 32'b11111111111111110101101101000110;
assign LUT_2[60563] = 32'b11111111111111110010100101011111;
assign LUT_2[60564] = 32'b11111111111111101011010001110010;
assign LUT_2[60565] = 32'b11111111111111101000001010001011;
assign LUT_2[60566] = 32'b11111111111111110010001010101110;
assign LUT_2[60567] = 32'b11111111111111101111000011000111;
assign LUT_2[60568] = 32'b11111111111111101001100101100111;
assign LUT_2[60569] = 32'b11111111111111100110011110000000;
assign LUT_2[60570] = 32'b11111111111111110000011110100011;
assign LUT_2[60571] = 32'b11111111111111101101010110111100;
assign LUT_2[60572] = 32'b11111111111111100110000011001111;
assign LUT_2[60573] = 32'b11111111111111100010111011101000;
assign LUT_2[60574] = 32'b11111111111111101100111100001011;
assign LUT_2[60575] = 32'b11111111111111101001110100100100;
assign LUT_2[60576] = 32'b11111111111111110100101011101001;
assign LUT_2[60577] = 32'b11111111111111110001100100000010;
assign LUT_2[60578] = 32'b11111111111111111011100100100101;
assign LUT_2[60579] = 32'b11111111111111111000011100111110;
assign LUT_2[60580] = 32'b11111111111111110001001001010001;
assign LUT_2[60581] = 32'b11111111111111101110000001101010;
assign LUT_2[60582] = 32'b11111111111111111000000010001101;
assign LUT_2[60583] = 32'b11111111111111110100111010100110;
assign LUT_2[60584] = 32'b11111111111111101111011101000110;
assign LUT_2[60585] = 32'b11111111111111101100010101011111;
assign LUT_2[60586] = 32'b11111111111111110110010110000010;
assign LUT_2[60587] = 32'b11111111111111110011001110011011;
assign LUT_2[60588] = 32'b11111111111111101011111010101110;
assign LUT_2[60589] = 32'b11111111111111101000110011000111;
assign LUT_2[60590] = 32'b11111111111111110010110011101010;
assign LUT_2[60591] = 32'b11111111111111101111101100000011;
assign LUT_2[60592] = 32'b11111111111111101111001111110011;
assign LUT_2[60593] = 32'b11111111111111101100001000001100;
assign LUT_2[60594] = 32'b11111111111111110110001000101111;
assign LUT_2[60595] = 32'b11111111111111110011000001001000;
assign LUT_2[60596] = 32'b11111111111111101011101101011011;
assign LUT_2[60597] = 32'b11111111111111101000100101110100;
assign LUT_2[60598] = 32'b11111111111111110010100110010111;
assign LUT_2[60599] = 32'b11111111111111101111011110110000;
assign LUT_2[60600] = 32'b11111111111111101010000001010000;
assign LUT_2[60601] = 32'b11111111111111100110111001101001;
assign LUT_2[60602] = 32'b11111111111111110000111010001100;
assign LUT_2[60603] = 32'b11111111111111101101110010100101;
assign LUT_2[60604] = 32'b11111111111111100110011110111000;
assign LUT_2[60605] = 32'b11111111111111100011010111010001;
assign LUT_2[60606] = 32'b11111111111111101101010111110100;
assign LUT_2[60607] = 32'b11111111111111101010010000001101;
assign LUT_2[60608] = 32'b11111111111111101100011000100011;
assign LUT_2[60609] = 32'b11111111111111101001010000111100;
assign LUT_2[60610] = 32'b11111111111111110011010001011111;
assign LUT_2[60611] = 32'b11111111111111110000001001111000;
assign LUT_2[60612] = 32'b11111111111111101000110110001011;
assign LUT_2[60613] = 32'b11111111111111100101101110100100;
assign LUT_2[60614] = 32'b11111111111111101111101111000111;
assign LUT_2[60615] = 32'b11111111111111101100100111100000;
assign LUT_2[60616] = 32'b11111111111111100111001010000000;
assign LUT_2[60617] = 32'b11111111111111100100000010011001;
assign LUT_2[60618] = 32'b11111111111111101110000010111100;
assign LUT_2[60619] = 32'b11111111111111101010111011010101;
assign LUT_2[60620] = 32'b11111111111111100011100111101000;
assign LUT_2[60621] = 32'b11111111111111100000100000000001;
assign LUT_2[60622] = 32'b11111111111111101010100000100100;
assign LUT_2[60623] = 32'b11111111111111100111011000111101;
assign LUT_2[60624] = 32'b11111111111111100110111100101101;
assign LUT_2[60625] = 32'b11111111111111100011110101000110;
assign LUT_2[60626] = 32'b11111111111111101101110101101001;
assign LUT_2[60627] = 32'b11111111111111101010101110000010;
assign LUT_2[60628] = 32'b11111111111111100011011010010101;
assign LUT_2[60629] = 32'b11111111111111100000010010101110;
assign LUT_2[60630] = 32'b11111111111111101010010011010001;
assign LUT_2[60631] = 32'b11111111111111100111001011101010;
assign LUT_2[60632] = 32'b11111111111111100001101110001010;
assign LUT_2[60633] = 32'b11111111111111011110100110100011;
assign LUT_2[60634] = 32'b11111111111111101000100111000110;
assign LUT_2[60635] = 32'b11111111111111100101011111011111;
assign LUT_2[60636] = 32'b11111111111111011110001011110010;
assign LUT_2[60637] = 32'b11111111111111011011000100001011;
assign LUT_2[60638] = 32'b11111111111111100101000100101110;
assign LUT_2[60639] = 32'b11111111111111100001111101000111;
assign LUT_2[60640] = 32'b11111111111111101100110100001100;
assign LUT_2[60641] = 32'b11111111111111101001101100100101;
assign LUT_2[60642] = 32'b11111111111111110011101101001000;
assign LUT_2[60643] = 32'b11111111111111110000100101100001;
assign LUT_2[60644] = 32'b11111111111111101001010001110100;
assign LUT_2[60645] = 32'b11111111111111100110001010001101;
assign LUT_2[60646] = 32'b11111111111111110000001010110000;
assign LUT_2[60647] = 32'b11111111111111101101000011001001;
assign LUT_2[60648] = 32'b11111111111111100111100101101001;
assign LUT_2[60649] = 32'b11111111111111100100011110000010;
assign LUT_2[60650] = 32'b11111111111111101110011110100101;
assign LUT_2[60651] = 32'b11111111111111101011010110111110;
assign LUT_2[60652] = 32'b11111111111111100100000011010001;
assign LUT_2[60653] = 32'b11111111111111100000111011101010;
assign LUT_2[60654] = 32'b11111111111111101010111100001101;
assign LUT_2[60655] = 32'b11111111111111100111110100100110;
assign LUT_2[60656] = 32'b11111111111111100111011000010110;
assign LUT_2[60657] = 32'b11111111111111100100010000101111;
assign LUT_2[60658] = 32'b11111111111111101110010001010010;
assign LUT_2[60659] = 32'b11111111111111101011001001101011;
assign LUT_2[60660] = 32'b11111111111111100011110101111110;
assign LUT_2[60661] = 32'b11111111111111100000101110010111;
assign LUT_2[60662] = 32'b11111111111111101010101110111010;
assign LUT_2[60663] = 32'b11111111111111100111100111010011;
assign LUT_2[60664] = 32'b11111111111111100010001001110011;
assign LUT_2[60665] = 32'b11111111111111011111000010001100;
assign LUT_2[60666] = 32'b11111111111111101001000010101111;
assign LUT_2[60667] = 32'b11111111111111100101111011001000;
assign LUT_2[60668] = 32'b11111111111111011110100111011011;
assign LUT_2[60669] = 32'b11111111111111011011011111110100;
assign LUT_2[60670] = 32'b11111111111111100101100000010111;
assign LUT_2[60671] = 32'b11111111111111100010011000110000;
assign LUT_2[60672] = 32'b11111111111111110011111010010111;
assign LUT_2[60673] = 32'b11111111111111110000110010110000;
assign LUT_2[60674] = 32'b11111111111111111010110011010011;
assign LUT_2[60675] = 32'b11111111111111110111101011101100;
assign LUT_2[60676] = 32'b11111111111111110000010111111111;
assign LUT_2[60677] = 32'b11111111111111101101010000011000;
assign LUT_2[60678] = 32'b11111111111111110111010000111011;
assign LUT_2[60679] = 32'b11111111111111110100001001010100;
assign LUT_2[60680] = 32'b11111111111111101110101011110100;
assign LUT_2[60681] = 32'b11111111111111101011100100001101;
assign LUT_2[60682] = 32'b11111111111111110101100100110000;
assign LUT_2[60683] = 32'b11111111111111110010011101001001;
assign LUT_2[60684] = 32'b11111111111111101011001001011100;
assign LUT_2[60685] = 32'b11111111111111101000000001110101;
assign LUT_2[60686] = 32'b11111111111111110010000010011000;
assign LUT_2[60687] = 32'b11111111111111101110111010110001;
assign LUT_2[60688] = 32'b11111111111111101110011110100001;
assign LUT_2[60689] = 32'b11111111111111101011010110111010;
assign LUT_2[60690] = 32'b11111111111111110101010111011101;
assign LUT_2[60691] = 32'b11111111111111110010001111110110;
assign LUT_2[60692] = 32'b11111111111111101010111100001001;
assign LUT_2[60693] = 32'b11111111111111100111110100100010;
assign LUT_2[60694] = 32'b11111111111111110001110101000101;
assign LUT_2[60695] = 32'b11111111111111101110101101011110;
assign LUT_2[60696] = 32'b11111111111111101001001111111110;
assign LUT_2[60697] = 32'b11111111111111100110001000010111;
assign LUT_2[60698] = 32'b11111111111111110000001000111010;
assign LUT_2[60699] = 32'b11111111111111101101000001010011;
assign LUT_2[60700] = 32'b11111111111111100101101101100110;
assign LUT_2[60701] = 32'b11111111111111100010100101111111;
assign LUT_2[60702] = 32'b11111111111111101100100110100010;
assign LUT_2[60703] = 32'b11111111111111101001011110111011;
assign LUT_2[60704] = 32'b11111111111111110100010110000000;
assign LUT_2[60705] = 32'b11111111111111110001001110011001;
assign LUT_2[60706] = 32'b11111111111111111011001110111100;
assign LUT_2[60707] = 32'b11111111111111111000000111010101;
assign LUT_2[60708] = 32'b11111111111111110000110011101000;
assign LUT_2[60709] = 32'b11111111111111101101101100000001;
assign LUT_2[60710] = 32'b11111111111111110111101100100100;
assign LUT_2[60711] = 32'b11111111111111110100100100111101;
assign LUT_2[60712] = 32'b11111111111111101111000111011101;
assign LUT_2[60713] = 32'b11111111111111101011111111110110;
assign LUT_2[60714] = 32'b11111111111111110110000000011001;
assign LUT_2[60715] = 32'b11111111111111110010111000110010;
assign LUT_2[60716] = 32'b11111111111111101011100101000101;
assign LUT_2[60717] = 32'b11111111111111101000011101011110;
assign LUT_2[60718] = 32'b11111111111111110010011110000001;
assign LUT_2[60719] = 32'b11111111111111101111010110011010;
assign LUT_2[60720] = 32'b11111111111111101110111010001010;
assign LUT_2[60721] = 32'b11111111111111101011110010100011;
assign LUT_2[60722] = 32'b11111111111111110101110011000110;
assign LUT_2[60723] = 32'b11111111111111110010101011011111;
assign LUT_2[60724] = 32'b11111111111111101011010111110010;
assign LUT_2[60725] = 32'b11111111111111101000010000001011;
assign LUT_2[60726] = 32'b11111111111111110010010000101110;
assign LUT_2[60727] = 32'b11111111111111101111001001000111;
assign LUT_2[60728] = 32'b11111111111111101001101011100111;
assign LUT_2[60729] = 32'b11111111111111100110100100000000;
assign LUT_2[60730] = 32'b11111111111111110000100100100011;
assign LUT_2[60731] = 32'b11111111111111101101011100111100;
assign LUT_2[60732] = 32'b11111111111111100110001001001111;
assign LUT_2[60733] = 32'b11111111111111100011000001101000;
assign LUT_2[60734] = 32'b11111111111111101101000010001011;
assign LUT_2[60735] = 32'b11111111111111101001111010100100;
assign LUT_2[60736] = 32'b11111111111111101100000010111010;
assign LUT_2[60737] = 32'b11111111111111101000111011010011;
assign LUT_2[60738] = 32'b11111111111111110010111011110110;
assign LUT_2[60739] = 32'b11111111111111101111110100001111;
assign LUT_2[60740] = 32'b11111111111111101000100000100010;
assign LUT_2[60741] = 32'b11111111111111100101011000111011;
assign LUT_2[60742] = 32'b11111111111111101111011001011110;
assign LUT_2[60743] = 32'b11111111111111101100010001110111;
assign LUT_2[60744] = 32'b11111111111111100110110100010111;
assign LUT_2[60745] = 32'b11111111111111100011101100110000;
assign LUT_2[60746] = 32'b11111111111111101101101101010011;
assign LUT_2[60747] = 32'b11111111111111101010100101101100;
assign LUT_2[60748] = 32'b11111111111111100011010001111111;
assign LUT_2[60749] = 32'b11111111111111100000001010011000;
assign LUT_2[60750] = 32'b11111111111111101010001010111011;
assign LUT_2[60751] = 32'b11111111111111100111000011010100;
assign LUT_2[60752] = 32'b11111111111111100110100111000100;
assign LUT_2[60753] = 32'b11111111111111100011011111011101;
assign LUT_2[60754] = 32'b11111111111111101101100000000000;
assign LUT_2[60755] = 32'b11111111111111101010011000011001;
assign LUT_2[60756] = 32'b11111111111111100011000100101100;
assign LUT_2[60757] = 32'b11111111111111011111111101000101;
assign LUT_2[60758] = 32'b11111111111111101001111101101000;
assign LUT_2[60759] = 32'b11111111111111100110110110000001;
assign LUT_2[60760] = 32'b11111111111111100001011000100001;
assign LUT_2[60761] = 32'b11111111111111011110010000111010;
assign LUT_2[60762] = 32'b11111111111111101000010001011101;
assign LUT_2[60763] = 32'b11111111111111100101001001110110;
assign LUT_2[60764] = 32'b11111111111111011101110110001001;
assign LUT_2[60765] = 32'b11111111111111011010101110100010;
assign LUT_2[60766] = 32'b11111111111111100100101111000101;
assign LUT_2[60767] = 32'b11111111111111100001100111011110;
assign LUT_2[60768] = 32'b11111111111111101100011110100011;
assign LUT_2[60769] = 32'b11111111111111101001010110111100;
assign LUT_2[60770] = 32'b11111111111111110011010111011111;
assign LUT_2[60771] = 32'b11111111111111110000001111111000;
assign LUT_2[60772] = 32'b11111111111111101000111100001011;
assign LUT_2[60773] = 32'b11111111111111100101110100100100;
assign LUT_2[60774] = 32'b11111111111111101111110101000111;
assign LUT_2[60775] = 32'b11111111111111101100101101100000;
assign LUT_2[60776] = 32'b11111111111111100111010000000000;
assign LUT_2[60777] = 32'b11111111111111100100001000011001;
assign LUT_2[60778] = 32'b11111111111111101110001000111100;
assign LUT_2[60779] = 32'b11111111111111101011000001010101;
assign LUT_2[60780] = 32'b11111111111111100011101101101000;
assign LUT_2[60781] = 32'b11111111111111100000100110000001;
assign LUT_2[60782] = 32'b11111111111111101010100110100100;
assign LUT_2[60783] = 32'b11111111111111100111011110111101;
assign LUT_2[60784] = 32'b11111111111111100111000010101101;
assign LUT_2[60785] = 32'b11111111111111100011111011000110;
assign LUT_2[60786] = 32'b11111111111111101101111011101001;
assign LUT_2[60787] = 32'b11111111111111101010110100000010;
assign LUT_2[60788] = 32'b11111111111111100011100000010101;
assign LUT_2[60789] = 32'b11111111111111100000011000101110;
assign LUT_2[60790] = 32'b11111111111111101010011001010001;
assign LUT_2[60791] = 32'b11111111111111100111010001101010;
assign LUT_2[60792] = 32'b11111111111111100001110100001010;
assign LUT_2[60793] = 32'b11111111111111011110101100100011;
assign LUT_2[60794] = 32'b11111111111111101000101101000110;
assign LUT_2[60795] = 32'b11111111111111100101100101011111;
assign LUT_2[60796] = 32'b11111111111111011110010001110010;
assign LUT_2[60797] = 32'b11111111111111011011001010001011;
assign LUT_2[60798] = 32'b11111111111111100101001010101110;
assign LUT_2[60799] = 32'b11111111111111100010000011000111;
assign LUT_2[60800] = 32'b11111111111111111000001110100110;
assign LUT_2[60801] = 32'b11111111111111110101000110111111;
assign LUT_2[60802] = 32'b11111111111111111111000111100010;
assign LUT_2[60803] = 32'b11111111111111111011111111111011;
assign LUT_2[60804] = 32'b11111111111111110100101100001110;
assign LUT_2[60805] = 32'b11111111111111110001100100100111;
assign LUT_2[60806] = 32'b11111111111111111011100101001010;
assign LUT_2[60807] = 32'b11111111111111111000011101100011;
assign LUT_2[60808] = 32'b11111111111111110011000000000011;
assign LUT_2[60809] = 32'b11111111111111101111111000011100;
assign LUT_2[60810] = 32'b11111111111111111001111000111111;
assign LUT_2[60811] = 32'b11111111111111110110110001011000;
assign LUT_2[60812] = 32'b11111111111111101111011101101011;
assign LUT_2[60813] = 32'b11111111111111101100010110000100;
assign LUT_2[60814] = 32'b11111111111111110110010110100111;
assign LUT_2[60815] = 32'b11111111111111110011001111000000;
assign LUT_2[60816] = 32'b11111111111111110010110010110000;
assign LUT_2[60817] = 32'b11111111111111101111101011001001;
assign LUT_2[60818] = 32'b11111111111111111001101011101100;
assign LUT_2[60819] = 32'b11111111111111110110100100000101;
assign LUT_2[60820] = 32'b11111111111111101111010000011000;
assign LUT_2[60821] = 32'b11111111111111101100001000110001;
assign LUT_2[60822] = 32'b11111111111111110110001001010100;
assign LUT_2[60823] = 32'b11111111111111110011000001101101;
assign LUT_2[60824] = 32'b11111111111111101101100100001101;
assign LUT_2[60825] = 32'b11111111111111101010011100100110;
assign LUT_2[60826] = 32'b11111111111111110100011101001001;
assign LUT_2[60827] = 32'b11111111111111110001010101100010;
assign LUT_2[60828] = 32'b11111111111111101010000001110101;
assign LUT_2[60829] = 32'b11111111111111100110111010001110;
assign LUT_2[60830] = 32'b11111111111111110000111010110001;
assign LUT_2[60831] = 32'b11111111111111101101110011001010;
assign LUT_2[60832] = 32'b11111111111111111000101010001111;
assign LUT_2[60833] = 32'b11111111111111110101100010101000;
assign LUT_2[60834] = 32'b11111111111111111111100011001011;
assign LUT_2[60835] = 32'b11111111111111111100011011100100;
assign LUT_2[60836] = 32'b11111111111111110101000111110111;
assign LUT_2[60837] = 32'b11111111111111110010000000010000;
assign LUT_2[60838] = 32'b11111111111111111100000000110011;
assign LUT_2[60839] = 32'b11111111111111111000111001001100;
assign LUT_2[60840] = 32'b11111111111111110011011011101100;
assign LUT_2[60841] = 32'b11111111111111110000010100000101;
assign LUT_2[60842] = 32'b11111111111111111010010100101000;
assign LUT_2[60843] = 32'b11111111111111110111001101000001;
assign LUT_2[60844] = 32'b11111111111111101111111001010100;
assign LUT_2[60845] = 32'b11111111111111101100110001101101;
assign LUT_2[60846] = 32'b11111111111111110110110010010000;
assign LUT_2[60847] = 32'b11111111111111110011101010101001;
assign LUT_2[60848] = 32'b11111111111111110011001110011001;
assign LUT_2[60849] = 32'b11111111111111110000000110110010;
assign LUT_2[60850] = 32'b11111111111111111010000111010101;
assign LUT_2[60851] = 32'b11111111111111110110111111101110;
assign LUT_2[60852] = 32'b11111111111111101111101100000001;
assign LUT_2[60853] = 32'b11111111111111101100100100011010;
assign LUT_2[60854] = 32'b11111111111111110110100100111101;
assign LUT_2[60855] = 32'b11111111111111110011011101010110;
assign LUT_2[60856] = 32'b11111111111111101101111111110110;
assign LUT_2[60857] = 32'b11111111111111101010111000001111;
assign LUT_2[60858] = 32'b11111111111111110100111000110010;
assign LUT_2[60859] = 32'b11111111111111110001110001001011;
assign LUT_2[60860] = 32'b11111111111111101010011101011110;
assign LUT_2[60861] = 32'b11111111111111100111010101110111;
assign LUT_2[60862] = 32'b11111111111111110001010110011010;
assign LUT_2[60863] = 32'b11111111111111101110001110110011;
assign LUT_2[60864] = 32'b11111111111111110000010111001001;
assign LUT_2[60865] = 32'b11111111111111101101001111100010;
assign LUT_2[60866] = 32'b11111111111111110111010000000101;
assign LUT_2[60867] = 32'b11111111111111110100001000011110;
assign LUT_2[60868] = 32'b11111111111111101100110100110001;
assign LUT_2[60869] = 32'b11111111111111101001101101001010;
assign LUT_2[60870] = 32'b11111111111111110011101101101101;
assign LUT_2[60871] = 32'b11111111111111110000100110000110;
assign LUT_2[60872] = 32'b11111111111111101011001000100110;
assign LUT_2[60873] = 32'b11111111111111101000000000111111;
assign LUT_2[60874] = 32'b11111111111111110010000001100010;
assign LUT_2[60875] = 32'b11111111111111101110111001111011;
assign LUT_2[60876] = 32'b11111111111111100111100110001110;
assign LUT_2[60877] = 32'b11111111111111100100011110100111;
assign LUT_2[60878] = 32'b11111111111111101110011111001010;
assign LUT_2[60879] = 32'b11111111111111101011010111100011;
assign LUT_2[60880] = 32'b11111111111111101010111011010011;
assign LUT_2[60881] = 32'b11111111111111100111110011101100;
assign LUT_2[60882] = 32'b11111111111111110001110100001111;
assign LUT_2[60883] = 32'b11111111111111101110101100101000;
assign LUT_2[60884] = 32'b11111111111111100111011000111011;
assign LUT_2[60885] = 32'b11111111111111100100010001010100;
assign LUT_2[60886] = 32'b11111111111111101110010001110111;
assign LUT_2[60887] = 32'b11111111111111101011001010010000;
assign LUT_2[60888] = 32'b11111111111111100101101100110000;
assign LUT_2[60889] = 32'b11111111111111100010100101001001;
assign LUT_2[60890] = 32'b11111111111111101100100101101100;
assign LUT_2[60891] = 32'b11111111111111101001011110000101;
assign LUT_2[60892] = 32'b11111111111111100010001010011000;
assign LUT_2[60893] = 32'b11111111111111011111000010110001;
assign LUT_2[60894] = 32'b11111111111111101001000011010100;
assign LUT_2[60895] = 32'b11111111111111100101111011101101;
assign LUT_2[60896] = 32'b11111111111111110000110010110010;
assign LUT_2[60897] = 32'b11111111111111101101101011001011;
assign LUT_2[60898] = 32'b11111111111111110111101011101110;
assign LUT_2[60899] = 32'b11111111111111110100100100000111;
assign LUT_2[60900] = 32'b11111111111111101101010000011010;
assign LUT_2[60901] = 32'b11111111111111101010001000110011;
assign LUT_2[60902] = 32'b11111111111111110100001001010110;
assign LUT_2[60903] = 32'b11111111111111110001000001101111;
assign LUT_2[60904] = 32'b11111111111111101011100100001111;
assign LUT_2[60905] = 32'b11111111111111101000011100101000;
assign LUT_2[60906] = 32'b11111111111111110010011101001011;
assign LUT_2[60907] = 32'b11111111111111101111010101100100;
assign LUT_2[60908] = 32'b11111111111111101000000001110111;
assign LUT_2[60909] = 32'b11111111111111100100111010010000;
assign LUT_2[60910] = 32'b11111111111111101110111010110011;
assign LUT_2[60911] = 32'b11111111111111101011110011001100;
assign LUT_2[60912] = 32'b11111111111111101011010110111100;
assign LUT_2[60913] = 32'b11111111111111101000001111010101;
assign LUT_2[60914] = 32'b11111111111111110010001111111000;
assign LUT_2[60915] = 32'b11111111111111101111001000010001;
assign LUT_2[60916] = 32'b11111111111111100111110100100100;
assign LUT_2[60917] = 32'b11111111111111100100101100111101;
assign LUT_2[60918] = 32'b11111111111111101110101101100000;
assign LUT_2[60919] = 32'b11111111111111101011100101111001;
assign LUT_2[60920] = 32'b11111111111111100110001000011001;
assign LUT_2[60921] = 32'b11111111111111100011000000110010;
assign LUT_2[60922] = 32'b11111111111111101101000001010101;
assign LUT_2[60923] = 32'b11111111111111101001111001101110;
assign LUT_2[60924] = 32'b11111111111111100010100110000001;
assign LUT_2[60925] = 32'b11111111111111011111011110011010;
assign LUT_2[60926] = 32'b11111111111111101001011110111101;
assign LUT_2[60927] = 32'b11111111111111100110010111010110;
assign LUT_2[60928] = 32'b11111111111111110100101101100011;
assign LUT_2[60929] = 32'b11111111111111110001100101111100;
assign LUT_2[60930] = 32'b11111111111111111011100110011111;
assign LUT_2[60931] = 32'b11111111111111111000011110111000;
assign LUT_2[60932] = 32'b11111111111111110001001011001011;
assign LUT_2[60933] = 32'b11111111111111101110000011100100;
assign LUT_2[60934] = 32'b11111111111111111000000100000111;
assign LUT_2[60935] = 32'b11111111111111110100111100100000;
assign LUT_2[60936] = 32'b11111111111111101111011111000000;
assign LUT_2[60937] = 32'b11111111111111101100010111011001;
assign LUT_2[60938] = 32'b11111111111111110110010111111100;
assign LUT_2[60939] = 32'b11111111111111110011010000010101;
assign LUT_2[60940] = 32'b11111111111111101011111100101000;
assign LUT_2[60941] = 32'b11111111111111101000110101000001;
assign LUT_2[60942] = 32'b11111111111111110010110101100100;
assign LUT_2[60943] = 32'b11111111111111101111101101111101;
assign LUT_2[60944] = 32'b11111111111111101111010001101101;
assign LUT_2[60945] = 32'b11111111111111101100001010000110;
assign LUT_2[60946] = 32'b11111111111111110110001010101001;
assign LUT_2[60947] = 32'b11111111111111110011000011000010;
assign LUT_2[60948] = 32'b11111111111111101011101111010101;
assign LUT_2[60949] = 32'b11111111111111101000100111101110;
assign LUT_2[60950] = 32'b11111111111111110010101000010001;
assign LUT_2[60951] = 32'b11111111111111101111100000101010;
assign LUT_2[60952] = 32'b11111111111111101010000011001010;
assign LUT_2[60953] = 32'b11111111111111100110111011100011;
assign LUT_2[60954] = 32'b11111111111111110000111100000110;
assign LUT_2[60955] = 32'b11111111111111101101110100011111;
assign LUT_2[60956] = 32'b11111111111111100110100000110010;
assign LUT_2[60957] = 32'b11111111111111100011011001001011;
assign LUT_2[60958] = 32'b11111111111111101101011001101110;
assign LUT_2[60959] = 32'b11111111111111101010010010000111;
assign LUT_2[60960] = 32'b11111111111111110101001001001100;
assign LUT_2[60961] = 32'b11111111111111110010000001100101;
assign LUT_2[60962] = 32'b11111111111111111100000010001000;
assign LUT_2[60963] = 32'b11111111111111111000111010100001;
assign LUT_2[60964] = 32'b11111111111111110001100110110100;
assign LUT_2[60965] = 32'b11111111111111101110011111001101;
assign LUT_2[60966] = 32'b11111111111111111000011111110000;
assign LUT_2[60967] = 32'b11111111111111110101011000001001;
assign LUT_2[60968] = 32'b11111111111111101111111010101001;
assign LUT_2[60969] = 32'b11111111111111101100110011000010;
assign LUT_2[60970] = 32'b11111111111111110110110011100101;
assign LUT_2[60971] = 32'b11111111111111110011101011111110;
assign LUT_2[60972] = 32'b11111111111111101100011000010001;
assign LUT_2[60973] = 32'b11111111111111101001010000101010;
assign LUT_2[60974] = 32'b11111111111111110011010001001101;
assign LUT_2[60975] = 32'b11111111111111110000001001100110;
assign LUT_2[60976] = 32'b11111111111111101111101101010110;
assign LUT_2[60977] = 32'b11111111111111101100100101101111;
assign LUT_2[60978] = 32'b11111111111111110110100110010010;
assign LUT_2[60979] = 32'b11111111111111110011011110101011;
assign LUT_2[60980] = 32'b11111111111111101100001010111110;
assign LUT_2[60981] = 32'b11111111111111101001000011010111;
assign LUT_2[60982] = 32'b11111111111111110011000011111010;
assign LUT_2[60983] = 32'b11111111111111101111111100010011;
assign LUT_2[60984] = 32'b11111111111111101010011110110011;
assign LUT_2[60985] = 32'b11111111111111100111010111001100;
assign LUT_2[60986] = 32'b11111111111111110001010111101111;
assign LUT_2[60987] = 32'b11111111111111101110010000001000;
assign LUT_2[60988] = 32'b11111111111111100110111100011011;
assign LUT_2[60989] = 32'b11111111111111100011110100110100;
assign LUT_2[60990] = 32'b11111111111111101101110101010111;
assign LUT_2[60991] = 32'b11111111111111101010101101110000;
assign LUT_2[60992] = 32'b11111111111111101100110110000110;
assign LUT_2[60993] = 32'b11111111111111101001101110011111;
assign LUT_2[60994] = 32'b11111111111111110011101111000010;
assign LUT_2[60995] = 32'b11111111111111110000100111011011;
assign LUT_2[60996] = 32'b11111111111111101001010011101110;
assign LUT_2[60997] = 32'b11111111111111100110001100000111;
assign LUT_2[60998] = 32'b11111111111111110000001100101010;
assign LUT_2[60999] = 32'b11111111111111101101000101000011;
assign LUT_2[61000] = 32'b11111111111111100111100111100011;
assign LUT_2[61001] = 32'b11111111111111100100011111111100;
assign LUT_2[61002] = 32'b11111111111111101110100000011111;
assign LUT_2[61003] = 32'b11111111111111101011011000111000;
assign LUT_2[61004] = 32'b11111111111111100100000101001011;
assign LUT_2[61005] = 32'b11111111111111100000111101100100;
assign LUT_2[61006] = 32'b11111111111111101010111110000111;
assign LUT_2[61007] = 32'b11111111111111100111110110100000;
assign LUT_2[61008] = 32'b11111111111111100111011010010000;
assign LUT_2[61009] = 32'b11111111111111100100010010101001;
assign LUT_2[61010] = 32'b11111111111111101110010011001100;
assign LUT_2[61011] = 32'b11111111111111101011001011100101;
assign LUT_2[61012] = 32'b11111111111111100011110111111000;
assign LUT_2[61013] = 32'b11111111111111100000110000010001;
assign LUT_2[61014] = 32'b11111111111111101010110000110100;
assign LUT_2[61015] = 32'b11111111111111100111101001001101;
assign LUT_2[61016] = 32'b11111111111111100010001011101101;
assign LUT_2[61017] = 32'b11111111111111011111000100000110;
assign LUT_2[61018] = 32'b11111111111111101001000100101001;
assign LUT_2[61019] = 32'b11111111111111100101111101000010;
assign LUT_2[61020] = 32'b11111111111111011110101001010101;
assign LUT_2[61021] = 32'b11111111111111011011100001101110;
assign LUT_2[61022] = 32'b11111111111111100101100010010001;
assign LUT_2[61023] = 32'b11111111111111100010011010101010;
assign LUT_2[61024] = 32'b11111111111111101101010001101111;
assign LUT_2[61025] = 32'b11111111111111101010001010001000;
assign LUT_2[61026] = 32'b11111111111111110100001010101011;
assign LUT_2[61027] = 32'b11111111111111110001000011000100;
assign LUT_2[61028] = 32'b11111111111111101001101111010111;
assign LUT_2[61029] = 32'b11111111111111100110100111110000;
assign LUT_2[61030] = 32'b11111111111111110000101000010011;
assign LUT_2[61031] = 32'b11111111111111101101100000101100;
assign LUT_2[61032] = 32'b11111111111111101000000011001100;
assign LUT_2[61033] = 32'b11111111111111100100111011100101;
assign LUT_2[61034] = 32'b11111111111111101110111100001000;
assign LUT_2[61035] = 32'b11111111111111101011110100100001;
assign LUT_2[61036] = 32'b11111111111111100100100000110100;
assign LUT_2[61037] = 32'b11111111111111100001011001001101;
assign LUT_2[61038] = 32'b11111111111111101011011001110000;
assign LUT_2[61039] = 32'b11111111111111101000010010001001;
assign LUT_2[61040] = 32'b11111111111111100111110101111001;
assign LUT_2[61041] = 32'b11111111111111100100101110010010;
assign LUT_2[61042] = 32'b11111111111111101110101110110101;
assign LUT_2[61043] = 32'b11111111111111101011100111001110;
assign LUT_2[61044] = 32'b11111111111111100100010011100001;
assign LUT_2[61045] = 32'b11111111111111100001001011111010;
assign LUT_2[61046] = 32'b11111111111111101011001100011101;
assign LUT_2[61047] = 32'b11111111111111101000000100110110;
assign LUT_2[61048] = 32'b11111111111111100010100111010110;
assign LUT_2[61049] = 32'b11111111111111011111011111101111;
assign LUT_2[61050] = 32'b11111111111111101001100000010010;
assign LUT_2[61051] = 32'b11111111111111100110011000101011;
assign LUT_2[61052] = 32'b11111111111111011111000100111110;
assign LUT_2[61053] = 32'b11111111111111011011111101010111;
assign LUT_2[61054] = 32'b11111111111111100101111101111010;
assign LUT_2[61055] = 32'b11111111111111100010110110010011;
assign LUT_2[61056] = 32'b11111111111111111001000001110010;
assign LUT_2[61057] = 32'b11111111111111110101111010001011;
assign LUT_2[61058] = 32'b11111111111111111111111010101110;
assign LUT_2[61059] = 32'b11111111111111111100110011000111;
assign LUT_2[61060] = 32'b11111111111111110101011111011010;
assign LUT_2[61061] = 32'b11111111111111110010010111110011;
assign LUT_2[61062] = 32'b11111111111111111100011000010110;
assign LUT_2[61063] = 32'b11111111111111111001010000101111;
assign LUT_2[61064] = 32'b11111111111111110011110011001111;
assign LUT_2[61065] = 32'b11111111111111110000101011101000;
assign LUT_2[61066] = 32'b11111111111111111010101100001011;
assign LUT_2[61067] = 32'b11111111111111110111100100100100;
assign LUT_2[61068] = 32'b11111111111111110000010000110111;
assign LUT_2[61069] = 32'b11111111111111101101001001010000;
assign LUT_2[61070] = 32'b11111111111111110111001001110011;
assign LUT_2[61071] = 32'b11111111111111110100000010001100;
assign LUT_2[61072] = 32'b11111111111111110011100101111100;
assign LUT_2[61073] = 32'b11111111111111110000011110010101;
assign LUT_2[61074] = 32'b11111111111111111010011110111000;
assign LUT_2[61075] = 32'b11111111111111110111010111010001;
assign LUT_2[61076] = 32'b11111111111111110000000011100100;
assign LUT_2[61077] = 32'b11111111111111101100111011111101;
assign LUT_2[61078] = 32'b11111111111111110110111100100000;
assign LUT_2[61079] = 32'b11111111111111110011110100111001;
assign LUT_2[61080] = 32'b11111111111111101110010111011001;
assign LUT_2[61081] = 32'b11111111111111101011001111110010;
assign LUT_2[61082] = 32'b11111111111111110101010000010101;
assign LUT_2[61083] = 32'b11111111111111110010001000101110;
assign LUT_2[61084] = 32'b11111111111111101010110101000001;
assign LUT_2[61085] = 32'b11111111111111100111101101011010;
assign LUT_2[61086] = 32'b11111111111111110001101101111101;
assign LUT_2[61087] = 32'b11111111111111101110100110010110;
assign LUT_2[61088] = 32'b11111111111111111001011101011011;
assign LUT_2[61089] = 32'b11111111111111110110010101110100;
assign LUT_2[61090] = 32'b00000000000000000000010110010111;
assign LUT_2[61091] = 32'b11111111111111111101001110110000;
assign LUT_2[61092] = 32'b11111111111111110101111011000011;
assign LUT_2[61093] = 32'b11111111111111110010110011011100;
assign LUT_2[61094] = 32'b11111111111111111100110011111111;
assign LUT_2[61095] = 32'b11111111111111111001101100011000;
assign LUT_2[61096] = 32'b11111111111111110100001110111000;
assign LUT_2[61097] = 32'b11111111111111110001000111010001;
assign LUT_2[61098] = 32'b11111111111111111011000111110100;
assign LUT_2[61099] = 32'b11111111111111111000000000001101;
assign LUT_2[61100] = 32'b11111111111111110000101100100000;
assign LUT_2[61101] = 32'b11111111111111101101100100111001;
assign LUT_2[61102] = 32'b11111111111111110111100101011100;
assign LUT_2[61103] = 32'b11111111111111110100011101110101;
assign LUT_2[61104] = 32'b11111111111111110100000001100101;
assign LUT_2[61105] = 32'b11111111111111110000111001111110;
assign LUT_2[61106] = 32'b11111111111111111010111010100001;
assign LUT_2[61107] = 32'b11111111111111110111110010111010;
assign LUT_2[61108] = 32'b11111111111111110000011111001101;
assign LUT_2[61109] = 32'b11111111111111101101010111100110;
assign LUT_2[61110] = 32'b11111111111111110111011000001001;
assign LUT_2[61111] = 32'b11111111111111110100010000100010;
assign LUT_2[61112] = 32'b11111111111111101110110011000010;
assign LUT_2[61113] = 32'b11111111111111101011101011011011;
assign LUT_2[61114] = 32'b11111111111111110101101011111110;
assign LUT_2[61115] = 32'b11111111111111110010100100010111;
assign LUT_2[61116] = 32'b11111111111111101011010000101010;
assign LUT_2[61117] = 32'b11111111111111101000001001000011;
assign LUT_2[61118] = 32'b11111111111111110010001001100110;
assign LUT_2[61119] = 32'b11111111111111101111000001111111;
assign LUT_2[61120] = 32'b11111111111111110001001010010101;
assign LUT_2[61121] = 32'b11111111111111101110000010101110;
assign LUT_2[61122] = 32'b11111111111111111000000011010001;
assign LUT_2[61123] = 32'b11111111111111110100111011101010;
assign LUT_2[61124] = 32'b11111111111111101101100111111101;
assign LUT_2[61125] = 32'b11111111111111101010100000010110;
assign LUT_2[61126] = 32'b11111111111111110100100000111001;
assign LUT_2[61127] = 32'b11111111111111110001011001010010;
assign LUT_2[61128] = 32'b11111111111111101011111011110010;
assign LUT_2[61129] = 32'b11111111111111101000110100001011;
assign LUT_2[61130] = 32'b11111111111111110010110100101110;
assign LUT_2[61131] = 32'b11111111111111101111101101000111;
assign LUT_2[61132] = 32'b11111111111111101000011001011010;
assign LUT_2[61133] = 32'b11111111111111100101010001110011;
assign LUT_2[61134] = 32'b11111111111111101111010010010110;
assign LUT_2[61135] = 32'b11111111111111101100001010101111;
assign LUT_2[61136] = 32'b11111111111111101011101110011111;
assign LUT_2[61137] = 32'b11111111111111101000100110111000;
assign LUT_2[61138] = 32'b11111111111111110010100111011011;
assign LUT_2[61139] = 32'b11111111111111101111011111110100;
assign LUT_2[61140] = 32'b11111111111111101000001100000111;
assign LUT_2[61141] = 32'b11111111111111100101000100100000;
assign LUT_2[61142] = 32'b11111111111111101111000101000011;
assign LUT_2[61143] = 32'b11111111111111101011111101011100;
assign LUT_2[61144] = 32'b11111111111111100110011111111100;
assign LUT_2[61145] = 32'b11111111111111100011011000010101;
assign LUT_2[61146] = 32'b11111111111111101101011000111000;
assign LUT_2[61147] = 32'b11111111111111101010010001010001;
assign LUT_2[61148] = 32'b11111111111111100010111101100100;
assign LUT_2[61149] = 32'b11111111111111011111110101111101;
assign LUT_2[61150] = 32'b11111111111111101001110110100000;
assign LUT_2[61151] = 32'b11111111111111100110101110111001;
assign LUT_2[61152] = 32'b11111111111111110001100101111110;
assign LUT_2[61153] = 32'b11111111111111101110011110010111;
assign LUT_2[61154] = 32'b11111111111111111000011110111010;
assign LUT_2[61155] = 32'b11111111111111110101010111010011;
assign LUT_2[61156] = 32'b11111111111111101110000011100110;
assign LUT_2[61157] = 32'b11111111111111101010111011111111;
assign LUT_2[61158] = 32'b11111111111111110100111100100010;
assign LUT_2[61159] = 32'b11111111111111110001110100111011;
assign LUT_2[61160] = 32'b11111111111111101100010111011011;
assign LUT_2[61161] = 32'b11111111111111101001001111110100;
assign LUT_2[61162] = 32'b11111111111111110011010000010111;
assign LUT_2[61163] = 32'b11111111111111110000001000110000;
assign LUT_2[61164] = 32'b11111111111111101000110101000011;
assign LUT_2[61165] = 32'b11111111111111100101101101011100;
assign LUT_2[61166] = 32'b11111111111111101111101101111111;
assign LUT_2[61167] = 32'b11111111111111101100100110011000;
assign LUT_2[61168] = 32'b11111111111111101100001010001000;
assign LUT_2[61169] = 32'b11111111111111101001000010100001;
assign LUT_2[61170] = 32'b11111111111111110011000011000100;
assign LUT_2[61171] = 32'b11111111111111101111111011011101;
assign LUT_2[61172] = 32'b11111111111111101000100111110000;
assign LUT_2[61173] = 32'b11111111111111100101100000001001;
assign LUT_2[61174] = 32'b11111111111111101111100000101100;
assign LUT_2[61175] = 32'b11111111111111101100011001000101;
assign LUT_2[61176] = 32'b11111111111111100110111011100101;
assign LUT_2[61177] = 32'b11111111111111100011110011111110;
assign LUT_2[61178] = 32'b11111111111111101101110100100001;
assign LUT_2[61179] = 32'b11111111111111101010101100111010;
assign LUT_2[61180] = 32'b11111111111111100011011001001101;
assign LUT_2[61181] = 32'b11111111111111100000010001100110;
assign LUT_2[61182] = 32'b11111111111111101010010010001001;
assign LUT_2[61183] = 32'b11111111111111100111001010100010;
assign LUT_2[61184] = 32'b11111111111111111000101100001001;
assign LUT_2[61185] = 32'b11111111111111110101100100100010;
assign LUT_2[61186] = 32'b11111111111111111111100101000101;
assign LUT_2[61187] = 32'b11111111111111111100011101011110;
assign LUT_2[61188] = 32'b11111111111111110101001001110001;
assign LUT_2[61189] = 32'b11111111111111110010000010001010;
assign LUT_2[61190] = 32'b11111111111111111100000010101101;
assign LUT_2[61191] = 32'b11111111111111111000111011000110;
assign LUT_2[61192] = 32'b11111111111111110011011101100110;
assign LUT_2[61193] = 32'b11111111111111110000010101111111;
assign LUT_2[61194] = 32'b11111111111111111010010110100010;
assign LUT_2[61195] = 32'b11111111111111110111001110111011;
assign LUT_2[61196] = 32'b11111111111111101111111011001110;
assign LUT_2[61197] = 32'b11111111111111101100110011100111;
assign LUT_2[61198] = 32'b11111111111111110110110100001010;
assign LUT_2[61199] = 32'b11111111111111110011101100100011;
assign LUT_2[61200] = 32'b11111111111111110011010000010011;
assign LUT_2[61201] = 32'b11111111111111110000001000101100;
assign LUT_2[61202] = 32'b11111111111111111010001001001111;
assign LUT_2[61203] = 32'b11111111111111110111000001101000;
assign LUT_2[61204] = 32'b11111111111111101111101101111011;
assign LUT_2[61205] = 32'b11111111111111101100100110010100;
assign LUT_2[61206] = 32'b11111111111111110110100110110111;
assign LUT_2[61207] = 32'b11111111111111110011011111010000;
assign LUT_2[61208] = 32'b11111111111111101110000001110000;
assign LUT_2[61209] = 32'b11111111111111101010111010001001;
assign LUT_2[61210] = 32'b11111111111111110100111010101100;
assign LUT_2[61211] = 32'b11111111111111110001110011000101;
assign LUT_2[61212] = 32'b11111111111111101010011111011000;
assign LUT_2[61213] = 32'b11111111111111100111010111110001;
assign LUT_2[61214] = 32'b11111111111111110001011000010100;
assign LUT_2[61215] = 32'b11111111111111101110010000101101;
assign LUT_2[61216] = 32'b11111111111111111001000111110010;
assign LUT_2[61217] = 32'b11111111111111110110000000001011;
assign LUT_2[61218] = 32'b00000000000000000000000000101110;
assign LUT_2[61219] = 32'b11111111111111111100111001000111;
assign LUT_2[61220] = 32'b11111111111111110101100101011010;
assign LUT_2[61221] = 32'b11111111111111110010011101110011;
assign LUT_2[61222] = 32'b11111111111111111100011110010110;
assign LUT_2[61223] = 32'b11111111111111111001010110101111;
assign LUT_2[61224] = 32'b11111111111111110011111001001111;
assign LUT_2[61225] = 32'b11111111111111110000110001101000;
assign LUT_2[61226] = 32'b11111111111111111010110010001011;
assign LUT_2[61227] = 32'b11111111111111110111101010100100;
assign LUT_2[61228] = 32'b11111111111111110000010110110111;
assign LUT_2[61229] = 32'b11111111111111101101001111010000;
assign LUT_2[61230] = 32'b11111111111111110111001111110011;
assign LUT_2[61231] = 32'b11111111111111110100001000001100;
assign LUT_2[61232] = 32'b11111111111111110011101011111100;
assign LUT_2[61233] = 32'b11111111111111110000100100010101;
assign LUT_2[61234] = 32'b11111111111111111010100100111000;
assign LUT_2[61235] = 32'b11111111111111110111011101010001;
assign LUT_2[61236] = 32'b11111111111111110000001001100100;
assign LUT_2[61237] = 32'b11111111111111101101000001111101;
assign LUT_2[61238] = 32'b11111111111111110111000010100000;
assign LUT_2[61239] = 32'b11111111111111110011111010111001;
assign LUT_2[61240] = 32'b11111111111111101110011101011001;
assign LUT_2[61241] = 32'b11111111111111101011010101110010;
assign LUT_2[61242] = 32'b11111111111111110101010110010101;
assign LUT_2[61243] = 32'b11111111111111110010001110101110;
assign LUT_2[61244] = 32'b11111111111111101010111011000001;
assign LUT_2[61245] = 32'b11111111111111100111110011011010;
assign LUT_2[61246] = 32'b11111111111111110001110011111101;
assign LUT_2[61247] = 32'b11111111111111101110101100010110;
assign LUT_2[61248] = 32'b11111111111111110000110100101100;
assign LUT_2[61249] = 32'b11111111111111101101101101000101;
assign LUT_2[61250] = 32'b11111111111111110111101101101000;
assign LUT_2[61251] = 32'b11111111111111110100100110000001;
assign LUT_2[61252] = 32'b11111111111111101101010010010100;
assign LUT_2[61253] = 32'b11111111111111101010001010101101;
assign LUT_2[61254] = 32'b11111111111111110100001011010000;
assign LUT_2[61255] = 32'b11111111111111110001000011101001;
assign LUT_2[61256] = 32'b11111111111111101011100110001001;
assign LUT_2[61257] = 32'b11111111111111101000011110100010;
assign LUT_2[61258] = 32'b11111111111111110010011111000101;
assign LUT_2[61259] = 32'b11111111111111101111010111011110;
assign LUT_2[61260] = 32'b11111111111111101000000011110001;
assign LUT_2[61261] = 32'b11111111111111100100111100001010;
assign LUT_2[61262] = 32'b11111111111111101110111100101101;
assign LUT_2[61263] = 32'b11111111111111101011110101000110;
assign LUT_2[61264] = 32'b11111111111111101011011000110110;
assign LUT_2[61265] = 32'b11111111111111101000010001001111;
assign LUT_2[61266] = 32'b11111111111111110010010001110010;
assign LUT_2[61267] = 32'b11111111111111101111001010001011;
assign LUT_2[61268] = 32'b11111111111111100111110110011110;
assign LUT_2[61269] = 32'b11111111111111100100101110110111;
assign LUT_2[61270] = 32'b11111111111111101110101111011010;
assign LUT_2[61271] = 32'b11111111111111101011100111110011;
assign LUT_2[61272] = 32'b11111111111111100110001010010011;
assign LUT_2[61273] = 32'b11111111111111100011000010101100;
assign LUT_2[61274] = 32'b11111111111111101101000011001111;
assign LUT_2[61275] = 32'b11111111111111101001111011101000;
assign LUT_2[61276] = 32'b11111111111111100010100111111011;
assign LUT_2[61277] = 32'b11111111111111011111100000010100;
assign LUT_2[61278] = 32'b11111111111111101001100000110111;
assign LUT_2[61279] = 32'b11111111111111100110011001010000;
assign LUT_2[61280] = 32'b11111111111111110001010000010101;
assign LUT_2[61281] = 32'b11111111111111101110001000101110;
assign LUT_2[61282] = 32'b11111111111111111000001001010001;
assign LUT_2[61283] = 32'b11111111111111110101000001101010;
assign LUT_2[61284] = 32'b11111111111111101101101101111101;
assign LUT_2[61285] = 32'b11111111111111101010100110010110;
assign LUT_2[61286] = 32'b11111111111111110100100110111001;
assign LUT_2[61287] = 32'b11111111111111110001011111010010;
assign LUT_2[61288] = 32'b11111111111111101100000001110010;
assign LUT_2[61289] = 32'b11111111111111101000111010001011;
assign LUT_2[61290] = 32'b11111111111111110010111010101110;
assign LUT_2[61291] = 32'b11111111111111101111110011000111;
assign LUT_2[61292] = 32'b11111111111111101000011111011010;
assign LUT_2[61293] = 32'b11111111111111100101010111110011;
assign LUT_2[61294] = 32'b11111111111111101111011000010110;
assign LUT_2[61295] = 32'b11111111111111101100010000101111;
assign LUT_2[61296] = 32'b11111111111111101011110100011111;
assign LUT_2[61297] = 32'b11111111111111101000101100111000;
assign LUT_2[61298] = 32'b11111111111111110010101101011011;
assign LUT_2[61299] = 32'b11111111111111101111100101110100;
assign LUT_2[61300] = 32'b11111111111111101000010010000111;
assign LUT_2[61301] = 32'b11111111111111100101001010100000;
assign LUT_2[61302] = 32'b11111111111111101111001011000011;
assign LUT_2[61303] = 32'b11111111111111101100000011011100;
assign LUT_2[61304] = 32'b11111111111111100110100101111100;
assign LUT_2[61305] = 32'b11111111111111100011011110010101;
assign LUT_2[61306] = 32'b11111111111111101101011110111000;
assign LUT_2[61307] = 32'b11111111111111101010010111010001;
assign LUT_2[61308] = 32'b11111111111111100011000011100100;
assign LUT_2[61309] = 32'b11111111111111011111111011111101;
assign LUT_2[61310] = 32'b11111111111111101001111100100000;
assign LUT_2[61311] = 32'b11111111111111100110110100111001;
assign LUT_2[61312] = 32'b11111111111111111101000000011000;
assign LUT_2[61313] = 32'b11111111111111111001111000110001;
assign LUT_2[61314] = 32'b00000000000000000011111001010100;
assign LUT_2[61315] = 32'b00000000000000000000110001101101;
assign LUT_2[61316] = 32'b11111111111111111001011110000000;
assign LUT_2[61317] = 32'b11111111111111110110010110011001;
assign LUT_2[61318] = 32'b00000000000000000000010110111100;
assign LUT_2[61319] = 32'b11111111111111111101001111010101;
assign LUT_2[61320] = 32'b11111111111111110111110001110101;
assign LUT_2[61321] = 32'b11111111111111110100101010001110;
assign LUT_2[61322] = 32'b11111111111111111110101010110001;
assign LUT_2[61323] = 32'b11111111111111111011100011001010;
assign LUT_2[61324] = 32'b11111111111111110100001111011101;
assign LUT_2[61325] = 32'b11111111111111110001000111110110;
assign LUT_2[61326] = 32'b11111111111111111011001000011001;
assign LUT_2[61327] = 32'b11111111111111111000000000110010;
assign LUT_2[61328] = 32'b11111111111111110111100100100010;
assign LUT_2[61329] = 32'b11111111111111110100011100111011;
assign LUT_2[61330] = 32'b11111111111111111110011101011110;
assign LUT_2[61331] = 32'b11111111111111111011010101110111;
assign LUT_2[61332] = 32'b11111111111111110100000010001010;
assign LUT_2[61333] = 32'b11111111111111110000111010100011;
assign LUT_2[61334] = 32'b11111111111111111010111011000110;
assign LUT_2[61335] = 32'b11111111111111110111110011011111;
assign LUT_2[61336] = 32'b11111111111111110010010101111111;
assign LUT_2[61337] = 32'b11111111111111101111001110011000;
assign LUT_2[61338] = 32'b11111111111111111001001110111011;
assign LUT_2[61339] = 32'b11111111111111110110000111010100;
assign LUT_2[61340] = 32'b11111111111111101110110011100111;
assign LUT_2[61341] = 32'b11111111111111101011101100000000;
assign LUT_2[61342] = 32'b11111111111111110101101100100011;
assign LUT_2[61343] = 32'b11111111111111110010100100111100;
assign LUT_2[61344] = 32'b11111111111111111101011100000001;
assign LUT_2[61345] = 32'b11111111111111111010010100011010;
assign LUT_2[61346] = 32'b00000000000000000100010100111101;
assign LUT_2[61347] = 32'b00000000000000000001001101010110;
assign LUT_2[61348] = 32'b11111111111111111001111001101001;
assign LUT_2[61349] = 32'b11111111111111110110110010000010;
assign LUT_2[61350] = 32'b00000000000000000000110010100101;
assign LUT_2[61351] = 32'b11111111111111111101101010111110;
assign LUT_2[61352] = 32'b11111111111111111000001101011110;
assign LUT_2[61353] = 32'b11111111111111110101000101110111;
assign LUT_2[61354] = 32'b11111111111111111111000110011010;
assign LUT_2[61355] = 32'b11111111111111111011111110110011;
assign LUT_2[61356] = 32'b11111111111111110100101011000110;
assign LUT_2[61357] = 32'b11111111111111110001100011011111;
assign LUT_2[61358] = 32'b11111111111111111011100100000010;
assign LUT_2[61359] = 32'b11111111111111111000011100011011;
assign LUT_2[61360] = 32'b11111111111111111000000000001011;
assign LUT_2[61361] = 32'b11111111111111110100111000100100;
assign LUT_2[61362] = 32'b11111111111111111110111001000111;
assign LUT_2[61363] = 32'b11111111111111111011110001100000;
assign LUT_2[61364] = 32'b11111111111111110100011101110011;
assign LUT_2[61365] = 32'b11111111111111110001010110001100;
assign LUT_2[61366] = 32'b11111111111111111011010110101111;
assign LUT_2[61367] = 32'b11111111111111111000001111001000;
assign LUT_2[61368] = 32'b11111111111111110010110001101000;
assign LUT_2[61369] = 32'b11111111111111101111101010000001;
assign LUT_2[61370] = 32'b11111111111111111001101010100100;
assign LUT_2[61371] = 32'b11111111111111110110100010111101;
assign LUT_2[61372] = 32'b11111111111111101111001111010000;
assign LUT_2[61373] = 32'b11111111111111101100000111101001;
assign LUT_2[61374] = 32'b11111111111111110110001000001100;
assign LUT_2[61375] = 32'b11111111111111110011000000100101;
assign LUT_2[61376] = 32'b11111111111111110101001000111011;
assign LUT_2[61377] = 32'b11111111111111110010000001010100;
assign LUT_2[61378] = 32'b11111111111111111100000001110111;
assign LUT_2[61379] = 32'b11111111111111111000111010010000;
assign LUT_2[61380] = 32'b11111111111111110001100110100011;
assign LUT_2[61381] = 32'b11111111111111101110011110111100;
assign LUT_2[61382] = 32'b11111111111111111000011111011111;
assign LUT_2[61383] = 32'b11111111111111110101010111111000;
assign LUT_2[61384] = 32'b11111111111111101111111010011000;
assign LUT_2[61385] = 32'b11111111111111101100110010110001;
assign LUT_2[61386] = 32'b11111111111111110110110011010100;
assign LUT_2[61387] = 32'b11111111111111110011101011101101;
assign LUT_2[61388] = 32'b11111111111111101100011000000000;
assign LUT_2[61389] = 32'b11111111111111101001010000011001;
assign LUT_2[61390] = 32'b11111111111111110011010000111100;
assign LUT_2[61391] = 32'b11111111111111110000001001010101;
assign LUT_2[61392] = 32'b11111111111111101111101101000101;
assign LUT_2[61393] = 32'b11111111111111101100100101011110;
assign LUT_2[61394] = 32'b11111111111111110110100110000001;
assign LUT_2[61395] = 32'b11111111111111110011011110011010;
assign LUT_2[61396] = 32'b11111111111111101100001010101101;
assign LUT_2[61397] = 32'b11111111111111101001000011000110;
assign LUT_2[61398] = 32'b11111111111111110011000011101001;
assign LUT_2[61399] = 32'b11111111111111101111111100000010;
assign LUT_2[61400] = 32'b11111111111111101010011110100010;
assign LUT_2[61401] = 32'b11111111111111100111010110111011;
assign LUT_2[61402] = 32'b11111111111111110001010111011110;
assign LUT_2[61403] = 32'b11111111111111101110001111110111;
assign LUT_2[61404] = 32'b11111111111111100110111100001010;
assign LUT_2[61405] = 32'b11111111111111100011110100100011;
assign LUT_2[61406] = 32'b11111111111111101101110101000110;
assign LUT_2[61407] = 32'b11111111111111101010101101011111;
assign LUT_2[61408] = 32'b11111111111111110101100100100100;
assign LUT_2[61409] = 32'b11111111111111110010011100111101;
assign LUT_2[61410] = 32'b11111111111111111100011101100000;
assign LUT_2[61411] = 32'b11111111111111111001010101111001;
assign LUT_2[61412] = 32'b11111111111111110010000010001100;
assign LUT_2[61413] = 32'b11111111111111101110111010100101;
assign LUT_2[61414] = 32'b11111111111111111000111011001000;
assign LUT_2[61415] = 32'b11111111111111110101110011100001;
assign LUT_2[61416] = 32'b11111111111111110000010110000001;
assign LUT_2[61417] = 32'b11111111111111101101001110011010;
assign LUT_2[61418] = 32'b11111111111111110111001110111101;
assign LUT_2[61419] = 32'b11111111111111110100000111010110;
assign LUT_2[61420] = 32'b11111111111111101100110011101001;
assign LUT_2[61421] = 32'b11111111111111101001101100000010;
assign LUT_2[61422] = 32'b11111111111111110011101100100101;
assign LUT_2[61423] = 32'b11111111111111110000100100111110;
assign LUT_2[61424] = 32'b11111111111111110000001000101110;
assign LUT_2[61425] = 32'b11111111111111101101000001000111;
assign LUT_2[61426] = 32'b11111111111111110111000001101010;
assign LUT_2[61427] = 32'b11111111111111110011111010000011;
assign LUT_2[61428] = 32'b11111111111111101100100110010110;
assign LUT_2[61429] = 32'b11111111111111101001011110101111;
assign LUT_2[61430] = 32'b11111111111111110011011111010010;
assign LUT_2[61431] = 32'b11111111111111110000010111101011;
assign LUT_2[61432] = 32'b11111111111111101010111010001011;
assign LUT_2[61433] = 32'b11111111111111100111110010100100;
assign LUT_2[61434] = 32'b11111111111111110001110011000111;
assign LUT_2[61435] = 32'b11111111111111101110101011100000;
assign LUT_2[61436] = 32'b11111111111111100111010111110011;
assign LUT_2[61437] = 32'b11111111111111100100010000001100;
assign LUT_2[61438] = 32'b11111111111111101110010000101111;
assign LUT_2[61439] = 32'b11111111111111101011001001001000;
assign LUT_2[61440] = 32'b11111111111111101100011101111011;
assign LUT_2[61441] = 32'b11111111111111101001010110010100;
assign LUT_2[61442] = 32'b11111111111111110011010110110111;
assign LUT_2[61443] = 32'b11111111111111110000001111010000;
assign LUT_2[61444] = 32'b11111111111111101000111011100011;
assign LUT_2[61445] = 32'b11111111111111100101110011111100;
assign LUT_2[61446] = 32'b11111111111111101111110100011111;
assign LUT_2[61447] = 32'b11111111111111101100101100111000;
assign LUT_2[61448] = 32'b11111111111111100111001111011000;
assign LUT_2[61449] = 32'b11111111111111100100000111110001;
assign LUT_2[61450] = 32'b11111111111111101110001000010100;
assign LUT_2[61451] = 32'b11111111111111101011000000101101;
assign LUT_2[61452] = 32'b11111111111111100011101101000000;
assign LUT_2[61453] = 32'b11111111111111100000100101011001;
assign LUT_2[61454] = 32'b11111111111111101010100101111100;
assign LUT_2[61455] = 32'b11111111111111100111011110010101;
assign LUT_2[61456] = 32'b11111111111111100111000010000101;
assign LUT_2[61457] = 32'b11111111111111100011111010011110;
assign LUT_2[61458] = 32'b11111111111111101101111011000001;
assign LUT_2[61459] = 32'b11111111111111101010110011011010;
assign LUT_2[61460] = 32'b11111111111111100011011111101101;
assign LUT_2[61461] = 32'b11111111111111100000011000000110;
assign LUT_2[61462] = 32'b11111111111111101010011000101001;
assign LUT_2[61463] = 32'b11111111111111100111010001000010;
assign LUT_2[61464] = 32'b11111111111111100001110011100010;
assign LUT_2[61465] = 32'b11111111111111011110101011111011;
assign LUT_2[61466] = 32'b11111111111111101000101100011110;
assign LUT_2[61467] = 32'b11111111111111100101100100110111;
assign LUT_2[61468] = 32'b11111111111111011110010001001010;
assign LUT_2[61469] = 32'b11111111111111011011001001100011;
assign LUT_2[61470] = 32'b11111111111111100101001010000110;
assign LUT_2[61471] = 32'b11111111111111100010000010011111;
assign LUT_2[61472] = 32'b11111111111111101100111001100100;
assign LUT_2[61473] = 32'b11111111111111101001110001111101;
assign LUT_2[61474] = 32'b11111111111111110011110010100000;
assign LUT_2[61475] = 32'b11111111111111110000101010111001;
assign LUT_2[61476] = 32'b11111111111111101001010111001100;
assign LUT_2[61477] = 32'b11111111111111100110001111100101;
assign LUT_2[61478] = 32'b11111111111111110000010000001000;
assign LUT_2[61479] = 32'b11111111111111101101001000100001;
assign LUT_2[61480] = 32'b11111111111111100111101011000001;
assign LUT_2[61481] = 32'b11111111111111100100100011011010;
assign LUT_2[61482] = 32'b11111111111111101110100011111101;
assign LUT_2[61483] = 32'b11111111111111101011011100010110;
assign LUT_2[61484] = 32'b11111111111111100100001000101001;
assign LUT_2[61485] = 32'b11111111111111100001000001000010;
assign LUT_2[61486] = 32'b11111111111111101011000001100101;
assign LUT_2[61487] = 32'b11111111111111100111111001111110;
assign LUT_2[61488] = 32'b11111111111111100111011101101110;
assign LUT_2[61489] = 32'b11111111111111100100010110000111;
assign LUT_2[61490] = 32'b11111111111111101110010110101010;
assign LUT_2[61491] = 32'b11111111111111101011001111000011;
assign LUT_2[61492] = 32'b11111111111111100011111011010110;
assign LUT_2[61493] = 32'b11111111111111100000110011101111;
assign LUT_2[61494] = 32'b11111111111111101010110100010010;
assign LUT_2[61495] = 32'b11111111111111100111101100101011;
assign LUT_2[61496] = 32'b11111111111111100010001111001011;
assign LUT_2[61497] = 32'b11111111111111011111000111100100;
assign LUT_2[61498] = 32'b11111111111111101001001000000111;
assign LUT_2[61499] = 32'b11111111111111100110000000100000;
assign LUT_2[61500] = 32'b11111111111111011110101100110011;
assign LUT_2[61501] = 32'b11111111111111011011100101001100;
assign LUT_2[61502] = 32'b11111111111111100101100101101111;
assign LUT_2[61503] = 32'b11111111111111100010011110001000;
assign LUT_2[61504] = 32'b11111111111111100100100110011110;
assign LUT_2[61505] = 32'b11111111111111100001011110110111;
assign LUT_2[61506] = 32'b11111111111111101011011111011010;
assign LUT_2[61507] = 32'b11111111111111101000010111110011;
assign LUT_2[61508] = 32'b11111111111111100001000100000110;
assign LUT_2[61509] = 32'b11111111111111011101111100011111;
assign LUT_2[61510] = 32'b11111111111111100111111101000010;
assign LUT_2[61511] = 32'b11111111111111100100110101011011;
assign LUT_2[61512] = 32'b11111111111111011111010111111011;
assign LUT_2[61513] = 32'b11111111111111011100010000010100;
assign LUT_2[61514] = 32'b11111111111111100110010000110111;
assign LUT_2[61515] = 32'b11111111111111100011001001010000;
assign LUT_2[61516] = 32'b11111111111111011011110101100011;
assign LUT_2[61517] = 32'b11111111111111011000101101111100;
assign LUT_2[61518] = 32'b11111111111111100010101110011111;
assign LUT_2[61519] = 32'b11111111111111011111100110111000;
assign LUT_2[61520] = 32'b11111111111111011111001010101000;
assign LUT_2[61521] = 32'b11111111111111011100000011000001;
assign LUT_2[61522] = 32'b11111111111111100110000011100100;
assign LUT_2[61523] = 32'b11111111111111100010111011111101;
assign LUT_2[61524] = 32'b11111111111111011011101000010000;
assign LUT_2[61525] = 32'b11111111111111011000100000101001;
assign LUT_2[61526] = 32'b11111111111111100010100001001100;
assign LUT_2[61527] = 32'b11111111111111011111011001100101;
assign LUT_2[61528] = 32'b11111111111111011001111100000101;
assign LUT_2[61529] = 32'b11111111111111010110110100011110;
assign LUT_2[61530] = 32'b11111111111111100000110101000001;
assign LUT_2[61531] = 32'b11111111111111011101101101011010;
assign LUT_2[61532] = 32'b11111111111111010110011001101101;
assign LUT_2[61533] = 32'b11111111111111010011010010000110;
assign LUT_2[61534] = 32'b11111111111111011101010010101001;
assign LUT_2[61535] = 32'b11111111111111011010001011000010;
assign LUT_2[61536] = 32'b11111111111111100101000010000111;
assign LUT_2[61537] = 32'b11111111111111100001111010100000;
assign LUT_2[61538] = 32'b11111111111111101011111011000011;
assign LUT_2[61539] = 32'b11111111111111101000110011011100;
assign LUT_2[61540] = 32'b11111111111111100001011111101111;
assign LUT_2[61541] = 32'b11111111111111011110011000001000;
assign LUT_2[61542] = 32'b11111111111111101000011000101011;
assign LUT_2[61543] = 32'b11111111111111100101010001000100;
assign LUT_2[61544] = 32'b11111111111111011111110011100100;
assign LUT_2[61545] = 32'b11111111111111011100101011111101;
assign LUT_2[61546] = 32'b11111111111111100110101100100000;
assign LUT_2[61547] = 32'b11111111111111100011100100111001;
assign LUT_2[61548] = 32'b11111111111111011100010001001100;
assign LUT_2[61549] = 32'b11111111111111011001001001100101;
assign LUT_2[61550] = 32'b11111111111111100011001010001000;
assign LUT_2[61551] = 32'b11111111111111100000000010100001;
assign LUT_2[61552] = 32'b11111111111111011111100110010001;
assign LUT_2[61553] = 32'b11111111111111011100011110101010;
assign LUT_2[61554] = 32'b11111111111111100110011111001101;
assign LUT_2[61555] = 32'b11111111111111100011010111100110;
assign LUT_2[61556] = 32'b11111111111111011100000011111001;
assign LUT_2[61557] = 32'b11111111111111011000111100010010;
assign LUT_2[61558] = 32'b11111111111111100010111100110101;
assign LUT_2[61559] = 32'b11111111111111011111110101001110;
assign LUT_2[61560] = 32'b11111111111111011010010111101110;
assign LUT_2[61561] = 32'b11111111111111010111010000000111;
assign LUT_2[61562] = 32'b11111111111111100001010000101010;
assign LUT_2[61563] = 32'b11111111111111011110001001000011;
assign LUT_2[61564] = 32'b11111111111111010110110101010110;
assign LUT_2[61565] = 32'b11111111111111010011101101101111;
assign LUT_2[61566] = 32'b11111111111111011101101110010010;
assign LUT_2[61567] = 32'b11111111111111011010100110101011;
assign LUT_2[61568] = 32'b11111111111111110000110010001010;
assign LUT_2[61569] = 32'b11111111111111101101101010100011;
assign LUT_2[61570] = 32'b11111111111111110111101011000110;
assign LUT_2[61571] = 32'b11111111111111110100100011011111;
assign LUT_2[61572] = 32'b11111111111111101101001111110010;
assign LUT_2[61573] = 32'b11111111111111101010001000001011;
assign LUT_2[61574] = 32'b11111111111111110100001000101110;
assign LUT_2[61575] = 32'b11111111111111110001000001000111;
assign LUT_2[61576] = 32'b11111111111111101011100011100111;
assign LUT_2[61577] = 32'b11111111111111101000011100000000;
assign LUT_2[61578] = 32'b11111111111111110010011100100011;
assign LUT_2[61579] = 32'b11111111111111101111010100111100;
assign LUT_2[61580] = 32'b11111111111111101000000001001111;
assign LUT_2[61581] = 32'b11111111111111100100111001101000;
assign LUT_2[61582] = 32'b11111111111111101110111010001011;
assign LUT_2[61583] = 32'b11111111111111101011110010100100;
assign LUT_2[61584] = 32'b11111111111111101011010110010100;
assign LUT_2[61585] = 32'b11111111111111101000001110101101;
assign LUT_2[61586] = 32'b11111111111111110010001111010000;
assign LUT_2[61587] = 32'b11111111111111101111000111101001;
assign LUT_2[61588] = 32'b11111111111111100111110011111100;
assign LUT_2[61589] = 32'b11111111111111100100101100010101;
assign LUT_2[61590] = 32'b11111111111111101110101100111000;
assign LUT_2[61591] = 32'b11111111111111101011100101010001;
assign LUT_2[61592] = 32'b11111111111111100110000111110001;
assign LUT_2[61593] = 32'b11111111111111100011000000001010;
assign LUT_2[61594] = 32'b11111111111111101101000000101101;
assign LUT_2[61595] = 32'b11111111111111101001111001000110;
assign LUT_2[61596] = 32'b11111111111111100010100101011001;
assign LUT_2[61597] = 32'b11111111111111011111011101110010;
assign LUT_2[61598] = 32'b11111111111111101001011110010101;
assign LUT_2[61599] = 32'b11111111111111100110010110101110;
assign LUT_2[61600] = 32'b11111111111111110001001101110011;
assign LUT_2[61601] = 32'b11111111111111101110000110001100;
assign LUT_2[61602] = 32'b11111111111111111000000110101111;
assign LUT_2[61603] = 32'b11111111111111110100111111001000;
assign LUT_2[61604] = 32'b11111111111111101101101011011011;
assign LUT_2[61605] = 32'b11111111111111101010100011110100;
assign LUT_2[61606] = 32'b11111111111111110100100100010111;
assign LUT_2[61607] = 32'b11111111111111110001011100110000;
assign LUT_2[61608] = 32'b11111111111111101011111111010000;
assign LUT_2[61609] = 32'b11111111111111101000110111101001;
assign LUT_2[61610] = 32'b11111111111111110010111000001100;
assign LUT_2[61611] = 32'b11111111111111101111110000100101;
assign LUT_2[61612] = 32'b11111111111111101000011100111000;
assign LUT_2[61613] = 32'b11111111111111100101010101010001;
assign LUT_2[61614] = 32'b11111111111111101111010101110100;
assign LUT_2[61615] = 32'b11111111111111101100001110001101;
assign LUT_2[61616] = 32'b11111111111111101011110001111101;
assign LUT_2[61617] = 32'b11111111111111101000101010010110;
assign LUT_2[61618] = 32'b11111111111111110010101010111001;
assign LUT_2[61619] = 32'b11111111111111101111100011010010;
assign LUT_2[61620] = 32'b11111111111111101000001111100101;
assign LUT_2[61621] = 32'b11111111111111100101000111111110;
assign LUT_2[61622] = 32'b11111111111111101111001000100001;
assign LUT_2[61623] = 32'b11111111111111101100000000111010;
assign LUT_2[61624] = 32'b11111111111111100110100011011010;
assign LUT_2[61625] = 32'b11111111111111100011011011110011;
assign LUT_2[61626] = 32'b11111111111111101101011100010110;
assign LUT_2[61627] = 32'b11111111111111101010010100101111;
assign LUT_2[61628] = 32'b11111111111111100011000001000010;
assign LUT_2[61629] = 32'b11111111111111011111111001011011;
assign LUT_2[61630] = 32'b11111111111111101001111001111110;
assign LUT_2[61631] = 32'b11111111111111100110110010010111;
assign LUT_2[61632] = 32'b11111111111111101000111010101101;
assign LUT_2[61633] = 32'b11111111111111100101110011000110;
assign LUT_2[61634] = 32'b11111111111111101111110011101001;
assign LUT_2[61635] = 32'b11111111111111101100101100000010;
assign LUT_2[61636] = 32'b11111111111111100101011000010101;
assign LUT_2[61637] = 32'b11111111111111100010010000101110;
assign LUT_2[61638] = 32'b11111111111111101100010001010001;
assign LUT_2[61639] = 32'b11111111111111101001001001101010;
assign LUT_2[61640] = 32'b11111111111111100011101100001010;
assign LUT_2[61641] = 32'b11111111111111100000100100100011;
assign LUT_2[61642] = 32'b11111111111111101010100101000110;
assign LUT_2[61643] = 32'b11111111111111100111011101011111;
assign LUT_2[61644] = 32'b11111111111111100000001001110010;
assign LUT_2[61645] = 32'b11111111111111011101000010001011;
assign LUT_2[61646] = 32'b11111111111111100111000010101110;
assign LUT_2[61647] = 32'b11111111111111100011111011000111;
assign LUT_2[61648] = 32'b11111111111111100011011110110111;
assign LUT_2[61649] = 32'b11111111111111100000010111010000;
assign LUT_2[61650] = 32'b11111111111111101010010111110011;
assign LUT_2[61651] = 32'b11111111111111100111010000001100;
assign LUT_2[61652] = 32'b11111111111111011111111100011111;
assign LUT_2[61653] = 32'b11111111111111011100110100111000;
assign LUT_2[61654] = 32'b11111111111111100110110101011011;
assign LUT_2[61655] = 32'b11111111111111100011101101110100;
assign LUT_2[61656] = 32'b11111111111111011110010000010100;
assign LUT_2[61657] = 32'b11111111111111011011001000101101;
assign LUT_2[61658] = 32'b11111111111111100101001001010000;
assign LUT_2[61659] = 32'b11111111111111100010000001101001;
assign LUT_2[61660] = 32'b11111111111111011010101101111100;
assign LUT_2[61661] = 32'b11111111111111010111100110010101;
assign LUT_2[61662] = 32'b11111111111111100001100110111000;
assign LUT_2[61663] = 32'b11111111111111011110011111010001;
assign LUT_2[61664] = 32'b11111111111111101001010110010110;
assign LUT_2[61665] = 32'b11111111111111100110001110101111;
assign LUT_2[61666] = 32'b11111111111111110000001111010010;
assign LUT_2[61667] = 32'b11111111111111101101000111101011;
assign LUT_2[61668] = 32'b11111111111111100101110011111110;
assign LUT_2[61669] = 32'b11111111111111100010101100010111;
assign LUT_2[61670] = 32'b11111111111111101100101100111010;
assign LUT_2[61671] = 32'b11111111111111101001100101010011;
assign LUT_2[61672] = 32'b11111111111111100100000111110011;
assign LUT_2[61673] = 32'b11111111111111100001000000001100;
assign LUT_2[61674] = 32'b11111111111111101011000000101111;
assign LUT_2[61675] = 32'b11111111111111100111111001001000;
assign LUT_2[61676] = 32'b11111111111111100000100101011011;
assign LUT_2[61677] = 32'b11111111111111011101011101110100;
assign LUT_2[61678] = 32'b11111111111111100111011110010111;
assign LUT_2[61679] = 32'b11111111111111100100010110110000;
assign LUT_2[61680] = 32'b11111111111111100011111010100000;
assign LUT_2[61681] = 32'b11111111111111100000110010111001;
assign LUT_2[61682] = 32'b11111111111111101010110011011100;
assign LUT_2[61683] = 32'b11111111111111100111101011110101;
assign LUT_2[61684] = 32'b11111111111111100000011000001000;
assign LUT_2[61685] = 32'b11111111111111011101010000100001;
assign LUT_2[61686] = 32'b11111111111111100111010001000100;
assign LUT_2[61687] = 32'b11111111111111100100001001011101;
assign LUT_2[61688] = 32'b11111111111111011110101011111101;
assign LUT_2[61689] = 32'b11111111111111011011100100010110;
assign LUT_2[61690] = 32'b11111111111111100101100100111001;
assign LUT_2[61691] = 32'b11111111111111100010011101010010;
assign LUT_2[61692] = 32'b11111111111111011011001001100101;
assign LUT_2[61693] = 32'b11111111111111011000000001111110;
assign LUT_2[61694] = 32'b11111111111111100010000010100001;
assign LUT_2[61695] = 32'b11111111111111011110111010111010;
assign LUT_2[61696] = 32'b11111111111111110000011100100001;
assign LUT_2[61697] = 32'b11111111111111101101010100111010;
assign LUT_2[61698] = 32'b11111111111111110111010101011101;
assign LUT_2[61699] = 32'b11111111111111110100001101110110;
assign LUT_2[61700] = 32'b11111111111111101100111010001001;
assign LUT_2[61701] = 32'b11111111111111101001110010100010;
assign LUT_2[61702] = 32'b11111111111111110011110011000101;
assign LUT_2[61703] = 32'b11111111111111110000101011011110;
assign LUT_2[61704] = 32'b11111111111111101011001101111110;
assign LUT_2[61705] = 32'b11111111111111101000000110010111;
assign LUT_2[61706] = 32'b11111111111111110010000110111010;
assign LUT_2[61707] = 32'b11111111111111101110111111010011;
assign LUT_2[61708] = 32'b11111111111111100111101011100110;
assign LUT_2[61709] = 32'b11111111111111100100100011111111;
assign LUT_2[61710] = 32'b11111111111111101110100100100010;
assign LUT_2[61711] = 32'b11111111111111101011011100111011;
assign LUT_2[61712] = 32'b11111111111111101011000000101011;
assign LUT_2[61713] = 32'b11111111111111100111111001000100;
assign LUT_2[61714] = 32'b11111111111111110001111001100111;
assign LUT_2[61715] = 32'b11111111111111101110110010000000;
assign LUT_2[61716] = 32'b11111111111111100111011110010011;
assign LUT_2[61717] = 32'b11111111111111100100010110101100;
assign LUT_2[61718] = 32'b11111111111111101110010111001111;
assign LUT_2[61719] = 32'b11111111111111101011001111101000;
assign LUT_2[61720] = 32'b11111111111111100101110010001000;
assign LUT_2[61721] = 32'b11111111111111100010101010100001;
assign LUT_2[61722] = 32'b11111111111111101100101011000100;
assign LUT_2[61723] = 32'b11111111111111101001100011011101;
assign LUT_2[61724] = 32'b11111111111111100010001111110000;
assign LUT_2[61725] = 32'b11111111111111011111001000001001;
assign LUT_2[61726] = 32'b11111111111111101001001000101100;
assign LUT_2[61727] = 32'b11111111111111100110000001000101;
assign LUT_2[61728] = 32'b11111111111111110000111000001010;
assign LUT_2[61729] = 32'b11111111111111101101110000100011;
assign LUT_2[61730] = 32'b11111111111111110111110001000110;
assign LUT_2[61731] = 32'b11111111111111110100101001011111;
assign LUT_2[61732] = 32'b11111111111111101101010101110010;
assign LUT_2[61733] = 32'b11111111111111101010001110001011;
assign LUT_2[61734] = 32'b11111111111111110100001110101110;
assign LUT_2[61735] = 32'b11111111111111110001000111000111;
assign LUT_2[61736] = 32'b11111111111111101011101001100111;
assign LUT_2[61737] = 32'b11111111111111101000100010000000;
assign LUT_2[61738] = 32'b11111111111111110010100010100011;
assign LUT_2[61739] = 32'b11111111111111101111011010111100;
assign LUT_2[61740] = 32'b11111111111111101000000111001111;
assign LUT_2[61741] = 32'b11111111111111100100111111101000;
assign LUT_2[61742] = 32'b11111111111111101111000000001011;
assign LUT_2[61743] = 32'b11111111111111101011111000100100;
assign LUT_2[61744] = 32'b11111111111111101011011100010100;
assign LUT_2[61745] = 32'b11111111111111101000010100101101;
assign LUT_2[61746] = 32'b11111111111111110010010101010000;
assign LUT_2[61747] = 32'b11111111111111101111001101101001;
assign LUT_2[61748] = 32'b11111111111111100111111001111100;
assign LUT_2[61749] = 32'b11111111111111100100110010010101;
assign LUT_2[61750] = 32'b11111111111111101110110010111000;
assign LUT_2[61751] = 32'b11111111111111101011101011010001;
assign LUT_2[61752] = 32'b11111111111111100110001101110001;
assign LUT_2[61753] = 32'b11111111111111100011000110001010;
assign LUT_2[61754] = 32'b11111111111111101101000110101101;
assign LUT_2[61755] = 32'b11111111111111101001111111000110;
assign LUT_2[61756] = 32'b11111111111111100010101011011001;
assign LUT_2[61757] = 32'b11111111111111011111100011110010;
assign LUT_2[61758] = 32'b11111111111111101001100100010101;
assign LUT_2[61759] = 32'b11111111111111100110011100101110;
assign LUT_2[61760] = 32'b11111111111111101000100101000100;
assign LUT_2[61761] = 32'b11111111111111100101011101011101;
assign LUT_2[61762] = 32'b11111111111111101111011110000000;
assign LUT_2[61763] = 32'b11111111111111101100010110011001;
assign LUT_2[61764] = 32'b11111111111111100101000010101100;
assign LUT_2[61765] = 32'b11111111111111100001111011000101;
assign LUT_2[61766] = 32'b11111111111111101011111011101000;
assign LUT_2[61767] = 32'b11111111111111101000110100000001;
assign LUT_2[61768] = 32'b11111111111111100011010110100001;
assign LUT_2[61769] = 32'b11111111111111100000001110111010;
assign LUT_2[61770] = 32'b11111111111111101010001111011101;
assign LUT_2[61771] = 32'b11111111111111100111000111110110;
assign LUT_2[61772] = 32'b11111111111111011111110100001001;
assign LUT_2[61773] = 32'b11111111111111011100101100100010;
assign LUT_2[61774] = 32'b11111111111111100110101101000101;
assign LUT_2[61775] = 32'b11111111111111100011100101011110;
assign LUT_2[61776] = 32'b11111111111111100011001001001110;
assign LUT_2[61777] = 32'b11111111111111100000000001100111;
assign LUT_2[61778] = 32'b11111111111111101010000010001010;
assign LUT_2[61779] = 32'b11111111111111100110111010100011;
assign LUT_2[61780] = 32'b11111111111111011111100110110110;
assign LUT_2[61781] = 32'b11111111111111011100011111001111;
assign LUT_2[61782] = 32'b11111111111111100110011111110010;
assign LUT_2[61783] = 32'b11111111111111100011011000001011;
assign LUT_2[61784] = 32'b11111111111111011101111010101011;
assign LUT_2[61785] = 32'b11111111111111011010110011000100;
assign LUT_2[61786] = 32'b11111111111111100100110011100111;
assign LUT_2[61787] = 32'b11111111111111100001101100000000;
assign LUT_2[61788] = 32'b11111111111111011010011000010011;
assign LUT_2[61789] = 32'b11111111111111010111010000101100;
assign LUT_2[61790] = 32'b11111111111111100001010001001111;
assign LUT_2[61791] = 32'b11111111111111011110001001101000;
assign LUT_2[61792] = 32'b11111111111111101001000000101101;
assign LUT_2[61793] = 32'b11111111111111100101111001000110;
assign LUT_2[61794] = 32'b11111111111111101111111001101001;
assign LUT_2[61795] = 32'b11111111111111101100110010000010;
assign LUT_2[61796] = 32'b11111111111111100101011110010101;
assign LUT_2[61797] = 32'b11111111111111100010010110101110;
assign LUT_2[61798] = 32'b11111111111111101100010111010001;
assign LUT_2[61799] = 32'b11111111111111101001001111101010;
assign LUT_2[61800] = 32'b11111111111111100011110010001010;
assign LUT_2[61801] = 32'b11111111111111100000101010100011;
assign LUT_2[61802] = 32'b11111111111111101010101011000110;
assign LUT_2[61803] = 32'b11111111111111100111100011011111;
assign LUT_2[61804] = 32'b11111111111111100000001111110010;
assign LUT_2[61805] = 32'b11111111111111011101001000001011;
assign LUT_2[61806] = 32'b11111111111111100111001000101110;
assign LUT_2[61807] = 32'b11111111111111100100000001000111;
assign LUT_2[61808] = 32'b11111111111111100011100100110111;
assign LUT_2[61809] = 32'b11111111111111100000011101010000;
assign LUT_2[61810] = 32'b11111111111111101010011101110011;
assign LUT_2[61811] = 32'b11111111111111100111010110001100;
assign LUT_2[61812] = 32'b11111111111111100000000010011111;
assign LUT_2[61813] = 32'b11111111111111011100111010111000;
assign LUT_2[61814] = 32'b11111111111111100110111011011011;
assign LUT_2[61815] = 32'b11111111111111100011110011110100;
assign LUT_2[61816] = 32'b11111111111111011110010110010100;
assign LUT_2[61817] = 32'b11111111111111011011001110101101;
assign LUT_2[61818] = 32'b11111111111111100101001111010000;
assign LUT_2[61819] = 32'b11111111111111100010000111101001;
assign LUT_2[61820] = 32'b11111111111111011010110011111100;
assign LUT_2[61821] = 32'b11111111111111010111101100010101;
assign LUT_2[61822] = 32'b11111111111111100001101100111000;
assign LUT_2[61823] = 32'b11111111111111011110100101010001;
assign LUT_2[61824] = 32'b11111111111111110100110000110000;
assign LUT_2[61825] = 32'b11111111111111110001101001001001;
assign LUT_2[61826] = 32'b11111111111111111011101001101100;
assign LUT_2[61827] = 32'b11111111111111111000100010000101;
assign LUT_2[61828] = 32'b11111111111111110001001110011000;
assign LUT_2[61829] = 32'b11111111111111101110000110110001;
assign LUT_2[61830] = 32'b11111111111111111000000111010100;
assign LUT_2[61831] = 32'b11111111111111110100111111101101;
assign LUT_2[61832] = 32'b11111111111111101111100010001101;
assign LUT_2[61833] = 32'b11111111111111101100011010100110;
assign LUT_2[61834] = 32'b11111111111111110110011011001001;
assign LUT_2[61835] = 32'b11111111111111110011010011100010;
assign LUT_2[61836] = 32'b11111111111111101011111111110101;
assign LUT_2[61837] = 32'b11111111111111101000111000001110;
assign LUT_2[61838] = 32'b11111111111111110010111000110001;
assign LUT_2[61839] = 32'b11111111111111101111110001001010;
assign LUT_2[61840] = 32'b11111111111111101111010100111010;
assign LUT_2[61841] = 32'b11111111111111101100001101010011;
assign LUT_2[61842] = 32'b11111111111111110110001101110110;
assign LUT_2[61843] = 32'b11111111111111110011000110001111;
assign LUT_2[61844] = 32'b11111111111111101011110010100010;
assign LUT_2[61845] = 32'b11111111111111101000101010111011;
assign LUT_2[61846] = 32'b11111111111111110010101011011110;
assign LUT_2[61847] = 32'b11111111111111101111100011110111;
assign LUT_2[61848] = 32'b11111111111111101010000110010111;
assign LUT_2[61849] = 32'b11111111111111100110111110110000;
assign LUT_2[61850] = 32'b11111111111111110000111111010011;
assign LUT_2[61851] = 32'b11111111111111101101110111101100;
assign LUT_2[61852] = 32'b11111111111111100110100011111111;
assign LUT_2[61853] = 32'b11111111111111100011011100011000;
assign LUT_2[61854] = 32'b11111111111111101101011100111011;
assign LUT_2[61855] = 32'b11111111111111101010010101010100;
assign LUT_2[61856] = 32'b11111111111111110101001100011001;
assign LUT_2[61857] = 32'b11111111111111110010000100110010;
assign LUT_2[61858] = 32'b11111111111111111100000101010101;
assign LUT_2[61859] = 32'b11111111111111111000111101101110;
assign LUT_2[61860] = 32'b11111111111111110001101010000001;
assign LUT_2[61861] = 32'b11111111111111101110100010011010;
assign LUT_2[61862] = 32'b11111111111111111000100010111101;
assign LUT_2[61863] = 32'b11111111111111110101011011010110;
assign LUT_2[61864] = 32'b11111111111111101111111101110110;
assign LUT_2[61865] = 32'b11111111111111101100110110001111;
assign LUT_2[61866] = 32'b11111111111111110110110110110010;
assign LUT_2[61867] = 32'b11111111111111110011101111001011;
assign LUT_2[61868] = 32'b11111111111111101100011011011110;
assign LUT_2[61869] = 32'b11111111111111101001010011110111;
assign LUT_2[61870] = 32'b11111111111111110011010100011010;
assign LUT_2[61871] = 32'b11111111111111110000001100110011;
assign LUT_2[61872] = 32'b11111111111111101111110000100011;
assign LUT_2[61873] = 32'b11111111111111101100101000111100;
assign LUT_2[61874] = 32'b11111111111111110110101001011111;
assign LUT_2[61875] = 32'b11111111111111110011100001111000;
assign LUT_2[61876] = 32'b11111111111111101100001110001011;
assign LUT_2[61877] = 32'b11111111111111101001000110100100;
assign LUT_2[61878] = 32'b11111111111111110011000111000111;
assign LUT_2[61879] = 32'b11111111111111101111111111100000;
assign LUT_2[61880] = 32'b11111111111111101010100010000000;
assign LUT_2[61881] = 32'b11111111111111100111011010011001;
assign LUT_2[61882] = 32'b11111111111111110001011010111100;
assign LUT_2[61883] = 32'b11111111111111101110010011010101;
assign LUT_2[61884] = 32'b11111111111111100110111111101000;
assign LUT_2[61885] = 32'b11111111111111100011111000000001;
assign LUT_2[61886] = 32'b11111111111111101101111000100100;
assign LUT_2[61887] = 32'b11111111111111101010110000111101;
assign LUT_2[61888] = 32'b11111111111111101100111001010011;
assign LUT_2[61889] = 32'b11111111111111101001110001101100;
assign LUT_2[61890] = 32'b11111111111111110011110010001111;
assign LUT_2[61891] = 32'b11111111111111110000101010101000;
assign LUT_2[61892] = 32'b11111111111111101001010110111011;
assign LUT_2[61893] = 32'b11111111111111100110001111010100;
assign LUT_2[61894] = 32'b11111111111111110000001111110111;
assign LUT_2[61895] = 32'b11111111111111101101001000010000;
assign LUT_2[61896] = 32'b11111111111111100111101010110000;
assign LUT_2[61897] = 32'b11111111111111100100100011001001;
assign LUT_2[61898] = 32'b11111111111111101110100011101100;
assign LUT_2[61899] = 32'b11111111111111101011011100000101;
assign LUT_2[61900] = 32'b11111111111111100100001000011000;
assign LUT_2[61901] = 32'b11111111111111100001000000110001;
assign LUT_2[61902] = 32'b11111111111111101011000001010100;
assign LUT_2[61903] = 32'b11111111111111100111111001101101;
assign LUT_2[61904] = 32'b11111111111111100111011101011101;
assign LUT_2[61905] = 32'b11111111111111100100010101110110;
assign LUT_2[61906] = 32'b11111111111111101110010110011001;
assign LUT_2[61907] = 32'b11111111111111101011001110110010;
assign LUT_2[61908] = 32'b11111111111111100011111011000101;
assign LUT_2[61909] = 32'b11111111111111100000110011011110;
assign LUT_2[61910] = 32'b11111111111111101010110100000001;
assign LUT_2[61911] = 32'b11111111111111100111101100011010;
assign LUT_2[61912] = 32'b11111111111111100010001110111010;
assign LUT_2[61913] = 32'b11111111111111011111000111010011;
assign LUT_2[61914] = 32'b11111111111111101001000111110110;
assign LUT_2[61915] = 32'b11111111111111100110000000001111;
assign LUT_2[61916] = 32'b11111111111111011110101100100010;
assign LUT_2[61917] = 32'b11111111111111011011100100111011;
assign LUT_2[61918] = 32'b11111111111111100101100101011110;
assign LUT_2[61919] = 32'b11111111111111100010011101110111;
assign LUT_2[61920] = 32'b11111111111111101101010100111100;
assign LUT_2[61921] = 32'b11111111111111101010001101010101;
assign LUT_2[61922] = 32'b11111111111111110100001101111000;
assign LUT_2[61923] = 32'b11111111111111110001000110010001;
assign LUT_2[61924] = 32'b11111111111111101001110010100100;
assign LUT_2[61925] = 32'b11111111111111100110101010111101;
assign LUT_2[61926] = 32'b11111111111111110000101011100000;
assign LUT_2[61927] = 32'b11111111111111101101100011111001;
assign LUT_2[61928] = 32'b11111111111111101000000110011001;
assign LUT_2[61929] = 32'b11111111111111100100111110110010;
assign LUT_2[61930] = 32'b11111111111111101110111111010101;
assign LUT_2[61931] = 32'b11111111111111101011110111101110;
assign LUT_2[61932] = 32'b11111111111111100100100100000001;
assign LUT_2[61933] = 32'b11111111111111100001011100011010;
assign LUT_2[61934] = 32'b11111111111111101011011100111101;
assign LUT_2[61935] = 32'b11111111111111101000010101010110;
assign LUT_2[61936] = 32'b11111111111111100111111001000110;
assign LUT_2[61937] = 32'b11111111111111100100110001011111;
assign LUT_2[61938] = 32'b11111111111111101110110010000010;
assign LUT_2[61939] = 32'b11111111111111101011101010011011;
assign LUT_2[61940] = 32'b11111111111111100100010110101110;
assign LUT_2[61941] = 32'b11111111111111100001001111000111;
assign LUT_2[61942] = 32'b11111111111111101011001111101010;
assign LUT_2[61943] = 32'b11111111111111101000001000000011;
assign LUT_2[61944] = 32'b11111111111111100010101010100011;
assign LUT_2[61945] = 32'b11111111111111011111100010111100;
assign LUT_2[61946] = 32'b11111111111111101001100011011111;
assign LUT_2[61947] = 32'b11111111111111100110011011111000;
assign LUT_2[61948] = 32'b11111111111111011111001000001011;
assign LUT_2[61949] = 32'b11111111111111011100000000100100;
assign LUT_2[61950] = 32'b11111111111111100110000001000111;
assign LUT_2[61951] = 32'b11111111111111100010111001100000;
assign LUT_2[61952] = 32'b11111111111111110001001111101101;
assign LUT_2[61953] = 32'b11111111111111101110001000000110;
assign LUT_2[61954] = 32'b11111111111111111000001000101001;
assign LUT_2[61955] = 32'b11111111111111110101000001000010;
assign LUT_2[61956] = 32'b11111111111111101101101101010101;
assign LUT_2[61957] = 32'b11111111111111101010100101101110;
assign LUT_2[61958] = 32'b11111111111111110100100110010001;
assign LUT_2[61959] = 32'b11111111111111110001011110101010;
assign LUT_2[61960] = 32'b11111111111111101100000001001010;
assign LUT_2[61961] = 32'b11111111111111101000111001100011;
assign LUT_2[61962] = 32'b11111111111111110010111010000110;
assign LUT_2[61963] = 32'b11111111111111101111110010011111;
assign LUT_2[61964] = 32'b11111111111111101000011110110010;
assign LUT_2[61965] = 32'b11111111111111100101010111001011;
assign LUT_2[61966] = 32'b11111111111111101111010111101110;
assign LUT_2[61967] = 32'b11111111111111101100010000000111;
assign LUT_2[61968] = 32'b11111111111111101011110011110111;
assign LUT_2[61969] = 32'b11111111111111101000101100010000;
assign LUT_2[61970] = 32'b11111111111111110010101100110011;
assign LUT_2[61971] = 32'b11111111111111101111100101001100;
assign LUT_2[61972] = 32'b11111111111111101000010001011111;
assign LUT_2[61973] = 32'b11111111111111100101001001111000;
assign LUT_2[61974] = 32'b11111111111111101111001010011011;
assign LUT_2[61975] = 32'b11111111111111101100000010110100;
assign LUT_2[61976] = 32'b11111111111111100110100101010100;
assign LUT_2[61977] = 32'b11111111111111100011011101101101;
assign LUT_2[61978] = 32'b11111111111111101101011110010000;
assign LUT_2[61979] = 32'b11111111111111101010010110101001;
assign LUT_2[61980] = 32'b11111111111111100011000010111100;
assign LUT_2[61981] = 32'b11111111111111011111111011010101;
assign LUT_2[61982] = 32'b11111111111111101001111011111000;
assign LUT_2[61983] = 32'b11111111111111100110110100010001;
assign LUT_2[61984] = 32'b11111111111111110001101011010110;
assign LUT_2[61985] = 32'b11111111111111101110100011101111;
assign LUT_2[61986] = 32'b11111111111111111000100100010010;
assign LUT_2[61987] = 32'b11111111111111110101011100101011;
assign LUT_2[61988] = 32'b11111111111111101110001000111110;
assign LUT_2[61989] = 32'b11111111111111101011000001010111;
assign LUT_2[61990] = 32'b11111111111111110101000001111010;
assign LUT_2[61991] = 32'b11111111111111110001111010010011;
assign LUT_2[61992] = 32'b11111111111111101100011100110011;
assign LUT_2[61993] = 32'b11111111111111101001010101001100;
assign LUT_2[61994] = 32'b11111111111111110011010101101111;
assign LUT_2[61995] = 32'b11111111111111110000001110001000;
assign LUT_2[61996] = 32'b11111111111111101000111010011011;
assign LUT_2[61997] = 32'b11111111111111100101110010110100;
assign LUT_2[61998] = 32'b11111111111111101111110011010111;
assign LUT_2[61999] = 32'b11111111111111101100101011110000;
assign LUT_2[62000] = 32'b11111111111111101100001111100000;
assign LUT_2[62001] = 32'b11111111111111101001000111111001;
assign LUT_2[62002] = 32'b11111111111111110011001000011100;
assign LUT_2[62003] = 32'b11111111111111110000000000110101;
assign LUT_2[62004] = 32'b11111111111111101000101101001000;
assign LUT_2[62005] = 32'b11111111111111100101100101100001;
assign LUT_2[62006] = 32'b11111111111111101111100110000100;
assign LUT_2[62007] = 32'b11111111111111101100011110011101;
assign LUT_2[62008] = 32'b11111111111111100111000000111101;
assign LUT_2[62009] = 32'b11111111111111100011111001010110;
assign LUT_2[62010] = 32'b11111111111111101101111001111001;
assign LUT_2[62011] = 32'b11111111111111101010110010010010;
assign LUT_2[62012] = 32'b11111111111111100011011110100101;
assign LUT_2[62013] = 32'b11111111111111100000010110111110;
assign LUT_2[62014] = 32'b11111111111111101010010111100001;
assign LUT_2[62015] = 32'b11111111111111100111001111111010;
assign LUT_2[62016] = 32'b11111111111111101001011000010000;
assign LUT_2[62017] = 32'b11111111111111100110010000101001;
assign LUT_2[62018] = 32'b11111111111111110000010001001100;
assign LUT_2[62019] = 32'b11111111111111101101001001100101;
assign LUT_2[62020] = 32'b11111111111111100101110101111000;
assign LUT_2[62021] = 32'b11111111111111100010101110010001;
assign LUT_2[62022] = 32'b11111111111111101100101110110100;
assign LUT_2[62023] = 32'b11111111111111101001100111001101;
assign LUT_2[62024] = 32'b11111111111111100100001001101101;
assign LUT_2[62025] = 32'b11111111111111100001000010000110;
assign LUT_2[62026] = 32'b11111111111111101011000010101001;
assign LUT_2[62027] = 32'b11111111111111100111111011000010;
assign LUT_2[62028] = 32'b11111111111111100000100111010101;
assign LUT_2[62029] = 32'b11111111111111011101011111101110;
assign LUT_2[62030] = 32'b11111111111111100111100000010001;
assign LUT_2[62031] = 32'b11111111111111100100011000101010;
assign LUT_2[62032] = 32'b11111111111111100011111100011010;
assign LUT_2[62033] = 32'b11111111111111100000110100110011;
assign LUT_2[62034] = 32'b11111111111111101010110101010110;
assign LUT_2[62035] = 32'b11111111111111100111101101101111;
assign LUT_2[62036] = 32'b11111111111111100000011010000010;
assign LUT_2[62037] = 32'b11111111111111011101010010011011;
assign LUT_2[62038] = 32'b11111111111111100111010010111110;
assign LUT_2[62039] = 32'b11111111111111100100001011010111;
assign LUT_2[62040] = 32'b11111111111111011110101101110111;
assign LUT_2[62041] = 32'b11111111111111011011100110010000;
assign LUT_2[62042] = 32'b11111111111111100101100110110011;
assign LUT_2[62043] = 32'b11111111111111100010011111001100;
assign LUT_2[62044] = 32'b11111111111111011011001011011111;
assign LUT_2[62045] = 32'b11111111111111011000000011111000;
assign LUT_2[62046] = 32'b11111111111111100010000100011011;
assign LUT_2[62047] = 32'b11111111111111011110111100110100;
assign LUT_2[62048] = 32'b11111111111111101001110011111001;
assign LUT_2[62049] = 32'b11111111111111100110101100010010;
assign LUT_2[62050] = 32'b11111111111111110000101100110101;
assign LUT_2[62051] = 32'b11111111111111101101100101001110;
assign LUT_2[62052] = 32'b11111111111111100110010001100001;
assign LUT_2[62053] = 32'b11111111111111100011001001111010;
assign LUT_2[62054] = 32'b11111111111111101101001010011101;
assign LUT_2[62055] = 32'b11111111111111101010000010110110;
assign LUT_2[62056] = 32'b11111111111111100100100101010110;
assign LUT_2[62057] = 32'b11111111111111100001011101101111;
assign LUT_2[62058] = 32'b11111111111111101011011110010010;
assign LUT_2[62059] = 32'b11111111111111101000010110101011;
assign LUT_2[62060] = 32'b11111111111111100001000010111110;
assign LUT_2[62061] = 32'b11111111111111011101111011010111;
assign LUT_2[62062] = 32'b11111111111111100111111011111010;
assign LUT_2[62063] = 32'b11111111111111100100110100010011;
assign LUT_2[62064] = 32'b11111111111111100100011000000011;
assign LUT_2[62065] = 32'b11111111111111100001010000011100;
assign LUT_2[62066] = 32'b11111111111111101011010000111111;
assign LUT_2[62067] = 32'b11111111111111101000001001011000;
assign LUT_2[62068] = 32'b11111111111111100000110101101011;
assign LUT_2[62069] = 32'b11111111111111011101101110000100;
assign LUT_2[62070] = 32'b11111111111111100111101110100111;
assign LUT_2[62071] = 32'b11111111111111100100100111000000;
assign LUT_2[62072] = 32'b11111111111111011111001001100000;
assign LUT_2[62073] = 32'b11111111111111011100000001111001;
assign LUT_2[62074] = 32'b11111111111111100110000010011100;
assign LUT_2[62075] = 32'b11111111111111100010111010110101;
assign LUT_2[62076] = 32'b11111111111111011011100111001000;
assign LUT_2[62077] = 32'b11111111111111011000011111100001;
assign LUT_2[62078] = 32'b11111111111111100010100000000100;
assign LUT_2[62079] = 32'b11111111111111011111011000011101;
assign LUT_2[62080] = 32'b11111111111111110101100011111100;
assign LUT_2[62081] = 32'b11111111111111110010011100010101;
assign LUT_2[62082] = 32'b11111111111111111100011100111000;
assign LUT_2[62083] = 32'b11111111111111111001010101010001;
assign LUT_2[62084] = 32'b11111111111111110010000001100100;
assign LUT_2[62085] = 32'b11111111111111101110111001111101;
assign LUT_2[62086] = 32'b11111111111111111000111010100000;
assign LUT_2[62087] = 32'b11111111111111110101110010111001;
assign LUT_2[62088] = 32'b11111111111111110000010101011001;
assign LUT_2[62089] = 32'b11111111111111101101001101110010;
assign LUT_2[62090] = 32'b11111111111111110111001110010101;
assign LUT_2[62091] = 32'b11111111111111110100000110101110;
assign LUT_2[62092] = 32'b11111111111111101100110011000001;
assign LUT_2[62093] = 32'b11111111111111101001101011011010;
assign LUT_2[62094] = 32'b11111111111111110011101011111101;
assign LUT_2[62095] = 32'b11111111111111110000100100010110;
assign LUT_2[62096] = 32'b11111111111111110000001000000110;
assign LUT_2[62097] = 32'b11111111111111101101000000011111;
assign LUT_2[62098] = 32'b11111111111111110111000001000010;
assign LUT_2[62099] = 32'b11111111111111110011111001011011;
assign LUT_2[62100] = 32'b11111111111111101100100101101110;
assign LUT_2[62101] = 32'b11111111111111101001011110000111;
assign LUT_2[62102] = 32'b11111111111111110011011110101010;
assign LUT_2[62103] = 32'b11111111111111110000010111000011;
assign LUT_2[62104] = 32'b11111111111111101010111001100011;
assign LUT_2[62105] = 32'b11111111111111100111110001111100;
assign LUT_2[62106] = 32'b11111111111111110001110010011111;
assign LUT_2[62107] = 32'b11111111111111101110101010111000;
assign LUT_2[62108] = 32'b11111111111111100111010111001011;
assign LUT_2[62109] = 32'b11111111111111100100001111100100;
assign LUT_2[62110] = 32'b11111111111111101110010000000111;
assign LUT_2[62111] = 32'b11111111111111101011001000100000;
assign LUT_2[62112] = 32'b11111111111111110101111111100101;
assign LUT_2[62113] = 32'b11111111111111110010110111111110;
assign LUT_2[62114] = 32'b11111111111111111100111000100001;
assign LUT_2[62115] = 32'b11111111111111111001110000111010;
assign LUT_2[62116] = 32'b11111111111111110010011101001101;
assign LUT_2[62117] = 32'b11111111111111101111010101100110;
assign LUT_2[62118] = 32'b11111111111111111001010110001001;
assign LUT_2[62119] = 32'b11111111111111110110001110100010;
assign LUT_2[62120] = 32'b11111111111111110000110001000010;
assign LUT_2[62121] = 32'b11111111111111101101101001011011;
assign LUT_2[62122] = 32'b11111111111111110111101001111110;
assign LUT_2[62123] = 32'b11111111111111110100100010010111;
assign LUT_2[62124] = 32'b11111111111111101101001110101010;
assign LUT_2[62125] = 32'b11111111111111101010000111000011;
assign LUT_2[62126] = 32'b11111111111111110100000111100110;
assign LUT_2[62127] = 32'b11111111111111110000111111111111;
assign LUT_2[62128] = 32'b11111111111111110000100011101111;
assign LUT_2[62129] = 32'b11111111111111101101011100001000;
assign LUT_2[62130] = 32'b11111111111111110111011100101011;
assign LUT_2[62131] = 32'b11111111111111110100010101000100;
assign LUT_2[62132] = 32'b11111111111111101101000001010111;
assign LUT_2[62133] = 32'b11111111111111101001111001110000;
assign LUT_2[62134] = 32'b11111111111111110011111010010011;
assign LUT_2[62135] = 32'b11111111111111110000110010101100;
assign LUT_2[62136] = 32'b11111111111111101011010101001100;
assign LUT_2[62137] = 32'b11111111111111101000001101100101;
assign LUT_2[62138] = 32'b11111111111111110010001110001000;
assign LUT_2[62139] = 32'b11111111111111101111000110100001;
assign LUT_2[62140] = 32'b11111111111111100111110010110100;
assign LUT_2[62141] = 32'b11111111111111100100101011001101;
assign LUT_2[62142] = 32'b11111111111111101110101011110000;
assign LUT_2[62143] = 32'b11111111111111101011100100001001;
assign LUT_2[62144] = 32'b11111111111111101101101100011111;
assign LUT_2[62145] = 32'b11111111111111101010100100111000;
assign LUT_2[62146] = 32'b11111111111111110100100101011011;
assign LUT_2[62147] = 32'b11111111111111110001011101110100;
assign LUT_2[62148] = 32'b11111111111111101010001010000111;
assign LUT_2[62149] = 32'b11111111111111100111000010100000;
assign LUT_2[62150] = 32'b11111111111111110001000011000011;
assign LUT_2[62151] = 32'b11111111111111101101111011011100;
assign LUT_2[62152] = 32'b11111111111111101000011101111100;
assign LUT_2[62153] = 32'b11111111111111100101010110010101;
assign LUT_2[62154] = 32'b11111111111111101111010110111000;
assign LUT_2[62155] = 32'b11111111111111101100001111010001;
assign LUT_2[62156] = 32'b11111111111111100100111011100100;
assign LUT_2[62157] = 32'b11111111111111100001110011111101;
assign LUT_2[62158] = 32'b11111111111111101011110100100000;
assign LUT_2[62159] = 32'b11111111111111101000101100111001;
assign LUT_2[62160] = 32'b11111111111111101000010000101001;
assign LUT_2[62161] = 32'b11111111111111100101001001000010;
assign LUT_2[62162] = 32'b11111111111111101111001001100101;
assign LUT_2[62163] = 32'b11111111111111101100000001111110;
assign LUT_2[62164] = 32'b11111111111111100100101110010001;
assign LUT_2[62165] = 32'b11111111111111100001100110101010;
assign LUT_2[62166] = 32'b11111111111111101011100111001101;
assign LUT_2[62167] = 32'b11111111111111101000011111100110;
assign LUT_2[62168] = 32'b11111111111111100011000010000110;
assign LUT_2[62169] = 32'b11111111111111011111111010011111;
assign LUT_2[62170] = 32'b11111111111111101001111011000010;
assign LUT_2[62171] = 32'b11111111111111100110110011011011;
assign LUT_2[62172] = 32'b11111111111111011111011111101110;
assign LUT_2[62173] = 32'b11111111111111011100011000000111;
assign LUT_2[62174] = 32'b11111111111111100110011000101010;
assign LUT_2[62175] = 32'b11111111111111100011010001000011;
assign LUT_2[62176] = 32'b11111111111111101110001000001000;
assign LUT_2[62177] = 32'b11111111111111101011000000100001;
assign LUT_2[62178] = 32'b11111111111111110101000001000100;
assign LUT_2[62179] = 32'b11111111111111110001111001011101;
assign LUT_2[62180] = 32'b11111111111111101010100101110000;
assign LUT_2[62181] = 32'b11111111111111100111011110001001;
assign LUT_2[62182] = 32'b11111111111111110001011110101100;
assign LUT_2[62183] = 32'b11111111111111101110010111000101;
assign LUT_2[62184] = 32'b11111111111111101000111001100101;
assign LUT_2[62185] = 32'b11111111111111100101110001111110;
assign LUT_2[62186] = 32'b11111111111111101111110010100001;
assign LUT_2[62187] = 32'b11111111111111101100101010111010;
assign LUT_2[62188] = 32'b11111111111111100101010111001101;
assign LUT_2[62189] = 32'b11111111111111100010001111100110;
assign LUT_2[62190] = 32'b11111111111111101100010000001001;
assign LUT_2[62191] = 32'b11111111111111101001001000100010;
assign LUT_2[62192] = 32'b11111111111111101000101100010010;
assign LUT_2[62193] = 32'b11111111111111100101100100101011;
assign LUT_2[62194] = 32'b11111111111111101111100101001110;
assign LUT_2[62195] = 32'b11111111111111101100011101100111;
assign LUT_2[62196] = 32'b11111111111111100101001001111010;
assign LUT_2[62197] = 32'b11111111111111100010000010010011;
assign LUT_2[62198] = 32'b11111111111111101100000010110110;
assign LUT_2[62199] = 32'b11111111111111101000111011001111;
assign LUT_2[62200] = 32'b11111111111111100011011101101111;
assign LUT_2[62201] = 32'b11111111111111100000010110001000;
assign LUT_2[62202] = 32'b11111111111111101010010110101011;
assign LUT_2[62203] = 32'b11111111111111100111001111000100;
assign LUT_2[62204] = 32'b11111111111111011111111011010111;
assign LUT_2[62205] = 32'b11111111111111011100110011110000;
assign LUT_2[62206] = 32'b11111111111111100110110100010011;
assign LUT_2[62207] = 32'b11111111111111100011101100101100;
assign LUT_2[62208] = 32'b11111111111111110101001110010011;
assign LUT_2[62209] = 32'b11111111111111110010000110101100;
assign LUT_2[62210] = 32'b11111111111111111100000111001111;
assign LUT_2[62211] = 32'b11111111111111111000111111101000;
assign LUT_2[62212] = 32'b11111111111111110001101011111011;
assign LUT_2[62213] = 32'b11111111111111101110100100010100;
assign LUT_2[62214] = 32'b11111111111111111000100100110111;
assign LUT_2[62215] = 32'b11111111111111110101011101010000;
assign LUT_2[62216] = 32'b11111111111111101111111111110000;
assign LUT_2[62217] = 32'b11111111111111101100111000001001;
assign LUT_2[62218] = 32'b11111111111111110110111000101100;
assign LUT_2[62219] = 32'b11111111111111110011110001000101;
assign LUT_2[62220] = 32'b11111111111111101100011101011000;
assign LUT_2[62221] = 32'b11111111111111101001010101110001;
assign LUT_2[62222] = 32'b11111111111111110011010110010100;
assign LUT_2[62223] = 32'b11111111111111110000001110101101;
assign LUT_2[62224] = 32'b11111111111111101111110010011101;
assign LUT_2[62225] = 32'b11111111111111101100101010110110;
assign LUT_2[62226] = 32'b11111111111111110110101011011001;
assign LUT_2[62227] = 32'b11111111111111110011100011110010;
assign LUT_2[62228] = 32'b11111111111111101100010000000101;
assign LUT_2[62229] = 32'b11111111111111101001001000011110;
assign LUT_2[62230] = 32'b11111111111111110011001001000001;
assign LUT_2[62231] = 32'b11111111111111110000000001011010;
assign LUT_2[62232] = 32'b11111111111111101010100011111010;
assign LUT_2[62233] = 32'b11111111111111100111011100010011;
assign LUT_2[62234] = 32'b11111111111111110001011100110110;
assign LUT_2[62235] = 32'b11111111111111101110010101001111;
assign LUT_2[62236] = 32'b11111111111111100111000001100010;
assign LUT_2[62237] = 32'b11111111111111100011111001111011;
assign LUT_2[62238] = 32'b11111111111111101101111010011110;
assign LUT_2[62239] = 32'b11111111111111101010110010110111;
assign LUT_2[62240] = 32'b11111111111111110101101001111100;
assign LUT_2[62241] = 32'b11111111111111110010100010010101;
assign LUT_2[62242] = 32'b11111111111111111100100010111000;
assign LUT_2[62243] = 32'b11111111111111111001011011010001;
assign LUT_2[62244] = 32'b11111111111111110010000111100100;
assign LUT_2[62245] = 32'b11111111111111101110111111111101;
assign LUT_2[62246] = 32'b11111111111111111001000000100000;
assign LUT_2[62247] = 32'b11111111111111110101111000111001;
assign LUT_2[62248] = 32'b11111111111111110000011011011001;
assign LUT_2[62249] = 32'b11111111111111101101010011110010;
assign LUT_2[62250] = 32'b11111111111111110111010100010101;
assign LUT_2[62251] = 32'b11111111111111110100001100101110;
assign LUT_2[62252] = 32'b11111111111111101100111001000001;
assign LUT_2[62253] = 32'b11111111111111101001110001011010;
assign LUT_2[62254] = 32'b11111111111111110011110001111101;
assign LUT_2[62255] = 32'b11111111111111110000101010010110;
assign LUT_2[62256] = 32'b11111111111111110000001110000110;
assign LUT_2[62257] = 32'b11111111111111101101000110011111;
assign LUT_2[62258] = 32'b11111111111111110111000111000010;
assign LUT_2[62259] = 32'b11111111111111110011111111011011;
assign LUT_2[62260] = 32'b11111111111111101100101011101110;
assign LUT_2[62261] = 32'b11111111111111101001100100000111;
assign LUT_2[62262] = 32'b11111111111111110011100100101010;
assign LUT_2[62263] = 32'b11111111111111110000011101000011;
assign LUT_2[62264] = 32'b11111111111111101010111111100011;
assign LUT_2[62265] = 32'b11111111111111100111110111111100;
assign LUT_2[62266] = 32'b11111111111111110001111000011111;
assign LUT_2[62267] = 32'b11111111111111101110110000111000;
assign LUT_2[62268] = 32'b11111111111111100111011101001011;
assign LUT_2[62269] = 32'b11111111111111100100010101100100;
assign LUT_2[62270] = 32'b11111111111111101110010110000111;
assign LUT_2[62271] = 32'b11111111111111101011001110100000;
assign LUT_2[62272] = 32'b11111111111111101101010110110110;
assign LUT_2[62273] = 32'b11111111111111101010001111001111;
assign LUT_2[62274] = 32'b11111111111111110100001111110010;
assign LUT_2[62275] = 32'b11111111111111110001001000001011;
assign LUT_2[62276] = 32'b11111111111111101001110100011110;
assign LUT_2[62277] = 32'b11111111111111100110101100110111;
assign LUT_2[62278] = 32'b11111111111111110000101101011010;
assign LUT_2[62279] = 32'b11111111111111101101100101110011;
assign LUT_2[62280] = 32'b11111111111111101000001000010011;
assign LUT_2[62281] = 32'b11111111111111100101000000101100;
assign LUT_2[62282] = 32'b11111111111111101111000001001111;
assign LUT_2[62283] = 32'b11111111111111101011111001101000;
assign LUT_2[62284] = 32'b11111111111111100100100101111011;
assign LUT_2[62285] = 32'b11111111111111100001011110010100;
assign LUT_2[62286] = 32'b11111111111111101011011110110111;
assign LUT_2[62287] = 32'b11111111111111101000010111010000;
assign LUT_2[62288] = 32'b11111111111111100111111011000000;
assign LUT_2[62289] = 32'b11111111111111100100110011011001;
assign LUT_2[62290] = 32'b11111111111111101110110011111100;
assign LUT_2[62291] = 32'b11111111111111101011101100010101;
assign LUT_2[62292] = 32'b11111111111111100100011000101000;
assign LUT_2[62293] = 32'b11111111111111100001010001000001;
assign LUT_2[62294] = 32'b11111111111111101011010001100100;
assign LUT_2[62295] = 32'b11111111111111101000001001111101;
assign LUT_2[62296] = 32'b11111111111111100010101100011101;
assign LUT_2[62297] = 32'b11111111111111011111100100110110;
assign LUT_2[62298] = 32'b11111111111111101001100101011001;
assign LUT_2[62299] = 32'b11111111111111100110011101110010;
assign LUT_2[62300] = 32'b11111111111111011111001010000101;
assign LUT_2[62301] = 32'b11111111111111011100000010011110;
assign LUT_2[62302] = 32'b11111111111111100110000011000001;
assign LUT_2[62303] = 32'b11111111111111100010111011011010;
assign LUT_2[62304] = 32'b11111111111111101101110010011111;
assign LUT_2[62305] = 32'b11111111111111101010101010111000;
assign LUT_2[62306] = 32'b11111111111111110100101011011011;
assign LUT_2[62307] = 32'b11111111111111110001100011110100;
assign LUT_2[62308] = 32'b11111111111111101010010000000111;
assign LUT_2[62309] = 32'b11111111111111100111001000100000;
assign LUT_2[62310] = 32'b11111111111111110001001001000011;
assign LUT_2[62311] = 32'b11111111111111101110000001011100;
assign LUT_2[62312] = 32'b11111111111111101000100011111100;
assign LUT_2[62313] = 32'b11111111111111100101011100010101;
assign LUT_2[62314] = 32'b11111111111111101111011100111000;
assign LUT_2[62315] = 32'b11111111111111101100010101010001;
assign LUT_2[62316] = 32'b11111111111111100101000001100100;
assign LUT_2[62317] = 32'b11111111111111100001111001111101;
assign LUT_2[62318] = 32'b11111111111111101011111010100000;
assign LUT_2[62319] = 32'b11111111111111101000110010111001;
assign LUT_2[62320] = 32'b11111111111111101000010110101001;
assign LUT_2[62321] = 32'b11111111111111100101001111000010;
assign LUT_2[62322] = 32'b11111111111111101111001111100101;
assign LUT_2[62323] = 32'b11111111111111101100000111111110;
assign LUT_2[62324] = 32'b11111111111111100100110100010001;
assign LUT_2[62325] = 32'b11111111111111100001101100101010;
assign LUT_2[62326] = 32'b11111111111111101011101101001101;
assign LUT_2[62327] = 32'b11111111111111101000100101100110;
assign LUT_2[62328] = 32'b11111111111111100011001000000110;
assign LUT_2[62329] = 32'b11111111111111100000000000011111;
assign LUT_2[62330] = 32'b11111111111111101010000001000010;
assign LUT_2[62331] = 32'b11111111111111100110111001011011;
assign LUT_2[62332] = 32'b11111111111111011111100101101110;
assign LUT_2[62333] = 32'b11111111111111011100011110000111;
assign LUT_2[62334] = 32'b11111111111111100110011110101010;
assign LUT_2[62335] = 32'b11111111111111100011010111000011;
assign LUT_2[62336] = 32'b11111111111111111001100010100010;
assign LUT_2[62337] = 32'b11111111111111110110011010111011;
assign LUT_2[62338] = 32'b00000000000000000000011011011110;
assign LUT_2[62339] = 32'b11111111111111111101010011110111;
assign LUT_2[62340] = 32'b11111111111111110110000000001010;
assign LUT_2[62341] = 32'b11111111111111110010111000100011;
assign LUT_2[62342] = 32'b11111111111111111100111001000110;
assign LUT_2[62343] = 32'b11111111111111111001110001011111;
assign LUT_2[62344] = 32'b11111111111111110100010011111111;
assign LUT_2[62345] = 32'b11111111111111110001001100011000;
assign LUT_2[62346] = 32'b11111111111111111011001100111011;
assign LUT_2[62347] = 32'b11111111111111111000000101010100;
assign LUT_2[62348] = 32'b11111111111111110000110001100111;
assign LUT_2[62349] = 32'b11111111111111101101101010000000;
assign LUT_2[62350] = 32'b11111111111111110111101010100011;
assign LUT_2[62351] = 32'b11111111111111110100100010111100;
assign LUT_2[62352] = 32'b11111111111111110100000110101100;
assign LUT_2[62353] = 32'b11111111111111110000111111000101;
assign LUT_2[62354] = 32'b11111111111111111010111111101000;
assign LUT_2[62355] = 32'b11111111111111110111111000000001;
assign LUT_2[62356] = 32'b11111111111111110000100100010100;
assign LUT_2[62357] = 32'b11111111111111101101011100101101;
assign LUT_2[62358] = 32'b11111111111111110111011101010000;
assign LUT_2[62359] = 32'b11111111111111110100010101101001;
assign LUT_2[62360] = 32'b11111111111111101110111000001001;
assign LUT_2[62361] = 32'b11111111111111101011110000100010;
assign LUT_2[62362] = 32'b11111111111111110101110001000101;
assign LUT_2[62363] = 32'b11111111111111110010101001011110;
assign LUT_2[62364] = 32'b11111111111111101011010101110001;
assign LUT_2[62365] = 32'b11111111111111101000001110001010;
assign LUT_2[62366] = 32'b11111111111111110010001110101101;
assign LUT_2[62367] = 32'b11111111111111101111000111000110;
assign LUT_2[62368] = 32'b11111111111111111001111110001011;
assign LUT_2[62369] = 32'b11111111111111110110110110100100;
assign LUT_2[62370] = 32'b00000000000000000000110111000111;
assign LUT_2[62371] = 32'b11111111111111111101101111100000;
assign LUT_2[62372] = 32'b11111111111111110110011011110011;
assign LUT_2[62373] = 32'b11111111111111110011010100001100;
assign LUT_2[62374] = 32'b11111111111111111101010100101111;
assign LUT_2[62375] = 32'b11111111111111111010001101001000;
assign LUT_2[62376] = 32'b11111111111111110100101111101000;
assign LUT_2[62377] = 32'b11111111111111110001101000000001;
assign LUT_2[62378] = 32'b11111111111111111011101000100100;
assign LUT_2[62379] = 32'b11111111111111111000100000111101;
assign LUT_2[62380] = 32'b11111111111111110001001101010000;
assign LUT_2[62381] = 32'b11111111111111101110000101101001;
assign LUT_2[62382] = 32'b11111111111111111000000110001100;
assign LUT_2[62383] = 32'b11111111111111110100111110100101;
assign LUT_2[62384] = 32'b11111111111111110100100010010101;
assign LUT_2[62385] = 32'b11111111111111110001011010101110;
assign LUT_2[62386] = 32'b11111111111111111011011011010001;
assign LUT_2[62387] = 32'b11111111111111111000010011101010;
assign LUT_2[62388] = 32'b11111111111111110000111111111101;
assign LUT_2[62389] = 32'b11111111111111101101111000010110;
assign LUT_2[62390] = 32'b11111111111111110111111000111001;
assign LUT_2[62391] = 32'b11111111111111110100110001010010;
assign LUT_2[62392] = 32'b11111111111111101111010011110010;
assign LUT_2[62393] = 32'b11111111111111101100001100001011;
assign LUT_2[62394] = 32'b11111111111111110110001100101110;
assign LUT_2[62395] = 32'b11111111111111110011000101000111;
assign LUT_2[62396] = 32'b11111111111111101011110001011010;
assign LUT_2[62397] = 32'b11111111111111101000101001110011;
assign LUT_2[62398] = 32'b11111111111111110010101010010110;
assign LUT_2[62399] = 32'b11111111111111101111100010101111;
assign LUT_2[62400] = 32'b11111111111111110001101011000101;
assign LUT_2[62401] = 32'b11111111111111101110100011011110;
assign LUT_2[62402] = 32'b11111111111111111000100100000001;
assign LUT_2[62403] = 32'b11111111111111110101011100011010;
assign LUT_2[62404] = 32'b11111111111111101110001000101101;
assign LUT_2[62405] = 32'b11111111111111101011000001000110;
assign LUT_2[62406] = 32'b11111111111111110101000001101001;
assign LUT_2[62407] = 32'b11111111111111110001111010000010;
assign LUT_2[62408] = 32'b11111111111111101100011100100010;
assign LUT_2[62409] = 32'b11111111111111101001010100111011;
assign LUT_2[62410] = 32'b11111111111111110011010101011110;
assign LUT_2[62411] = 32'b11111111111111110000001101110111;
assign LUT_2[62412] = 32'b11111111111111101000111010001010;
assign LUT_2[62413] = 32'b11111111111111100101110010100011;
assign LUT_2[62414] = 32'b11111111111111101111110011000110;
assign LUT_2[62415] = 32'b11111111111111101100101011011111;
assign LUT_2[62416] = 32'b11111111111111101100001111001111;
assign LUT_2[62417] = 32'b11111111111111101001000111101000;
assign LUT_2[62418] = 32'b11111111111111110011001000001011;
assign LUT_2[62419] = 32'b11111111111111110000000000100100;
assign LUT_2[62420] = 32'b11111111111111101000101100110111;
assign LUT_2[62421] = 32'b11111111111111100101100101010000;
assign LUT_2[62422] = 32'b11111111111111101111100101110011;
assign LUT_2[62423] = 32'b11111111111111101100011110001100;
assign LUT_2[62424] = 32'b11111111111111100111000000101100;
assign LUT_2[62425] = 32'b11111111111111100011111001000101;
assign LUT_2[62426] = 32'b11111111111111101101111001101000;
assign LUT_2[62427] = 32'b11111111111111101010110010000001;
assign LUT_2[62428] = 32'b11111111111111100011011110010100;
assign LUT_2[62429] = 32'b11111111111111100000010110101101;
assign LUT_2[62430] = 32'b11111111111111101010010111010000;
assign LUT_2[62431] = 32'b11111111111111100111001111101001;
assign LUT_2[62432] = 32'b11111111111111110010000110101110;
assign LUT_2[62433] = 32'b11111111111111101110111111000111;
assign LUT_2[62434] = 32'b11111111111111111000111111101010;
assign LUT_2[62435] = 32'b11111111111111110101111000000011;
assign LUT_2[62436] = 32'b11111111111111101110100100010110;
assign LUT_2[62437] = 32'b11111111111111101011011100101111;
assign LUT_2[62438] = 32'b11111111111111110101011101010010;
assign LUT_2[62439] = 32'b11111111111111110010010101101011;
assign LUT_2[62440] = 32'b11111111111111101100111000001011;
assign LUT_2[62441] = 32'b11111111111111101001110000100100;
assign LUT_2[62442] = 32'b11111111111111110011110001000111;
assign LUT_2[62443] = 32'b11111111111111110000101001100000;
assign LUT_2[62444] = 32'b11111111111111101001010101110011;
assign LUT_2[62445] = 32'b11111111111111100110001110001100;
assign LUT_2[62446] = 32'b11111111111111110000001110101111;
assign LUT_2[62447] = 32'b11111111111111101101000111001000;
assign LUT_2[62448] = 32'b11111111111111101100101010111000;
assign LUT_2[62449] = 32'b11111111111111101001100011010001;
assign LUT_2[62450] = 32'b11111111111111110011100011110100;
assign LUT_2[62451] = 32'b11111111111111110000011100001101;
assign LUT_2[62452] = 32'b11111111111111101001001000100000;
assign LUT_2[62453] = 32'b11111111111111100110000000111001;
assign LUT_2[62454] = 32'b11111111111111110000000001011100;
assign LUT_2[62455] = 32'b11111111111111101100111001110101;
assign LUT_2[62456] = 32'b11111111111111100111011100010101;
assign LUT_2[62457] = 32'b11111111111111100100010100101110;
assign LUT_2[62458] = 32'b11111111111111101110010101010001;
assign LUT_2[62459] = 32'b11111111111111101011001101101010;
assign LUT_2[62460] = 32'b11111111111111100011111001111101;
assign LUT_2[62461] = 32'b11111111111111100000110010010110;
assign LUT_2[62462] = 32'b11111111111111101010110010111001;
assign LUT_2[62463] = 32'b11111111111111100111101011010010;
assign LUT_2[62464] = 32'b11111111111111110011001010000000;
assign LUT_2[62465] = 32'b11111111111111110000000010011001;
assign LUT_2[62466] = 32'b11111111111111111010000010111100;
assign LUT_2[62467] = 32'b11111111111111110110111011010101;
assign LUT_2[62468] = 32'b11111111111111101111100111101000;
assign LUT_2[62469] = 32'b11111111111111101100100000000001;
assign LUT_2[62470] = 32'b11111111111111110110100000100100;
assign LUT_2[62471] = 32'b11111111111111110011011000111101;
assign LUT_2[62472] = 32'b11111111111111101101111011011101;
assign LUT_2[62473] = 32'b11111111111111101010110011110110;
assign LUT_2[62474] = 32'b11111111111111110100110100011001;
assign LUT_2[62475] = 32'b11111111111111110001101100110010;
assign LUT_2[62476] = 32'b11111111111111101010011001000101;
assign LUT_2[62477] = 32'b11111111111111100111010001011110;
assign LUT_2[62478] = 32'b11111111111111110001010010000001;
assign LUT_2[62479] = 32'b11111111111111101110001010011010;
assign LUT_2[62480] = 32'b11111111111111101101101110001010;
assign LUT_2[62481] = 32'b11111111111111101010100110100011;
assign LUT_2[62482] = 32'b11111111111111110100100111000110;
assign LUT_2[62483] = 32'b11111111111111110001011111011111;
assign LUT_2[62484] = 32'b11111111111111101010001011110010;
assign LUT_2[62485] = 32'b11111111111111100111000100001011;
assign LUT_2[62486] = 32'b11111111111111110001000100101110;
assign LUT_2[62487] = 32'b11111111111111101101111101000111;
assign LUT_2[62488] = 32'b11111111111111101000011111100111;
assign LUT_2[62489] = 32'b11111111111111100101011000000000;
assign LUT_2[62490] = 32'b11111111111111101111011000100011;
assign LUT_2[62491] = 32'b11111111111111101100010000111100;
assign LUT_2[62492] = 32'b11111111111111100100111101001111;
assign LUT_2[62493] = 32'b11111111111111100001110101101000;
assign LUT_2[62494] = 32'b11111111111111101011110110001011;
assign LUT_2[62495] = 32'b11111111111111101000101110100100;
assign LUT_2[62496] = 32'b11111111111111110011100101101001;
assign LUT_2[62497] = 32'b11111111111111110000011110000010;
assign LUT_2[62498] = 32'b11111111111111111010011110100101;
assign LUT_2[62499] = 32'b11111111111111110111010110111110;
assign LUT_2[62500] = 32'b11111111111111110000000011010001;
assign LUT_2[62501] = 32'b11111111111111101100111011101010;
assign LUT_2[62502] = 32'b11111111111111110110111100001101;
assign LUT_2[62503] = 32'b11111111111111110011110100100110;
assign LUT_2[62504] = 32'b11111111111111101110010111000110;
assign LUT_2[62505] = 32'b11111111111111101011001111011111;
assign LUT_2[62506] = 32'b11111111111111110101010000000010;
assign LUT_2[62507] = 32'b11111111111111110010001000011011;
assign LUT_2[62508] = 32'b11111111111111101010110100101110;
assign LUT_2[62509] = 32'b11111111111111100111101101000111;
assign LUT_2[62510] = 32'b11111111111111110001101101101010;
assign LUT_2[62511] = 32'b11111111111111101110100110000011;
assign LUT_2[62512] = 32'b11111111111111101110001001110011;
assign LUT_2[62513] = 32'b11111111111111101011000010001100;
assign LUT_2[62514] = 32'b11111111111111110101000010101111;
assign LUT_2[62515] = 32'b11111111111111110001111011001000;
assign LUT_2[62516] = 32'b11111111111111101010100111011011;
assign LUT_2[62517] = 32'b11111111111111100111011111110100;
assign LUT_2[62518] = 32'b11111111111111110001100000010111;
assign LUT_2[62519] = 32'b11111111111111101110011000110000;
assign LUT_2[62520] = 32'b11111111111111101000111011010000;
assign LUT_2[62521] = 32'b11111111111111100101110011101001;
assign LUT_2[62522] = 32'b11111111111111101111110100001100;
assign LUT_2[62523] = 32'b11111111111111101100101100100101;
assign LUT_2[62524] = 32'b11111111111111100101011000111000;
assign LUT_2[62525] = 32'b11111111111111100010010001010001;
assign LUT_2[62526] = 32'b11111111111111101100010001110100;
assign LUT_2[62527] = 32'b11111111111111101001001010001101;
assign LUT_2[62528] = 32'b11111111111111101011010010100011;
assign LUT_2[62529] = 32'b11111111111111101000001010111100;
assign LUT_2[62530] = 32'b11111111111111110010001011011111;
assign LUT_2[62531] = 32'b11111111111111101111000011111000;
assign LUT_2[62532] = 32'b11111111111111100111110000001011;
assign LUT_2[62533] = 32'b11111111111111100100101000100100;
assign LUT_2[62534] = 32'b11111111111111101110101001000111;
assign LUT_2[62535] = 32'b11111111111111101011100001100000;
assign LUT_2[62536] = 32'b11111111111111100110000100000000;
assign LUT_2[62537] = 32'b11111111111111100010111100011001;
assign LUT_2[62538] = 32'b11111111111111101100111100111100;
assign LUT_2[62539] = 32'b11111111111111101001110101010101;
assign LUT_2[62540] = 32'b11111111111111100010100001101000;
assign LUT_2[62541] = 32'b11111111111111011111011010000001;
assign LUT_2[62542] = 32'b11111111111111101001011010100100;
assign LUT_2[62543] = 32'b11111111111111100110010010111101;
assign LUT_2[62544] = 32'b11111111111111100101110110101101;
assign LUT_2[62545] = 32'b11111111111111100010101111000110;
assign LUT_2[62546] = 32'b11111111111111101100101111101001;
assign LUT_2[62547] = 32'b11111111111111101001101000000010;
assign LUT_2[62548] = 32'b11111111111111100010010100010101;
assign LUT_2[62549] = 32'b11111111111111011111001100101110;
assign LUT_2[62550] = 32'b11111111111111101001001101010001;
assign LUT_2[62551] = 32'b11111111111111100110000101101010;
assign LUT_2[62552] = 32'b11111111111111100000101000001010;
assign LUT_2[62553] = 32'b11111111111111011101100000100011;
assign LUT_2[62554] = 32'b11111111111111100111100001000110;
assign LUT_2[62555] = 32'b11111111111111100100011001011111;
assign LUT_2[62556] = 32'b11111111111111011101000101110010;
assign LUT_2[62557] = 32'b11111111111111011001111110001011;
assign LUT_2[62558] = 32'b11111111111111100011111110101110;
assign LUT_2[62559] = 32'b11111111111111100000110111000111;
assign LUT_2[62560] = 32'b11111111111111101011101110001100;
assign LUT_2[62561] = 32'b11111111111111101000100110100101;
assign LUT_2[62562] = 32'b11111111111111110010100111001000;
assign LUT_2[62563] = 32'b11111111111111101111011111100001;
assign LUT_2[62564] = 32'b11111111111111101000001011110100;
assign LUT_2[62565] = 32'b11111111111111100101000100001101;
assign LUT_2[62566] = 32'b11111111111111101111000100110000;
assign LUT_2[62567] = 32'b11111111111111101011111101001001;
assign LUT_2[62568] = 32'b11111111111111100110011111101001;
assign LUT_2[62569] = 32'b11111111111111100011011000000010;
assign LUT_2[62570] = 32'b11111111111111101101011000100101;
assign LUT_2[62571] = 32'b11111111111111101010010000111110;
assign LUT_2[62572] = 32'b11111111111111100010111101010001;
assign LUT_2[62573] = 32'b11111111111111011111110101101010;
assign LUT_2[62574] = 32'b11111111111111101001110110001101;
assign LUT_2[62575] = 32'b11111111111111100110101110100110;
assign LUT_2[62576] = 32'b11111111111111100110010010010110;
assign LUT_2[62577] = 32'b11111111111111100011001010101111;
assign LUT_2[62578] = 32'b11111111111111101101001011010010;
assign LUT_2[62579] = 32'b11111111111111101010000011101011;
assign LUT_2[62580] = 32'b11111111111111100010101111111110;
assign LUT_2[62581] = 32'b11111111111111011111101000010111;
assign LUT_2[62582] = 32'b11111111111111101001101000111010;
assign LUT_2[62583] = 32'b11111111111111100110100001010011;
assign LUT_2[62584] = 32'b11111111111111100001000011110011;
assign LUT_2[62585] = 32'b11111111111111011101111100001100;
assign LUT_2[62586] = 32'b11111111111111100111111100101111;
assign LUT_2[62587] = 32'b11111111111111100100110101001000;
assign LUT_2[62588] = 32'b11111111111111011101100001011011;
assign LUT_2[62589] = 32'b11111111111111011010011001110100;
assign LUT_2[62590] = 32'b11111111111111100100011010010111;
assign LUT_2[62591] = 32'b11111111111111100001010010110000;
assign LUT_2[62592] = 32'b11111111111111110111011110001111;
assign LUT_2[62593] = 32'b11111111111111110100010110101000;
assign LUT_2[62594] = 32'b11111111111111111110010111001011;
assign LUT_2[62595] = 32'b11111111111111111011001111100100;
assign LUT_2[62596] = 32'b11111111111111110011111011110111;
assign LUT_2[62597] = 32'b11111111111111110000110100010000;
assign LUT_2[62598] = 32'b11111111111111111010110100110011;
assign LUT_2[62599] = 32'b11111111111111110111101101001100;
assign LUT_2[62600] = 32'b11111111111111110010001111101100;
assign LUT_2[62601] = 32'b11111111111111101111001000000101;
assign LUT_2[62602] = 32'b11111111111111111001001000101000;
assign LUT_2[62603] = 32'b11111111111111110110000001000001;
assign LUT_2[62604] = 32'b11111111111111101110101101010100;
assign LUT_2[62605] = 32'b11111111111111101011100101101101;
assign LUT_2[62606] = 32'b11111111111111110101100110010000;
assign LUT_2[62607] = 32'b11111111111111110010011110101001;
assign LUT_2[62608] = 32'b11111111111111110010000010011001;
assign LUT_2[62609] = 32'b11111111111111101110111010110010;
assign LUT_2[62610] = 32'b11111111111111111000111011010101;
assign LUT_2[62611] = 32'b11111111111111110101110011101110;
assign LUT_2[62612] = 32'b11111111111111101110100000000001;
assign LUT_2[62613] = 32'b11111111111111101011011000011010;
assign LUT_2[62614] = 32'b11111111111111110101011000111101;
assign LUT_2[62615] = 32'b11111111111111110010010001010110;
assign LUT_2[62616] = 32'b11111111111111101100110011110110;
assign LUT_2[62617] = 32'b11111111111111101001101100001111;
assign LUT_2[62618] = 32'b11111111111111110011101100110010;
assign LUT_2[62619] = 32'b11111111111111110000100101001011;
assign LUT_2[62620] = 32'b11111111111111101001010001011110;
assign LUT_2[62621] = 32'b11111111111111100110001001110111;
assign LUT_2[62622] = 32'b11111111111111110000001010011010;
assign LUT_2[62623] = 32'b11111111111111101101000010110011;
assign LUT_2[62624] = 32'b11111111111111110111111001111000;
assign LUT_2[62625] = 32'b11111111111111110100110010010001;
assign LUT_2[62626] = 32'b11111111111111111110110010110100;
assign LUT_2[62627] = 32'b11111111111111111011101011001101;
assign LUT_2[62628] = 32'b11111111111111110100010111100000;
assign LUT_2[62629] = 32'b11111111111111110001001111111001;
assign LUT_2[62630] = 32'b11111111111111111011010000011100;
assign LUT_2[62631] = 32'b11111111111111111000001000110101;
assign LUT_2[62632] = 32'b11111111111111110010101011010101;
assign LUT_2[62633] = 32'b11111111111111101111100011101110;
assign LUT_2[62634] = 32'b11111111111111111001100100010001;
assign LUT_2[62635] = 32'b11111111111111110110011100101010;
assign LUT_2[62636] = 32'b11111111111111101111001000111101;
assign LUT_2[62637] = 32'b11111111111111101100000001010110;
assign LUT_2[62638] = 32'b11111111111111110110000001111001;
assign LUT_2[62639] = 32'b11111111111111110010111010010010;
assign LUT_2[62640] = 32'b11111111111111110010011110000010;
assign LUT_2[62641] = 32'b11111111111111101111010110011011;
assign LUT_2[62642] = 32'b11111111111111111001010110111110;
assign LUT_2[62643] = 32'b11111111111111110110001111010111;
assign LUT_2[62644] = 32'b11111111111111101110111011101010;
assign LUT_2[62645] = 32'b11111111111111101011110100000011;
assign LUT_2[62646] = 32'b11111111111111110101110100100110;
assign LUT_2[62647] = 32'b11111111111111110010101100111111;
assign LUT_2[62648] = 32'b11111111111111101101001111011111;
assign LUT_2[62649] = 32'b11111111111111101010000111111000;
assign LUT_2[62650] = 32'b11111111111111110100001000011011;
assign LUT_2[62651] = 32'b11111111111111110001000000110100;
assign LUT_2[62652] = 32'b11111111111111101001101101000111;
assign LUT_2[62653] = 32'b11111111111111100110100101100000;
assign LUT_2[62654] = 32'b11111111111111110000100110000011;
assign LUT_2[62655] = 32'b11111111111111101101011110011100;
assign LUT_2[62656] = 32'b11111111111111101111100110110010;
assign LUT_2[62657] = 32'b11111111111111101100011111001011;
assign LUT_2[62658] = 32'b11111111111111110110011111101110;
assign LUT_2[62659] = 32'b11111111111111110011011000000111;
assign LUT_2[62660] = 32'b11111111111111101100000100011010;
assign LUT_2[62661] = 32'b11111111111111101000111100110011;
assign LUT_2[62662] = 32'b11111111111111110010111101010110;
assign LUT_2[62663] = 32'b11111111111111101111110101101111;
assign LUT_2[62664] = 32'b11111111111111101010011000001111;
assign LUT_2[62665] = 32'b11111111111111100111010000101000;
assign LUT_2[62666] = 32'b11111111111111110001010001001011;
assign LUT_2[62667] = 32'b11111111111111101110001001100100;
assign LUT_2[62668] = 32'b11111111111111100110110101110111;
assign LUT_2[62669] = 32'b11111111111111100011101110010000;
assign LUT_2[62670] = 32'b11111111111111101101101110110011;
assign LUT_2[62671] = 32'b11111111111111101010100111001100;
assign LUT_2[62672] = 32'b11111111111111101010001010111100;
assign LUT_2[62673] = 32'b11111111111111100111000011010101;
assign LUT_2[62674] = 32'b11111111111111110001000011111000;
assign LUT_2[62675] = 32'b11111111111111101101111100010001;
assign LUT_2[62676] = 32'b11111111111111100110101000100100;
assign LUT_2[62677] = 32'b11111111111111100011100000111101;
assign LUT_2[62678] = 32'b11111111111111101101100001100000;
assign LUT_2[62679] = 32'b11111111111111101010011001111001;
assign LUT_2[62680] = 32'b11111111111111100100111100011001;
assign LUT_2[62681] = 32'b11111111111111100001110100110010;
assign LUT_2[62682] = 32'b11111111111111101011110101010101;
assign LUT_2[62683] = 32'b11111111111111101000101101101110;
assign LUT_2[62684] = 32'b11111111111111100001011010000001;
assign LUT_2[62685] = 32'b11111111111111011110010010011010;
assign LUT_2[62686] = 32'b11111111111111101000010010111101;
assign LUT_2[62687] = 32'b11111111111111100101001011010110;
assign LUT_2[62688] = 32'b11111111111111110000000010011011;
assign LUT_2[62689] = 32'b11111111111111101100111010110100;
assign LUT_2[62690] = 32'b11111111111111110110111011010111;
assign LUT_2[62691] = 32'b11111111111111110011110011110000;
assign LUT_2[62692] = 32'b11111111111111101100100000000011;
assign LUT_2[62693] = 32'b11111111111111101001011000011100;
assign LUT_2[62694] = 32'b11111111111111110011011000111111;
assign LUT_2[62695] = 32'b11111111111111110000010001011000;
assign LUT_2[62696] = 32'b11111111111111101010110011111000;
assign LUT_2[62697] = 32'b11111111111111100111101100010001;
assign LUT_2[62698] = 32'b11111111111111110001101100110100;
assign LUT_2[62699] = 32'b11111111111111101110100101001101;
assign LUT_2[62700] = 32'b11111111111111100111010001100000;
assign LUT_2[62701] = 32'b11111111111111100100001001111001;
assign LUT_2[62702] = 32'b11111111111111101110001010011100;
assign LUT_2[62703] = 32'b11111111111111101011000010110101;
assign LUT_2[62704] = 32'b11111111111111101010100110100101;
assign LUT_2[62705] = 32'b11111111111111100111011110111110;
assign LUT_2[62706] = 32'b11111111111111110001011111100001;
assign LUT_2[62707] = 32'b11111111111111101110010111111010;
assign LUT_2[62708] = 32'b11111111111111100111000100001101;
assign LUT_2[62709] = 32'b11111111111111100011111100100110;
assign LUT_2[62710] = 32'b11111111111111101101111101001001;
assign LUT_2[62711] = 32'b11111111111111101010110101100010;
assign LUT_2[62712] = 32'b11111111111111100101011000000010;
assign LUT_2[62713] = 32'b11111111111111100010010000011011;
assign LUT_2[62714] = 32'b11111111111111101100010000111110;
assign LUT_2[62715] = 32'b11111111111111101001001001010111;
assign LUT_2[62716] = 32'b11111111111111100001110101101010;
assign LUT_2[62717] = 32'b11111111111111011110101110000011;
assign LUT_2[62718] = 32'b11111111111111101000101110100110;
assign LUT_2[62719] = 32'b11111111111111100101100110111111;
assign LUT_2[62720] = 32'b11111111111111110111001000100110;
assign LUT_2[62721] = 32'b11111111111111110100000000111111;
assign LUT_2[62722] = 32'b11111111111111111110000001100010;
assign LUT_2[62723] = 32'b11111111111111111010111001111011;
assign LUT_2[62724] = 32'b11111111111111110011100110001110;
assign LUT_2[62725] = 32'b11111111111111110000011110100111;
assign LUT_2[62726] = 32'b11111111111111111010011111001010;
assign LUT_2[62727] = 32'b11111111111111110111010111100011;
assign LUT_2[62728] = 32'b11111111111111110001111010000011;
assign LUT_2[62729] = 32'b11111111111111101110110010011100;
assign LUT_2[62730] = 32'b11111111111111111000110010111111;
assign LUT_2[62731] = 32'b11111111111111110101101011011000;
assign LUT_2[62732] = 32'b11111111111111101110010111101011;
assign LUT_2[62733] = 32'b11111111111111101011010000000100;
assign LUT_2[62734] = 32'b11111111111111110101010000100111;
assign LUT_2[62735] = 32'b11111111111111110010001001000000;
assign LUT_2[62736] = 32'b11111111111111110001101100110000;
assign LUT_2[62737] = 32'b11111111111111101110100101001001;
assign LUT_2[62738] = 32'b11111111111111111000100101101100;
assign LUT_2[62739] = 32'b11111111111111110101011110000101;
assign LUT_2[62740] = 32'b11111111111111101110001010011000;
assign LUT_2[62741] = 32'b11111111111111101011000010110001;
assign LUT_2[62742] = 32'b11111111111111110101000011010100;
assign LUT_2[62743] = 32'b11111111111111110001111011101101;
assign LUT_2[62744] = 32'b11111111111111101100011110001101;
assign LUT_2[62745] = 32'b11111111111111101001010110100110;
assign LUT_2[62746] = 32'b11111111111111110011010111001001;
assign LUT_2[62747] = 32'b11111111111111110000001111100010;
assign LUT_2[62748] = 32'b11111111111111101000111011110101;
assign LUT_2[62749] = 32'b11111111111111100101110100001110;
assign LUT_2[62750] = 32'b11111111111111101111110100110001;
assign LUT_2[62751] = 32'b11111111111111101100101101001010;
assign LUT_2[62752] = 32'b11111111111111110111100100001111;
assign LUT_2[62753] = 32'b11111111111111110100011100101000;
assign LUT_2[62754] = 32'b11111111111111111110011101001011;
assign LUT_2[62755] = 32'b11111111111111111011010101100100;
assign LUT_2[62756] = 32'b11111111111111110100000001110111;
assign LUT_2[62757] = 32'b11111111111111110000111010010000;
assign LUT_2[62758] = 32'b11111111111111111010111010110011;
assign LUT_2[62759] = 32'b11111111111111110111110011001100;
assign LUT_2[62760] = 32'b11111111111111110010010101101100;
assign LUT_2[62761] = 32'b11111111111111101111001110000101;
assign LUT_2[62762] = 32'b11111111111111111001001110101000;
assign LUT_2[62763] = 32'b11111111111111110110000111000001;
assign LUT_2[62764] = 32'b11111111111111101110110011010100;
assign LUT_2[62765] = 32'b11111111111111101011101011101101;
assign LUT_2[62766] = 32'b11111111111111110101101100010000;
assign LUT_2[62767] = 32'b11111111111111110010100100101001;
assign LUT_2[62768] = 32'b11111111111111110010001000011001;
assign LUT_2[62769] = 32'b11111111111111101111000000110010;
assign LUT_2[62770] = 32'b11111111111111111001000001010101;
assign LUT_2[62771] = 32'b11111111111111110101111001101110;
assign LUT_2[62772] = 32'b11111111111111101110100110000001;
assign LUT_2[62773] = 32'b11111111111111101011011110011010;
assign LUT_2[62774] = 32'b11111111111111110101011110111101;
assign LUT_2[62775] = 32'b11111111111111110010010111010110;
assign LUT_2[62776] = 32'b11111111111111101100111001110110;
assign LUT_2[62777] = 32'b11111111111111101001110010001111;
assign LUT_2[62778] = 32'b11111111111111110011110010110010;
assign LUT_2[62779] = 32'b11111111111111110000101011001011;
assign LUT_2[62780] = 32'b11111111111111101001010111011110;
assign LUT_2[62781] = 32'b11111111111111100110001111110111;
assign LUT_2[62782] = 32'b11111111111111110000010000011010;
assign LUT_2[62783] = 32'b11111111111111101101001000110011;
assign LUT_2[62784] = 32'b11111111111111101111010001001001;
assign LUT_2[62785] = 32'b11111111111111101100001001100010;
assign LUT_2[62786] = 32'b11111111111111110110001010000101;
assign LUT_2[62787] = 32'b11111111111111110011000010011110;
assign LUT_2[62788] = 32'b11111111111111101011101110110001;
assign LUT_2[62789] = 32'b11111111111111101000100111001010;
assign LUT_2[62790] = 32'b11111111111111110010100111101101;
assign LUT_2[62791] = 32'b11111111111111101111100000000110;
assign LUT_2[62792] = 32'b11111111111111101010000010100110;
assign LUT_2[62793] = 32'b11111111111111100110111010111111;
assign LUT_2[62794] = 32'b11111111111111110000111011100010;
assign LUT_2[62795] = 32'b11111111111111101101110011111011;
assign LUT_2[62796] = 32'b11111111111111100110100000001110;
assign LUT_2[62797] = 32'b11111111111111100011011000100111;
assign LUT_2[62798] = 32'b11111111111111101101011001001010;
assign LUT_2[62799] = 32'b11111111111111101010010001100011;
assign LUT_2[62800] = 32'b11111111111111101001110101010011;
assign LUT_2[62801] = 32'b11111111111111100110101101101100;
assign LUT_2[62802] = 32'b11111111111111110000101110001111;
assign LUT_2[62803] = 32'b11111111111111101101100110101000;
assign LUT_2[62804] = 32'b11111111111111100110010010111011;
assign LUT_2[62805] = 32'b11111111111111100011001011010100;
assign LUT_2[62806] = 32'b11111111111111101101001011110111;
assign LUT_2[62807] = 32'b11111111111111101010000100010000;
assign LUT_2[62808] = 32'b11111111111111100100100110110000;
assign LUT_2[62809] = 32'b11111111111111100001011111001001;
assign LUT_2[62810] = 32'b11111111111111101011011111101100;
assign LUT_2[62811] = 32'b11111111111111101000011000000101;
assign LUT_2[62812] = 32'b11111111111111100001000100011000;
assign LUT_2[62813] = 32'b11111111111111011101111100110001;
assign LUT_2[62814] = 32'b11111111111111100111111101010100;
assign LUT_2[62815] = 32'b11111111111111100100110101101101;
assign LUT_2[62816] = 32'b11111111111111101111101100110010;
assign LUT_2[62817] = 32'b11111111111111101100100101001011;
assign LUT_2[62818] = 32'b11111111111111110110100101101110;
assign LUT_2[62819] = 32'b11111111111111110011011110000111;
assign LUT_2[62820] = 32'b11111111111111101100001010011010;
assign LUT_2[62821] = 32'b11111111111111101001000010110011;
assign LUT_2[62822] = 32'b11111111111111110011000011010110;
assign LUT_2[62823] = 32'b11111111111111101111111011101111;
assign LUT_2[62824] = 32'b11111111111111101010011110001111;
assign LUT_2[62825] = 32'b11111111111111100111010110101000;
assign LUT_2[62826] = 32'b11111111111111110001010111001011;
assign LUT_2[62827] = 32'b11111111111111101110001111100100;
assign LUT_2[62828] = 32'b11111111111111100110111011110111;
assign LUT_2[62829] = 32'b11111111111111100011110100010000;
assign LUT_2[62830] = 32'b11111111111111101101110100110011;
assign LUT_2[62831] = 32'b11111111111111101010101101001100;
assign LUT_2[62832] = 32'b11111111111111101010010000111100;
assign LUT_2[62833] = 32'b11111111111111100111001001010101;
assign LUT_2[62834] = 32'b11111111111111110001001001111000;
assign LUT_2[62835] = 32'b11111111111111101110000010010001;
assign LUT_2[62836] = 32'b11111111111111100110101110100100;
assign LUT_2[62837] = 32'b11111111111111100011100110111101;
assign LUT_2[62838] = 32'b11111111111111101101100111100000;
assign LUT_2[62839] = 32'b11111111111111101010011111111001;
assign LUT_2[62840] = 32'b11111111111111100101000010011001;
assign LUT_2[62841] = 32'b11111111111111100001111010110010;
assign LUT_2[62842] = 32'b11111111111111101011111011010101;
assign LUT_2[62843] = 32'b11111111111111101000110011101110;
assign LUT_2[62844] = 32'b11111111111111100001100000000001;
assign LUT_2[62845] = 32'b11111111111111011110011000011010;
assign LUT_2[62846] = 32'b11111111111111101000011000111101;
assign LUT_2[62847] = 32'b11111111111111100101010001010110;
assign LUT_2[62848] = 32'b11111111111111111011011100110101;
assign LUT_2[62849] = 32'b11111111111111111000010101001110;
assign LUT_2[62850] = 32'b00000000000000000010010101110001;
assign LUT_2[62851] = 32'b11111111111111111111001110001010;
assign LUT_2[62852] = 32'b11111111111111110111111010011101;
assign LUT_2[62853] = 32'b11111111111111110100110010110110;
assign LUT_2[62854] = 32'b11111111111111111110110011011001;
assign LUT_2[62855] = 32'b11111111111111111011101011110010;
assign LUT_2[62856] = 32'b11111111111111110110001110010010;
assign LUT_2[62857] = 32'b11111111111111110011000110101011;
assign LUT_2[62858] = 32'b11111111111111111101000111001110;
assign LUT_2[62859] = 32'b11111111111111111001111111100111;
assign LUT_2[62860] = 32'b11111111111111110010101011111010;
assign LUT_2[62861] = 32'b11111111111111101111100100010011;
assign LUT_2[62862] = 32'b11111111111111111001100100110110;
assign LUT_2[62863] = 32'b11111111111111110110011101001111;
assign LUT_2[62864] = 32'b11111111111111110110000000111111;
assign LUT_2[62865] = 32'b11111111111111110010111001011000;
assign LUT_2[62866] = 32'b11111111111111111100111001111011;
assign LUT_2[62867] = 32'b11111111111111111001110010010100;
assign LUT_2[62868] = 32'b11111111111111110010011110100111;
assign LUT_2[62869] = 32'b11111111111111101111010111000000;
assign LUT_2[62870] = 32'b11111111111111111001010111100011;
assign LUT_2[62871] = 32'b11111111111111110110001111111100;
assign LUT_2[62872] = 32'b11111111111111110000110010011100;
assign LUT_2[62873] = 32'b11111111111111101101101010110101;
assign LUT_2[62874] = 32'b11111111111111110111101011011000;
assign LUT_2[62875] = 32'b11111111111111110100100011110001;
assign LUT_2[62876] = 32'b11111111111111101101010000000100;
assign LUT_2[62877] = 32'b11111111111111101010001000011101;
assign LUT_2[62878] = 32'b11111111111111110100001001000000;
assign LUT_2[62879] = 32'b11111111111111110001000001011001;
assign LUT_2[62880] = 32'b11111111111111111011111000011110;
assign LUT_2[62881] = 32'b11111111111111111000110000110111;
assign LUT_2[62882] = 32'b00000000000000000010110001011010;
assign LUT_2[62883] = 32'b11111111111111111111101001110011;
assign LUT_2[62884] = 32'b11111111111111111000010110000110;
assign LUT_2[62885] = 32'b11111111111111110101001110011111;
assign LUT_2[62886] = 32'b11111111111111111111001111000010;
assign LUT_2[62887] = 32'b11111111111111111100000111011011;
assign LUT_2[62888] = 32'b11111111111111110110101001111011;
assign LUT_2[62889] = 32'b11111111111111110011100010010100;
assign LUT_2[62890] = 32'b11111111111111111101100010110111;
assign LUT_2[62891] = 32'b11111111111111111010011011010000;
assign LUT_2[62892] = 32'b11111111111111110011000111100011;
assign LUT_2[62893] = 32'b11111111111111101111111111111100;
assign LUT_2[62894] = 32'b11111111111111111010000000011111;
assign LUT_2[62895] = 32'b11111111111111110110111000111000;
assign LUT_2[62896] = 32'b11111111111111110110011100101000;
assign LUT_2[62897] = 32'b11111111111111110011010101000001;
assign LUT_2[62898] = 32'b11111111111111111101010101100100;
assign LUT_2[62899] = 32'b11111111111111111010001101111101;
assign LUT_2[62900] = 32'b11111111111111110010111010010000;
assign LUT_2[62901] = 32'b11111111111111101111110010101001;
assign LUT_2[62902] = 32'b11111111111111111001110011001100;
assign LUT_2[62903] = 32'b11111111111111110110101011100101;
assign LUT_2[62904] = 32'b11111111111111110001001110000101;
assign LUT_2[62905] = 32'b11111111111111101110000110011110;
assign LUT_2[62906] = 32'b11111111111111111000000111000001;
assign LUT_2[62907] = 32'b11111111111111110100111111011010;
assign LUT_2[62908] = 32'b11111111111111101101101011101101;
assign LUT_2[62909] = 32'b11111111111111101010100100000110;
assign LUT_2[62910] = 32'b11111111111111110100100100101001;
assign LUT_2[62911] = 32'b11111111111111110001011101000010;
assign LUT_2[62912] = 32'b11111111111111110011100101011000;
assign LUT_2[62913] = 32'b11111111111111110000011101110001;
assign LUT_2[62914] = 32'b11111111111111111010011110010100;
assign LUT_2[62915] = 32'b11111111111111110111010110101101;
assign LUT_2[62916] = 32'b11111111111111110000000011000000;
assign LUT_2[62917] = 32'b11111111111111101100111011011001;
assign LUT_2[62918] = 32'b11111111111111110110111011111100;
assign LUT_2[62919] = 32'b11111111111111110011110100010101;
assign LUT_2[62920] = 32'b11111111111111101110010110110101;
assign LUT_2[62921] = 32'b11111111111111101011001111001110;
assign LUT_2[62922] = 32'b11111111111111110101001111110001;
assign LUT_2[62923] = 32'b11111111111111110010001000001010;
assign LUT_2[62924] = 32'b11111111111111101010110100011101;
assign LUT_2[62925] = 32'b11111111111111100111101100110110;
assign LUT_2[62926] = 32'b11111111111111110001101101011001;
assign LUT_2[62927] = 32'b11111111111111101110100101110010;
assign LUT_2[62928] = 32'b11111111111111101110001001100010;
assign LUT_2[62929] = 32'b11111111111111101011000001111011;
assign LUT_2[62930] = 32'b11111111111111110101000010011110;
assign LUT_2[62931] = 32'b11111111111111110001111010110111;
assign LUT_2[62932] = 32'b11111111111111101010100111001010;
assign LUT_2[62933] = 32'b11111111111111100111011111100011;
assign LUT_2[62934] = 32'b11111111111111110001100000000110;
assign LUT_2[62935] = 32'b11111111111111101110011000011111;
assign LUT_2[62936] = 32'b11111111111111101000111010111111;
assign LUT_2[62937] = 32'b11111111111111100101110011011000;
assign LUT_2[62938] = 32'b11111111111111101111110011111011;
assign LUT_2[62939] = 32'b11111111111111101100101100010100;
assign LUT_2[62940] = 32'b11111111111111100101011000100111;
assign LUT_2[62941] = 32'b11111111111111100010010001000000;
assign LUT_2[62942] = 32'b11111111111111101100010001100011;
assign LUT_2[62943] = 32'b11111111111111101001001001111100;
assign LUT_2[62944] = 32'b11111111111111110100000001000001;
assign LUT_2[62945] = 32'b11111111111111110000111001011010;
assign LUT_2[62946] = 32'b11111111111111111010111001111101;
assign LUT_2[62947] = 32'b11111111111111110111110010010110;
assign LUT_2[62948] = 32'b11111111111111110000011110101001;
assign LUT_2[62949] = 32'b11111111111111101101010111000010;
assign LUT_2[62950] = 32'b11111111111111110111010111100101;
assign LUT_2[62951] = 32'b11111111111111110100001111111110;
assign LUT_2[62952] = 32'b11111111111111101110110010011110;
assign LUT_2[62953] = 32'b11111111111111101011101010110111;
assign LUT_2[62954] = 32'b11111111111111110101101011011010;
assign LUT_2[62955] = 32'b11111111111111110010100011110011;
assign LUT_2[62956] = 32'b11111111111111101011010000000110;
assign LUT_2[62957] = 32'b11111111111111101000001000011111;
assign LUT_2[62958] = 32'b11111111111111110010001001000010;
assign LUT_2[62959] = 32'b11111111111111101111000001011011;
assign LUT_2[62960] = 32'b11111111111111101110100101001011;
assign LUT_2[62961] = 32'b11111111111111101011011101100100;
assign LUT_2[62962] = 32'b11111111111111110101011110000111;
assign LUT_2[62963] = 32'b11111111111111110010010110100000;
assign LUT_2[62964] = 32'b11111111111111101011000010110011;
assign LUT_2[62965] = 32'b11111111111111100111111011001100;
assign LUT_2[62966] = 32'b11111111111111110001111011101111;
assign LUT_2[62967] = 32'b11111111111111101110110100001000;
assign LUT_2[62968] = 32'b11111111111111101001010110101000;
assign LUT_2[62969] = 32'b11111111111111100110001111000001;
assign LUT_2[62970] = 32'b11111111111111110000001111100100;
assign LUT_2[62971] = 32'b11111111111111101101000111111101;
assign LUT_2[62972] = 32'b11111111111111100101110100010000;
assign LUT_2[62973] = 32'b11111111111111100010101100101001;
assign LUT_2[62974] = 32'b11111111111111101100101101001100;
assign LUT_2[62975] = 32'b11111111111111101001100101100101;
assign LUT_2[62976] = 32'b11111111111111110111111011110010;
assign LUT_2[62977] = 32'b11111111111111110100110100001011;
assign LUT_2[62978] = 32'b11111111111111111110110100101110;
assign LUT_2[62979] = 32'b11111111111111111011101101000111;
assign LUT_2[62980] = 32'b11111111111111110100011001011010;
assign LUT_2[62981] = 32'b11111111111111110001010001110011;
assign LUT_2[62982] = 32'b11111111111111111011010010010110;
assign LUT_2[62983] = 32'b11111111111111111000001010101111;
assign LUT_2[62984] = 32'b11111111111111110010101101001111;
assign LUT_2[62985] = 32'b11111111111111101111100101101000;
assign LUT_2[62986] = 32'b11111111111111111001100110001011;
assign LUT_2[62987] = 32'b11111111111111110110011110100100;
assign LUT_2[62988] = 32'b11111111111111101111001010110111;
assign LUT_2[62989] = 32'b11111111111111101100000011010000;
assign LUT_2[62990] = 32'b11111111111111110110000011110011;
assign LUT_2[62991] = 32'b11111111111111110010111100001100;
assign LUT_2[62992] = 32'b11111111111111110010011111111100;
assign LUT_2[62993] = 32'b11111111111111101111011000010101;
assign LUT_2[62994] = 32'b11111111111111111001011000111000;
assign LUT_2[62995] = 32'b11111111111111110110010001010001;
assign LUT_2[62996] = 32'b11111111111111101110111101100100;
assign LUT_2[62997] = 32'b11111111111111101011110101111101;
assign LUT_2[62998] = 32'b11111111111111110101110110100000;
assign LUT_2[62999] = 32'b11111111111111110010101110111001;
assign LUT_2[63000] = 32'b11111111111111101101010001011001;
assign LUT_2[63001] = 32'b11111111111111101010001001110010;
assign LUT_2[63002] = 32'b11111111111111110100001010010101;
assign LUT_2[63003] = 32'b11111111111111110001000010101110;
assign LUT_2[63004] = 32'b11111111111111101001101111000001;
assign LUT_2[63005] = 32'b11111111111111100110100111011010;
assign LUT_2[63006] = 32'b11111111111111110000100111111101;
assign LUT_2[63007] = 32'b11111111111111101101100000010110;
assign LUT_2[63008] = 32'b11111111111111111000010111011011;
assign LUT_2[63009] = 32'b11111111111111110101001111110100;
assign LUT_2[63010] = 32'b11111111111111111111010000010111;
assign LUT_2[63011] = 32'b11111111111111111100001000110000;
assign LUT_2[63012] = 32'b11111111111111110100110101000011;
assign LUT_2[63013] = 32'b11111111111111110001101101011100;
assign LUT_2[63014] = 32'b11111111111111111011101101111111;
assign LUT_2[63015] = 32'b11111111111111111000100110011000;
assign LUT_2[63016] = 32'b11111111111111110011001000111000;
assign LUT_2[63017] = 32'b11111111111111110000000001010001;
assign LUT_2[63018] = 32'b11111111111111111010000001110100;
assign LUT_2[63019] = 32'b11111111111111110110111010001101;
assign LUT_2[63020] = 32'b11111111111111101111100110100000;
assign LUT_2[63021] = 32'b11111111111111101100011110111001;
assign LUT_2[63022] = 32'b11111111111111110110011111011100;
assign LUT_2[63023] = 32'b11111111111111110011010111110101;
assign LUT_2[63024] = 32'b11111111111111110010111011100101;
assign LUT_2[63025] = 32'b11111111111111101111110011111110;
assign LUT_2[63026] = 32'b11111111111111111001110100100001;
assign LUT_2[63027] = 32'b11111111111111110110101100111010;
assign LUT_2[63028] = 32'b11111111111111101111011001001101;
assign LUT_2[63029] = 32'b11111111111111101100010001100110;
assign LUT_2[63030] = 32'b11111111111111110110010010001001;
assign LUT_2[63031] = 32'b11111111111111110011001010100010;
assign LUT_2[63032] = 32'b11111111111111101101101101000010;
assign LUT_2[63033] = 32'b11111111111111101010100101011011;
assign LUT_2[63034] = 32'b11111111111111110100100101111110;
assign LUT_2[63035] = 32'b11111111111111110001011110010111;
assign LUT_2[63036] = 32'b11111111111111101010001010101010;
assign LUT_2[63037] = 32'b11111111111111100111000011000011;
assign LUT_2[63038] = 32'b11111111111111110001000011100110;
assign LUT_2[63039] = 32'b11111111111111101101111011111111;
assign LUT_2[63040] = 32'b11111111111111110000000100010101;
assign LUT_2[63041] = 32'b11111111111111101100111100101110;
assign LUT_2[63042] = 32'b11111111111111110110111101010001;
assign LUT_2[63043] = 32'b11111111111111110011110101101010;
assign LUT_2[63044] = 32'b11111111111111101100100001111101;
assign LUT_2[63045] = 32'b11111111111111101001011010010110;
assign LUT_2[63046] = 32'b11111111111111110011011010111001;
assign LUT_2[63047] = 32'b11111111111111110000010011010010;
assign LUT_2[63048] = 32'b11111111111111101010110101110010;
assign LUT_2[63049] = 32'b11111111111111100111101110001011;
assign LUT_2[63050] = 32'b11111111111111110001101110101110;
assign LUT_2[63051] = 32'b11111111111111101110100111000111;
assign LUT_2[63052] = 32'b11111111111111100111010011011010;
assign LUT_2[63053] = 32'b11111111111111100100001011110011;
assign LUT_2[63054] = 32'b11111111111111101110001100010110;
assign LUT_2[63055] = 32'b11111111111111101011000100101111;
assign LUT_2[63056] = 32'b11111111111111101010101000011111;
assign LUT_2[63057] = 32'b11111111111111100111100000111000;
assign LUT_2[63058] = 32'b11111111111111110001100001011011;
assign LUT_2[63059] = 32'b11111111111111101110011001110100;
assign LUT_2[63060] = 32'b11111111111111100111000110000111;
assign LUT_2[63061] = 32'b11111111111111100011111110100000;
assign LUT_2[63062] = 32'b11111111111111101101111111000011;
assign LUT_2[63063] = 32'b11111111111111101010110111011100;
assign LUT_2[63064] = 32'b11111111111111100101011001111100;
assign LUT_2[63065] = 32'b11111111111111100010010010010101;
assign LUT_2[63066] = 32'b11111111111111101100010010111000;
assign LUT_2[63067] = 32'b11111111111111101001001011010001;
assign LUT_2[63068] = 32'b11111111111111100001110111100100;
assign LUT_2[63069] = 32'b11111111111111011110101111111101;
assign LUT_2[63070] = 32'b11111111111111101000110000100000;
assign LUT_2[63071] = 32'b11111111111111100101101000111001;
assign LUT_2[63072] = 32'b11111111111111110000011111111110;
assign LUT_2[63073] = 32'b11111111111111101101011000010111;
assign LUT_2[63074] = 32'b11111111111111110111011000111010;
assign LUT_2[63075] = 32'b11111111111111110100010001010011;
assign LUT_2[63076] = 32'b11111111111111101100111101100110;
assign LUT_2[63077] = 32'b11111111111111101001110101111111;
assign LUT_2[63078] = 32'b11111111111111110011110110100010;
assign LUT_2[63079] = 32'b11111111111111110000101110111011;
assign LUT_2[63080] = 32'b11111111111111101011010001011011;
assign LUT_2[63081] = 32'b11111111111111101000001001110100;
assign LUT_2[63082] = 32'b11111111111111110010001010010111;
assign LUT_2[63083] = 32'b11111111111111101111000010110000;
assign LUT_2[63084] = 32'b11111111111111100111101111000011;
assign LUT_2[63085] = 32'b11111111111111100100100111011100;
assign LUT_2[63086] = 32'b11111111111111101110100111111111;
assign LUT_2[63087] = 32'b11111111111111101011100000011000;
assign LUT_2[63088] = 32'b11111111111111101011000100001000;
assign LUT_2[63089] = 32'b11111111111111100111111100100001;
assign LUT_2[63090] = 32'b11111111111111110001111101000100;
assign LUT_2[63091] = 32'b11111111111111101110110101011101;
assign LUT_2[63092] = 32'b11111111111111100111100001110000;
assign LUT_2[63093] = 32'b11111111111111100100011010001001;
assign LUT_2[63094] = 32'b11111111111111101110011010101100;
assign LUT_2[63095] = 32'b11111111111111101011010011000101;
assign LUT_2[63096] = 32'b11111111111111100101110101100101;
assign LUT_2[63097] = 32'b11111111111111100010101101111110;
assign LUT_2[63098] = 32'b11111111111111101100101110100001;
assign LUT_2[63099] = 32'b11111111111111101001100110111010;
assign LUT_2[63100] = 32'b11111111111111100010010011001101;
assign LUT_2[63101] = 32'b11111111111111011111001011100110;
assign LUT_2[63102] = 32'b11111111111111101001001100001001;
assign LUT_2[63103] = 32'b11111111111111100110000100100010;
assign LUT_2[63104] = 32'b11111111111111111100010000000001;
assign LUT_2[63105] = 32'b11111111111111111001001000011010;
assign LUT_2[63106] = 32'b00000000000000000011001000111101;
assign LUT_2[63107] = 32'b00000000000000000000000001010110;
assign LUT_2[63108] = 32'b11111111111111111000101101101001;
assign LUT_2[63109] = 32'b11111111111111110101100110000010;
assign LUT_2[63110] = 32'b11111111111111111111100110100101;
assign LUT_2[63111] = 32'b11111111111111111100011110111110;
assign LUT_2[63112] = 32'b11111111111111110111000001011110;
assign LUT_2[63113] = 32'b11111111111111110011111001110111;
assign LUT_2[63114] = 32'b11111111111111111101111010011010;
assign LUT_2[63115] = 32'b11111111111111111010110010110011;
assign LUT_2[63116] = 32'b11111111111111110011011111000110;
assign LUT_2[63117] = 32'b11111111111111110000010111011111;
assign LUT_2[63118] = 32'b11111111111111111010011000000010;
assign LUT_2[63119] = 32'b11111111111111110111010000011011;
assign LUT_2[63120] = 32'b11111111111111110110110100001011;
assign LUT_2[63121] = 32'b11111111111111110011101100100100;
assign LUT_2[63122] = 32'b11111111111111111101101101000111;
assign LUT_2[63123] = 32'b11111111111111111010100101100000;
assign LUT_2[63124] = 32'b11111111111111110011010001110011;
assign LUT_2[63125] = 32'b11111111111111110000001010001100;
assign LUT_2[63126] = 32'b11111111111111111010001010101111;
assign LUT_2[63127] = 32'b11111111111111110111000011001000;
assign LUT_2[63128] = 32'b11111111111111110001100101101000;
assign LUT_2[63129] = 32'b11111111111111101110011110000001;
assign LUT_2[63130] = 32'b11111111111111111000011110100100;
assign LUT_2[63131] = 32'b11111111111111110101010110111101;
assign LUT_2[63132] = 32'b11111111111111101110000011010000;
assign LUT_2[63133] = 32'b11111111111111101010111011101001;
assign LUT_2[63134] = 32'b11111111111111110100111100001100;
assign LUT_2[63135] = 32'b11111111111111110001110100100101;
assign LUT_2[63136] = 32'b11111111111111111100101011101010;
assign LUT_2[63137] = 32'b11111111111111111001100100000011;
assign LUT_2[63138] = 32'b00000000000000000011100100100110;
assign LUT_2[63139] = 32'b00000000000000000000011100111111;
assign LUT_2[63140] = 32'b11111111111111111001001001010010;
assign LUT_2[63141] = 32'b11111111111111110110000001101011;
assign LUT_2[63142] = 32'b00000000000000000000000010001110;
assign LUT_2[63143] = 32'b11111111111111111100111010100111;
assign LUT_2[63144] = 32'b11111111111111110111011101000111;
assign LUT_2[63145] = 32'b11111111111111110100010101100000;
assign LUT_2[63146] = 32'b11111111111111111110010110000011;
assign LUT_2[63147] = 32'b11111111111111111011001110011100;
assign LUT_2[63148] = 32'b11111111111111110011111010101111;
assign LUT_2[63149] = 32'b11111111111111110000110011001000;
assign LUT_2[63150] = 32'b11111111111111111010110011101011;
assign LUT_2[63151] = 32'b11111111111111110111101100000100;
assign LUT_2[63152] = 32'b11111111111111110111001111110100;
assign LUT_2[63153] = 32'b11111111111111110100001000001101;
assign LUT_2[63154] = 32'b11111111111111111110001000110000;
assign LUT_2[63155] = 32'b11111111111111111011000001001001;
assign LUT_2[63156] = 32'b11111111111111110011101101011100;
assign LUT_2[63157] = 32'b11111111111111110000100101110101;
assign LUT_2[63158] = 32'b11111111111111111010100110011000;
assign LUT_2[63159] = 32'b11111111111111110111011110110001;
assign LUT_2[63160] = 32'b11111111111111110010000001010001;
assign LUT_2[63161] = 32'b11111111111111101110111001101010;
assign LUT_2[63162] = 32'b11111111111111111000111010001101;
assign LUT_2[63163] = 32'b11111111111111110101110010100110;
assign LUT_2[63164] = 32'b11111111111111101110011110111001;
assign LUT_2[63165] = 32'b11111111111111101011010111010010;
assign LUT_2[63166] = 32'b11111111111111110101010111110101;
assign LUT_2[63167] = 32'b11111111111111110010010000001110;
assign LUT_2[63168] = 32'b11111111111111110100011000100100;
assign LUT_2[63169] = 32'b11111111111111110001010000111101;
assign LUT_2[63170] = 32'b11111111111111111011010001100000;
assign LUT_2[63171] = 32'b11111111111111111000001001111001;
assign LUT_2[63172] = 32'b11111111111111110000110110001100;
assign LUT_2[63173] = 32'b11111111111111101101101110100101;
assign LUT_2[63174] = 32'b11111111111111110111101111001000;
assign LUT_2[63175] = 32'b11111111111111110100100111100001;
assign LUT_2[63176] = 32'b11111111111111101111001010000001;
assign LUT_2[63177] = 32'b11111111111111101100000010011010;
assign LUT_2[63178] = 32'b11111111111111110110000010111101;
assign LUT_2[63179] = 32'b11111111111111110010111011010110;
assign LUT_2[63180] = 32'b11111111111111101011100111101001;
assign LUT_2[63181] = 32'b11111111111111101000100000000010;
assign LUT_2[63182] = 32'b11111111111111110010100000100101;
assign LUT_2[63183] = 32'b11111111111111101111011000111110;
assign LUT_2[63184] = 32'b11111111111111101110111100101110;
assign LUT_2[63185] = 32'b11111111111111101011110101000111;
assign LUT_2[63186] = 32'b11111111111111110101110101101010;
assign LUT_2[63187] = 32'b11111111111111110010101110000011;
assign LUT_2[63188] = 32'b11111111111111101011011010010110;
assign LUT_2[63189] = 32'b11111111111111101000010010101111;
assign LUT_2[63190] = 32'b11111111111111110010010011010010;
assign LUT_2[63191] = 32'b11111111111111101111001011101011;
assign LUT_2[63192] = 32'b11111111111111101001101110001011;
assign LUT_2[63193] = 32'b11111111111111100110100110100100;
assign LUT_2[63194] = 32'b11111111111111110000100111000111;
assign LUT_2[63195] = 32'b11111111111111101101011111100000;
assign LUT_2[63196] = 32'b11111111111111100110001011110011;
assign LUT_2[63197] = 32'b11111111111111100011000100001100;
assign LUT_2[63198] = 32'b11111111111111101101000100101111;
assign LUT_2[63199] = 32'b11111111111111101001111101001000;
assign LUT_2[63200] = 32'b11111111111111110100110100001101;
assign LUT_2[63201] = 32'b11111111111111110001101100100110;
assign LUT_2[63202] = 32'b11111111111111111011101101001001;
assign LUT_2[63203] = 32'b11111111111111111000100101100010;
assign LUT_2[63204] = 32'b11111111111111110001010001110101;
assign LUT_2[63205] = 32'b11111111111111101110001010001110;
assign LUT_2[63206] = 32'b11111111111111111000001010110001;
assign LUT_2[63207] = 32'b11111111111111110101000011001010;
assign LUT_2[63208] = 32'b11111111111111101111100101101010;
assign LUT_2[63209] = 32'b11111111111111101100011110000011;
assign LUT_2[63210] = 32'b11111111111111110110011110100110;
assign LUT_2[63211] = 32'b11111111111111110011010110111111;
assign LUT_2[63212] = 32'b11111111111111101100000011010010;
assign LUT_2[63213] = 32'b11111111111111101000111011101011;
assign LUT_2[63214] = 32'b11111111111111110010111100001110;
assign LUT_2[63215] = 32'b11111111111111101111110100100111;
assign LUT_2[63216] = 32'b11111111111111101111011000010111;
assign LUT_2[63217] = 32'b11111111111111101100010000110000;
assign LUT_2[63218] = 32'b11111111111111110110010001010011;
assign LUT_2[63219] = 32'b11111111111111110011001001101100;
assign LUT_2[63220] = 32'b11111111111111101011110101111111;
assign LUT_2[63221] = 32'b11111111111111101000101110011000;
assign LUT_2[63222] = 32'b11111111111111110010101110111011;
assign LUT_2[63223] = 32'b11111111111111101111100111010100;
assign LUT_2[63224] = 32'b11111111111111101010001001110100;
assign LUT_2[63225] = 32'b11111111111111100111000010001101;
assign LUT_2[63226] = 32'b11111111111111110001000010110000;
assign LUT_2[63227] = 32'b11111111111111101101111011001001;
assign LUT_2[63228] = 32'b11111111111111100110100111011100;
assign LUT_2[63229] = 32'b11111111111111100011011111110101;
assign LUT_2[63230] = 32'b11111111111111101101100000011000;
assign LUT_2[63231] = 32'b11111111111111101010011000110001;
assign LUT_2[63232] = 32'b11111111111111111011111010011000;
assign LUT_2[63233] = 32'b11111111111111111000110010110001;
assign LUT_2[63234] = 32'b00000000000000000010110011010100;
assign LUT_2[63235] = 32'b11111111111111111111101011101101;
assign LUT_2[63236] = 32'b11111111111111111000011000000000;
assign LUT_2[63237] = 32'b11111111111111110101010000011001;
assign LUT_2[63238] = 32'b11111111111111111111010000111100;
assign LUT_2[63239] = 32'b11111111111111111100001001010101;
assign LUT_2[63240] = 32'b11111111111111110110101011110101;
assign LUT_2[63241] = 32'b11111111111111110011100100001110;
assign LUT_2[63242] = 32'b11111111111111111101100100110001;
assign LUT_2[63243] = 32'b11111111111111111010011101001010;
assign LUT_2[63244] = 32'b11111111111111110011001001011101;
assign LUT_2[63245] = 32'b11111111111111110000000001110110;
assign LUT_2[63246] = 32'b11111111111111111010000010011001;
assign LUT_2[63247] = 32'b11111111111111110110111010110010;
assign LUT_2[63248] = 32'b11111111111111110110011110100010;
assign LUT_2[63249] = 32'b11111111111111110011010110111011;
assign LUT_2[63250] = 32'b11111111111111111101010111011110;
assign LUT_2[63251] = 32'b11111111111111111010001111110111;
assign LUT_2[63252] = 32'b11111111111111110010111100001010;
assign LUT_2[63253] = 32'b11111111111111101111110100100011;
assign LUT_2[63254] = 32'b11111111111111111001110101000110;
assign LUT_2[63255] = 32'b11111111111111110110101101011111;
assign LUT_2[63256] = 32'b11111111111111110001001111111111;
assign LUT_2[63257] = 32'b11111111111111101110001000011000;
assign LUT_2[63258] = 32'b11111111111111111000001000111011;
assign LUT_2[63259] = 32'b11111111111111110101000001010100;
assign LUT_2[63260] = 32'b11111111111111101101101101100111;
assign LUT_2[63261] = 32'b11111111111111101010100110000000;
assign LUT_2[63262] = 32'b11111111111111110100100110100011;
assign LUT_2[63263] = 32'b11111111111111110001011110111100;
assign LUT_2[63264] = 32'b11111111111111111100010110000001;
assign LUT_2[63265] = 32'b11111111111111111001001110011010;
assign LUT_2[63266] = 32'b00000000000000000011001110111101;
assign LUT_2[63267] = 32'b00000000000000000000000111010110;
assign LUT_2[63268] = 32'b11111111111111111000110011101001;
assign LUT_2[63269] = 32'b11111111111111110101101100000010;
assign LUT_2[63270] = 32'b11111111111111111111101100100101;
assign LUT_2[63271] = 32'b11111111111111111100100100111110;
assign LUT_2[63272] = 32'b11111111111111110111000111011110;
assign LUT_2[63273] = 32'b11111111111111110011111111110111;
assign LUT_2[63274] = 32'b11111111111111111110000000011010;
assign LUT_2[63275] = 32'b11111111111111111010111000110011;
assign LUT_2[63276] = 32'b11111111111111110011100101000110;
assign LUT_2[63277] = 32'b11111111111111110000011101011111;
assign LUT_2[63278] = 32'b11111111111111111010011110000010;
assign LUT_2[63279] = 32'b11111111111111110111010110011011;
assign LUT_2[63280] = 32'b11111111111111110110111010001011;
assign LUT_2[63281] = 32'b11111111111111110011110010100100;
assign LUT_2[63282] = 32'b11111111111111111101110011000111;
assign LUT_2[63283] = 32'b11111111111111111010101011100000;
assign LUT_2[63284] = 32'b11111111111111110011010111110011;
assign LUT_2[63285] = 32'b11111111111111110000010000001100;
assign LUT_2[63286] = 32'b11111111111111111010010000101111;
assign LUT_2[63287] = 32'b11111111111111110111001001001000;
assign LUT_2[63288] = 32'b11111111111111110001101011101000;
assign LUT_2[63289] = 32'b11111111111111101110100100000001;
assign LUT_2[63290] = 32'b11111111111111111000100100100100;
assign LUT_2[63291] = 32'b11111111111111110101011100111101;
assign LUT_2[63292] = 32'b11111111111111101110001001010000;
assign LUT_2[63293] = 32'b11111111111111101011000001101001;
assign LUT_2[63294] = 32'b11111111111111110101000010001100;
assign LUT_2[63295] = 32'b11111111111111110001111010100101;
assign LUT_2[63296] = 32'b11111111111111110100000010111011;
assign LUT_2[63297] = 32'b11111111111111110000111011010100;
assign LUT_2[63298] = 32'b11111111111111111010111011110111;
assign LUT_2[63299] = 32'b11111111111111110111110100010000;
assign LUT_2[63300] = 32'b11111111111111110000100000100011;
assign LUT_2[63301] = 32'b11111111111111101101011000111100;
assign LUT_2[63302] = 32'b11111111111111110111011001011111;
assign LUT_2[63303] = 32'b11111111111111110100010001111000;
assign LUT_2[63304] = 32'b11111111111111101110110100011000;
assign LUT_2[63305] = 32'b11111111111111101011101100110001;
assign LUT_2[63306] = 32'b11111111111111110101101101010100;
assign LUT_2[63307] = 32'b11111111111111110010100101101101;
assign LUT_2[63308] = 32'b11111111111111101011010010000000;
assign LUT_2[63309] = 32'b11111111111111101000001010011001;
assign LUT_2[63310] = 32'b11111111111111110010001010111100;
assign LUT_2[63311] = 32'b11111111111111101111000011010101;
assign LUT_2[63312] = 32'b11111111111111101110100111000101;
assign LUT_2[63313] = 32'b11111111111111101011011111011110;
assign LUT_2[63314] = 32'b11111111111111110101100000000001;
assign LUT_2[63315] = 32'b11111111111111110010011000011010;
assign LUT_2[63316] = 32'b11111111111111101011000100101101;
assign LUT_2[63317] = 32'b11111111111111100111111101000110;
assign LUT_2[63318] = 32'b11111111111111110001111101101001;
assign LUT_2[63319] = 32'b11111111111111101110110110000010;
assign LUT_2[63320] = 32'b11111111111111101001011000100010;
assign LUT_2[63321] = 32'b11111111111111100110010000111011;
assign LUT_2[63322] = 32'b11111111111111110000010001011110;
assign LUT_2[63323] = 32'b11111111111111101101001001110111;
assign LUT_2[63324] = 32'b11111111111111100101110110001010;
assign LUT_2[63325] = 32'b11111111111111100010101110100011;
assign LUT_2[63326] = 32'b11111111111111101100101111000110;
assign LUT_2[63327] = 32'b11111111111111101001100111011111;
assign LUT_2[63328] = 32'b11111111111111110100011110100100;
assign LUT_2[63329] = 32'b11111111111111110001010110111101;
assign LUT_2[63330] = 32'b11111111111111111011010111100000;
assign LUT_2[63331] = 32'b11111111111111111000001111111001;
assign LUT_2[63332] = 32'b11111111111111110000111100001100;
assign LUT_2[63333] = 32'b11111111111111101101110100100101;
assign LUT_2[63334] = 32'b11111111111111110111110101001000;
assign LUT_2[63335] = 32'b11111111111111110100101101100001;
assign LUT_2[63336] = 32'b11111111111111101111010000000001;
assign LUT_2[63337] = 32'b11111111111111101100001000011010;
assign LUT_2[63338] = 32'b11111111111111110110001000111101;
assign LUT_2[63339] = 32'b11111111111111110011000001010110;
assign LUT_2[63340] = 32'b11111111111111101011101101101001;
assign LUT_2[63341] = 32'b11111111111111101000100110000010;
assign LUT_2[63342] = 32'b11111111111111110010100110100101;
assign LUT_2[63343] = 32'b11111111111111101111011110111110;
assign LUT_2[63344] = 32'b11111111111111101111000010101110;
assign LUT_2[63345] = 32'b11111111111111101011111011000111;
assign LUT_2[63346] = 32'b11111111111111110101111011101010;
assign LUT_2[63347] = 32'b11111111111111110010110100000011;
assign LUT_2[63348] = 32'b11111111111111101011100000010110;
assign LUT_2[63349] = 32'b11111111111111101000011000101111;
assign LUT_2[63350] = 32'b11111111111111110010011001010010;
assign LUT_2[63351] = 32'b11111111111111101111010001101011;
assign LUT_2[63352] = 32'b11111111111111101001110100001011;
assign LUT_2[63353] = 32'b11111111111111100110101100100100;
assign LUT_2[63354] = 32'b11111111111111110000101101000111;
assign LUT_2[63355] = 32'b11111111111111101101100101100000;
assign LUT_2[63356] = 32'b11111111111111100110010001110011;
assign LUT_2[63357] = 32'b11111111111111100011001010001100;
assign LUT_2[63358] = 32'b11111111111111101101001010101111;
assign LUT_2[63359] = 32'b11111111111111101010000011001000;
assign LUT_2[63360] = 32'b00000000000000000000001110100111;
assign LUT_2[63361] = 32'b11111111111111111101000111000000;
assign LUT_2[63362] = 32'b00000000000000000111000111100011;
assign LUT_2[63363] = 32'b00000000000000000011111111111100;
assign LUT_2[63364] = 32'b11111111111111111100101100001111;
assign LUT_2[63365] = 32'b11111111111111111001100100101000;
assign LUT_2[63366] = 32'b00000000000000000011100101001011;
assign LUT_2[63367] = 32'b00000000000000000000011101100100;
assign LUT_2[63368] = 32'b11111111111111111011000000000100;
assign LUT_2[63369] = 32'b11111111111111110111111000011101;
assign LUT_2[63370] = 32'b00000000000000000001111001000000;
assign LUT_2[63371] = 32'b11111111111111111110110001011001;
assign LUT_2[63372] = 32'b11111111111111110111011101101100;
assign LUT_2[63373] = 32'b11111111111111110100010110000101;
assign LUT_2[63374] = 32'b11111111111111111110010110101000;
assign LUT_2[63375] = 32'b11111111111111111011001111000001;
assign LUT_2[63376] = 32'b11111111111111111010110010110001;
assign LUT_2[63377] = 32'b11111111111111110111101011001010;
assign LUT_2[63378] = 32'b00000000000000000001101011101101;
assign LUT_2[63379] = 32'b11111111111111111110100100000110;
assign LUT_2[63380] = 32'b11111111111111110111010000011001;
assign LUT_2[63381] = 32'b11111111111111110100001000110010;
assign LUT_2[63382] = 32'b11111111111111111110001001010101;
assign LUT_2[63383] = 32'b11111111111111111011000001101110;
assign LUT_2[63384] = 32'b11111111111111110101100100001110;
assign LUT_2[63385] = 32'b11111111111111110010011100100111;
assign LUT_2[63386] = 32'b11111111111111111100011101001010;
assign LUT_2[63387] = 32'b11111111111111111001010101100011;
assign LUT_2[63388] = 32'b11111111111111110010000001110110;
assign LUT_2[63389] = 32'b11111111111111101110111010001111;
assign LUT_2[63390] = 32'b11111111111111111000111010110010;
assign LUT_2[63391] = 32'b11111111111111110101110011001011;
assign LUT_2[63392] = 32'b00000000000000000000101010010000;
assign LUT_2[63393] = 32'b11111111111111111101100010101001;
assign LUT_2[63394] = 32'b00000000000000000111100011001100;
assign LUT_2[63395] = 32'b00000000000000000100011011100101;
assign LUT_2[63396] = 32'b11111111111111111101000111111000;
assign LUT_2[63397] = 32'b11111111111111111010000000010001;
assign LUT_2[63398] = 32'b00000000000000000100000000110100;
assign LUT_2[63399] = 32'b00000000000000000000111001001101;
assign LUT_2[63400] = 32'b11111111111111111011011011101101;
assign LUT_2[63401] = 32'b11111111111111111000010100000110;
assign LUT_2[63402] = 32'b00000000000000000010010100101001;
assign LUT_2[63403] = 32'b11111111111111111111001101000010;
assign LUT_2[63404] = 32'b11111111111111110111111001010101;
assign LUT_2[63405] = 32'b11111111111111110100110001101110;
assign LUT_2[63406] = 32'b11111111111111111110110010010001;
assign LUT_2[63407] = 32'b11111111111111111011101010101010;
assign LUT_2[63408] = 32'b11111111111111111011001110011010;
assign LUT_2[63409] = 32'b11111111111111111000000110110011;
assign LUT_2[63410] = 32'b00000000000000000010000111010110;
assign LUT_2[63411] = 32'b11111111111111111110111111101111;
assign LUT_2[63412] = 32'b11111111111111110111101100000010;
assign LUT_2[63413] = 32'b11111111111111110100100100011011;
assign LUT_2[63414] = 32'b11111111111111111110100100111110;
assign LUT_2[63415] = 32'b11111111111111111011011101010111;
assign LUT_2[63416] = 32'b11111111111111110101111111110111;
assign LUT_2[63417] = 32'b11111111111111110010111000010000;
assign LUT_2[63418] = 32'b11111111111111111100111000110011;
assign LUT_2[63419] = 32'b11111111111111111001110001001100;
assign LUT_2[63420] = 32'b11111111111111110010011101011111;
assign LUT_2[63421] = 32'b11111111111111101111010101111000;
assign LUT_2[63422] = 32'b11111111111111111001010110011011;
assign LUT_2[63423] = 32'b11111111111111110110001110110100;
assign LUT_2[63424] = 32'b11111111111111111000010111001010;
assign LUT_2[63425] = 32'b11111111111111110101001111100011;
assign LUT_2[63426] = 32'b11111111111111111111010000000110;
assign LUT_2[63427] = 32'b11111111111111111100001000011111;
assign LUT_2[63428] = 32'b11111111111111110100110100110010;
assign LUT_2[63429] = 32'b11111111111111110001101101001011;
assign LUT_2[63430] = 32'b11111111111111111011101101101110;
assign LUT_2[63431] = 32'b11111111111111111000100110000111;
assign LUT_2[63432] = 32'b11111111111111110011001000100111;
assign LUT_2[63433] = 32'b11111111111111110000000001000000;
assign LUT_2[63434] = 32'b11111111111111111010000001100011;
assign LUT_2[63435] = 32'b11111111111111110110111001111100;
assign LUT_2[63436] = 32'b11111111111111101111100110001111;
assign LUT_2[63437] = 32'b11111111111111101100011110101000;
assign LUT_2[63438] = 32'b11111111111111110110011111001011;
assign LUT_2[63439] = 32'b11111111111111110011010111100100;
assign LUT_2[63440] = 32'b11111111111111110010111011010100;
assign LUT_2[63441] = 32'b11111111111111101111110011101101;
assign LUT_2[63442] = 32'b11111111111111111001110100010000;
assign LUT_2[63443] = 32'b11111111111111110110101100101001;
assign LUT_2[63444] = 32'b11111111111111101111011000111100;
assign LUT_2[63445] = 32'b11111111111111101100010001010101;
assign LUT_2[63446] = 32'b11111111111111110110010001111000;
assign LUT_2[63447] = 32'b11111111111111110011001010010001;
assign LUT_2[63448] = 32'b11111111111111101101101100110001;
assign LUT_2[63449] = 32'b11111111111111101010100101001010;
assign LUT_2[63450] = 32'b11111111111111110100100101101101;
assign LUT_2[63451] = 32'b11111111111111110001011110000110;
assign LUT_2[63452] = 32'b11111111111111101010001010011001;
assign LUT_2[63453] = 32'b11111111111111100111000010110010;
assign LUT_2[63454] = 32'b11111111111111110001000011010101;
assign LUT_2[63455] = 32'b11111111111111101101111011101110;
assign LUT_2[63456] = 32'b11111111111111111000110010110011;
assign LUT_2[63457] = 32'b11111111111111110101101011001100;
assign LUT_2[63458] = 32'b11111111111111111111101011101111;
assign LUT_2[63459] = 32'b11111111111111111100100100001000;
assign LUT_2[63460] = 32'b11111111111111110101010000011011;
assign LUT_2[63461] = 32'b11111111111111110010001000110100;
assign LUT_2[63462] = 32'b11111111111111111100001001010111;
assign LUT_2[63463] = 32'b11111111111111111001000001110000;
assign LUT_2[63464] = 32'b11111111111111110011100100010000;
assign LUT_2[63465] = 32'b11111111111111110000011100101001;
assign LUT_2[63466] = 32'b11111111111111111010011101001100;
assign LUT_2[63467] = 32'b11111111111111110111010101100101;
assign LUT_2[63468] = 32'b11111111111111110000000001111000;
assign LUT_2[63469] = 32'b11111111111111101100111010010001;
assign LUT_2[63470] = 32'b11111111111111110110111010110100;
assign LUT_2[63471] = 32'b11111111111111110011110011001101;
assign LUT_2[63472] = 32'b11111111111111110011010110111101;
assign LUT_2[63473] = 32'b11111111111111110000001111010110;
assign LUT_2[63474] = 32'b11111111111111111010001111111001;
assign LUT_2[63475] = 32'b11111111111111110111001000010010;
assign LUT_2[63476] = 32'b11111111111111101111110100100101;
assign LUT_2[63477] = 32'b11111111111111101100101100111110;
assign LUT_2[63478] = 32'b11111111111111110110101101100001;
assign LUT_2[63479] = 32'b11111111111111110011100101111010;
assign LUT_2[63480] = 32'b11111111111111101110001000011010;
assign LUT_2[63481] = 32'b11111111111111101011000000110011;
assign LUT_2[63482] = 32'b11111111111111110101000001010110;
assign LUT_2[63483] = 32'b11111111111111110001111001101111;
assign LUT_2[63484] = 32'b11111111111111101010100110000010;
assign LUT_2[63485] = 32'b11111111111111100111011110011011;
assign LUT_2[63486] = 32'b11111111111111110001011110111110;
assign LUT_2[63487] = 32'b11111111111111101110010111010111;
assign LUT_2[63488] = 32'b11111111111111101000010011110111;
assign LUT_2[63489] = 32'b11111111111111100101001100010000;
assign LUT_2[63490] = 32'b11111111111111101111001100110011;
assign LUT_2[63491] = 32'b11111111111111101100000101001100;
assign LUT_2[63492] = 32'b11111111111111100100110001011111;
assign LUT_2[63493] = 32'b11111111111111100001101001111000;
assign LUT_2[63494] = 32'b11111111111111101011101010011011;
assign LUT_2[63495] = 32'b11111111111111101000100010110100;
assign LUT_2[63496] = 32'b11111111111111100011000101010100;
assign LUT_2[63497] = 32'b11111111111111011111111101101101;
assign LUT_2[63498] = 32'b11111111111111101001111110010000;
assign LUT_2[63499] = 32'b11111111111111100110110110101001;
assign LUT_2[63500] = 32'b11111111111111011111100010111100;
assign LUT_2[63501] = 32'b11111111111111011100011011010101;
assign LUT_2[63502] = 32'b11111111111111100110011011111000;
assign LUT_2[63503] = 32'b11111111111111100011010100010001;
assign LUT_2[63504] = 32'b11111111111111100010111000000001;
assign LUT_2[63505] = 32'b11111111111111011111110000011010;
assign LUT_2[63506] = 32'b11111111111111101001110000111101;
assign LUT_2[63507] = 32'b11111111111111100110101001010110;
assign LUT_2[63508] = 32'b11111111111111011111010101101001;
assign LUT_2[63509] = 32'b11111111111111011100001110000010;
assign LUT_2[63510] = 32'b11111111111111100110001110100101;
assign LUT_2[63511] = 32'b11111111111111100011000110111110;
assign LUT_2[63512] = 32'b11111111111111011101101001011110;
assign LUT_2[63513] = 32'b11111111111111011010100001110111;
assign LUT_2[63514] = 32'b11111111111111100100100010011010;
assign LUT_2[63515] = 32'b11111111111111100001011010110011;
assign LUT_2[63516] = 32'b11111111111111011010000111000110;
assign LUT_2[63517] = 32'b11111111111111010110111111011111;
assign LUT_2[63518] = 32'b11111111111111100001000000000010;
assign LUT_2[63519] = 32'b11111111111111011101111000011011;
assign LUT_2[63520] = 32'b11111111111111101000101111100000;
assign LUT_2[63521] = 32'b11111111111111100101100111111001;
assign LUT_2[63522] = 32'b11111111111111101111101000011100;
assign LUT_2[63523] = 32'b11111111111111101100100000110101;
assign LUT_2[63524] = 32'b11111111111111100101001101001000;
assign LUT_2[63525] = 32'b11111111111111100010000101100001;
assign LUT_2[63526] = 32'b11111111111111101100000110000100;
assign LUT_2[63527] = 32'b11111111111111101000111110011101;
assign LUT_2[63528] = 32'b11111111111111100011100000111101;
assign LUT_2[63529] = 32'b11111111111111100000011001010110;
assign LUT_2[63530] = 32'b11111111111111101010011001111001;
assign LUT_2[63531] = 32'b11111111111111100111010010010010;
assign LUT_2[63532] = 32'b11111111111111011111111110100101;
assign LUT_2[63533] = 32'b11111111111111011100110110111110;
assign LUT_2[63534] = 32'b11111111111111100110110111100001;
assign LUT_2[63535] = 32'b11111111111111100011101111111010;
assign LUT_2[63536] = 32'b11111111111111100011010011101010;
assign LUT_2[63537] = 32'b11111111111111100000001100000011;
assign LUT_2[63538] = 32'b11111111111111101010001100100110;
assign LUT_2[63539] = 32'b11111111111111100111000100111111;
assign LUT_2[63540] = 32'b11111111111111011111110001010010;
assign LUT_2[63541] = 32'b11111111111111011100101001101011;
assign LUT_2[63542] = 32'b11111111111111100110101010001110;
assign LUT_2[63543] = 32'b11111111111111100011100010100111;
assign LUT_2[63544] = 32'b11111111111111011110000101000111;
assign LUT_2[63545] = 32'b11111111111111011010111101100000;
assign LUT_2[63546] = 32'b11111111111111100100111110000011;
assign LUT_2[63547] = 32'b11111111111111100001110110011100;
assign LUT_2[63548] = 32'b11111111111111011010100010101111;
assign LUT_2[63549] = 32'b11111111111111010111011011001000;
assign LUT_2[63550] = 32'b11111111111111100001011011101011;
assign LUT_2[63551] = 32'b11111111111111011110010100000100;
assign LUT_2[63552] = 32'b11111111111111100000011100011010;
assign LUT_2[63553] = 32'b11111111111111011101010100110011;
assign LUT_2[63554] = 32'b11111111111111100111010101010110;
assign LUT_2[63555] = 32'b11111111111111100100001101101111;
assign LUT_2[63556] = 32'b11111111111111011100111010000010;
assign LUT_2[63557] = 32'b11111111111111011001110010011011;
assign LUT_2[63558] = 32'b11111111111111100011110010111110;
assign LUT_2[63559] = 32'b11111111111111100000101011010111;
assign LUT_2[63560] = 32'b11111111111111011011001101110111;
assign LUT_2[63561] = 32'b11111111111111011000000110010000;
assign LUT_2[63562] = 32'b11111111111111100010000110110011;
assign LUT_2[63563] = 32'b11111111111111011110111111001100;
assign LUT_2[63564] = 32'b11111111111111010111101011011111;
assign LUT_2[63565] = 32'b11111111111111010100100011111000;
assign LUT_2[63566] = 32'b11111111111111011110100100011011;
assign LUT_2[63567] = 32'b11111111111111011011011100110100;
assign LUT_2[63568] = 32'b11111111111111011011000000100100;
assign LUT_2[63569] = 32'b11111111111111010111111000111101;
assign LUT_2[63570] = 32'b11111111111111100001111001100000;
assign LUT_2[63571] = 32'b11111111111111011110110001111001;
assign LUT_2[63572] = 32'b11111111111111010111011110001100;
assign LUT_2[63573] = 32'b11111111111111010100010110100101;
assign LUT_2[63574] = 32'b11111111111111011110010111001000;
assign LUT_2[63575] = 32'b11111111111111011011001111100001;
assign LUT_2[63576] = 32'b11111111111111010101110010000001;
assign LUT_2[63577] = 32'b11111111111111010010101010011010;
assign LUT_2[63578] = 32'b11111111111111011100101010111101;
assign LUT_2[63579] = 32'b11111111111111011001100011010110;
assign LUT_2[63580] = 32'b11111111111111010010001111101001;
assign LUT_2[63581] = 32'b11111111111111001111001000000010;
assign LUT_2[63582] = 32'b11111111111111011001001000100101;
assign LUT_2[63583] = 32'b11111111111111010110000000111110;
assign LUT_2[63584] = 32'b11111111111111100000111000000011;
assign LUT_2[63585] = 32'b11111111111111011101110000011100;
assign LUT_2[63586] = 32'b11111111111111100111110000111111;
assign LUT_2[63587] = 32'b11111111111111100100101001011000;
assign LUT_2[63588] = 32'b11111111111111011101010101101011;
assign LUT_2[63589] = 32'b11111111111111011010001110000100;
assign LUT_2[63590] = 32'b11111111111111100100001110100111;
assign LUT_2[63591] = 32'b11111111111111100001000111000000;
assign LUT_2[63592] = 32'b11111111111111011011101001100000;
assign LUT_2[63593] = 32'b11111111111111011000100001111001;
assign LUT_2[63594] = 32'b11111111111111100010100010011100;
assign LUT_2[63595] = 32'b11111111111111011111011010110101;
assign LUT_2[63596] = 32'b11111111111111011000000111001000;
assign LUT_2[63597] = 32'b11111111111111010100111111100001;
assign LUT_2[63598] = 32'b11111111111111011111000000000100;
assign LUT_2[63599] = 32'b11111111111111011011111000011101;
assign LUT_2[63600] = 32'b11111111111111011011011100001101;
assign LUT_2[63601] = 32'b11111111111111011000010100100110;
assign LUT_2[63602] = 32'b11111111111111100010010101001001;
assign LUT_2[63603] = 32'b11111111111111011111001101100010;
assign LUT_2[63604] = 32'b11111111111111010111111001110101;
assign LUT_2[63605] = 32'b11111111111111010100110010001110;
assign LUT_2[63606] = 32'b11111111111111011110110010110001;
assign LUT_2[63607] = 32'b11111111111111011011101011001010;
assign LUT_2[63608] = 32'b11111111111111010110001101101010;
assign LUT_2[63609] = 32'b11111111111111010011000110000011;
assign LUT_2[63610] = 32'b11111111111111011101000110100110;
assign LUT_2[63611] = 32'b11111111111111011001111110111111;
assign LUT_2[63612] = 32'b11111111111111010010101011010010;
assign LUT_2[63613] = 32'b11111111111111001111100011101011;
assign LUT_2[63614] = 32'b11111111111111011001100100001110;
assign LUT_2[63615] = 32'b11111111111111010110011100100111;
assign LUT_2[63616] = 32'b11111111111111101100101000000110;
assign LUT_2[63617] = 32'b11111111111111101001100000011111;
assign LUT_2[63618] = 32'b11111111111111110011100001000010;
assign LUT_2[63619] = 32'b11111111111111110000011001011011;
assign LUT_2[63620] = 32'b11111111111111101001000101101110;
assign LUT_2[63621] = 32'b11111111111111100101111110000111;
assign LUT_2[63622] = 32'b11111111111111101111111110101010;
assign LUT_2[63623] = 32'b11111111111111101100110111000011;
assign LUT_2[63624] = 32'b11111111111111100111011001100011;
assign LUT_2[63625] = 32'b11111111111111100100010001111100;
assign LUT_2[63626] = 32'b11111111111111101110010010011111;
assign LUT_2[63627] = 32'b11111111111111101011001010111000;
assign LUT_2[63628] = 32'b11111111111111100011110111001011;
assign LUT_2[63629] = 32'b11111111111111100000101111100100;
assign LUT_2[63630] = 32'b11111111111111101010110000000111;
assign LUT_2[63631] = 32'b11111111111111100111101000100000;
assign LUT_2[63632] = 32'b11111111111111100111001100010000;
assign LUT_2[63633] = 32'b11111111111111100100000100101001;
assign LUT_2[63634] = 32'b11111111111111101110000101001100;
assign LUT_2[63635] = 32'b11111111111111101010111101100101;
assign LUT_2[63636] = 32'b11111111111111100011101001111000;
assign LUT_2[63637] = 32'b11111111111111100000100010010001;
assign LUT_2[63638] = 32'b11111111111111101010100010110100;
assign LUT_2[63639] = 32'b11111111111111100111011011001101;
assign LUT_2[63640] = 32'b11111111111111100001111101101101;
assign LUT_2[63641] = 32'b11111111111111011110110110000110;
assign LUT_2[63642] = 32'b11111111111111101000110110101001;
assign LUT_2[63643] = 32'b11111111111111100101101111000010;
assign LUT_2[63644] = 32'b11111111111111011110011011010101;
assign LUT_2[63645] = 32'b11111111111111011011010011101110;
assign LUT_2[63646] = 32'b11111111111111100101010100010001;
assign LUT_2[63647] = 32'b11111111111111100010001100101010;
assign LUT_2[63648] = 32'b11111111111111101101000011101111;
assign LUT_2[63649] = 32'b11111111111111101001111100001000;
assign LUT_2[63650] = 32'b11111111111111110011111100101011;
assign LUT_2[63651] = 32'b11111111111111110000110101000100;
assign LUT_2[63652] = 32'b11111111111111101001100001010111;
assign LUT_2[63653] = 32'b11111111111111100110011001110000;
assign LUT_2[63654] = 32'b11111111111111110000011010010011;
assign LUT_2[63655] = 32'b11111111111111101101010010101100;
assign LUT_2[63656] = 32'b11111111111111100111110101001100;
assign LUT_2[63657] = 32'b11111111111111100100101101100101;
assign LUT_2[63658] = 32'b11111111111111101110101110001000;
assign LUT_2[63659] = 32'b11111111111111101011100110100001;
assign LUT_2[63660] = 32'b11111111111111100100010010110100;
assign LUT_2[63661] = 32'b11111111111111100001001011001101;
assign LUT_2[63662] = 32'b11111111111111101011001011110000;
assign LUT_2[63663] = 32'b11111111111111101000000100001001;
assign LUT_2[63664] = 32'b11111111111111100111100111111001;
assign LUT_2[63665] = 32'b11111111111111100100100000010010;
assign LUT_2[63666] = 32'b11111111111111101110100000110101;
assign LUT_2[63667] = 32'b11111111111111101011011001001110;
assign LUT_2[63668] = 32'b11111111111111100100000101100001;
assign LUT_2[63669] = 32'b11111111111111100000111101111010;
assign LUT_2[63670] = 32'b11111111111111101010111110011101;
assign LUT_2[63671] = 32'b11111111111111100111110110110110;
assign LUT_2[63672] = 32'b11111111111111100010011001010110;
assign LUT_2[63673] = 32'b11111111111111011111010001101111;
assign LUT_2[63674] = 32'b11111111111111101001010010010010;
assign LUT_2[63675] = 32'b11111111111111100110001010101011;
assign LUT_2[63676] = 32'b11111111111111011110110110111110;
assign LUT_2[63677] = 32'b11111111111111011011101111010111;
assign LUT_2[63678] = 32'b11111111111111100101101111111010;
assign LUT_2[63679] = 32'b11111111111111100010101000010011;
assign LUT_2[63680] = 32'b11111111111111100100110000101001;
assign LUT_2[63681] = 32'b11111111111111100001101001000010;
assign LUT_2[63682] = 32'b11111111111111101011101001100101;
assign LUT_2[63683] = 32'b11111111111111101000100001111110;
assign LUT_2[63684] = 32'b11111111111111100001001110010001;
assign LUT_2[63685] = 32'b11111111111111011110000110101010;
assign LUT_2[63686] = 32'b11111111111111101000000111001101;
assign LUT_2[63687] = 32'b11111111111111100100111111100110;
assign LUT_2[63688] = 32'b11111111111111011111100010000110;
assign LUT_2[63689] = 32'b11111111111111011100011010011111;
assign LUT_2[63690] = 32'b11111111111111100110011011000010;
assign LUT_2[63691] = 32'b11111111111111100011010011011011;
assign LUT_2[63692] = 32'b11111111111111011011111111101110;
assign LUT_2[63693] = 32'b11111111111111011000111000000111;
assign LUT_2[63694] = 32'b11111111111111100010111000101010;
assign LUT_2[63695] = 32'b11111111111111011111110001000011;
assign LUT_2[63696] = 32'b11111111111111011111010100110011;
assign LUT_2[63697] = 32'b11111111111111011100001101001100;
assign LUT_2[63698] = 32'b11111111111111100110001101101111;
assign LUT_2[63699] = 32'b11111111111111100011000110001000;
assign LUT_2[63700] = 32'b11111111111111011011110010011011;
assign LUT_2[63701] = 32'b11111111111111011000101010110100;
assign LUT_2[63702] = 32'b11111111111111100010101011010111;
assign LUT_2[63703] = 32'b11111111111111011111100011110000;
assign LUT_2[63704] = 32'b11111111111111011010000110010000;
assign LUT_2[63705] = 32'b11111111111111010110111110101001;
assign LUT_2[63706] = 32'b11111111111111100000111111001100;
assign LUT_2[63707] = 32'b11111111111111011101110111100101;
assign LUT_2[63708] = 32'b11111111111111010110100011111000;
assign LUT_2[63709] = 32'b11111111111111010011011100010001;
assign LUT_2[63710] = 32'b11111111111111011101011100110100;
assign LUT_2[63711] = 32'b11111111111111011010010101001101;
assign LUT_2[63712] = 32'b11111111111111100101001100010010;
assign LUT_2[63713] = 32'b11111111111111100010000100101011;
assign LUT_2[63714] = 32'b11111111111111101100000101001110;
assign LUT_2[63715] = 32'b11111111111111101000111101100111;
assign LUT_2[63716] = 32'b11111111111111100001101001111010;
assign LUT_2[63717] = 32'b11111111111111011110100010010011;
assign LUT_2[63718] = 32'b11111111111111101000100010110110;
assign LUT_2[63719] = 32'b11111111111111100101011011001111;
assign LUT_2[63720] = 32'b11111111111111011111111101101111;
assign LUT_2[63721] = 32'b11111111111111011100110110001000;
assign LUT_2[63722] = 32'b11111111111111100110110110101011;
assign LUT_2[63723] = 32'b11111111111111100011101111000100;
assign LUT_2[63724] = 32'b11111111111111011100011011010111;
assign LUT_2[63725] = 32'b11111111111111011001010011110000;
assign LUT_2[63726] = 32'b11111111111111100011010100010011;
assign LUT_2[63727] = 32'b11111111111111100000001100101100;
assign LUT_2[63728] = 32'b11111111111111011111110000011100;
assign LUT_2[63729] = 32'b11111111111111011100101000110101;
assign LUT_2[63730] = 32'b11111111111111100110101001011000;
assign LUT_2[63731] = 32'b11111111111111100011100001110001;
assign LUT_2[63732] = 32'b11111111111111011100001110000100;
assign LUT_2[63733] = 32'b11111111111111011001000110011101;
assign LUT_2[63734] = 32'b11111111111111100011000111000000;
assign LUT_2[63735] = 32'b11111111111111011111111111011001;
assign LUT_2[63736] = 32'b11111111111111011010100001111001;
assign LUT_2[63737] = 32'b11111111111111010111011010010010;
assign LUT_2[63738] = 32'b11111111111111100001011010110101;
assign LUT_2[63739] = 32'b11111111111111011110010011001110;
assign LUT_2[63740] = 32'b11111111111111010110111111100001;
assign LUT_2[63741] = 32'b11111111111111010011110111111010;
assign LUT_2[63742] = 32'b11111111111111011101111000011101;
assign LUT_2[63743] = 32'b11111111111111011010110000110110;
assign LUT_2[63744] = 32'b11111111111111101100010010011101;
assign LUT_2[63745] = 32'b11111111111111101001001010110110;
assign LUT_2[63746] = 32'b11111111111111110011001011011001;
assign LUT_2[63747] = 32'b11111111111111110000000011110010;
assign LUT_2[63748] = 32'b11111111111111101000110000000101;
assign LUT_2[63749] = 32'b11111111111111100101101000011110;
assign LUT_2[63750] = 32'b11111111111111101111101001000001;
assign LUT_2[63751] = 32'b11111111111111101100100001011010;
assign LUT_2[63752] = 32'b11111111111111100111000011111010;
assign LUT_2[63753] = 32'b11111111111111100011111100010011;
assign LUT_2[63754] = 32'b11111111111111101101111100110110;
assign LUT_2[63755] = 32'b11111111111111101010110101001111;
assign LUT_2[63756] = 32'b11111111111111100011100001100010;
assign LUT_2[63757] = 32'b11111111111111100000011001111011;
assign LUT_2[63758] = 32'b11111111111111101010011010011110;
assign LUT_2[63759] = 32'b11111111111111100111010010110111;
assign LUT_2[63760] = 32'b11111111111111100110110110100111;
assign LUT_2[63761] = 32'b11111111111111100011101111000000;
assign LUT_2[63762] = 32'b11111111111111101101101111100011;
assign LUT_2[63763] = 32'b11111111111111101010100111111100;
assign LUT_2[63764] = 32'b11111111111111100011010100001111;
assign LUT_2[63765] = 32'b11111111111111100000001100101000;
assign LUT_2[63766] = 32'b11111111111111101010001101001011;
assign LUT_2[63767] = 32'b11111111111111100111000101100100;
assign LUT_2[63768] = 32'b11111111111111100001101000000100;
assign LUT_2[63769] = 32'b11111111111111011110100000011101;
assign LUT_2[63770] = 32'b11111111111111101000100001000000;
assign LUT_2[63771] = 32'b11111111111111100101011001011001;
assign LUT_2[63772] = 32'b11111111111111011110000101101100;
assign LUT_2[63773] = 32'b11111111111111011010111110000101;
assign LUT_2[63774] = 32'b11111111111111100100111110101000;
assign LUT_2[63775] = 32'b11111111111111100001110111000001;
assign LUT_2[63776] = 32'b11111111111111101100101110000110;
assign LUT_2[63777] = 32'b11111111111111101001100110011111;
assign LUT_2[63778] = 32'b11111111111111110011100111000010;
assign LUT_2[63779] = 32'b11111111111111110000011111011011;
assign LUT_2[63780] = 32'b11111111111111101001001011101110;
assign LUT_2[63781] = 32'b11111111111111100110000100000111;
assign LUT_2[63782] = 32'b11111111111111110000000100101010;
assign LUT_2[63783] = 32'b11111111111111101100111101000011;
assign LUT_2[63784] = 32'b11111111111111100111011111100011;
assign LUT_2[63785] = 32'b11111111111111100100010111111100;
assign LUT_2[63786] = 32'b11111111111111101110011000011111;
assign LUT_2[63787] = 32'b11111111111111101011010000111000;
assign LUT_2[63788] = 32'b11111111111111100011111101001011;
assign LUT_2[63789] = 32'b11111111111111100000110101100100;
assign LUT_2[63790] = 32'b11111111111111101010110110000111;
assign LUT_2[63791] = 32'b11111111111111100111101110100000;
assign LUT_2[63792] = 32'b11111111111111100111010010010000;
assign LUT_2[63793] = 32'b11111111111111100100001010101001;
assign LUT_2[63794] = 32'b11111111111111101110001011001100;
assign LUT_2[63795] = 32'b11111111111111101011000011100101;
assign LUT_2[63796] = 32'b11111111111111100011101111111000;
assign LUT_2[63797] = 32'b11111111111111100000101000010001;
assign LUT_2[63798] = 32'b11111111111111101010101000110100;
assign LUT_2[63799] = 32'b11111111111111100111100001001101;
assign LUT_2[63800] = 32'b11111111111111100010000011101101;
assign LUT_2[63801] = 32'b11111111111111011110111100000110;
assign LUT_2[63802] = 32'b11111111111111101000111100101001;
assign LUT_2[63803] = 32'b11111111111111100101110101000010;
assign LUT_2[63804] = 32'b11111111111111011110100001010101;
assign LUT_2[63805] = 32'b11111111111111011011011001101110;
assign LUT_2[63806] = 32'b11111111111111100101011010010001;
assign LUT_2[63807] = 32'b11111111111111100010010010101010;
assign LUT_2[63808] = 32'b11111111111111100100011011000000;
assign LUT_2[63809] = 32'b11111111111111100001010011011001;
assign LUT_2[63810] = 32'b11111111111111101011010011111100;
assign LUT_2[63811] = 32'b11111111111111101000001100010101;
assign LUT_2[63812] = 32'b11111111111111100000111000101000;
assign LUT_2[63813] = 32'b11111111111111011101110001000001;
assign LUT_2[63814] = 32'b11111111111111100111110001100100;
assign LUT_2[63815] = 32'b11111111111111100100101001111101;
assign LUT_2[63816] = 32'b11111111111111011111001100011101;
assign LUT_2[63817] = 32'b11111111111111011100000100110110;
assign LUT_2[63818] = 32'b11111111111111100110000101011001;
assign LUT_2[63819] = 32'b11111111111111100010111101110010;
assign LUT_2[63820] = 32'b11111111111111011011101010000101;
assign LUT_2[63821] = 32'b11111111111111011000100010011110;
assign LUT_2[63822] = 32'b11111111111111100010100011000001;
assign LUT_2[63823] = 32'b11111111111111011111011011011010;
assign LUT_2[63824] = 32'b11111111111111011110111111001010;
assign LUT_2[63825] = 32'b11111111111111011011110111100011;
assign LUT_2[63826] = 32'b11111111111111100101111000000110;
assign LUT_2[63827] = 32'b11111111111111100010110000011111;
assign LUT_2[63828] = 32'b11111111111111011011011100110010;
assign LUT_2[63829] = 32'b11111111111111011000010101001011;
assign LUT_2[63830] = 32'b11111111111111100010010101101110;
assign LUT_2[63831] = 32'b11111111111111011111001110000111;
assign LUT_2[63832] = 32'b11111111111111011001110000100111;
assign LUT_2[63833] = 32'b11111111111111010110101001000000;
assign LUT_2[63834] = 32'b11111111111111100000101001100011;
assign LUT_2[63835] = 32'b11111111111111011101100001111100;
assign LUT_2[63836] = 32'b11111111111111010110001110001111;
assign LUT_2[63837] = 32'b11111111111111010011000110101000;
assign LUT_2[63838] = 32'b11111111111111011101000111001011;
assign LUT_2[63839] = 32'b11111111111111011001111111100100;
assign LUT_2[63840] = 32'b11111111111111100100110110101001;
assign LUT_2[63841] = 32'b11111111111111100001101111000010;
assign LUT_2[63842] = 32'b11111111111111101011101111100101;
assign LUT_2[63843] = 32'b11111111111111101000100111111110;
assign LUT_2[63844] = 32'b11111111111111100001010100010001;
assign LUT_2[63845] = 32'b11111111111111011110001100101010;
assign LUT_2[63846] = 32'b11111111111111101000001101001101;
assign LUT_2[63847] = 32'b11111111111111100101000101100110;
assign LUT_2[63848] = 32'b11111111111111011111101000000110;
assign LUT_2[63849] = 32'b11111111111111011100100000011111;
assign LUT_2[63850] = 32'b11111111111111100110100001000010;
assign LUT_2[63851] = 32'b11111111111111100011011001011011;
assign LUT_2[63852] = 32'b11111111111111011100000101101110;
assign LUT_2[63853] = 32'b11111111111111011000111110000111;
assign LUT_2[63854] = 32'b11111111111111100010111110101010;
assign LUT_2[63855] = 32'b11111111111111011111110111000011;
assign LUT_2[63856] = 32'b11111111111111011111011010110011;
assign LUT_2[63857] = 32'b11111111111111011100010011001100;
assign LUT_2[63858] = 32'b11111111111111100110010011101111;
assign LUT_2[63859] = 32'b11111111111111100011001100001000;
assign LUT_2[63860] = 32'b11111111111111011011111000011011;
assign LUT_2[63861] = 32'b11111111111111011000110000110100;
assign LUT_2[63862] = 32'b11111111111111100010110001010111;
assign LUT_2[63863] = 32'b11111111111111011111101001110000;
assign LUT_2[63864] = 32'b11111111111111011010001100010000;
assign LUT_2[63865] = 32'b11111111111111010111000100101001;
assign LUT_2[63866] = 32'b11111111111111100001000101001100;
assign LUT_2[63867] = 32'b11111111111111011101111101100101;
assign LUT_2[63868] = 32'b11111111111111010110101001111000;
assign LUT_2[63869] = 32'b11111111111111010011100010010001;
assign LUT_2[63870] = 32'b11111111111111011101100010110100;
assign LUT_2[63871] = 32'b11111111111111011010011011001101;
assign LUT_2[63872] = 32'b11111111111111110000100110101100;
assign LUT_2[63873] = 32'b11111111111111101101011111000101;
assign LUT_2[63874] = 32'b11111111111111110111011111101000;
assign LUT_2[63875] = 32'b11111111111111110100011000000001;
assign LUT_2[63876] = 32'b11111111111111101101000100010100;
assign LUT_2[63877] = 32'b11111111111111101001111100101101;
assign LUT_2[63878] = 32'b11111111111111110011111101010000;
assign LUT_2[63879] = 32'b11111111111111110000110101101001;
assign LUT_2[63880] = 32'b11111111111111101011011000001001;
assign LUT_2[63881] = 32'b11111111111111101000010000100010;
assign LUT_2[63882] = 32'b11111111111111110010010001000101;
assign LUT_2[63883] = 32'b11111111111111101111001001011110;
assign LUT_2[63884] = 32'b11111111111111100111110101110001;
assign LUT_2[63885] = 32'b11111111111111100100101110001010;
assign LUT_2[63886] = 32'b11111111111111101110101110101101;
assign LUT_2[63887] = 32'b11111111111111101011100111000110;
assign LUT_2[63888] = 32'b11111111111111101011001010110110;
assign LUT_2[63889] = 32'b11111111111111101000000011001111;
assign LUT_2[63890] = 32'b11111111111111110010000011110010;
assign LUT_2[63891] = 32'b11111111111111101110111100001011;
assign LUT_2[63892] = 32'b11111111111111100111101000011110;
assign LUT_2[63893] = 32'b11111111111111100100100000110111;
assign LUT_2[63894] = 32'b11111111111111101110100001011010;
assign LUT_2[63895] = 32'b11111111111111101011011001110011;
assign LUT_2[63896] = 32'b11111111111111100101111100010011;
assign LUT_2[63897] = 32'b11111111111111100010110100101100;
assign LUT_2[63898] = 32'b11111111111111101100110101001111;
assign LUT_2[63899] = 32'b11111111111111101001101101101000;
assign LUT_2[63900] = 32'b11111111111111100010011001111011;
assign LUT_2[63901] = 32'b11111111111111011111010010010100;
assign LUT_2[63902] = 32'b11111111111111101001010010110111;
assign LUT_2[63903] = 32'b11111111111111100110001011010000;
assign LUT_2[63904] = 32'b11111111111111110001000010010101;
assign LUT_2[63905] = 32'b11111111111111101101111010101110;
assign LUT_2[63906] = 32'b11111111111111110111111011010001;
assign LUT_2[63907] = 32'b11111111111111110100110011101010;
assign LUT_2[63908] = 32'b11111111111111101101011111111101;
assign LUT_2[63909] = 32'b11111111111111101010011000010110;
assign LUT_2[63910] = 32'b11111111111111110100011000111001;
assign LUT_2[63911] = 32'b11111111111111110001010001010010;
assign LUT_2[63912] = 32'b11111111111111101011110011110010;
assign LUT_2[63913] = 32'b11111111111111101000101100001011;
assign LUT_2[63914] = 32'b11111111111111110010101100101110;
assign LUT_2[63915] = 32'b11111111111111101111100101000111;
assign LUT_2[63916] = 32'b11111111111111101000010001011010;
assign LUT_2[63917] = 32'b11111111111111100101001001110011;
assign LUT_2[63918] = 32'b11111111111111101111001010010110;
assign LUT_2[63919] = 32'b11111111111111101100000010101111;
assign LUT_2[63920] = 32'b11111111111111101011100110011111;
assign LUT_2[63921] = 32'b11111111111111101000011110111000;
assign LUT_2[63922] = 32'b11111111111111110010011111011011;
assign LUT_2[63923] = 32'b11111111111111101111010111110100;
assign LUT_2[63924] = 32'b11111111111111101000000100000111;
assign LUT_2[63925] = 32'b11111111111111100100111100100000;
assign LUT_2[63926] = 32'b11111111111111101110111101000011;
assign LUT_2[63927] = 32'b11111111111111101011110101011100;
assign LUT_2[63928] = 32'b11111111111111100110010111111100;
assign LUT_2[63929] = 32'b11111111111111100011010000010101;
assign LUT_2[63930] = 32'b11111111111111101101010000111000;
assign LUT_2[63931] = 32'b11111111111111101010001001010001;
assign LUT_2[63932] = 32'b11111111111111100010110101100100;
assign LUT_2[63933] = 32'b11111111111111011111101101111101;
assign LUT_2[63934] = 32'b11111111111111101001101110100000;
assign LUT_2[63935] = 32'b11111111111111100110100110111001;
assign LUT_2[63936] = 32'b11111111111111101000101111001111;
assign LUT_2[63937] = 32'b11111111111111100101100111101000;
assign LUT_2[63938] = 32'b11111111111111101111101000001011;
assign LUT_2[63939] = 32'b11111111111111101100100000100100;
assign LUT_2[63940] = 32'b11111111111111100101001100110111;
assign LUT_2[63941] = 32'b11111111111111100010000101010000;
assign LUT_2[63942] = 32'b11111111111111101100000101110011;
assign LUT_2[63943] = 32'b11111111111111101000111110001100;
assign LUT_2[63944] = 32'b11111111111111100011100000101100;
assign LUT_2[63945] = 32'b11111111111111100000011001000101;
assign LUT_2[63946] = 32'b11111111111111101010011001101000;
assign LUT_2[63947] = 32'b11111111111111100111010010000001;
assign LUT_2[63948] = 32'b11111111111111011111111110010100;
assign LUT_2[63949] = 32'b11111111111111011100110110101101;
assign LUT_2[63950] = 32'b11111111111111100110110111010000;
assign LUT_2[63951] = 32'b11111111111111100011101111101001;
assign LUT_2[63952] = 32'b11111111111111100011010011011001;
assign LUT_2[63953] = 32'b11111111111111100000001011110010;
assign LUT_2[63954] = 32'b11111111111111101010001100010101;
assign LUT_2[63955] = 32'b11111111111111100111000100101110;
assign LUT_2[63956] = 32'b11111111111111011111110001000001;
assign LUT_2[63957] = 32'b11111111111111011100101001011010;
assign LUT_2[63958] = 32'b11111111111111100110101001111101;
assign LUT_2[63959] = 32'b11111111111111100011100010010110;
assign LUT_2[63960] = 32'b11111111111111011110000100110110;
assign LUT_2[63961] = 32'b11111111111111011010111101001111;
assign LUT_2[63962] = 32'b11111111111111100100111101110010;
assign LUT_2[63963] = 32'b11111111111111100001110110001011;
assign LUT_2[63964] = 32'b11111111111111011010100010011110;
assign LUT_2[63965] = 32'b11111111111111010111011010110111;
assign LUT_2[63966] = 32'b11111111111111100001011011011010;
assign LUT_2[63967] = 32'b11111111111111011110010011110011;
assign LUT_2[63968] = 32'b11111111111111101001001010111000;
assign LUT_2[63969] = 32'b11111111111111100110000011010001;
assign LUT_2[63970] = 32'b11111111111111110000000011110100;
assign LUT_2[63971] = 32'b11111111111111101100111100001101;
assign LUT_2[63972] = 32'b11111111111111100101101000100000;
assign LUT_2[63973] = 32'b11111111111111100010100000111001;
assign LUT_2[63974] = 32'b11111111111111101100100001011100;
assign LUT_2[63975] = 32'b11111111111111101001011001110101;
assign LUT_2[63976] = 32'b11111111111111100011111100010101;
assign LUT_2[63977] = 32'b11111111111111100000110100101110;
assign LUT_2[63978] = 32'b11111111111111101010110101010001;
assign LUT_2[63979] = 32'b11111111111111100111101101101010;
assign LUT_2[63980] = 32'b11111111111111100000011001111101;
assign LUT_2[63981] = 32'b11111111111111011101010010010110;
assign LUT_2[63982] = 32'b11111111111111100111010010111001;
assign LUT_2[63983] = 32'b11111111111111100100001011010010;
assign LUT_2[63984] = 32'b11111111111111100011101111000010;
assign LUT_2[63985] = 32'b11111111111111100000100111011011;
assign LUT_2[63986] = 32'b11111111111111101010100111111110;
assign LUT_2[63987] = 32'b11111111111111100111100000010111;
assign LUT_2[63988] = 32'b11111111111111100000001100101010;
assign LUT_2[63989] = 32'b11111111111111011101000101000011;
assign LUT_2[63990] = 32'b11111111111111100111000101100110;
assign LUT_2[63991] = 32'b11111111111111100011111101111111;
assign LUT_2[63992] = 32'b11111111111111011110100000011111;
assign LUT_2[63993] = 32'b11111111111111011011011000111000;
assign LUT_2[63994] = 32'b11111111111111100101011001011011;
assign LUT_2[63995] = 32'b11111111111111100010010001110100;
assign LUT_2[63996] = 32'b11111111111111011010111110000111;
assign LUT_2[63997] = 32'b11111111111111010111110110100000;
assign LUT_2[63998] = 32'b11111111111111100001110111000011;
assign LUT_2[63999] = 32'b11111111111111011110101111011100;
assign LUT_2[64000] = 32'b11111111111111101101000101101001;
assign LUT_2[64001] = 32'b11111111111111101001111110000010;
assign LUT_2[64002] = 32'b11111111111111110011111110100101;
assign LUT_2[64003] = 32'b11111111111111110000110110111110;
assign LUT_2[64004] = 32'b11111111111111101001100011010001;
assign LUT_2[64005] = 32'b11111111111111100110011011101010;
assign LUT_2[64006] = 32'b11111111111111110000011100001101;
assign LUT_2[64007] = 32'b11111111111111101101010100100110;
assign LUT_2[64008] = 32'b11111111111111100111110111000110;
assign LUT_2[64009] = 32'b11111111111111100100101111011111;
assign LUT_2[64010] = 32'b11111111111111101110110000000010;
assign LUT_2[64011] = 32'b11111111111111101011101000011011;
assign LUT_2[64012] = 32'b11111111111111100100010100101110;
assign LUT_2[64013] = 32'b11111111111111100001001101000111;
assign LUT_2[64014] = 32'b11111111111111101011001101101010;
assign LUT_2[64015] = 32'b11111111111111101000000110000011;
assign LUT_2[64016] = 32'b11111111111111100111101001110011;
assign LUT_2[64017] = 32'b11111111111111100100100010001100;
assign LUT_2[64018] = 32'b11111111111111101110100010101111;
assign LUT_2[64019] = 32'b11111111111111101011011011001000;
assign LUT_2[64020] = 32'b11111111111111100100000111011011;
assign LUT_2[64021] = 32'b11111111111111100000111111110100;
assign LUT_2[64022] = 32'b11111111111111101011000000010111;
assign LUT_2[64023] = 32'b11111111111111100111111000110000;
assign LUT_2[64024] = 32'b11111111111111100010011011010000;
assign LUT_2[64025] = 32'b11111111111111011111010011101001;
assign LUT_2[64026] = 32'b11111111111111101001010100001100;
assign LUT_2[64027] = 32'b11111111111111100110001100100101;
assign LUT_2[64028] = 32'b11111111111111011110111000111000;
assign LUT_2[64029] = 32'b11111111111111011011110001010001;
assign LUT_2[64030] = 32'b11111111111111100101110001110100;
assign LUT_2[64031] = 32'b11111111111111100010101010001101;
assign LUT_2[64032] = 32'b11111111111111101101100001010010;
assign LUT_2[64033] = 32'b11111111111111101010011001101011;
assign LUT_2[64034] = 32'b11111111111111110100011010001110;
assign LUT_2[64035] = 32'b11111111111111110001010010100111;
assign LUT_2[64036] = 32'b11111111111111101001111110111010;
assign LUT_2[64037] = 32'b11111111111111100110110111010011;
assign LUT_2[64038] = 32'b11111111111111110000110111110110;
assign LUT_2[64039] = 32'b11111111111111101101110000001111;
assign LUT_2[64040] = 32'b11111111111111101000010010101111;
assign LUT_2[64041] = 32'b11111111111111100101001011001000;
assign LUT_2[64042] = 32'b11111111111111101111001011101011;
assign LUT_2[64043] = 32'b11111111111111101100000100000100;
assign LUT_2[64044] = 32'b11111111111111100100110000010111;
assign LUT_2[64045] = 32'b11111111111111100001101000110000;
assign LUT_2[64046] = 32'b11111111111111101011101001010011;
assign LUT_2[64047] = 32'b11111111111111101000100001101100;
assign LUT_2[64048] = 32'b11111111111111101000000101011100;
assign LUT_2[64049] = 32'b11111111111111100100111101110101;
assign LUT_2[64050] = 32'b11111111111111101110111110011000;
assign LUT_2[64051] = 32'b11111111111111101011110110110001;
assign LUT_2[64052] = 32'b11111111111111100100100011000100;
assign LUT_2[64053] = 32'b11111111111111100001011011011101;
assign LUT_2[64054] = 32'b11111111111111101011011100000000;
assign LUT_2[64055] = 32'b11111111111111101000010100011001;
assign LUT_2[64056] = 32'b11111111111111100010110110111001;
assign LUT_2[64057] = 32'b11111111111111011111101111010010;
assign LUT_2[64058] = 32'b11111111111111101001101111110101;
assign LUT_2[64059] = 32'b11111111111111100110101000001110;
assign LUT_2[64060] = 32'b11111111111111011111010100100001;
assign LUT_2[64061] = 32'b11111111111111011100001100111010;
assign LUT_2[64062] = 32'b11111111111111100110001101011101;
assign LUT_2[64063] = 32'b11111111111111100011000101110110;
assign LUT_2[64064] = 32'b11111111111111100101001110001100;
assign LUT_2[64065] = 32'b11111111111111100010000110100101;
assign LUT_2[64066] = 32'b11111111111111101100000111001000;
assign LUT_2[64067] = 32'b11111111111111101000111111100001;
assign LUT_2[64068] = 32'b11111111111111100001101011110100;
assign LUT_2[64069] = 32'b11111111111111011110100100001101;
assign LUT_2[64070] = 32'b11111111111111101000100100110000;
assign LUT_2[64071] = 32'b11111111111111100101011101001001;
assign LUT_2[64072] = 32'b11111111111111011111111111101001;
assign LUT_2[64073] = 32'b11111111111111011100111000000010;
assign LUT_2[64074] = 32'b11111111111111100110111000100101;
assign LUT_2[64075] = 32'b11111111111111100011110000111110;
assign LUT_2[64076] = 32'b11111111111111011100011101010001;
assign LUT_2[64077] = 32'b11111111111111011001010101101010;
assign LUT_2[64078] = 32'b11111111111111100011010110001101;
assign LUT_2[64079] = 32'b11111111111111100000001110100110;
assign LUT_2[64080] = 32'b11111111111111011111110010010110;
assign LUT_2[64081] = 32'b11111111111111011100101010101111;
assign LUT_2[64082] = 32'b11111111111111100110101011010010;
assign LUT_2[64083] = 32'b11111111111111100011100011101011;
assign LUT_2[64084] = 32'b11111111111111011100001111111110;
assign LUT_2[64085] = 32'b11111111111111011001001000010111;
assign LUT_2[64086] = 32'b11111111111111100011001000111010;
assign LUT_2[64087] = 32'b11111111111111100000000001010011;
assign LUT_2[64088] = 32'b11111111111111011010100011110011;
assign LUT_2[64089] = 32'b11111111111111010111011100001100;
assign LUT_2[64090] = 32'b11111111111111100001011100101111;
assign LUT_2[64091] = 32'b11111111111111011110010101001000;
assign LUT_2[64092] = 32'b11111111111111010111000001011011;
assign LUT_2[64093] = 32'b11111111111111010011111001110100;
assign LUT_2[64094] = 32'b11111111111111011101111010010111;
assign LUT_2[64095] = 32'b11111111111111011010110010110000;
assign LUT_2[64096] = 32'b11111111111111100101101001110101;
assign LUT_2[64097] = 32'b11111111111111100010100010001110;
assign LUT_2[64098] = 32'b11111111111111101100100010110001;
assign LUT_2[64099] = 32'b11111111111111101001011011001010;
assign LUT_2[64100] = 32'b11111111111111100010000111011101;
assign LUT_2[64101] = 32'b11111111111111011110111111110110;
assign LUT_2[64102] = 32'b11111111111111101001000000011001;
assign LUT_2[64103] = 32'b11111111111111100101111000110010;
assign LUT_2[64104] = 32'b11111111111111100000011011010010;
assign LUT_2[64105] = 32'b11111111111111011101010011101011;
assign LUT_2[64106] = 32'b11111111111111100111010100001110;
assign LUT_2[64107] = 32'b11111111111111100100001100100111;
assign LUT_2[64108] = 32'b11111111111111011100111000111010;
assign LUT_2[64109] = 32'b11111111111111011001110001010011;
assign LUT_2[64110] = 32'b11111111111111100011110001110110;
assign LUT_2[64111] = 32'b11111111111111100000101010001111;
assign LUT_2[64112] = 32'b11111111111111100000001101111111;
assign LUT_2[64113] = 32'b11111111111111011101000110011000;
assign LUT_2[64114] = 32'b11111111111111100111000110111011;
assign LUT_2[64115] = 32'b11111111111111100011111111010100;
assign LUT_2[64116] = 32'b11111111111111011100101011100111;
assign LUT_2[64117] = 32'b11111111111111011001100100000000;
assign LUT_2[64118] = 32'b11111111111111100011100100100011;
assign LUT_2[64119] = 32'b11111111111111100000011100111100;
assign LUT_2[64120] = 32'b11111111111111011010111111011100;
assign LUT_2[64121] = 32'b11111111111111010111110111110101;
assign LUT_2[64122] = 32'b11111111111111100001111000011000;
assign LUT_2[64123] = 32'b11111111111111011110110000110001;
assign LUT_2[64124] = 32'b11111111111111010111011101000100;
assign LUT_2[64125] = 32'b11111111111111010100010101011101;
assign LUT_2[64126] = 32'b11111111111111011110010110000000;
assign LUT_2[64127] = 32'b11111111111111011011001110011001;
assign LUT_2[64128] = 32'b11111111111111110001011001111000;
assign LUT_2[64129] = 32'b11111111111111101110010010010001;
assign LUT_2[64130] = 32'b11111111111111111000010010110100;
assign LUT_2[64131] = 32'b11111111111111110101001011001101;
assign LUT_2[64132] = 32'b11111111111111101101110111100000;
assign LUT_2[64133] = 32'b11111111111111101010101111111001;
assign LUT_2[64134] = 32'b11111111111111110100110000011100;
assign LUT_2[64135] = 32'b11111111111111110001101000110101;
assign LUT_2[64136] = 32'b11111111111111101100001011010101;
assign LUT_2[64137] = 32'b11111111111111101001000011101110;
assign LUT_2[64138] = 32'b11111111111111110011000100010001;
assign LUT_2[64139] = 32'b11111111111111101111111100101010;
assign LUT_2[64140] = 32'b11111111111111101000101000111101;
assign LUT_2[64141] = 32'b11111111111111100101100001010110;
assign LUT_2[64142] = 32'b11111111111111101111100001111001;
assign LUT_2[64143] = 32'b11111111111111101100011010010010;
assign LUT_2[64144] = 32'b11111111111111101011111110000010;
assign LUT_2[64145] = 32'b11111111111111101000110110011011;
assign LUT_2[64146] = 32'b11111111111111110010110110111110;
assign LUT_2[64147] = 32'b11111111111111101111101111010111;
assign LUT_2[64148] = 32'b11111111111111101000011011101010;
assign LUT_2[64149] = 32'b11111111111111100101010100000011;
assign LUT_2[64150] = 32'b11111111111111101111010100100110;
assign LUT_2[64151] = 32'b11111111111111101100001100111111;
assign LUT_2[64152] = 32'b11111111111111100110101111011111;
assign LUT_2[64153] = 32'b11111111111111100011100111111000;
assign LUT_2[64154] = 32'b11111111111111101101101000011011;
assign LUT_2[64155] = 32'b11111111111111101010100000110100;
assign LUT_2[64156] = 32'b11111111111111100011001101000111;
assign LUT_2[64157] = 32'b11111111111111100000000101100000;
assign LUT_2[64158] = 32'b11111111111111101010000110000011;
assign LUT_2[64159] = 32'b11111111111111100110111110011100;
assign LUT_2[64160] = 32'b11111111111111110001110101100001;
assign LUT_2[64161] = 32'b11111111111111101110101101111010;
assign LUT_2[64162] = 32'b11111111111111111000101110011101;
assign LUT_2[64163] = 32'b11111111111111110101100110110110;
assign LUT_2[64164] = 32'b11111111111111101110010011001001;
assign LUT_2[64165] = 32'b11111111111111101011001011100010;
assign LUT_2[64166] = 32'b11111111111111110101001100000101;
assign LUT_2[64167] = 32'b11111111111111110010000100011110;
assign LUT_2[64168] = 32'b11111111111111101100100110111110;
assign LUT_2[64169] = 32'b11111111111111101001011111010111;
assign LUT_2[64170] = 32'b11111111111111110011011111111010;
assign LUT_2[64171] = 32'b11111111111111110000011000010011;
assign LUT_2[64172] = 32'b11111111111111101001000100100110;
assign LUT_2[64173] = 32'b11111111111111100101111100111111;
assign LUT_2[64174] = 32'b11111111111111101111111101100010;
assign LUT_2[64175] = 32'b11111111111111101100110101111011;
assign LUT_2[64176] = 32'b11111111111111101100011001101011;
assign LUT_2[64177] = 32'b11111111111111101001010010000100;
assign LUT_2[64178] = 32'b11111111111111110011010010100111;
assign LUT_2[64179] = 32'b11111111111111110000001011000000;
assign LUT_2[64180] = 32'b11111111111111101000110111010011;
assign LUT_2[64181] = 32'b11111111111111100101101111101100;
assign LUT_2[64182] = 32'b11111111111111101111110000001111;
assign LUT_2[64183] = 32'b11111111111111101100101000101000;
assign LUT_2[64184] = 32'b11111111111111100111001011001000;
assign LUT_2[64185] = 32'b11111111111111100100000011100001;
assign LUT_2[64186] = 32'b11111111111111101110000100000100;
assign LUT_2[64187] = 32'b11111111111111101010111100011101;
assign LUT_2[64188] = 32'b11111111111111100011101000110000;
assign LUT_2[64189] = 32'b11111111111111100000100001001001;
assign LUT_2[64190] = 32'b11111111111111101010100001101100;
assign LUT_2[64191] = 32'b11111111111111100111011010000101;
assign LUT_2[64192] = 32'b11111111111111101001100010011011;
assign LUT_2[64193] = 32'b11111111111111100110011010110100;
assign LUT_2[64194] = 32'b11111111111111110000011011010111;
assign LUT_2[64195] = 32'b11111111111111101101010011110000;
assign LUT_2[64196] = 32'b11111111111111100110000000000011;
assign LUT_2[64197] = 32'b11111111111111100010111000011100;
assign LUT_2[64198] = 32'b11111111111111101100111000111111;
assign LUT_2[64199] = 32'b11111111111111101001110001011000;
assign LUT_2[64200] = 32'b11111111111111100100010011111000;
assign LUT_2[64201] = 32'b11111111111111100001001100010001;
assign LUT_2[64202] = 32'b11111111111111101011001100110100;
assign LUT_2[64203] = 32'b11111111111111101000000101001101;
assign LUT_2[64204] = 32'b11111111111111100000110001100000;
assign LUT_2[64205] = 32'b11111111111111011101101001111001;
assign LUT_2[64206] = 32'b11111111111111100111101010011100;
assign LUT_2[64207] = 32'b11111111111111100100100010110101;
assign LUT_2[64208] = 32'b11111111111111100100000110100101;
assign LUT_2[64209] = 32'b11111111111111100000111110111110;
assign LUT_2[64210] = 32'b11111111111111101010111111100001;
assign LUT_2[64211] = 32'b11111111111111100111110111111010;
assign LUT_2[64212] = 32'b11111111111111100000100100001101;
assign LUT_2[64213] = 32'b11111111111111011101011100100110;
assign LUT_2[64214] = 32'b11111111111111100111011101001001;
assign LUT_2[64215] = 32'b11111111111111100100010101100010;
assign LUT_2[64216] = 32'b11111111111111011110111000000010;
assign LUT_2[64217] = 32'b11111111111111011011110000011011;
assign LUT_2[64218] = 32'b11111111111111100101110000111110;
assign LUT_2[64219] = 32'b11111111111111100010101001010111;
assign LUT_2[64220] = 32'b11111111111111011011010101101010;
assign LUT_2[64221] = 32'b11111111111111011000001110000011;
assign LUT_2[64222] = 32'b11111111111111100010001110100110;
assign LUT_2[64223] = 32'b11111111111111011111000110111111;
assign LUT_2[64224] = 32'b11111111111111101001111110000100;
assign LUT_2[64225] = 32'b11111111111111100110110110011101;
assign LUT_2[64226] = 32'b11111111111111110000110111000000;
assign LUT_2[64227] = 32'b11111111111111101101101111011001;
assign LUT_2[64228] = 32'b11111111111111100110011011101100;
assign LUT_2[64229] = 32'b11111111111111100011010100000101;
assign LUT_2[64230] = 32'b11111111111111101101010100101000;
assign LUT_2[64231] = 32'b11111111111111101010001101000001;
assign LUT_2[64232] = 32'b11111111111111100100101111100001;
assign LUT_2[64233] = 32'b11111111111111100001100111111010;
assign LUT_2[64234] = 32'b11111111111111101011101000011101;
assign LUT_2[64235] = 32'b11111111111111101000100000110110;
assign LUT_2[64236] = 32'b11111111111111100001001101001001;
assign LUT_2[64237] = 32'b11111111111111011110000101100010;
assign LUT_2[64238] = 32'b11111111111111101000000110000101;
assign LUT_2[64239] = 32'b11111111111111100100111110011110;
assign LUT_2[64240] = 32'b11111111111111100100100010001110;
assign LUT_2[64241] = 32'b11111111111111100001011010100111;
assign LUT_2[64242] = 32'b11111111111111101011011011001010;
assign LUT_2[64243] = 32'b11111111111111101000010011100011;
assign LUT_2[64244] = 32'b11111111111111100000111111110110;
assign LUT_2[64245] = 32'b11111111111111011101111000001111;
assign LUT_2[64246] = 32'b11111111111111100111111000110010;
assign LUT_2[64247] = 32'b11111111111111100100110001001011;
assign LUT_2[64248] = 32'b11111111111111011111010011101011;
assign LUT_2[64249] = 32'b11111111111111011100001100000100;
assign LUT_2[64250] = 32'b11111111111111100110001100100111;
assign LUT_2[64251] = 32'b11111111111111100011000101000000;
assign LUT_2[64252] = 32'b11111111111111011011110001010011;
assign LUT_2[64253] = 32'b11111111111111011000101001101100;
assign LUT_2[64254] = 32'b11111111111111100010101010001111;
assign LUT_2[64255] = 32'b11111111111111011111100010101000;
assign LUT_2[64256] = 32'b11111111111111110001000100001111;
assign LUT_2[64257] = 32'b11111111111111101101111100101000;
assign LUT_2[64258] = 32'b11111111111111110111111101001011;
assign LUT_2[64259] = 32'b11111111111111110100110101100100;
assign LUT_2[64260] = 32'b11111111111111101101100001110111;
assign LUT_2[64261] = 32'b11111111111111101010011010010000;
assign LUT_2[64262] = 32'b11111111111111110100011010110011;
assign LUT_2[64263] = 32'b11111111111111110001010011001100;
assign LUT_2[64264] = 32'b11111111111111101011110101101100;
assign LUT_2[64265] = 32'b11111111111111101000101110000101;
assign LUT_2[64266] = 32'b11111111111111110010101110101000;
assign LUT_2[64267] = 32'b11111111111111101111100111000001;
assign LUT_2[64268] = 32'b11111111111111101000010011010100;
assign LUT_2[64269] = 32'b11111111111111100101001011101101;
assign LUT_2[64270] = 32'b11111111111111101111001100010000;
assign LUT_2[64271] = 32'b11111111111111101100000100101001;
assign LUT_2[64272] = 32'b11111111111111101011101000011001;
assign LUT_2[64273] = 32'b11111111111111101000100000110010;
assign LUT_2[64274] = 32'b11111111111111110010100001010101;
assign LUT_2[64275] = 32'b11111111111111101111011001101110;
assign LUT_2[64276] = 32'b11111111111111101000000110000001;
assign LUT_2[64277] = 32'b11111111111111100100111110011010;
assign LUT_2[64278] = 32'b11111111111111101110111110111101;
assign LUT_2[64279] = 32'b11111111111111101011110111010110;
assign LUT_2[64280] = 32'b11111111111111100110011001110110;
assign LUT_2[64281] = 32'b11111111111111100011010010001111;
assign LUT_2[64282] = 32'b11111111111111101101010010110010;
assign LUT_2[64283] = 32'b11111111111111101010001011001011;
assign LUT_2[64284] = 32'b11111111111111100010110111011110;
assign LUT_2[64285] = 32'b11111111111111011111101111110111;
assign LUT_2[64286] = 32'b11111111111111101001110000011010;
assign LUT_2[64287] = 32'b11111111111111100110101000110011;
assign LUT_2[64288] = 32'b11111111111111110001011111111000;
assign LUT_2[64289] = 32'b11111111111111101110011000010001;
assign LUT_2[64290] = 32'b11111111111111111000011000110100;
assign LUT_2[64291] = 32'b11111111111111110101010001001101;
assign LUT_2[64292] = 32'b11111111111111101101111101100000;
assign LUT_2[64293] = 32'b11111111111111101010110101111001;
assign LUT_2[64294] = 32'b11111111111111110100110110011100;
assign LUT_2[64295] = 32'b11111111111111110001101110110101;
assign LUT_2[64296] = 32'b11111111111111101100010001010101;
assign LUT_2[64297] = 32'b11111111111111101001001001101110;
assign LUT_2[64298] = 32'b11111111111111110011001010010001;
assign LUT_2[64299] = 32'b11111111111111110000000010101010;
assign LUT_2[64300] = 32'b11111111111111101000101110111101;
assign LUT_2[64301] = 32'b11111111111111100101100111010110;
assign LUT_2[64302] = 32'b11111111111111101111100111111001;
assign LUT_2[64303] = 32'b11111111111111101100100000010010;
assign LUT_2[64304] = 32'b11111111111111101100000100000010;
assign LUT_2[64305] = 32'b11111111111111101000111100011011;
assign LUT_2[64306] = 32'b11111111111111110010111100111110;
assign LUT_2[64307] = 32'b11111111111111101111110101010111;
assign LUT_2[64308] = 32'b11111111111111101000100001101010;
assign LUT_2[64309] = 32'b11111111111111100101011010000011;
assign LUT_2[64310] = 32'b11111111111111101111011010100110;
assign LUT_2[64311] = 32'b11111111111111101100010010111111;
assign LUT_2[64312] = 32'b11111111111111100110110101011111;
assign LUT_2[64313] = 32'b11111111111111100011101101111000;
assign LUT_2[64314] = 32'b11111111111111101101101110011011;
assign LUT_2[64315] = 32'b11111111111111101010100110110100;
assign LUT_2[64316] = 32'b11111111111111100011010011000111;
assign LUT_2[64317] = 32'b11111111111111100000001011100000;
assign LUT_2[64318] = 32'b11111111111111101010001100000011;
assign LUT_2[64319] = 32'b11111111111111100111000100011100;
assign LUT_2[64320] = 32'b11111111111111101001001100110010;
assign LUT_2[64321] = 32'b11111111111111100110000101001011;
assign LUT_2[64322] = 32'b11111111111111110000000101101110;
assign LUT_2[64323] = 32'b11111111111111101100111110000111;
assign LUT_2[64324] = 32'b11111111111111100101101010011010;
assign LUT_2[64325] = 32'b11111111111111100010100010110011;
assign LUT_2[64326] = 32'b11111111111111101100100011010110;
assign LUT_2[64327] = 32'b11111111111111101001011011101111;
assign LUT_2[64328] = 32'b11111111111111100011111110001111;
assign LUT_2[64329] = 32'b11111111111111100000110110101000;
assign LUT_2[64330] = 32'b11111111111111101010110111001011;
assign LUT_2[64331] = 32'b11111111111111100111101111100100;
assign LUT_2[64332] = 32'b11111111111111100000011011110111;
assign LUT_2[64333] = 32'b11111111111111011101010100010000;
assign LUT_2[64334] = 32'b11111111111111100111010100110011;
assign LUT_2[64335] = 32'b11111111111111100100001101001100;
assign LUT_2[64336] = 32'b11111111111111100011110000111100;
assign LUT_2[64337] = 32'b11111111111111100000101001010101;
assign LUT_2[64338] = 32'b11111111111111101010101001111000;
assign LUT_2[64339] = 32'b11111111111111100111100010010001;
assign LUT_2[64340] = 32'b11111111111111100000001110100100;
assign LUT_2[64341] = 32'b11111111111111011101000110111101;
assign LUT_2[64342] = 32'b11111111111111100111000111100000;
assign LUT_2[64343] = 32'b11111111111111100011111111111001;
assign LUT_2[64344] = 32'b11111111111111011110100010011001;
assign LUT_2[64345] = 32'b11111111111111011011011010110010;
assign LUT_2[64346] = 32'b11111111111111100101011011010101;
assign LUT_2[64347] = 32'b11111111111111100010010011101110;
assign LUT_2[64348] = 32'b11111111111111011011000000000001;
assign LUT_2[64349] = 32'b11111111111111010111111000011010;
assign LUT_2[64350] = 32'b11111111111111100001111000111101;
assign LUT_2[64351] = 32'b11111111111111011110110001010110;
assign LUT_2[64352] = 32'b11111111111111101001101000011011;
assign LUT_2[64353] = 32'b11111111111111100110100000110100;
assign LUT_2[64354] = 32'b11111111111111110000100001010111;
assign LUT_2[64355] = 32'b11111111111111101101011001110000;
assign LUT_2[64356] = 32'b11111111111111100110000110000011;
assign LUT_2[64357] = 32'b11111111111111100010111110011100;
assign LUT_2[64358] = 32'b11111111111111101100111110111111;
assign LUT_2[64359] = 32'b11111111111111101001110111011000;
assign LUT_2[64360] = 32'b11111111111111100100011001111000;
assign LUT_2[64361] = 32'b11111111111111100001010010010001;
assign LUT_2[64362] = 32'b11111111111111101011010010110100;
assign LUT_2[64363] = 32'b11111111111111101000001011001101;
assign LUT_2[64364] = 32'b11111111111111100000110111100000;
assign LUT_2[64365] = 32'b11111111111111011101101111111001;
assign LUT_2[64366] = 32'b11111111111111100111110000011100;
assign LUT_2[64367] = 32'b11111111111111100100101000110101;
assign LUT_2[64368] = 32'b11111111111111100100001100100101;
assign LUT_2[64369] = 32'b11111111111111100001000100111110;
assign LUT_2[64370] = 32'b11111111111111101011000101100001;
assign LUT_2[64371] = 32'b11111111111111100111111101111010;
assign LUT_2[64372] = 32'b11111111111111100000101010001101;
assign LUT_2[64373] = 32'b11111111111111011101100010100110;
assign LUT_2[64374] = 32'b11111111111111100111100011001001;
assign LUT_2[64375] = 32'b11111111111111100100011011100010;
assign LUT_2[64376] = 32'b11111111111111011110111110000010;
assign LUT_2[64377] = 32'b11111111111111011011110110011011;
assign LUT_2[64378] = 32'b11111111111111100101110110111110;
assign LUT_2[64379] = 32'b11111111111111100010101111010111;
assign LUT_2[64380] = 32'b11111111111111011011011011101010;
assign LUT_2[64381] = 32'b11111111111111011000010100000011;
assign LUT_2[64382] = 32'b11111111111111100010010100100110;
assign LUT_2[64383] = 32'b11111111111111011111001100111111;
assign LUT_2[64384] = 32'b11111111111111110101011000011110;
assign LUT_2[64385] = 32'b11111111111111110010010000110111;
assign LUT_2[64386] = 32'b11111111111111111100010001011010;
assign LUT_2[64387] = 32'b11111111111111111001001001110011;
assign LUT_2[64388] = 32'b11111111111111110001110110000110;
assign LUT_2[64389] = 32'b11111111111111101110101110011111;
assign LUT_2[64390] = 32'b11111111111111111000101111000010;
assign LUT_2[64391] = 32'b11111111111111110101100111011011;
assign LUT_2[64392] = 32'b11111111111111110000001001111011;
assign LUT_2[64393] = 32'b11111111111111101101000010010100;
assign LUT_2[64394] = 32'b11111111111111110111000010110111;
assign LUT_2[64395] = 32'b11111111111111110011111011010000;
assign LUT_2[64396] = 32'b11111111111111101100100111100011;
assign LUT_2[64397] = 32'b11111111111111101001011111111100;
assign LUT_2[64398] = 32'b11111111111111110011100000011111;
assign LUT_2[64399] = 32'b11111111111111110000011000111000;
assign LUT_2[64400] = 32'b11111111111111101111111100101000;
assign LUT_2[64401] = 32'b11111111111111101100110101000001;
assign LUT_2[64402] = 32'b11111111111111110110110101100100;
assign LUT_2[64403] = 32'b11111111111111110011101101111101;
assign LUT_2[64404] = 32'b11111111111111101100011010010000;
assign LUT_2[64405] = 32'b11111111111111101001010010101001;
assign LUT_2[64406] = 32'b11111111111111110011010011001100;
assign LUT_2[64407] = 32'b11111111111111110000001011100101;
assign LUT_2[64408] = 32'b11111111111111101010101110000101;
assign LUT_2[64409] = 32'b11111111111111100111100110011110;
assign LUT_2[64410] = 32'b11111111111111110001100111000001;
assign LUT_2[64411] = 32'b11111111111111101110011111011010;
assign LUT_2[64412] = 32'b11111111111111100111001011101101;
assign LUT_2[64413] = 32'b11111111111111100100000100000110;
assign LUT_2[64414] = 32'b11111111111111101110000100101001;
assign LUT_2[64415] = 32'b11111111111111101010111101000010;
assign LUT_2[64416] = 32'b11111111111111110101110100000111;
assign LUT_2[64417] = 32'b11111111111111110010101100100000;
assign LUT_2[64418] = 32'b11111111111111111100101101000011;
assign LUT_2[64419] = 32'b11111111111111111001100101011100;
assign LUT_2[64420] = 32'b11111111111111110010010001101111;
assign LUT_2[64421] = 32'b11111111111111101111001010001000;
assign LUT_2[64422] = 32'b11111111111111111001001010101011;
assign LUT_2[64423] = 32'b11111111111111110110000011000100;
assign LUT_2[64424] = 32'b11111111111111110000100101100100;
assign LUT_2[64425] = 32'b11111111111111101101011101111101;
assign LUT_2[64426] = 32'b11111111111111110111011110100000;
assign LUT_2[64427] = 32'b11111111111111110100010110111001;
assign LUT_2[64428] = 32'b11111111111111101101000011001100;
assign LUT_2[64429] = 32'b11111111111111101001111011100101;
assign LUT_2[64430] = 32'b11111111111111110011111100001000;
assign LUT_2[64431] = 32'b11111111111111110000110100100001;
assign LUT_2[64432] = 32'b11111111111111110000011000010001;
assign LUT_2[64433] = 32'b11111111111111101101010000101010;
assign LUT_2[64434] = 32'b11111111111111110111010001001101;
assign LUT_2[64435] = 32'b11111111111111110100001001100110;
assign LUT_2[64436] = 32'b11111111111111101100110101111001;
assign LUT_2[64437] = 32'b11111111111111101001101110010010;
assign LUT_2[64438] = 32'b11111111111111110011101110110101;
assign LUT_2[64439] = 32'b11111111111111110000100111001110;
assign LUT_2[64440] = 32'b11111111111111101011001001101110;
assign LUT_2[64441] = 32'b11111111111111101000000010000111;
assign LUT_2[64442] = 32'b11111111111111110010000010101010;
assign LUT_2[64443] = 32'b11111111111111101110111011000011;
assign LUT_2[64444] = 32'b11111111111111100111100111010110;
assign LUT_2[64445] = 32'b11111111111111100100011111101111;
assign LUT_2[64446] = 32'b11111111111111101110100000010010;
assign LUT_2[64447] = 32'b11111111111111101011011000101011;
assign LUT_2[64448] = 32'b11111111111111101101100001000001;
assign LUT_2[64449] = 32'b11111111111111101010011001011010;
assign LUT_2[64450] = 32'b11111111111111110100011001111101;
assign LUT_2[64451] = 32'b11111111111111110001010010010110;
assign LUT_2[64452] = 32'b11111111111111101001111110101001;
assign LUT_2[64453] = 32'b11111111111111100110110111000010;
assign LUT_2[64454] = 32'b11111111111111110000110111100101;
assign LUT_2[64455] = 32'b11111111111111101101101111111110;
assign LUT_2[64456] = 32'b11111111111111101000010010011110;
assign LUT_2[64457] = 32'b11111111111111100101001010110111;
assign LUT_2[64458] = 32'b11111111111111101111001011011010;
assign LUT_2[64459] = 32'b11111111111111101100000011110011;
assign LUT_2[64460] = 32'b11111111111111100100110000000110;
assign LUT_2[64461] = 32'b11111111111111100001101000011111;
assign LUT_2[64462] = 32'b11111111111111101011101001000010;
assign LUT_2[64463] = 32'b11111111111111101000100001011011;
assign LUT_2[64464] = 32'b11111111111111101000000101001011;
assign LUT_2[64465] = 32'b11111111111111100100111101100100;
assign LUT_2[64466] = 32'b11111111111111101110111110000111;
assign LUT_2[64467] = 32'b11111111111111101011110110100000;
assign LUT_2[64468] = 32'b11111111111111100100100010110011;
assign LUT_2[64469] = 32'b11111111111111100001011011001100;
assign LUT_2[64470] = 32'b11111111111111101011011011101111;
assign LUT_2[64471] = 32'b11111111111111101000010100001000;
assign LUT_2[64472] = 32'b11111111111111100010110110101000;
assign LUT_2[64473] = 32'b11111111111111011111101111000001;
assign LUT_2[64474] = 32'b11111111111111101001101111100100;
assign LUT_2[64475] = 32'b11111111111111100110100111111101;
assign LUT_2[64476] = 32'b11111111111111011111010100010000;
assign LUT_2[64477] = 32'b11111111111111011100001100101001;
assign LUT_2[64478] = 32'b11111111111111100110001101001100;
assign LUT_2[64479] = 32'b11111111111111100011000101100101;
assign LUT_2[64480] = 32'b11111111111111101101111100101010;
assign LUT_2[64481] = 32'b11111111111111101010110101000011;
assign LUT_2[64482] = 32'b11111111111111110100110101100110;
assign LUT_2[64483] = 32'b11111111111111110001101101111111;
assign LUT_2[64484] = 32'b11111111111111101010011010010010;
assign LUT_2[64485] = 32'b11111111111111100111010010101011;
assign LUT_2[64486] = 32'b11111111111111110001010011001110;
assign LUT_2[64487] = 32'b11111111111111101110001011100111;
assign LUT_2[64488] = 32'b11111111111111101000101110000111;
assign LUT_2[64489] = 32'b11111111111111100101100110100000;
assign LUT_2[64490] = 32'b11111111111111101111100111000011;
assign LUT_2[64491] = 32'b11111111111111101100011111011100;
assign LUT_2[64492] = 32'b11111111111111100101001011101111;
assign LUT_2[64493] = 32'b11111111111111100010000100001000;
assign LUT_2[64494] = 32'b11111111111111101100000100101011;
assign LUT_2[64495] = 32'b11111111111111101000111101000100;
assign LUT_2[64496] = 32'b11111111111111101000100000110100;
assign LUT_2[64497] = 32'b11111111111111100101011001001101;
assign LUT_2[64498] = 32'b11111111111111101111011001110000;
assign LUT_2[64499] = 32'b11111111111111101100010010001001;
assign LUT_2[64500] = 32'b11111111111111100100111110011100;
assign LUT_2[64501] = 32'b11111111111111100001110110110101;
assign LUT_2[64502] = 32'b11111111111111101011110111011000;
assign LUT_2[64503] = 32'b11111111111111101000101111110001;
assign LUT_2[64504] = 32'b11111111111111100011010010010001;
assign LUT_2[64505] = 32'b11111111111111100000001010101010;
assign LUT_2[64506] = 32'b11111111111111101010001011001101;
assign LUT_2[64507] = 32'b11111111111111100111000011100110;
assign LUT_2[64508] = 32'b11111111111111011111101111111001;
assign LUT_2[64509] = 32'b11111111111111011100101000010010;
assign LUT_2[64510] = 32'b11111111111111100110101000110101;
assign LUT_2[64511] = 32'b11111111111111100011100001001110;
assign LUT_2[64512] = 32'b11111111111111101110111111111100;
assign LUT_2[64513] = 32'b11111111111111101011111000010101;
assign LUT_2[64514] = 32'b11111111111111110101111000111000;
assign LUT_2[64515] = 32'b11111111111111110010110001010001;
assign LUT_2[64516] = 32'b11111111111111101011011101100100;
assign LUT_2[64517] = 32'b11111111111111101000010101111101;
assign LUT_2[64518] = 32'b11111111111111110010010110100000;
assign LUT_2[64519] = 32'b11111111111111101111001110111001;
assign LUT_2[64520] = 32'b11111111111111101001110001011001;
assign LUT_2[64521] = 32'b11111111111111100110101001110010;
assign LUT_2[64522] = 32'b11111111111111110000101010010101;
assign LUT_2[64523] = 32'b11111111111111101101100010101110;
assign LUT_2[64524] = 32'b11111111111111100110001111000001;
assign LUT_2[64525] = 32'b11111111111111100011000111011010;
assign LUT_2[64526] = 32'b11111111111111101101000111111101;
assign LUT_2[64527] = 32'b11111111111111101010000000010110;
assign LUT_2[64528] = 32'b11111111111111101001100100000110;
assign LUT_2[64529] = 32'b11111111111111100110011100011111;
assign LUT_2[64530] = 32'b11111111111111110000011101000010;
assign LUT_2[64531] = 32'b11111111111111101101010101011011;
assign LUT_2[64532] = 32'b11111111111111100110000001101110;
assign LUT_2[64533] = 32'b11111111111111100010111010000111;
assign LUT_2[64534] = 32'b11111111111111101100111010101010;
assign LUT_2[64535] = 32'b11111111111111101001110011000011;
assign LUT_2[64536] = 32'b11111111111111100100010101100011;
assign LUT_2[64537] = 32'b11111111111111100001001101111100;
assign LUT_2[64538] = 32'b11111111111111101011001110011111;
assign LUT_2[64539] = 32'b11111111111111101000000110111000;
assign LUT_2[64540] = 32'b11111111111111100000110011001011;
assign LUT_2[64541] = 32'b11111111111111011101101011100100;
assign LUT_2[64542] = 32'b11111111111111100111101100000111;
assign LUT_2[64543] = 32'b11111111111111100100100100100000;
assign LUT_2[64544] = 32'b11111111111111101111011011100101;
assign LUT_2[64545] = 32'b11111111111111101100010011111110;
assign LUT_2[64546] = 32'b11111111111111110110010100100001;
assign LUT_2[64547] = 32'b11111111111111110011001100111010;
assign LUT_2[64548] = 32'b11111111111111101011111001001101;
assign LUT_2[64549] = 32'b11111111111111101000110001100110;
assign LUT_2[64550] = 32'b11111111111111110010110010001001;
assign LUT_2[64551] = 32'b11111111111111101111101010100010;
assign LUT_2[64552] = 32'b11111111111111101010001101000010;
assign LUT_2[64553] = 32'b11111111111111100111000101011011;
assign LUT_2[64554] = 32'b11111111111111110001000101111110;
assign LUT_2[64555] = 32'b11111111111111101101111110010111;
assign LUT_2[64556] = 32'b11111111111111100110101010101010;
assign LUT_2[64557] = 32'b11111111111111100011100011000011;
assign LUT_2[64558] = 32'b11111111111111101101100011100110;
assign LUT_2[64559] = 32'b11111111111111101010011011111111;
assign LUT_2[64560] = 32'b11111111111111101001111111101111;
assign LUT_2[64561] = 32'b11111111111111100110111000001000;
assign LUT_2[64562] = 32'b11111111111111110000111000101011;
assign LUT_2[64563] = 32'b11111111111111101101110001000100;
assign LUT_2[64564] = 32'b11111111111111100110011101010111;
assign LUT_2[64565] = 32'b11111111111111100011010101110000;
assign LUT_2[64566] = 32'b11111111111111101101010110010011;
assign LUT_2[64567] = 32'b11111111111111101010001110101100;
assign LUT_2[64568] = 32'b11111111111111100100110001001100;
assign LUT_2[64569] = 32'b11111111111111100001101001100101;
assign LUT_2[64570] = 32'b11111111111111101011101010001000;
assign LUT_2[64571] = 32'b11111111111111101000100010100001;
assign LUT_2[64572] = 32'b11111111111111100001001110110100;
assign LUT_2[64573] = 32'b11111111111111011110000111001101;
assign LUT_2[64574] = 32'b11111111111111101000000111110000;
assign LUT_2[64575] = 32'b11111111111111100101000000001001;
assign LUT_2[64576] = 32'b11111111111111100111001000011111;
assign LUT_2[64577] = 32'b11111111111111100100000000111000;
assign LUT_2[64578] = 32'b11111111111111101110000001011011;
assign LUT_2[64579] = 32'b11111111111111101010111001110100;
assign LUT_2[64580] = 32'b11111111111111100011100110000111;
assign LUT_2[64581] = 32'b11111111111111100000011110100000;
assign LUT_2[64582] = 32'b11111111111111101010011111000011;
assign LUT_2[64583] = 32'b11111111111111100111010111011100;
assign LUT_2[64584] = 32'b11111111111111100001111001111100;
assign LUT_2[64585] = 32'b11111111111111011110110010010101;
assign LUT_2[64586] = 32'b11111111111111101000110010111000;
assign LUT_2[64587] = 32'b11111111111111100101101011010001;
assign LUT_2[64588] = 32'b11111111111111011110010111100100;
assign LUT_2[64589] = 32'b11111111111111011011001111111101;
assign LUT_2[64590] = 32'b11111111111111100101010000100000;
assign LUT_2[64591] = 32'b11111111111111100010001000111001;
assign LUT_2[64592] = 32'b11111111111111100001101100101001;
assign LUT_2[64593] = 32'b11111111111111011110100101000010;
assign LUT_2[64594] = 32'b11111111111111101000100101100101;
assign LUT_2[64595] = 32'b11111111111111100101011101111110;
assign LUT_2[64596] = 32'b11111111111111011110001010010001;
assign LUT_2[64597] = 32'b11111111111111011011000010101010;
assign LUT_2[64598] = 32'b11111111111111100101000011001101;
assign LUT_2[64599] = 32'b11111111111111100001111011100110;
assign LUT_2[64600] = 32'b11111111111111011100011110000110;
assign LUT_2[64601] = 32'b11111111111111011001010110011111;
assign LUT_2[64602] = 32'b11111111111111100011010111000010;
assign LUT_2[64603] = 32'b11111111111111100000001111011011;
assign LUT_2[64604] = 32'b11111111111111011000111011101110;
assign LUT_2[64605] = 32'b11111111111111010101110100000111;
assign LUT_2[64606] = 32'b11111111111111011111110100101010;
assign LUT_2[64607] = 32'b11111111111111011100101101000011;
assign LUT_2[64608] = 32'b11111111111111100111100100001000;
assign LUT_2[64609] = 32'b11111111111111100100011100100001;
assign LUT_2[64610] = 32'b11111111111111101110011101000100;
assign LUT_2[64611] = 32'b11111111111111101011010101011101;
assign LUT_2[64612] = 32'b11111111111111100100000001110000;
assign LUT_2[64613] = 32'b11111111111111100000111010001001;
assign LUT_2[64614] = 32'b11111111111111101010111010101100;
assign LUT_2[64615] = 32'b11111111111111100111110011000101;
assign LUT_2[64616] = 32'b11111111111111100010010101100101;
assign LUT_2[64617] = 32'b11111111111111011111001101111110;
assign LUT_2[64618] = 32'b11111111111111101001001110100001;
assign LUT_2[64619] = 32'b11111111111111100110000110111010;
assign LUT_2[64620] = 32'b11111111111111011110110011001101;
assign LUT_2[64621] = 32'b11111111111111011011101011100110;
assign LUT_2[64622] = 32'b11111111111111100101101100001001;
assign LUT_2[64623] = 32'b11111111111111100010100100100010;
assign LUT_2[64624] = 32'b11111111111111100010001000010010;
assign LUT_2[64625] = 32'b11111111111111011111000000101011;
assign LUT_2[64626] = 32'b11111111111111101001000001001110;
assign LUT_2[64627] = 32'b11111111111111100101111001100111;
assign LUT_2[64628] = 32'b11111111111111011110100101111010;
assign LUT_2[64629] = 32'b11111111111111011011011110010011;
assign LUT_2[64630] = 32'b11111111111111100101011110110110;
assign LUT_2[64631] = 32'b11111111111111100010010111001111;
assign LUT_2[64632] = 32'b11111111111111011100111001101111;
assign LUT_2[64633] = 32'b11111111111111011001110010001000;
assign LUT_2[64634] = 32'b11111111111111100011110010101011;
assign LUT_2[64635] = 32'b11111111111111100000101011000100;
assign LUT_2[64636] = 32'b11111111111111011001010111010111;
assign LUT_2[64637] = 32'b11111111111111010110001111110000;
assign LUT_2[64638] = 32'b11111111111111100000010000010011;
assign LUT_2[64639] = 32'b11111111111111011101001000101100;
assign LUT_2[64640] = 32'b11111111111111110011010100001011;
assign LUT_2[64641] = 32'b11111111111111110000001100100100;
assign LUT_2[64642] = 32'b11111111111111111010001101000111;
assign LUT_2[64643] = 32'b11111111111111110111000101100000;
assign LUT_2[64644] = 32'b11111111111111101111110001110011;
assign LUT_2[64645] = 32'b11111111111111101100101010001100;
assign LUT_2[64646] = 32'b11111111111111110110101010101111;
assign LUT_2[64647] = 32'b11111111111111110011100011001000;
assign LUT_2[64648] = 32'b11111111111111101110000101101000;
assign LUT_2[64649] = 32'b11111111111111101010111110000001;
assign LUT_2[64650] = 32'b11111111111111110100111110100100;
assign LUT_2[64651] = 32'b11111111111111110001110110111101;
assign LUT_2[64652] = 32'b11111111111111101010100011010000;
assign LUT_2[64653] = 32'b11111111111111100111011011101001;
assign LUT_2[64654] = 32'b11111111111111110001011100001100;
assign LUT_2[64655] = 32'b11111111111111101110010100100101;
assign LUT_2[64656] = 32'b11111111111111101101111000010101;
assign LUT_2[64657] = 32'b11111111111111101010110000101110;
assign LUT_2[64658] = 32'b11111111111111110100110001010001;
assign LUT_2[64659] = 32'b11111111111111110001101001101010;
assign LUT_2[64660] = 32'b11111111111111101010010101111101;
assign LUT_2[64661] = 32'b11111111111111100111001110010110;
assign LUT_2[64662] = 32'b11111111111111110001001110111001;
assign LUT_2[64663] = 32'b11111111111111101110000111010010;
assign LUT_2[64664] = 32'b11111111111111101000101001110010;
assign LUT_2[64665] = 32'b11111111111111100101100010001011;
assign LUT_2[64666] = 32'b11111111111111101111100010101110;
assign LUT_2[64667] = 32'b11111111111111101100011011000111;
assign LUT_2[64668] = 32'b11111111111111100101000111011010;
assign LUT_2[64669] = 32'b11111111111111100001111111110011;
assign LUT_2[64670] = 32'b11111111111111101100000000010110;
assign LUT_2[64671] = 32'b11111111111111101000111000101111;
assign LUT_2[64672] = 32'b11111111111111110011101111110100;
assign LUT_2[64673] = 32'b11111111111111110000101000001101;
assign LUT_2[64674] = 32'b11111111111111111010101000110000;
assign LUT_2[64675] = 32'b11111111111111110111100001001001;
assign LUT_2[64676] = 32'b11111111111111110000001101011100;
assign LUT_2[64677] = 32'b11111111111111101101000101110101;
assign LUT_2[64678] = 32'b11111111111111110111000110011000;
assign LUT_2[64679] = 32'b11111111111111110011111110110001;
assign LUT_2[64680] = 32'b11111111111111101110100001010001;
assign LUT_2[64681] = 32'b11111111111111101011011001101010;
assign LUT_2[64682] = 32'b11111111111111110101011010001101;
assign LUT_2[64683] = 32'b11111111111111110010010010100110;
assign LUT_2[64684] = 32'b11111111111111101010111110111001;
assign LUT_2[64685] = 32'b11111111111111100111110111010010;
assign LUT_2[64686] = 32'b11111111111111110001110111110101;
assign LUT_2[64687] = 32'b11111111111111101110110000001110;
assign LUT_2[64688] = 32'b11111111111111101110010011111110;
assign LUT_2[64689] = 32'b11111111111111101011001100010111;
assign LUT_2[64690] = 32'b11111111111111110101001100111010;
assign LUT_2[64691] = 32'b11111111111111110010000101010011;
assign LUT_2[64692] = 32'b11111111111111101010110001100110;
assign LUT_2[64693] = 32'b11111111111111100111101001111111;
assign LUT_2[64694] = 32'b11111111111111110001101010100010;
assign LUT_2[64695] = 32'b11111111111111101110100010111011;
assign LUT_2[64696] = 32'b11111111111111101001000101011011;
assign LUT_2[64697] = 32'b11111111111111100101111101110100;
assign LUT_2[64698] = 32'b11111111111111101111111110010111;
assign LUT_2[64699] = 32'b11111111111111101100110110110000;
assign LUT_2[64700] = 32'b11111111111111100101100011000011;
assign LUT_2[64701] = 32'b11111111111111100010011011011100;
assign LUT_2[64702] = 32'b11111111111111101100011011111111;
assign LUT_2[64703] = 32'b11111111111111101001010100011000;
assign LUT_2[64704] = 32'b11111111111111101011011100101110;
assign LUT_2[64705] = 32'b11111111111111101000010101000111;
assign LUT_2[64706] = 32'b11111111111111110010010101101010;
assign LUT_2[64707] = 32'b11111111111111101111001110000011;
assign LUT_2[64708] = 32'b11111111111111100111111010010110;
assign LUT_2[64709] = 32'b11111111111111100100110010101111;
assign LUT_2[64710] = 32'b11111111111111101110110011010010;
assign LUT_2[64711] = 32'b11111111111111101011101011101011;
assign LUT_2[64712] = 32'b11111111111111100110001110001011;
assign LUT_2[64713] = 32'b11111111111111100011000110100100;
assign LUT_2[64714] = 32'b11111111111111101101000111000111;
assign LUT_2[64715] = 32'b11111111111111101001111111100000;
assign LUT_2[64716] = 32'b11111111111111100010101011110011;
assign LUT_2[64717] = 32'b11111111111111011111100100001100;
assign LUT_2[64718] = 32'b11111111111111101001100100101111;
assign LUT_2[64719] = 32'b11111111111111100110011101001000;
assign LUT_2[64720] = 32'b11111111111111100110000000111000;
assign LUT_2[64721] = 32'b11111111111111100010111001010001;
assign LUT_2[64722] = 32'b11111111111111101100111001110100;
assign LUT_2[64723] = 32'b11111111111111101001110010001101;
assign LUT_2[64724] = 32'b11111111111111100010011110100000;
assign LUT_2[64725] = 32'b11111111111111011111010110111001;
assign LUT_2[64726] = 32'b11111111111111101001010111011100;
assign LUT_2[64727] = 32'b11111111111111100110001111110101;
assign LUT_2[64728] = 32'b11111111111111100000110010010101;
assign LUT_2[64729] = 32'b11111111111111011101101010101110;
assign LUT_2[64730] = 32'b11111111111111100111101011010001;
assign LUT_2[64731] = 32'b11111111111111100100100011101010;
assign LUT_2[64732] = 32'b11111111111111011101001111111101;
assign LUT_2[64733] = 32'b11111111111111011010001000010110;
assign LUT_2[64734] = 32'b11111111111111100100001000111001;
assign LUT_2[64735] = 32'b11111111111111100001000001010010;
assign LUT_2[64736] = 32'b11111111111111101011111000010111;
assign LUT_2[64737] = 32'b11111111111111101000110000110000;
assign LUT_2[64738] = 32'b11111111111111110010110001010011;
assign LUT_2[64739] = 32'b11111111111111101111101001101100;
assign LUT_2[64740] = 32'b11111111111111101000010101111111;
assign LUT_2[64741] = 32'b11111111111111100101001110011000;
assign LUT_2[64742] = 32'b11111111111111101111001110111011;
assign LUT_2[64743] = 32'b11111111111111101100000111010100;
assign LUT_2[64744] = 32'b11111111111111100110101001110100;
assign LUT_2[64745] = 32'b11111111111111100011100010001101;
assign LUT_2[64746] = 32'b11111111111111101101100010110000;
assign LUT_2[64747] = 32'b11111111111111101010011011001001;
assign LUT_2[64748] = 32'b11111111111111100011000111011100;
assign LUT_2[64749] = 32'b11111111111111011111111111110101;
assign LUT_2[64750] = 32'b11111111111111101010000000011000;
assign LUT_2[64751] = 32'b11111111111111100110111000110001;
assign LUT_2[64752] = 32'b11111111111111100110011100100001;
assign LUT_2[64753] = 32'b11111111111111100011010100111010;
assign LUT_2[64754] = 32'b11111111111111101101010101011101;
assign LUT_2[64755] = 32'b11111111111111101010001101110110;
assign LUT_2[64756] = 32'b11111111111111100010111010001001;
assign LUT_2[64757] = 32'b11111111111111011111110010100010;
assign LUT_2[64758] = 32'b11111111111111101001110011000101;
assign LUT_2[64759] = 32'b11111111111111100110101011011110;
assign LUT_2[64760] = 32'b11111111111111100001001101111110;
assign LUT_2[64761] = 32'b11111111111111011110000110010111;
assign LUT_2[64762] = 32'b11111111111111101000000110111010;
assign LUT_2[64763] = 32'b11111111111111100100111111010011;
assign LUT_2[64764] = 32'b11111111111111011101101011100110;
assign LUT_2[64765] = 32'b11111111111111011010100011111111;
assign LUT_2[64766] = 32'b11111111111111100100100100100010;
assign LUT_2[64767] = 32'b11111111111111100001011100111011;
assign LUT_2[64768] = 32'b11111111111111110010111110100010;
assign LUT_2[64769] = 32'b11111111111111101111110110111011;
assign LUT_2[64770] = 32'b11111111111111111001110111011110;
assign LUT_2[64771] = 32'b11111111111111110110101111110111;
assign LUT_2[64772] = 32'b11111111111111101111011100001010;
assign LUT_2[64773] = 32'b11111111111111101100010100100011;
assign LUT_2[64774] = 32'b11111111111111110110010101000110;
assign LUT_2[64775] = 32'b11111111111111110011001101011111;
assign LUT_2[64776] = 32'b11111111111111101101101111111111;
assign LUT_2[64777] = 32'b11111111111111101010101000011000;
assign LUT_2[64778] = 32'b11111111111111110100101000111011;
assign LUT_2[64779] = 32'b11111111111111110001100001010100;
assign LUT_2[64780] = 32'b11111111111111101010001101100111;
assign LUT_2[64781] = 32'b11111111111111100111000110000000;
assign LUT_2[64782] = 32'b11111111111111110001000110100011;
assign LUT_2[64783] = 32'b11111111111111101101111110111100;
assign LUT_2[64784] = 32'b11111111111111101101100010101100;
assign LUT_2[64785] = 32'b11111111111111101010011011000101;
assign LUT_2[64786] = 32'b11111111111111110100011011101000;
assign LUT_2[64787] = 32'b11111111111111110001010100000001;
assign LUT_2[64788] = 32'b11111111111111101010000000010100;
assign LUT_2[64789] = 32'b11111111111111100110111000101101;
assign LUT_2[64790] = 32'b11111111111111110000111001010000;
assign LUT_2[64791] = 32'b11111111111111101101110001101001;
assign LUT_2[64792] = 32'b11111111111111101000010100001001;
assign LUT_2[64793] = 32'b11111111111111100101001100100010;
assign LUT_2[64794] = 32'b11111111111111101111001101000101;
assign LUT_2[64795] = 32'b11111111111111101100000101011110;
assign LUT_2[64796] = 32'b11111111111111100100110001110001;
assign LUT_2[64797] = 32'b11111111111111100001101010001010;
assign LUT_2[64798] = 32'b11111111111111101011101010101101;
assign LUT_2[64799] = 32'b11111111111111101000100011000110;
assign LUT_2[64800] = 32'b11111111111111110011011010001011;
assign LUT_2[64801] = 32'b11111111111111110000010010100100;
assign LUT_2[64802] = 32'b11111111111111111010010011000111;
assign LUT_2[64803] = 32'b11111111111111110111001011100000;
assign LUT_2[64804] = 32'b11111111111111101111110111110011;
assign LUT_2[64805] = 32'b11111111111111101100110000001100;
assign LUT_2[64806] = 32'b11111111111111110110110000101111;
assign LUT_2[64807] = 32'b11111111111111110011101001001000;
assign LUT_2[64808] = 32'b11111111111111101110001011101000;
assign LUT_2[64809] = 32'b11111111111111101011000100000001;
assign LUT_2[64810] = 32'b11111111111111110101000100100100;
assign LUT_2[64811] = 32'b11111111111111110001111100111101;
assign LUT_2[64812] = 32'b11111111111111101010101001010000;
assign LUT_2[64813] = 32'b11111111111111100111100001101001;
assign LUT_2[64814] = 32'b11111111111111110001100010001100;
assign LUT_2[64815] = 32'b11111111111111101110011010100101;
assign LUT_2[64816] = 32'b11111111111111101101111110010101;
assign LUT_2[64817] = 32'b11111111111111101010110110101110;
assign LUT_2[64818] = 32'b11111111111111110100110111010001;
assign LUT_2[64819] = 32'b11111111111111110001101111101010;
assign LUT_2[64820] = 32'b11111111111111101010011011111101;
assign LUT_2[64821] = 32'b11111111111111100111010100010110;
assign LUT_2[64822] = 32'b11111111111111110001010100111001;
assign LUT_2[64823] = 32'b11111111111111101110001101010010;
assign LUT_2[64824] = 32'b11111111111111101000101111110010;
assign LUT_2[64825] = 32'b11111111111111100101101000001011;
assign LUT_2[64826] = 32'b11111111111111101111101000101110;
assign LUT_2[64827] = 32'b11111111111111101100100001000111;
assign LUT_2[64828] = 32'b11111111111111100101001101011010;
assign LUT_2[64829] = 32'b11111111111111100010000101110011;
assign LUT_2[64830] = 32'b11111111111111101100000110010110;
assign LUT_2[64831] = 32'b11111111111111101000111110101111;
assign LUT_2[64832] = 32'b11111111111111101011000111000101;
assign LUT_2[64833] = 32'b11111111111111100111111111011110;
assign LUT_2[64834] = 32'b11111111111111110010000000000001;
assign LUT_2[64835] = 32'b11111111111111101110111000011010;
assign LUT_2[64836] = 32'b11111111111111100111100100101101;
assign LUT_2[64837] = 32'b11111111111111100100011101000110;
assign LUT_2[64838] = 32'b11111111111111101110011101101001;
assign LUT_2[64839] = 32'b11111111111111101011010110000010;
assign LUT_2[64840] = 32'b11111111111111100101111000100010;
assign LUT_2[64841] = 32'b11111111111111100010110000111011;
assign LUT_2[64842] = 32'b11111111111111101100110001011110;
assign LUT_2[64843] = 32'b11111111111111101001101001110111;
assign LUT_2[64844] = 32'b11111111111111100010010110001010;
assign LUT_2[64845] = 32'b11111111111111011111001110100011;
assign LUT_2[64846] = 32'b11111111111111101001001111000110;
assign LUT_2[64847] = 32'b11111111111111100110000111011111;
assign LUT_2[64848] = 32'b11111111111111100101101011001111;
assign LUT_2[64849] = 32'b11111111111111100010100011101000;
assign LUT_2[64850] = 32'b11111111111111101100100100001011;
assign LUT_2[64851] = 32'b11111111111111101001011100100100;
assign LUT_2[64852] = 32'b11111111111111100010001000110111;
assign LUT_2[64853] = 32'b11111111111111011111000001010000;
assign LUT_2[64854] = 32'b11111111111111101001000001110011;
assign LUT_2[64855] = 32'b11111111111111100101111010001100;
assign LUT_2[64856] = 32'b11111111111111100000011100101100;
assign LUT_2[64857] = 32'b11111111111111011101010101000101;
assign LUT_2[64858] = 32'b11111111111111100111010101101000;
assign LUT_2[64859] = 32'b11111111111111100100001110000001;
assign LUT_2[64860] = 32'b11111111111111011100111010010100;
assign LUT_2[64861] = 32'b11111111111111011001110010101101;
assign LUT_2[64862] = 32'b11111111111111100011110011010000;
assign LUT_2[64863] = 32'b11111111111111100000101011101001;
assign LUT_2[64864] = 32'b11111111111111101011100010101110;
assign LUT_2[64865] = 32'b11111111111111101000011011000111;
assign LUT_2[64866] = 32'b11111111111111110010011011101010;
assign LUT_2[64867] = 32'b11111111111111101111010100000011;
assign LUT_2[64868] = 32'b11111111111111101000000000010110;
assign LUT_2[64869] = 32'b11111111111111100100111000101111;
assign LUT_2[64870] = 32'b11111111111111101110111001010010;
assign LUT_2[64871] = 32'b11111111111111101011110001101011;
assign LUT_2[64872] = 32'b11111111111111100110010100001011;
assign LUT_2[64873] = 32'b11111111111111100011001100100100;
assign LUT_2[64874] = 32'b11111111111111101101001101000111;
assign LUT_2[64875] = 32'b11111111111111101010000101100000;
assign LUT_2[64876] = 32'b11111111111111100010110001110011;
assign LUT_2[64877] = 32'b11111111111111011111101010001100;
assign LUT_2[64878] = 32'b11111111111111101001101010101111;
assign LUT_2[64879] = 32'b11111111111111100110100011001000;
assign LUT_2[64880] = 32'b11111111111111100110000110111000;
assign LUT_2[64881] = 32'b11111111111111100010111111010001;
assign LUT_2[64882] = 32'b11111111111111101100111111110100;
assign LUT_2[64883] = 32'b11111111111111101001111000001101;
assign LUT_2[64884] = 32'b11111111111111100010100100100000;
assign LUT_2[64885] = 32'b11111111111111011111011100111001;
assign LUT_2[64886] = 32'b11111111111111101001011101011100;
assign LUT_2[64887] = 32'b11111111111111100110010101110101;
assign LUT_2[64888] = 32'b11111111111111100000111000010101;
assign LUT_2[64889] = 32'b11111111111111011101110000101110;
assign LUT_2[64890] = 32'b11111111111111100111110001010001;
assign LUT_2[64891] = 32'b11111111111111100100101001101010;
assign LUT_2[64892] = 32'b11111111111111011101010101111101;
assign LUT_2[64893] = 32'b11111111111111011010001110010110;
assign LUT_2[64894] = 32'b11111111111111100100001110111001;
assign LUT_2[64895] = 32'b11111111111111100001000111010010;
assign LUT_2[64896] = 32'b11111111111111110111010010110001;
assign LUT_2[64897] = 32'b11111111111111110100001011001010;
assign LUT_2[64898] = 32'b11111111111111111110001011101101;
assign LUT_2[64899] = 32'b11111111111111111011000100000110;
assign LUT_2[64900] = 32'b11111111111111110011110000011001;
assign LUT_2[64901] = 32'b11111111111111110000101000110010;
assign LUT_2[64902] = 32'b11111111111111111010101001010101;
assign LUT_2[64903] = 32'b11111111111111110111100001101110;
assign LUT_2[64904] = 32'b11111111111111110010000100001110;
assign LUT_2[64905] = 32'b11111111111111101110111100100111;
assign LUT_2[64906] = 32'b11111111111111111000111101001010;
assign LUT_2[64907] = 32'b11111111111111110101110101100011;
assign LUT_2[64908] = 32'b11111111111111101110100001110110;
assign LUT_2[64909] = 32'b11111111111111101011011010001111;
assign LUT_2[64910] = 32'b11111111111111110101011010110010;
assign LUT_2[64911] = 32'b11111111111111110010010011001011;
assign LUT_2[64912] = 32'b11111111111111110001110110111011;
assign LUT_2[64913] = 32'b11111111111111101110101111010100;
assign LUT_2[64914] = 32'b11111111111111111000101111110111;
assign LUT_2[64915] = 32'b11111111111111110101101000010000;
assign LUT_2[64916] = 32'b11111111111111101110010100100011;
assign LUT_2[64917] = 32'b11111111111111101011001100111100;
assign LUT_2[64918] = 32'b11111111111111110101001101011111;
assign LUT_2[64919] = 32'b11111111111111110010000101111000;
assign LUT_2[64920] = 32'b11111111111111101100101000011000;
assign LUT_2[64921] = 32'b11111111111111101001100000110001;
assign LUT_2[64922] = 32'b11111111111111110011100001010100;
assign LUT_2[64923] = 32'b11111111111111110000011001101101;
assign LUT_2[64924] = 32'b11111111111111101001000110000000;
assign LUT_2[64925] = 32'b11111111111111100101111110011001;
assign LUT_2[64926] = 32'b11111111111111101111111110111100;
assign LUT_2[64927] = 32'b11111111111111101100110111010101;
assign LUT_2[64928] = 32'b11111111111111110111101110011010;
assign LUT_2[64929] = 32'b11111111111111110100100110110011;
assign LUT_2[64930] = 32'b11111111111111111110100111010110;
assign LUT_2[64931] = 32'b11111111111111111011011111101111;
assign LUT_2[64932] = 32'b11111111111111110100001100000010;
assign LUT_2[64933] = 32'b11111111111111110001000100011011;
assign LUT_2[64934] = 32'b11111111111111111011000100111110;
assign LUT_2[64935] = 32'b11111111111111110111111101010111;
assign LUT_2[64936] = 32'b11111111111111110010011111110111;
assign LUT_2[64937] = 32'b11111111111111101111011000010000;
assign LUT_2[64938] = 32'b11111111111111111001011000110011;
assign LUT_2[64939] = 32'b11111111111111110110010001001100;
assign LUT_2[64940] = 32'b11111111111111101110111101011111;
assign LUT_2[64941] = 32'b11111111111111101011110101111000;
assign LUT_2[64942] = 32'b11111111111111110101110110011011;
assign LUT_2[64943] = 32'b11111111111111110010101110110100;
assign LUT_2[64944] = 32'b11111111111111110010010010100100;
assign LUT_2[64945] = 32'b11111111111111101111001010111101;
assign LUT_2[64946] = 32'b11111111111111111001001011100000;
assign LUT_2[64947] = 32'b11111111111111110110000011111001;
assign LUT_2[64948] = 32'b11111111111111101110110000001100;
assign LUT_2[64949] = 32'b11111111111111101011101000100101;
assign LUT_2[64950] = 32'b11111111111111110101101001001000;
assign LUT_2[64951] = 32'b11111111111111110010100001100001;
assign LUT_2[64952] = 32'b11111111111111101101000100000001;
assign LUT_2[64953] = 32'b11111111111111101001111100011010;
assign LUT_2[64954] = 32'b11111111111111110011111100111101;
assign LUT_2[64955] = 32'b11111111111111110000110101010110;
assign LUT_2[64956] = 32'b11111111111111101001100001101001;
assign LUT_2[64957] = 32'b11111111111111100110011010000010;
assign LUT_2[64958] = 32'b11111111111111110000011010100101;
assign LUT_2[64959] = 32'b11111111111111101101010010111110;
assign LUT_2[64960] = 32'b11111111111111101111011011010100;
assign LUT_2[64961] = 32'b11111111111111101100010011101101;
assign LUT_2[64962] = 32'b11111111111111110110010100010000;
assign LUT_2[64963] = 32'b11111111111111110011001100101001;
assign LUT_2[64964] = 32'b11111111111111101011111000111100;
assign LUT_2[64965] = 32'b11111111111111101000110001010101;
assign LUT_2[64966] = 32'b11111111111111110010110001111000;
assign LUT_2[64967] = 32'b11111111111111101111101010010001;
assign LUT_2[64968] = 32'b11111111111111101010001100110001;
assign LUT_2[64969] = 32'b11111111111111100111000101001010;
assign LUT_2[64970] = 32'b11111111111111110001000101101101;
assign LUT_2[64971] = 32'b11111111111111101101111110000110;
assign LUT_2[64972] = 32'b11111111111111100110101010011001;
assign LUT_2[64973] = 32'b11111111111111100011100010110010;
assign LUT_2[64974] = 32'b11111111111111101101100011010101;
assign LUT_2[64975] = 32'b11111111111111101010011011101110;
assign LUT_2[64976] = 32'b11111111111111101001111111011110;
assign LUT_2[64977] = 32'b11111111111111100110110111110111;
assign LUT_2[64978] = 32'b11111111111111110000111000011010;
assign LUT_2[64979] = 32'b11111111111111101101110000110011;
assign LUT_2[64980] = 32'b11111111111111100110011101000110;
assign LUT_2[64981] = 32'b11111111111111100011010101011111;
assign LUT_2[64982] = 32'b11111111111111101101010110000010;
assign LUT_2[64983] = 32'b11111111111111101010001110011011;
assign LUT_2[64984] = 32'b11111111111111100100110000111011;
assign LUT_2[64985] = 32'b11111111111111100001101001010100;
assign LUT_2[64986] = 32'b11111111111111101011101001110111;
assign LUT_2[64987] = 32'b11111111111111101000100010010000;
assign LUT_2[64988] = 32'b11111111111111100001001110100011;
assign LUT_2[64989] = 32'b11111111111111011110000110111100;
assign LUT_2[64990] = 32'b11111111111111101000000111011111;
assign LUT_2[64991] = 32'b11111111111111100100111111111000;
assign LUT_2[64992] = 32'b11111111111111101111110110111101;
assign LUT_2[64993] = 32'b11111111111111101100101111010110;
assign LUT_2[64994] = 32'b11111111111111110110101111111001;
assign LUT_2[64995] = 32'b11111111111111110011101000010010;
assign LUT_2[64996] = 32'b11111111111111101100010100100101;
assign LUT_2[64997] = 32'b11111111111111101001001100111110;
assign LUT_2[64998] = 32'b11111111111111110011001101100001;
assign LUT_2[64999] = 32'b11111111111111110000000101111010;
assign LUT_2[65000] = 32'b11111111111111101010101000011010;
assign LUT_2[65001] = 32'b11111111111111100111100000110011;
assign LUT_2[65002] = 32'b11111111111111110001100001010110;
assign LUT_2[65003] = 32'b11111111111111101110011001101111;
assign LUT_2[65004] = 32'b11111111111111100111000110000010;
assign LUT_2[65005] = 32'b11111111111111100011111110011011;
assign LUT_2[65006] = 32'b11111111111111101101111110111110;
assign LUT_2[65007] = 32'b11111111111111101010110111010111;
assign LUT_2[65008] = 32'b11111111111111101010011011000111;
assign LUT_2[65009] = 32'b11111111111111100111010011100000;
assign LUT_2[65010] = 32'b11111111111111110001010100000011;
assign LUT_2[65011] = 32'b11111111111111101110001100011100;
assign LUT_2[65012] = 32'b11111111111111100110111000101111;
assign LUT_2[65013] = 32'b11111111111111100011110001001000;
assign LUT_2[65014] = 32'b11111111111111101101110001101011;
assign LUT_2[65015] = 32'b11111111111111101010101010000100;
assign LUT_2[65016] = 32'b11111111111111100101001100100100;
assign LUT_2[65017] = 32'b11111111111111100010000100111101;
assign LUT_2[65018] = 32'b11111111111111101100000101100000;
assign LUT_2[65019] = 32'b11111111111111101000111101111001;
assign LUT_2[65020] = 32'b11111111111111100001101010001100;
assign LUT_2[65021] = 32'b11111111111111011110100010100101;
assign LUT_2[65022] = 32'b11111111111111101000100011001000;
assign LUT_2[65023] = 32'b11111111111111100101011011100001;
assign LUT_2[65024] = 32'b11111111111111110011110001101110;
assign LUT_2[65025] = 32'b11111111111111110000101010000111;
assign LUT_2[65026] = 32'b11111111111111111010101010101010;
assign LUT_2[65027] = 32'b11111111111111110111100011000011;
assign LUT_2[65028] = 32'b11111111111111110000001111010110;
assign LUT_2[65029] = 32'b11111111111111101101000111101111;
assign LUT_2[65030] = 32'b11111111111111110111001000010010;
assign LUT_2[65031] = 32'b11111111111111110100000000101011;
assign LUT_2[65032] = 32'b11111111111111101110100011001011;
assign LUT_2[65033] = 32'b11111111111111101011011011100100;
assign LUT_2[65034] = 32'b11111111111111110101011100000111;
assign LUT_2[65035] = 32'b11111111111111110010010100100000;
assign LUT_2[65036] = 32'b11111111111111101011000000110011;
assign LUT_2[65037] = 32'b11111111111111100111111001001100;
assign LUT_2[65038] = 32'b11111111111111110001111001101111;
assign LUT_2[65039] = 32'b11111111111111101110110010001000;
assign LUT_2[65040] = 32'b11111111111111101110010101111000;
assign LUT_2[65041] = 32'b11111111111111101011001110010001;
assign LUT_2[65042] = 32'b11111111111111110101001110110100;
assign LUT_2[65043] = 32'b11111111111111110010000111001101;
assign LUT_2[65044] = 32'b11111111111111101010110011100000;
assign LUT_2[65045] = 32'b11111111111111100111101011111001;
assign LUT_2[65046] = 32'b11111111111111110001101100011100;
assign LUT_2[65047] = 32'b11111111111111101110100100110101;
assign LUT_2[65048] = 32'b11111111111111101001000111010101;
assign LUT_2[65049] = 32'b11111111111111100101111111101110;
assign LUT_2[65050] = 32'b11111111111111110000000000010001;
assign LUT_2[65051] = 32'b11111111111111101100111000101010;
assign LUT_2[65052] = 32'b11111111111111100101100100111101;
assign LUT_2[65053] = 32'b11111111111111100010011101010110;
assign LUT_2[65054] = 32'b11111111111111101100011101111001;
assign LUT_2[65055] = 32'b11111111111111101001010110010010;
assign LUT_2[65056] = 32'b11111111111111110100001101010111;
assign LUT_2[65057] = 32'b11111111111111110001000101110000;
assign LUT_2[65058] = 32'b11111111111111111011000110010011;
assign LUT_2[65059] = 32'b11111111111111110111111110101100;
assign LUT_2[65060] = 32'b11111111111111110000101010111111;
assign LUT_2[65061] = 32'b11111111111111101101100011011000;
assign LUT_2[65062] = 32'b11111111111111110111100011111011;
assign LUT_2[65063] = 32'b11111111111111110100011100010100;
assign LUT_2[65064] = 32'b11111111111111101110111110110100;
assign LUT_2[65065] = 32'b11111111111111101011110111001101;
assign LUT_2[65066] = 32'b11111111111111110101110111110000;
assign LUT_2[65067] = 32'b11111111111111110010110000001001;
assign LUT_2[65068] = 32'b11111111111111101011011100011100;
assign LUT_2[65069] = 32'b11111111111111101000010100110101;
assign LUT_2[65070] = 32'b11111111111111110010010101011000;
assign LUT_2[65071] = 32'b11111111111111101111001101110001;
assign LUT_2[65072] = 32'b11111111111111101110110001100001;
assign LUT_2[65073] = 32'b11111111111111101011101001111010;
assign LUT_2[65074] = 32'b11111111111111110101101010011101;
assign LUT_2[65075] = 32'b11111111111111110010100010110110;
assign LUT_2[65076] = 32'b11111111111111101011001111001001;
assign LUT_2[65077] = 32'b11111111111111101000000111100010;
assign LUT_2[65078] = 32'b11111111111111110010001000000101;
assign LUT_2[65079] = 32'b11111111111111101111000000011110;
assign LUT_2[65080] = 32'b11111111111111101001100010111110;
assign LUT_2[65081] = 32'b11111111111111100110011011010111;
assign LUT_2[65082] = 32'b11111111111111110000011011111010;
assign LUT_2[65083] = 32'b11111111111111101101010100010011;
assign LUT_2[65084] = 32'b11111111111111100110000000100110;
assign LUT_2[65085] = 32'b11111111111111100010111000111111;
assign LUT_2[65086] = 32'b11111111111111101100111001100010;
assign LUT_2[65087] = 32'b11111111111111101001110001111011;
assign LUT_2[65088] = 32'b11111111111111101011111010010001;
assign LUT_2[65089] = 32'b11111111111111101000110010101010;
assign LUT_2[65090] = 32'b11111111111111110010110011001101;
assign LUT_2[65091] = 32'b11111111111111101111101011100110;
assign LUT_2[65092] = 32'b11111111111111101000010111111001;
assign LUT_2[65093] = 32'b11111111111111100101010000010010;
assign LUT_2[65094] = 32'b11111111111111101111010000110101;
assign LUT_2[65095] = 32'b11111111111111101100001001001110;
assign LUT_2[65096] = 32'b11111111111111100110101011101110;
assign LUT_2[65097] = 32'b11111111111111100011100100000111;
assign LUT_2[65098] = 32'b11111111111111101101100100101010;
assign LUT_2[65099] = 32'b11111111111111101010011101000011;
assign LUT_2[65100] = 32'b11111111111111100011001001010110;
assign LUT_2[65101] = 32'b11111111111111100000000001101111;
assign LUT_2[65102] = 32'b11111111111111101010000010010010;
assign LUT_2[65103] = 32'b11111111111111100110111010101011;
assign LUT_2[65104] = 32'b11111111111111100110011110011011;
assign LUT_2[65105] = 32'b11111111111111100011010110110100;
assign LUT_2[65106] = 32'b11111111111111101101010111010111;
assign LUT_2[65107] = 32'b11111111111111101010001111110000;
assign LUT_2[65108] = 32'b11111111111111100010111100000011;
assign LUT_2[65109] = 32'b11111111111111011111110100011100;
assign LUT_2[65110] = 32'b11111111111111101001110100111111;
assign LUT_2[65111] = 32'b11111111111111100110101101011000;
assign LUT_2[65112] = 32'b11111111111111100001001111111000;
assign LUT_2[65113] = 32'b11111111111111011110001000010001;
assign LUT_2[65114] = 32'b11111111111111101000001000110100;
assign LUT_2[65115] = 32'b11111111111111100101000001001101;
assign LUT_2[65116] = 32'b11111111111111011101101101100000;
assign LUT_2[65117] = 32'b11111111111111011010100101111001;
assign LUT_2[65118] = 32'b11111111111111100100100110011100;
assign LUT_2[65119] = 32'b11111111111111100001011110110101;
assign LUT_2[65120] = 32'b11111111111111101100010101111010;
assign LUT_2[65121] = 32'b11111111111111101001001110010011;
assign LUT_2[65122] = 32'b11111111111111110011001110110110;
assign LUT_2[65123] = 32'b11111111111111110000000111001111;
assign LUT_2[65124] = 32'b11111111111111101000110011100010;
assign LUT_2[65125] = 32'b11111111111111100101101011111011;
assign LUT_2[65126] = 32'b11111111111111101111101100011110;
assign LUT_2[65127] = 32'b11111111111111101100100100110111;
assign LUT_2[65128] = 32'b11111111111111100111000111010111;
assign LUT_2[65129] = 32'b11111111111111100011111111110000;
assign LUT_2[65130] = 32'b11111111111111101110000000010011;
assign LUT_2[65131] = 32'b11111111111111101010111000101100;
assign LUT_2[65132] = 32'b11111111111111100011100100111111;
assign LUT_2[65133] = 32'b11111111111111100000011101011000;
assign LUT_2[65134] = 32'b11111111111111101010011101111011;
assign LUT_2[65135] = 32'b11111111111111100111010110010100;
assign LUT_2[65136] = 32'b11111111111111100110111010000100;
assign LUT_2[65137] = 32'b11111111111111100011110010011101;
assign LUT_2[65138] = 32'b11111111111111101101110011000000;
assign LUT_2[65139] = 32'b11111111111111101010101011011001;
assign LUT_2[65140] = 32'b11111111111111100011010111101100;
assign LUT_2[65141] = 32'b11111111111111100000010000000101;
assign LUT_2[65142] = 32'b11111111111111101010010000101000;
assign LUT_2[65143] = 32'b11111111111111100111001001000001;
assign LUT_2[65144] = 32'b11111111111111100001101011100001;
assign LUT_2[65145] = 32'b11111111111111011110100011111010;
assign LUT_2[65146] = 32'b11111111111111101000100100011101;
assign LUT_2[65147] = 32'b11111111111111100101011100110110;
assign LUT_2[65148] = 32'b11111111111111011110001001001001;
assign LUT_2[65149] = 32'b11111111111111011011000001100010;
assign LUT_2[65150] = 32'b11111111111111100101000010000101;
assign LUT_2[65151] = 32'b11111111111111100001111010011110;
assign LUT_2[65152] = 32'b11111111111111111000000101111101;
assign LUT_2[65153] = 32'b11111111111111110100111110010110;
assign LUT_2[65154] = 32'b11111111111111111110111110111001;
assign LUT_2[65155] = 32'b11111111111111111011110111010010;
assign LUT_2[65156] = 32'b11111111111111110100100011100101;
assign LUT_2[65157] = 32'b11111111111111110001011011111110;
assign LUT_2[65158] = 32'b11111111111111111011011100100001;
assign LUT_2[65159] = 32'b11111111111111111000010100111010;
assign LUT_2[65160] = 32'b11111111111111110010110111011010;
assign LUT_2[65161] = 32'b11111111111111101111101111110011;
assign LUT_2[65162] = 32'b11111111111111111001110000010110;
assign LUT_2[65163] = 32'b11111111111111110110101000101111;
assign LUT_2[65164] = 32'b11111111111111101111010101000010;
assign LUT_2[65165] = 32'b11111111111111101100001101011011;
assign LUT_2[65166] = 32'b11111111111111110110001101111110;
assign LUT_2[65167] = 32'b11111111111111110011000110010111;
assign LUT_2[65168] = 32'b11111111111111110010101010000111;
assign LUT_2[65169] = 32'b11111111111111101111100010100000;
assign LUT_2[65170] = 32'b11111111111111111001100011000011;
assign LUT_2[65171] = 32'b11111111111111110110011011011100;
assign LUT_2[65172] = 32'b11111111111111101111000111101111;
assign LUT_2[65173] = 32'b11111111111111101100000000001000;
assign LUT_2[65174] = 32'b11111111111111110110000000101011;
assign LUT_2[65175] = 32'b11111111111111110010111001000100;
assign LUT_2[65176] = 32'b11111111111111101101011011100100;
assign LUT_2[65177] = 32'b11111111111111101010010011111101;
assign LUT_2[65178] = 32'b11111111111111110100010100100000;
assign LUT_2[65179] = 32'b11111111111111110001001100111001;
assign LUT_2[65180] = 32'b11111111111111101001111001001100;
assign LUT_2[65181] = 32'b11111111111111100110110001100101;
assign LUT_2[65182] = 32'b11111111111111110000110010001000;
assign LUT_2[65183] = 32'b11111111111111101101101010100001;
assign LUT_2[65184] = 32'b11111111111111111000100001100110;
assign LUT_2[65185] = 32'b11111111111111110101011001111111;
assign LUT_2[65186] = 32'b11111111111111111111011010100010;
assign LUT_2[65187] = 32'b11111111111111111100010010111011;
assign LUT_2[65188] = 32'b11111111111111110100111111001110;
assign LUT_2[65189] = 32'b11111111111111110001110111100111;
assign LUT_2[65190] = 32'b11111111111111111011111000001010;
assign LUT_2[65191] = 32'b11111111111111111000110000100011;
assign LUT_2[65192] = 32'b11111111111111110011010011000011;
assign LUT_2[65193] = 32'b11111111111111110000001011011100;
assign LUT_2[65194] = 32'b11111111111111111010001011111111;
assign LUT_2[65195] = 32'b11111111111111110111000100011000;
assign LUT_2[65196] = 32'b11111111111111101111110000101011;
assign LUT_2[65197] = 32'b11111111111111101100101001000100;
assign LUT_2[65198] = 32'b11111111111111110110101001100111;
assign LUT_2[65199] = 32'b11111111111111110011100010000000;
assign LUT_2[65200] = 32'b11111111111111110011000101110000;
assign LUT_2[65201] = 32'b11111111111111101111111110001001;
assign LUT_2[65202] = 32'b11111111111111111001111110101100;
assign LUT_2[65203] = 32'b11111111111111110110110111000101;
assign LUT_2[65204] = 32'b11111111111111101111100011011000;
assign LUT_2[65205] = 32'b11111111111111101100011011110001;
assign LUT_2[65206] = 32'b11111111111111110110011100010100;
assign LUT_2[65207] = 32'b11111111111111110011010100101101;
assign LUT_2[65208] = 32'b11111111111111101101110111001101;
assign LUT_2[65209] = 32'b11111111111111101010101111100110;
assign LUT_2[65210] = 32'b11111111111111110100110000001001;
assign LUT_2[65211] = 32'b11111111111111110001101000100010;
assign LUT_2[65212] = 32'b11111111111111101010010100110101;
assign LUT_2[65213] = 32'b11111111111111100111001101001110;
assign LUT_2[65214] = 32'b11111111111111110001001101110001;
assign LUT_2[65215] = 32'b11111111111111101110000110001010;
assign LUT_2[65216] = 32'b11111111111111110000001110100000;
assign LUT_2[65217] = 32'b11111111111111101101000110111001;
assign LUT_2[65218] = 32'b11111111111111110111000111011100;
assign LUT_2[65219] = 32'b11111111111111110011111111110101;
assign LUT_2[65220] = 32'b11111111111111101100101100001000;
assign LUT_2[65221] = 32'b11111111111111101001100100100001;
assign LUT_2[65222] = 32'b11111111111111110011100101000100;
assign LUT_2[65223] = 32'b11111111111111110000011101011101;
assign LUT_2[65224] = 32'b11111111111111101010111111111101;
assign LUT_2[65225] = 32'b11111111111111100111111000010110;
assign LUT_2[65226] = 32'b11111111111111110001111000111001;
assign LUT_2[65227] = 32'b11111111111111101110110001010010;
assign LUT_2[65228] = 32'b11111111111111100111011101100101;
assign LUT_2[65229] = 32'b11111111111111100100010101111110;
assign LUT_2[65230] = 32'b11111111111111101110010110100001;
assign LUT_2[65231] = 32'b11111111111111101011001110111010;
assign LUT_2[65232] = 32'b11111111111111101010110010101010;
assign LUT_2[65233] = 32'b11111111111111100111101011000011;
assign LUT_2[65234] = 32'b11111111111111110001101011100110;
assign LUT_2[65235] = 32'b11111111111111101110100011111111;
assign LUT_2[65236] = 32'b11111111111111100111010000010010;
assign LUT_2[65237] = 32'b11111111111111100100001000101011;
assign LUT_2[65238] = 32'b11111111111111101110001001001110;
assign LUT_2[65239] = 32'b11111111111111101011000001100111;
assign LUT_2[65240] = 32'b11111111111111100101100100000111;
assign LUT_2[65241] = 32'b11111111111111100010011100100000;
assign LUT_2[65242] = 32'b11111111111111101100011101000011;
assign LUT_2[65243] = 32'b11111111111111101001010101011100;
assign LUT_2[65244] = 32'b11111111111111100010000001101111;
assign LUT_2[65245] = 32'b11111111111111011110111010001000;
assign LUT_2[65246] = 32'b11111111111111101000111010101011;
assign LUT_2[65247] = 32'b11111111111111100101110011000100;
assign LUT_2[65248] = 32'b11111111111111110000101010001001;
assign LUT_2[65249] = 32'b11111111111111101101100010100010;
assign LUT_2[65250] = 32'b11111111111111110111100011000101;
assign LUT_2[65251] = 32'b11111111111111110100011011011110;
assign LUT_2[65252] = 32'b11111111111111101101000111110001;
assign LUT_2[65253] = 32'b11111111111111101010000000001010;
assign LUT_2[65254] = 32'b11111111111111110100000000101101;
assign LUT_2[65255] = 32'b11111111111111110000111001000110;
assign LUT_2[65256] = 32'b11111111111111101011011011100110;
assign LUT_2[65257] = 32'b11111111111111101000010011111111;
assign LUT_2[65258] = 32'b11111111111111110010010100100010;
assign LUT_2[65259] = 32'b11111111111111101111001100111011;
assign LUT_2[65260] = 32'b11111111111111100111111001001110;
assign LUT_2[65261] = 32'b11111111111111100100110001100111;
assign LUT_2[65262] = 32'b11111111111111101110110010001010;
assign LUT_2[65263] = 32'b11111111111111101011101010100011;
assign LUT_2[65264] = 32'b11111111111111101011001110010011;
assign LUT_2[65265] = 32'b11111111111111101000000110101100;
assign LUT_2[65266] = 32'b11111111111111110010000111001111;
assign LUT_2[65267] = 32'b11111111111111101110111111101000;
assign LUT_2[65268] = 32'b11111111111111100111101011111011;
assign LUT_2[65269] = 32'b11111111111111100100100100010100;
assign LUT_2[65270] = 32'b11111111111111101110100100110111;
assign LUT_2[65271] = 32'b11111111111111101011011101010000;
assign LUT_2[65272] = 32'b11111111111111100101111111110000;
assign LUT_2[65273] = 32'b11111111111111100010111000001001;
assign LUT_2[65274] = 32'b11111111111111101100111000101100;
assign LUT_2[65275] = 32'b11111111111111101001110001000101;
assign LUT_2[65276] = 32'b11111111111111100010011101011000;
assign LUT_2[65277] = 32'b11111111111111011111010101110001;
assign LUT_2[65278] = 32'b11111111111111101001010110010100;
assign LUT_2[65279] = 32'b11111111111111100110001110101101;
assign LUT_2[65280] = 32'b11111111111111110111110000010100;
assign LUT_2[65281] = 32'b11111111111111110100101000101101;
assign LUT_2[65282] = 32'b11111111111111111110101001010000;
assign LUT_2[65283] = 32'b11111111111111111011100001101001;
assign LUT_2[65284] = 32'b11111111111111110100001101111100;
assign LUT_2[65285] = 32'b11111111111111110001000110010101;
assign LUT_2[65286] = 32'b11111111111111111011000110111000;
assign LUT_2[65287] = 32'b11111111111111110111111111010001;
assign LUT_2[65288] = 32'b11111111111111110010100001110001;
assign LUT_2[65289] = 32'b11111111111111101111011010001010;
assign LUT_2[65290] = 32'b11111111111111111001011010101101;
assign LUT_2[65291] = 32'b11111111111111110110010011000110;
assign LUT_2[65292] = 32'b11111111111111101110111111011001;
assign LUT_2[65293] = 32'b11111111111111101011110111110010;
assign LUT_2[65294] = 32'b11111111111111110101111000010101;
assign LUT_2[65295] = 32'b11111111111111110010110000101110;
assign LUT_2[65296] = 32'b11111111111111110010010100011110;
assign LUT_2[65297] = 32'b11111111111111101111001100110111;
assign LUT_2[65298] = 32'b11111111111111111001001101011010;
assign LUT_2[65299] = 32'b11111111111111110110000101110011;
assign LUT_2[65300] = 32'b11111111111111101110110010000110;
assign LUT_2[65301] = 32'b11111111111111101011101010011111;
assign LUT_2[65302] = 32'b11111111111111110101101011000010;
assign LUT_2[65303] = 32'b11111111111111110010100011011011;
assign LUT_2[65304] = 32'b11111111111111101101000101111011;
assign LUT_2[65305] = 32'b11111111111111101001111110010100;
assign LUT_2[65306] = 32'b11111111111111110011111110110111;
assign LUT_2[65307] = 32'b11111111111111110000110111010000;
assign LUT_2[65308] = 32'b11111111111111101001100011100011;
assign LUT_2[65309] = 32'b11111111111111100110011011111100;
assign LUT_2[65310] = 32'b11111111111111110000011100011111;
assign LUT_2[65311] = 32'b11111111111111101101010100111000;
assign LUT_2[65312] = 32'b11111111111111111000001011111101;
assign LUT_2[65313] = 32'b11111111111111110101000100010110;
assign LUT_2[65314] = 32'b11111111111111111111000100111001;
assign LUT_2[65315] = 32'b11111111111111111011111101010010;
assign LUT_2[65316] = 32'b11111111111111110100101001100101;
assign LUT_2[65317] = 32'b11111111111111110001100001111110;
assign LUT_2[65318] = 32'b11111111111111111011100010100001;
assign LUT_2[65319] = 32'b11111111111111111000011010111010;
assign LUT_2[65320] = 32'b11111111111111110010111101011010;
assign LUT_2[65321] = 32'b11111111111111101111110101110011;
assign LUT_2[65322] = 32'b11111111111111111001110110010110;
assign LUT_2[65323] = 32'b11111111111111110110101110101111;
assign LUT_2[65324] = 32'b11111111111111101111011011000010;
assign LUT_2[65325] = 32'b11111111111111101100010011011011;
assign LUT_2[65326] = 32'b11111111111111110110010011111110;
assign LUT_2[65327] = 32'b11111111111111110011001100010111;
assign LUT_2[65328] = 32'b11111111111111110010110000000111;
assign LUT_2[65329] = 32'b11111111111111101111101000100000;
assign LUT_2[65330] = 32'b11111111111111111001101001000011;
assign LUT_2[65331] = 32'b11111111111111110110100001011100;
assign LUT_2[65332] = 32'b11111111111111101111001101101111;
assign LUT_2[65333] = 32'b11111111111111101100000110001000;
assign LUT_2[65334] = 32'b11111111111111110110000110101011;
assign LUT_2[65335] = 32'b11111111111111110010111111000100;
assign LUT_2[65336] = 32'b11111111111111101101100001100100;
assign LUT_2[65337] = 32'b11111111111111101010011001111101;
assign LUT_2[65338] = 32'b11111111111111110100011010100000;
assign LUT_2[65339] = 32'b11111111111111110001010010111001;
assign LUT_2[65340] = 32'b11111111111111101001111111001100;
assign LUT_2[65341] = 32'b11111111111111100110110111100101;
assign LUT_2[65342] = 32'b11111111111111110000111000001000;
assign LUT_2[65343] = 32'b11111111111111101101110000100001;
assign LUT_2[65344] = 32'b11111111111111101111111000110111;
assign LUT_2[65345] = 32'b11111111111111101100110001010000;
assign LUT_2[65346] = 32'b11111111111111110110110001110011;
assign LUT_2[65347] = 32'b11111111111111110011101010001100;
assign LUT_2[65348] = 32'b11111111111111101100010110011111;
assign LUT_2[65349] = 32'b11111111111111101001001110111000;
assign LUT_2[65350] = 32'b11111111111111110011001111011011;
assign LUT_2[65351] = 32'b11111111111111110000000111110100;
assign LUT_2[65352] = 32'b11111111111111101010101010010100;
assign LUT_2[65353] = 32'b11111111111111100111100010101101;
assign LUT_2[65354] = 32'b11111111111111110001100011010000;
assign LUT_2[65355] = 32'b11111111111111101110011011101001;
assign LUT_2[65356] = 32'b11111111111111100111000111111100;
assign LUT_2[65357] = 32'b11111111111111100100000000010101;
assign LUT_2[65358] = 32'b11111111111111101110000000111000;
assign LUT_2[65359] = 32'b11111111111111101010111001010001;
assign LUT_2[65360] = 32'b11111111111111101010011101000001;
assign LUT_2[65361] = 32'b11111111111111100111010101011010;
assign LUT_2[65362] = 32'b11111111111111110001010101111101;
assign LUT_2[65363] = 32'b11111111111111101110001110010110;
assign LUT_2[65364] = 32'b11111111111111100110111010101001;
assign LUT_2[65365] = 32'b11111111111111100011110011000010;
assign LUT_2[65366] = 32'b11111111111111101101110011100101;
assign LUT_2[65367] = 32'b11111111111111101010101011111110;
assign LUT_2[65368] = 32'b11111111111111100101001110011110;
assign LUT_2[65369] = 32'b11111111111111100010000110110111;
assign LUT_2[65370] = 32'b11111111111111101100000111011010;
assign LUT_2[65371] = 32'b11111111111111101000111111110011;
assign LUT_2[65372] = 32'b11111111111111100001101100000110;
assign LUT_2[65373] = 32'b11111111111111011110100100011111;
assign LUT_2[65374] = 32'b11111111111111101000100101000010;
assign LUT_2[65375] = 32'b11111111111111100101011101011011;
assign LUT_2[65376] = 32'b11111111111111110000010100100000;
assign LUT_2[65377] = 32'b11111111111111101101001100111001;
assign LUT_2[65378] = 32'b11111111111111110111001101011100;
assign LUT_2[65379] = 32'b11111111111111110100000101110101;
assign LUT_2[65380] = 32'b11111111111111101100110010001000;
assign LUT_2[65381] = 32'b11111111111111101001101010100001;
assign LUT_2[65382] = 32'b11111111111111110011101011000100;
assign LUT_2[65383] = 32'b11111111111111110000100011011101;
assign LUT_2[65384] = 32'b11111111111111101011000101111101;
assign LUT_2[65385] = 32'b11111111111111100111111110010110;
assign LUT_2[65386] = 32'b11111111111111110001111110111001;
assign LUT_2[65387] = 32'b11111111111111101110110111010010;
assign LUT_2[65388] = 32'b11111111111111100111100011100101;
assign LUT_2[65389] = 32'b11111111111111100100011011111110;
assign LUT_2[65390] = 32'b11111111111111101110011100100001;
assign LUT_2[65391] = 32'b11111111111111101011010100111010;
assign LUT_2[65392] = 32'b11111111111111101010111000101010;
assign LUT_2[65393] = 32'b11111111111111100111110001000011;
assign LUT_2[65394] = 32'b11111111111111110001110001100110;
assign LUT_2[65395] = 32'b11111111111111101110101001111111;
assign LUT_2[65396] = 32'b11111111111111100111010110010010;
assign LUT_2[65397] = 32'b11111111111111100100001110101011;
assign LUT_2[65398] = 32'b11111111111111101110001111001110;
assign LUT_2[65399] = 32'b11111111111111101011000111100111;
assign LUT_2[65400] = 32'b11111111111111100101101010000111;
assign LUT_2[65401] = 32'b11111111111111100010100010100000;
assign LUT_2[65402] = 32'b11111111111111101100100011000011;
assign LUT_2[65403] = 32'b11111111111111101001011011011100;
assign LUT_2[65404] = 32'b11111111111111100010000111101111;
assign LUT_2[65405] = 32'b11111111111111011111000000001000;
assign LUT_2[65406] = 32'b11111111111111101001000000101011;
assign LUT_2[65407] = 32'b11111111111111100101111001000100;
assign LUT_2[65408] = 32'b11111111111111111100000100100011;
assign LUT_2[65409] = 32'b11111111111111111000111100111100;
assign LUT_2[65410] = 32'b00000000000000000010111101011111;
assign LUT_2[65411] = 32'b11111111111111111111110101111000;
assign LUT_2[65412] = 32'b11111111111111111000100010001011;
assign LUT_2[65413] = 32'b11111111111111110101011010100100;
assign LUT_2[65414] = 32'b11111111111111111111011011000111;
assign LUT_2[65415] = 32'b11111111111111111100010011100000;
assign LUT_2[65416] = 32'b11111111111111110110110110000000;
assign LUT_2[65417] = 32'b11111111111111110011101110011001;
assign LUT_2[65418] = 32'b11111111111111111101101110111100;
assign LUT_2[65419] = 32'b11111111111111111010100111010101;
assign LUT_2[65420] = 32'b11111111111111110011010011101000;
assign LUT_2[65421] = 32'b11111111111111110000001100000001;
assign LUT_2[65422] = 32'b11111111111111111010001100100100;
assign LUT_2[65423] = 32'b11111111111111110111000100111101;
assign LUT_2[65424] = 32'b11111111111111110110101000101101;
assign LUT_2[65425] = 32'b11111111111111110011100001000110;
assign LUT_2[65426] = 32'b11111111111111111101100001101001;
assign LUT_2[65427] = 32'b11111111111111111010011010000010;
assign LUT_2[65428] = 32'b11111111111111110011000110010101;
assign LUT_2[65429] = 32'b11111111111111101111111110101110;
assign LUT_2[65430] = 32'b11111111111111111001111111010001;
assign LUT_2[65431] = 32'b11111111111111110110110111101010;
assign LUT_2[65432] = 32'b11111111111111110001011010001010;
assign LUT_2[65433] = 32'b11111111111111101110010010100011;
assign LUT_2[65434] = 32'b11111111111111111000010011000110;
assign LUT_2[65435] = 32'b11111111111111110101001011011111;
assign LUT_2[65436] = 32'b11111111111111101101110111110010;
assign LUT_2[65437] = 32'b11111111111111101010110000001011;
assign LUT_2[65438] = 32'b11111111111111110100110000101110;
assign LUT_2[65439] = 32'b11111111111111110001101001000111;
assign LUT_2[65440] = 32'b11111111111111111100100000001100;
assign LUT_2[65441] = 32'b11111111111111111001011000100101;
assign LUT_2[65442] = 32'b00000000000000000011011001001000;
assign LUT_2[65443] = 32'b00000000000000000000010001100001;
assign LUT_2[65444] = 32'b11111111111111111000111101110100;
assign LUT_2[65445] = 32'b11111111111111110101110110001101;
assign LUT_2[65446] = 32'b11111111111111111111110110110000;
assign LUT_2[65447] = 32'b11111111111111111100101111001001;
assign LUT_2[65448] = 32'b11111111111111110111010001101001;
assign LUT_2[65449] = 32'b11111111111111110100001010000010;
assign LUT_2[65450] = 32'b11111111111111111110001010100101;
assign LUT_2[65451] = 32'b11111111111111111011000010111110;
assign LUT_2[65452] = 32'b11111111111111110011101111010001;
assign LUT_2[65453] = 32'b11111111111111110000100111101010;
assign LUT_2[65454] = 32'b11111111111111111010101000001101;
assign LUT_2[65455] = 32'b11111111111111110111100000100110;
assign LUT_2[65456] = 32'b11111111111111110111000100010110;
assign LUT_2[65457] = 32'b11111111111111110011111100101111;
assign LUT_2[65458] = 32'b11111111111111111101111101010010;
assign LUT_2[65459] = 32'b11111111111111111010110101101011;
assign LUT_2[65460] = 32'b11111111111111110011100001111110;
assign LUT_2[65461] = 32'b11111111111111110000011010010111;
assign LUT_2[65462] = 32'b11111111111111111010011010111010;
assign LUT_2[65463] = 32'b11111111111111110111010011010011;
assign LUT_2[65464] = 32'b11111111111111110001110101110011;
assign LUT_2[65465] = 32'b11111111111111101110101110001100;
assign LUT_2[65466] = 32'b11111111111111111000101110101111;
assign LUT_2[65467] = 32'b11111111111111110101100111001000;
assign LUT_2[65468] = 32'b11111111111111101110010011011011;
assign LUT_2[65469] = 32'b11111111111111101011001011110100;
assign LUT_2[65470] = 32'b11111111111111110101001100010111;
assign LUT_2[65471] = 32'b11111111111111110010000100110000;
assign LUT_2[65472] = 32'b11111111111111110100001101000110;
assign LUT_2[65473] = 32'b11111111111111110001000101011111;
assign LUT_2[65474] = 32'b11111111111111111011000110000010;
assign LUT_2[65475] = 32'b11111111111111110111111110011011;
assign LUT_2[65476] = 32'b11111111111111110000101010101110;
assign LUT_2[65477] = 32'b11111111111111101101100011000111;
assign LUT_2[65478] = 32'b11111111111111110111100011101010;
assign LUT_2[65479] = 32'b11111111111111110100011100000011;
assign LUT_2[65480] = 32'b11111111111111101110111110100011;
assign LUT_2[65481] = 32'b11111111111111101011110110111100;
assign LUT_2[65482] = 32'b11111111111111110101110111011111;
assign LUT_2[65483] = 32'b11111111111111110010101111111000;
assign LUT_2[65484] = 32'b11111111111111101011011100001011;
assign LUT_2[65485] = 32'b11111111111111101000010100100100;
assign LUT_2[65486] = 32'b11111111111111110010010101000111;
assign LUT_2[65487] = 32'b11111111111111101111001101100000;
assign LUT_2[65488] = 32'b11111111111111101110110001010000;
assign LUT_2[65489] = 32'b11111111111111101011101001101001;
assign LUT_2[65490] = 32'b11111111111111110101101010001100;
assign LUT_2[65491] = 32'b11111111111111110010100010100101;
assign LUT_2[65492] = 32'b11111111111111101011001110111000;
assign LUT_2[65493] = 32'b11111111111111101000000111010001;
assign LUT_2[65494] = 32'b11111111111111110010000111110100;
assign LUT_2[65495] = 32'b11111111111111101111000000001101;
assign LUT_2[65496] = 32'b11111111111111101001100010101101;
assign LUT_2[65497] = 32'b11111111111111100110011011000110;
assign LUT_2[65498] = 32'b11111111111111110000011011101001;
assign LUT_2[65499] = 32'b11111111111111101101010100000010;
assign LUT_2[65500] = 32'b11111111111111100110000000010101;
assign LUT_2[65501] = 32'b11111111111111100010111000101110;
assign LUT_2[65502] = 32'b11111111111111101100111001010001;
assign LUT_2[65503] = 32'b11111111111111101001110001101010;
assign LUT_2[65504] = 32'b11111111111111110100101000101111;
assign LUT_2[65505] = 32'b11111111111111110001100001001000;
assign LUT_2[65506] = 32'b11111111111111111011100001101011;
assign LUT_2[65507] = 32'b11111111111111111000011010000100;
assign LUT_2[65508] = 32'b11111111111111110001000110010111;
assign LUT_2[65509] = 32'b11111111111111101101111110110000;
assign LUT_2[65510] = 32'b11111111111111110111111111010011;
assign LUT_2[65511] = 32'b11111111111111110100110111101100;
assign LUT_2[65512] = 32'b11111111111111101111011010001100;
assign LUT_2[65513] = 32'b11111111111111101100010010100101;
assign LUT_2[65514] = 32'b11111111111111110110010011001000;
assign LUT_2[65515] = 32'b11111111111111110011001011100001;
assign LUT_2[65516] = 32'b11111111111111101011110111110100;
assign LUT_2[65517] = 32'b11111111111111101000110000001101;
assign LUT_2[65518] = 32'b11111111111111110010110000110000;
assign LUT_2[65519] = 32'b11111111111111101111101001001001;
assign LUT_2[65520] = 32'b11111111111111101111001100111001;
assign LUT_2[65521] = 32'b11111111111111101100000101010010;
assign LUT_2[65522] = 32'b11111111111111110110000101110101;
assign LUT_2[65523] = 32'b11111111111111110010111110001110;
assign LUT_2[65524] = 32'b11111111111111101011101010100001;
assign LUT_2[65525] = 32'b11111111111111101000100010111010;
assign LUT_2[65526] = 32'b11111111111111110010100011011101;
assign LUT_2[65527] = 32'b11111111111111101111011011110110;
assign LUT_2[65528] = 32'b11111111111111101001111110010110;
assign LUT_2[65529] = 32'b11111111111111100110110110101111;
assign LUT_2[65530] = 32'b11111111111111110000110111010010;
assign LUT_2[65531] = 32'b11111111111111101101101111101011;
assign LUT_2[65532] = 32'b11111111111111100110011011111110;
assign LUT_2[65533] = 32'b11111111111111100011010100010111;
assign LUT_2[65534] = 32'b11111111111111101101010100111010;
assign LUT_2[65535] = 32'b11111111111111101010001101010011;
endmodule
