module DA_table_4(table_in_4 , table_out_4);
input unsigned [15:0]table_in_4;
output [31:0]table_out_4;
wire  [31:0]LUT_4[65535:0]; 
wire [31:0]table_out_4; 
assign table_out_4 = LUT_4[table_in_4];
assign LUT_4[0] = 32'b00000000000000000000000000000000;
assign LUT_4[1] = 32'b11111111111111111001001011111000;
assign LUT_4[2] = 32'b11111111111111111111011010100100;
assign LUT_4[3] = 32'b11111111111111111000100110011100;
assign LUT_4[4] = 32'b11111111111111111101000000011100;
assign LUT_4[5] = 32'b11111111111111110110001100010100;
assign LUT_4[6] = 32'b11111111111111111100011011000000;
assign LUT_4[7] = 32'b11111111111111110101100110111000;
assign LUT_4[8] = 32'b11111111111111111001001100010101;
assign LUT_4[9] = 32'b11111111111111110010011000001101;
assign LUT_4[10] = 32'b11111111111111111000100110111001;
assign LUT_4[11] = 32'b11111111111111110001110010110001;
assign LUT_4[12] = 32'b11111111111111110110001100110001;
assign LUT_4[13] = 32'b11111111111111101111011000101001;
assign LUT_4[14] = 32'b11111111111111110101100111010101;
assign LUT_4[15] = 32'b11111111111111101110110011001101;
assign LUT_4[16] = 32'b11111111111111111101110001101110;
assign LUT_4[17] = 32'b11111111111111110110111101100110;
assign LUT_4[18] = 32'b11111111111111111101001100010010;
assign LUT_4[19] = 32'b11111111111111110110011000001010;
assign LUT_4[20] = 32'b11111111111111111010110010001010;
assign LUT_4[21] = 32'b11111111111111110011111110000010;
assign LUT_4[22] = 32'b11111111111111111010001100101110;
assign LUT_4[23] = 32'b11111111111111110011011000100110;
assign LUT_4[24] = 32'b11111111111111110110111110000011;
assign LUT_4[25] = 32'b11111111111111110000001001111011;
assign LUT_4[26] = 32'b11111111111111110110011000100111;
assign LUT_4[27] = 32'b11111111111111101111100100011111;
assign LUT_4[28] = 32'b11111111111111110011111110011111;
assign LUT_4[29] = 32'b11111111111111101101001010010111;
assign LUT_4[30] = 32'b11111111111111110011011001000011;
assign LUT_4[31] = 32'b11111111111111101100100100111011;
assign LUT_4[32] = 32'b11111111111111111110011011000111;
assign LUT_4[33] = 32'b11111111111111110111100110111111;
assign LUT_4[34] = 32'b11111111111111111101110101101011;
assign LUT_4[35] = 32'b11111111111111110111000001100011;
assign LUT_4[36] = 32'b11111111111111111011011011100011;
assign LUT_4[37] = 32'b11111111111111110100100111011011;
assign LUT_4[38] = 32'b11111111111111111010110110000111;
assign LUT_4[39] = 32'b11111111111111110100000001111111;
assign LUT_4[40] = 32'b11111111111111110111100111011100;
assign LUT_4[41] = 32'b11111111111111110000110011010100;
assign LUT_4[42] = 32'b11111111111111110111000010000000;
assign LUT_4[43] = 32'b11111111111111110000001101111000;
assign LUT_4[44] = 32'b11111111111111110100100111111000;
assign LUT_4[45] = 32'b11111111111111101101110011110000;
assign LUT_4[46] = 32'b11111111111111110100000010011100;
assign LUT_4[47] = 32'b11111111111111101101001110010100;
assign LUT_4[48] = 32'b11111111111111111100001100110101;
assign LUT_4[49] = 32'b11111111111111110101011000101101;
assign LUT_4[50] = 32'b11111111111111111011100111011001;
assign LUT_4[51] = 32'b11111111111111110100110011010001;
assign LUT_4[52] = 32'b11111111111111111001001101010001;
assign LUT_4[53] = 32'b11111111111111110010011001001001;
assign LUT_4[54] = 32'b11111111111111111000100111110101;
assign LUT_4[55] = 32'b11111111111111110001110011101101;
assign LUT_4[56] = 32'b11111111111111110101011001001010;
assign LUT_4[57] = 32'b11111111111111101110100101000010;
assign LUT_4[58] = 32'b11111111111111110100110011101110;
assign LUT_4[59] = 32'b11111111111111101101111111100110;
assign LUT_4[60] = 32'b11111111111111110010011001100110;
assign LUT_4[61] = 32'b11111111111111101011100101011110;
assign LUT_4[62] = 32'b11111111111111110001110100001010;
assign LUT_4[63] = 32'b11111111111111101011000000000010;
assign LUT_4[64] = 32'b00000000000000000001010111010100;
assign LUT_4[65] = 32'b11111111111111111010100011001100;
assign LUT_4[66] = 32'b00000000000000000000110001111000;
assign LUT_4[67] = 32'b11111111111111111001111101110000;
assign LUT_4[68] = 32'b11111111111111111110010111110000;
assign LUT_4[69] = 32'b11111111111111110111100011101000;
assign LUT_4[70] = 32'b11111111111111111101110010010100;
assign LUT_4[71] = 32'b11111111111111110110111110001100;
assign LUT_4[72] = 32'b11111111111111111010100011101001;
assign LUT_4[73] = 32'b11111111111111110011101111100001;
assign LUT_4[74] = 32'b11111111111111111001111110001101;
assign LUT_4[75] = 32'b11111111111111110011001010000101;
assign LUT_4[76] = 32'b11111111111111110111100100000101;
assign LUT_4[77] = 32'b11111111111111110000101111111101;
assign LUT_4[78] = 32'b11111111111111110110111110101001;
assign LUT_4[79] = 32'b11111111111111110000001010100001;
assign LUT_4[80] = 32'b11111111111111111111001001000010;
assign LUT_4[81] = 32'b11111111111111111000010100111010;
assign LUT_4[82] = 32'b11111111111111111110100011100110;
assign LUT_4[83] = 32'b11111111111111110111101111011110;
assign LUT_4[84] = 32'b11111111111111111100001001011110;
assign LUT_4[85] = 32'b11111111111111110101010101010110;
assign LUT_4[86] = 32'b11111111111111111011100100000010;
assign LUT_4[87] = 32'b11111111111111110100101111111010;
assign LUT_4[88] = 32'b11111111111111111000010101010111;
assign LUT_4[89] = 32'b11111111111111110001100001001111;
assign LUT_4[90] = 32'b11111111111111110111101111111011;
assign LUT_4[91] = 32'b11111111111111110000111011110011;
assign LUT_4[92] = 32'b11111111111111110101010101110011;
assign LUT_4[93] = 32'b11111111111111101110100001101011;
assign LUT_4[94] = 32'b11111111111111110100110000010111;
assign LUT_4[95] = 32'b11111111111111101101111100001111;
assign LUT_4[96] = 32'b11111111111111111111110010011011;
assign LUT_4[97] = 32'b11111111111111111000111110010011;
assign LUT_4[98] = 32'b11111111111111111111001100111111;
assign LUT_4[99] = 32'b11111111111111111000011000110111;
assign LUT_4[100] = 32'b11111111111111111100110010110111;
assign LUT_4[101] = 32'b11111111111111110101111110101111;
assign LUT_4[102] = 32'b11111111111111111100001101011011;
assign LUT_4[103] = 32'b11111111111111110101011001010011;
assign LUT_4[104] = 32'b11111111111111111000111110110000;
assign LUT_4[105] = 32'b11111111111111110010001010101000;
assign LUT_4[106] = 32'b11111111111111111000011001010100;
assign LUT_4[107] = 32'b11111111111111110001100101001100;
assign LUT_4[108] = 32'b11111111111111110101111111001100;
assign LUT_4[109] = 32'b11111111111111101111001011000100;
assign LUT_4[110] = 32'b11111111111111110101011001110000;
assign LUT_4[111] = 32'b11111111111111101110100101101000;
assign LUT_4[112] = 32'b11111111111111111101100100001001;
assign LUT_4[113] = 32'b11111111111111110110110000000001;
assign LUT_4[114] = 32'b11111111111111111100111110101101;
assign LUT_4[115] = 32'b11111111111111110110001010100101;
assign LUT_4[116] = 32'b11111111111111111010100100100101;
assign LUT_4[117] = 32'b11111111111111110011110000011101;
assign LUT_4[118] = 32'b11111111111111111001111111001001;
assign LUT_4[119] = 32'b11111111111111110011001011000001;
assign LUT_4[120] = 32'b11111111111111110110110000011110;
assign LUT_4[121] = 32'b11111111111111101111111100010110;
assign LUT_4[122] = 32'b11111111111111110110001011000010;
assign LUT_4[123] = 32'b11111111111111101111010110111010;
assign LUT_4[124] = 32'b11111111111111110011110000111010;
assign LUT_4[125] = 32'b11111111111111101100111100110010;
assign LUT_4[126] = 32'b11111111111111110011001011011110;
assign LUT_4[127] = 32'b11111111111111101100010111010110;
assign LUT_4[128] = 32'b00000000000000000010100110001000;
assign LUT_4[129] = 32'b11111111111111111011110010000000;
assign LUT_4[130] = 32'b00000000000000000010000000101100;
assign LUT_4[131] = 32'b11111111111111111011001100100100;
assign LUT_4[132] = 32'b11111111111111111111100110100100;
assign LUT_4[133] = 32'b11111111111111111000110010011100;
assign LUT_4[134] = 32'b11111111111111111111000001001000;
assign LUT_4[135] = 32'b11111111111111111000001101000000;
assign LUT_4[136] = 32'b11111111111111111011110010011101;
assign LUT_4[137] = 32'b11111111111111110100111110010101;
assign LUT_4[138] = 32'b11111111111111111011001101000001;
assign LUT_4[139] = 32'b11111111111111110100011000111001;
assign LUT_4[140] = 32'b11111111111111111000110010111001;
assign LUT_4[141] = 32'b11111111111111110001111110110001;
assign LUT_4[142] = 32'b11111111111111111000001101011101;
assign LUT_4[143] = 32'b11111111111111110001011001010101;
assign LUT_4[144] = 32'b00000000000000000000010111110110;
assign LUT_4[145] = 32'b11111111111111111001100011101110;
assign LUT_4[146] = 32'b11111111111111111111110010011010;
assign LUT_4[147] = 32'b11111111111111111000111110010010;
assign LUT_4[148] = 32'b11111111111111111101011000010010;
assign LUT_4[149] = 32'b11111111111111110110100100001010;
assign LUT_4[150] = 32'b11111111111111111100110010110110;
assign LUT_4[151] = 32'b11111111111111110101111110101110;
assign LUT_4[152] = 32'b11111111111111111001100100001011;
assign LUT_4[153] = 32'b11111111111111110010110000000011;
assign LUT_4[154] = 32'b11111111111111111000111110101111;
assign LUT_4[155] = 32'b11111111111111110010001010100111;
assign LUT_4[156] = 32'b11111111111111110110100100100111;
assign LUT_4[157] = 32'b11111111111111101111110000011111;
assign LUT_4[158] = 32'b11111111111111110101111111001011;
assign LUT_4[159] = 32'b11111111111111101111001011000011;
assign LUT_4[160] = 32'b00000000000000000001000001001111;
assign LUT_4[161] = 32'b11111111111111111010001101000111;
assign LUT_4[162] = 32'b00000000000000000000011011110011;
assign LUT_4[163] = 32'b11111111111111111001100111101011;
assign LUT_4[164] = 32'b11111111111111111110000001101011;
assign LUT_4[165] = 32'b11111111111111110111001101100011;
assign LUT_4[166] = 32'b11111111111111111101011100001111;
assign LUT_4[167] = 32'b11111111111111110110101000000111;
assign LUT_4[168] = 32'b11111111111111111010001101100100;
assign LUT_4[169] = 32'b11111111111111110011011001011100;
assign LUT_4[170] = 32'b11111111111111111001101000001000;
assign LUT_4[171] = 32'b11111111111111110010110100000000;
assign LUT_4[172] = 32'b11111111111111110111001110000000;
assign LUT_4[173] = 32'b11111111111111110000011001111000;
assign LUT_4[174] = 32'b11111111111111110110101000100100;
assign LUT_4[175] = 32'b11111111111111101111110100011100;
assign LUT_4[176] = 32'b11111111111111111110110010111101;
assign LUT_4[177] = 32'b11111111111111110111111110110101;
assign LUT_4[178] = 32'b11111111111111111110001101100001;
assign LUT_4[179] = 32'b11111111111111110111011001011001;
assign LUT_4[180] = 32'b11111111111111111011110011011001;
assign LUT_4[181] = 32'b11111111111111110100111111010001;
assign LUT_4[182] = 32'b11111111111111111011001101111101;
assign LUT_4[183] = 32'b11111111111111110100011001110101;
assign LUT_4[184] = 32'b11111111111111110111111111010010;
assign LUT_4[185] = 32'b11111111111111110001001011001010;
assign LUT_4[186] = 32'b11111111111111110111011001110110;
assign LUT_4[187] = 32'b11111111111111110000100101101110;
assign LUT_4[188] = 32'b11111111111111110100111111101110;
assign LUT_4[189] = 32'b11111111111111101110001011100110;
assign LUT_4[190] = 32'b11111111111111110100011010010010;
assign LUT_4[191] = 32'b11111111111111101101100110001010;
assign LUT_4[192] = 32'b00000000000000000011111101011100;
assign LUT_4[193] = 32'b11111111111111111101001001010100;
assign LUT_4[194] = 32'b00000000000000000011011000000000;
assign LUT_4[195] = 32'b11111111111111111100100011111000;
assign LUT_4[196] = 32'b00000000000000000000111101111000;
assign LUT_4[197] = 32'b11111111111111111010001001110000;
assign LUT_4[198] = 32'b00000000000000000000011000011100;
assign LUT_4[199] = 32'b11111111111111111001100100010100;
assign LUT_4[200] = 32'b11111111111111111101001001110001;
assign LUT_4[201] = 32'b11111111111111110110010101101001;
assign LUT_4[202] = 32'b11111111111111111100100100010101;
assign LUT_4[203] = 32'b11111111111111110101110000001101;
assign LUT_4[204] = 32'b11111111111111111010001010001101;
assign LUT_4[205] = 32'b11111111111111110011010110000101;
assign LUT_4[206] = 32'b11111111111111111001100100110001;
assign LUT_4[207] = 32'b11111111111111110010110000101001;
assign LUT_4[208] = 32'b00000000000000000001101111001010;
assign LUT_4[209] = 32'b11111111111111111010111011000010;
assign LUT_4[210] = 32'b00000000000000000001001001101110;
assign LUT_4[211] = 32'b11111111111111111010010101100110;
assign LUT_4[212] = 32'b11111111111111111110101111100110;
assign LUT_4[213] = 32'b11111111111111110111111011011110;
assign LUT_4[214] = 32'b11111111111111111110001010001010;
assign LUT_4[215] = 32'b11111111111111110111010110000010;
assign LUT_4[216] = 32'b11111111111111111010111011011111;
assign LUT_4[217] = 32'b11111111111111110100000111010111;
assign LUT_4[218] = 32'b11111111111111111010010110000011;
assign LUT_4[219] = 32'b11111111111111110011100001111011;
assign LUT_4[220] = 32'b11111111111111110111111011111011;
assign LUT_4[221] = 32'b11111111111111110001000111110011;
assign LUT_4[222] = 32'b11111111111111110111010110011111;
assign LUT_4[223] = 32'b11111111111111110000100010010111;
assign LUT_4[224] = 32'b00000000000000000010011000100011;
assign LUT_4[225] = 32'b11111111111111111011100100011011;
assign LUT_4[226] = 32'b00000000000000000001110011000111;
assign LUT_4[227] = 32'b11111111111111111010111110111111;
assign LUT_4[228] = 32'b11111111111111111111011000111111;
assign LUT_4[229] = 32'b11111111111111111000100100110111;
assign LUT_4[230] = 32'b11111111111111111110110011100011;
assign LUT_4[231] = 32'b11111111111111110111111111011011;
assign LUT_4[232] = 32'b11111111111111111011100100111000;
assign LUT_4[233] = 32'b11111111111111110100110000110000;
assign LUT_4[234] = 32'b11111111111111111010111111011100;
assign LUT_4[235] = 32'b11111111111111110100001011010100;
assign LUT_4[236] = 32'b11111111111111111000100101010100;
assign LUT_4[237] = 32'b11111111111111110001110001001100;
assign LUT_4[238] = 32'b11111111111111110111111111111000;
assign LUT_4[239] = 32'b11111111111111110001001011110000;
assign LUT_4[240] = 32'b00000000000000000000001010010001;
assign LUT_4[241] = 32'b11111111111111111001010110001001;
assign LUT_4[242] = 32'b11111111111111111111100100110101;
assign LUT_4[243] = 32'b11111111111111111000110000101101;
assign LUT_4[244] = 32'b11111111111111111101001010101101;
assign LUT_4[245] = 32'b11111111111111110110010110100101;
assign LUT_4[246] = 32'b11111111111111111100100101010001;
assign LUT_4[247] = 32'b11111111111111110101110001001001;
assign LUT_4[248] = 32'b11111111111111111001010110100110;
assign LUT_4[249] = 32'b11111111111111110010100010011110;
assign LUT_4[250] = 32'b11111111111111111000110001001010;
assign LUT_4[251] = 32'b11111111111111110001111101000010;
assign LUT_4[252] = 32'b11111111111111110110010111000010;
assign LUT_4[253] = 32'b11111111111111101111100010111010;
assign LUT_4[254] = 32'b11111111111111110101110001100110;
assign LUT_4[255] = 32'b11111111111111101110111101011110;
assign LUT_4[256] = 32'b00000000000000000100111011100011;
assign LUT_4[257] = 32'b11111111111111111110000111011011;
assign LUT_4[258] = 32'b00000000000000000100010110000111;
assign LUT_4[259] = 32'b11111111111111111101100001111111;
assign LUT_4[260] = 32'b00000000000000000001111011111111;
assign LUT_4[261] = 32'b11111111111111111011000111110111;
assign LUT_4[262] = 32'b00000000000000000001010110100011;
assign LUT_4[263] = 32'b11111111111111111010100010011011;
assign LUT_4[264] = 32'b11111111111111111110000111111000;
assign LUT_4[265] = 32'b11111111111111110111010011110000;
assign LUT_4[266] = 32'b11111111111111111101100010011100;
assign LUT_4[267] = 32'b11111111111111110110101110010100;
assign LUT_4[268] = 32'b11111111111111111011001000010100;
assign LUT_4[269] = 32'b11111111111111110100010100001100;
assign LUT_4[270] = 32'b11111111111111111010100010111000;
assign LUT_4[271] = 32'b11111111111111110011101110110000;
assign LUT_4[272] = 32'b00000000000000000010101101010001;
assign LUT_4[273] = 32'b11111111111111111011111001001001;
assign LUT_4[274] = 32'b00000000000000000010000111110101;
assign LUT_4[275] = 32'b11111111111111111011010011101101;
assign LUT_4[276] = 32'b11111111111111111111101101101101;
assign LUT_4[277] = 32'b11111111111111111000111001100101;
assign LUT_4[278] = 32'b11111111111111111111001000010001;
assign LUT_4[279] = 32'b11111111111111111000010100001001;
assign LUT_4[280] = 32'b11111111111111111011111001100110;
assign LUT_4[281] = 32'b11111111111111110101000101011110;
assign LUT_4[282] = 32'b11111111111111111011010100001010;
assign LUT_4[283] = 32'b11111111111111110100100000000010;
assign LUT_4[284] = 32'b11111111111111111000111010000010;
assign LUT_4[285] = 32'b11111111111111110010000101111010;
assign LUT_4[286] = 32'b11111111111111111000010100100110;
assign LUT_4[287] = 32'b11111111111111110001100000011110;
assign LUT_4[288] = 32'b00000000000000000011010110101010;
assign LUT_4[289] = 32'b11111111111111111100100010100010;
assign LUT_4[290] = 32'b00000000000000000010110001001110;
assign LUT_4[291] = 32'b11111111111111111011111101000110;
assign LUT_4[292] = 32'b00000000000000000000010111000110;
assign LUT_4[293] = 32'b11111111111111111001100010111110;
assign LUT_4[294] = 32'b11111111111111111111110001101010;
assign LUT_4[295] = 32'b11111111111111111000111101100010;
assign LUT_4[296] = 32'b11111111111111111100100010111111;
assign LUT_4[297] = 32'b11111111111111110101101110110111;
assign LUT_4[298] = 32'b11111111111111111011111101100011;
assign LUT_4[299] = 32'b11111111111111110101001001011011;
assign LUT_4[300] = 32'b11111111111111111001100011011011;
assign LUT_4[301] = 32'b11111111111111110010101111010011;
assign LUT_4[302] = 32'b11111111111111111000111101111111;
assign LUT_4[303] = 32'b11111111111111110010001001110111;
assign LUT_4[304] = 32'b00000000000000000001001000011000;
assign LUT_4[305] = 32'b11111111111111111010010100010000;
assign LUT_4[306] = 32'b00000000000000000000100010111100;
assign LUT_4[307] = 32'b11111111111111111001101110110100;
assign LUT_4[308] = 32'b11111111111111111110001000110100;
assign LUT_4[309] = 32'b11111111111111110111010100101100;
assign LUT_4[310] = 32'b11111111111111111101100011011000;
assign LUT_4[311] = 32'b11111111111111110110101111010000;
assign LUT_4[312] = 32'b11111111111111111010010100101101;
assign LUT_4[313] = 32'b11111111111111110011100000100101;
assign LUT_4[314] = 32'b11111111111111111001101111010001;
assign LUT_4[315] = 32'b11111111111111110010111011001001;
assign LUT_4[316] = 32'b11111111111111110111010101001001;
assign LUT_4[317] = 32'b11111111111111110000100001000001;
assign LUT_4[318] = 32'b11111111111111110110101111101101;
assign LUT_4[319] = 32'b11111111111111101111111011100101;
assign LUT_4[320] = 32'b00000000000000000110010010110111;
assign LUT_4[321] = 32'b11111111111111111111011110101111;
assign LUT_4[322] = 32'b00000000000000000101101101011011;
assign LUT_4[323] = 32'b11111111111111111110111001010011;
assign LUT_4[324] = 32'b00000000000000000011010011010011;
assign LUT_4[325] = 32'b11111111111111111100011111001011;
assign LUT_4[326] = 32'b00000000000000000010101101110111;
assign LUT_4[327] = 32'b11111111111111111011111001101111;
assign LUT_4[328] = 32'b11111111111111111111011111001100;
assign LUT_4[329] = 32'b11111111111111111000101011000100;
assign LUT_4[330] = 32'b11111111111111111110111001110000;
assign LUT_4[331] = 32'b11111111111111111000000101101000;
assign LUT_4[332] = 32'b11111111111111111100011111101000;
assign LUT_4[333] = 32'b11111111111111110101101011100000;
assign LUT_4[334] = 32'b11111111111111111011111010001100;
assign LUT_4[335] = 32'b11111111111111110101000110000100;
assign LUT_4[336] = 32'b00000000000000000100000100100101;
assign LUT_4[337] = 32'b11111111111111111101010000011101;
assign LUT_4[338] = 32'b00000000000000000011011111001001;
assign LUT_4[339] = 32'b11111111111111111100101011000001;
assign LUT_4[340] = 32'b00000000000000000001000101000001;
assign LUT_4[341] = 32'b11111111111111111010010000111001;
assign LUT_4[342] = 32'b00000000000000000000011111100101;
assign LUT_4[343] = 32'b11111111111111111001101011011101;
assign LUT_4[344] = 32'b11111111111111111101010000111010;
assign LUT_4[345] = 32'b11111111111111110110011100110010;
assign LUT_4[346] = 32'b11111111111111111100101011011110;
assign LUT_4[347] = 32'b11111111111111110101110111010110;
assign LUT_4[348] = 32'b11111111111111111010010001010110;
assign LUT_4[349] = 32'b11111111111111110011011101001110;
assign LUT_4[350] = 32'b11111111111111111001101011111010;
assign LUT_4[351] = 32'b11111111111111110010110111110010;
assign LUT_4[352] = 32'b00000000000000000100101101111110;
assign LUT_4[353] = 32'b11111111111111111101111001110110;
assign LUT_4[354] = 32'b00000000000000000100001000100010;
assign LUT_4[355] = 32'b11111111111111111101010100011010;
assign LUT_4[356] = 32'b00000000000000000001101110011010;
assign LUT_4[357] = 32'b11111111111111111010111010010010;
assign LUT_4[358] = 32'b00000000000000000001001000111110;
assign LUT_4[359] = 32'b11111111111111111010010100110110;
assign LUT_4[360] = 32'b11111111111111111101111010010011;
assign LUT_4[361] = 32'b11111111111111110111000110001011;
assign LUT_4[362] = 32'b11111111111111111101010100110111;
assign LUT_4[363] = 32'b11111111111111110110100000101111;
assign LUT_4[364] = 32'b11111111111111111010111010101111;
assign LUT_4[365] = 32'b11111111111111110100000110100111;
assign LUT_4[366] = 32'b11111111111111111010010101010011;
assign LUT_4[367] = 32'b11111111111111110011100001001011;
assign LUT_4[368] = 32'b00000000000000000010011111101100;
assign LUT_4[369] = 32'b11111111111111111011101011100100;
assign LUT_4[370] = 32'b00000000000000000001111010010000;
assign LUT_4[371] = 32'b11111111111111111011000110001000;
assign LUT_4[372] = 32'b11111111111111111111100000001000;
assign LUT_4[373] = 32'b11111111111111111000101100000000;
assign LUT_4[374] = 32'b11111111111111111110111010101100;
assign LUT_4[375] = 32'b11111111111111111000000110100100;
assign LUT_4[376] = 32'b11111111111111111011101100000001;
assign LUT_4[377] = 32'b11111111111111110100110111111001;
assign LUT_4[378] = 32'b11111111111111111011000110100101;
assign LUT_4[379] = 32'b11111111111111110100010010011101;
assign LUT_4[380] = 32'b11111111111111111000101100011101;
assign LUT_4[381] = 32'b11111111111111110001111000010101;
assign LUT_4[382] = 32'b11111111111111111000000111000001;
assign LUT_4[383] = 32'b11111111111111110001010010111001;
assign LUT_4[384] = 32'b00000000000000000111100001101011;
assign LUT_4[385] = 32'b00000000000000000000101101100011;
assign LUT_4[386] = 32'b00000000000000000110111100001111;
assign LUT_4[387] = 32'b00000000000000000000001000000111;
assign LUT_4[388] = 32'b00000000000000000100100010000111;
assign LUT_4[389] = 32'b11111111111111111101101101111111;
assign LUT_4[390] = 32'b00000000000000000011111100101011;
assign LUT_4[391] = 32'b11111111111111111101001000100011;
assign LUT_4[392] = 32'b00000000000000000000101110000000;
assign LUT_4[393] = 32'b11111111111111111001111001111000;
assign LUT_4[394] = 32'b00000000000000000000001000100100;
assign LUT_4[395] = 32'b11111111111111111001010100011100;
assign LUT_4[396] = 32'b11111111111111111101101110011100;
assign LUT_4[397] = 32'b11111111111111110110111010010100;
assign LUT_4[398] = 32'b11111111111111111101001001000000;
assign LUT_4[399] = 32'b11111111111111110110010100111000;
assign LUT_4[400] = 32'b00000000000000000101010011011001;
assign LUT_4[401] = 32'b11111111111111111110011111010001;
assign LUT_4[402] = 32'b00000000000000000100101101111101;
assign LUT_4[403] = 32'b11111111111111111101111001110101;
assign LUT_4[404] = 32'b00000000000000000010010011110101;
assign LUT_4[405] = 32'b11111111111111111011011111101101;
assign LUT_4[406] = 32'b00000000000000000001101110011001;
assign LUT_4[407] = 32'b11111111111111111010111010010001;
assign LUT_4[408] = 32'b11111111111111111110011111101110;
assign LUT_4[409] = 32'b11111111111111110111101011100110;
assign LUT_4[410] = 32'b11111111111111111101111010010010;
assign LUT_4[411] = 32'b11111111111111110111000110001010;
assign LUT_4[412] = 32'b11111111111111111011100000001010;
assign LUT_4[413] = 32'b11111111111111110100101100000010;
assign LUT_4[414] = 32'b11111111111111111010111010101110;
assign LUT_4[415] = 32'b11111111111111110100000110100110;
assign LUT_4[416] = 32'b00000000000000000101111100110010;
assign LUT_4[417] = 32'b11111111111111111111001000101010;
assign LUT_4[418] = 32'b00000000000000000101010111010110;
assign LUT_4[419] = 32'b11111111111111111110100011001110;
assign LUT_4[420] = 32'b00000000000000000010111101001110;
assign LUT_4[421] = 32'b11111111111111111100001001000110;
assign LUT_4[422] = 32'b00000000000000000010010111110010;
assign LUT_4[423] = 32'b11111111111111111011100011101010;
assign LUT_4[424] = 32'b11111111111111111111001001000111;
assign LUT_4[425] = 32'b11111111111111111000010100111111;
assign LUT_4[426] = 32'b11111111111111111110100011101011;
assign LUT_4[427] = 32'b11111111111111110111101111100011;
assign LUT_4[428] = 32'b11111111111111111100001001100011;
assign LUT_4[429] = 32'b11111111111111110101010101011011;
assign LUT_4[430] = 32'b11111111111111111011100100000111;
assign LUT_4[431] = 32'b11111111111111110100101111111111;
assign LUT_4[432] = 32'b00000000000000000011101110100000;
assign LUT_4[433] = 32'b11111111111111111100111010011000;
assign LUT_4[434] = 32'b00000000000000000011001001000100;
assign LUT_4[435] = 32'b11111111111111111100010100111100;
assign LUT_4[436] = 32'b00000000000000000000101110111100;
assign LUT_4[437] = 32'b11111111111111111001111010110100;
assign LUT_4[438] = 32'b00000000000000000000001001100000;
assign LUT_4[439] = 32'b11111111111111111001010101011000;
assign LUT_4[440] = 32'b11111111111111111100111010110101;
assign LUT_4[441] = 32'b11111111111111110110000110101101;
assign LUT_4[442] = 32'b11111111111111111100010101011001;
assign LUT_4[443] = 32'b11111111111111110101100001010001;
assign LUT_4[444] = 32'b11111111111111111001111011010001;
assign LUT_4[445] = 32'b11111111111111110011000111001001;
assign LUT_4[446] = 32'b11111111111111111001010101110101;
assign LUT_4[447] = 32'b11111111111111110010100001101101;
assign LUT_4[448] = 32'b00000000000000001000111000111111;
assign LUT_4[449] = 32'b00000000000000000010000100110111;
assign LUT_4[450] = 32'b00000000000000001000010011100011;
assign LUT_4[451] = 32'b00000000000000000001011111011011;
assign LUT_4[452] = 32'b00000000000000000101111001011011;
assign LUT_4[453] = 32'b11111111111111111111000101010011;
assign LUT_4[454] = 32'b00000000000000000101010011111111;
assign LUT_4[455] = 32'b11111111111111111110011111110111;
assign LUT_4[456] = 32'b00000000000000000010000101010100;
assign LUT_4[457] = 32'b11111111111111111011010001001100;
assign LUT_4[458] = 32'b00000000000000000001011111111000;
assign LUT_4[459] = 32'b11111111111111111010101011110000;
assign LUT_4[460] = 32'b11111111111111111111000101110000;
assign LUT_4[461] = 32'b11111111111111111000010001101000;
assign LUT_4[462] = 32'b11111111111111111110100000010100;
assign LUT_4[463] = 32'b11111111111111110111101100001100;
assign LUT_4[464] = 32'b00000000000000000110101010101101;
assign LUT_4[465] = 32'b11111111111111111111110110100101;
assign LUT_4[466] = 32'b00000000000000000110000101010001;
assign LUT_4[467] = 32'b11111111111111111111010001001001;
assign LUT_4[468] = 32'b00000000000000000011101011001001;
assign LUT_4[469] = 32'b11111111111111111100110111000001;
assign LUT_4[470] = 32'b00000000000000000011000101101101;
assign LUT_4[471] = 32'b11111111111111111100010001100101;
assign LUT_4[472] = 32'b11111111111111111111110111000010;
assign LUT_4[473] = 32'b11111111111111111001000010111010;
assign LUT_4[474] = 32'b11111111111111111111010001100110;
assign LUT_4[475] = 32'b11111111111111111000011101011110;
assign LUT_4[476] = 32'b11111111111111111100110111011110;
assign LUT_4[477] = 32'b11111111111111110110000011010110;
assign LUT_4[478] = 32'b11111111111111111100010010000010;
assign LUT_4[479] = 32'b11111111111111110101011101111010;
assign LUT_4[480] = 32'b00000000000000000111010100000110;
assign LUT_4[481] = 32'b00000000000000000000011111111110;
assign LUT_4[482] = 32'b00000000000000000110101110101010;
assign LUT_4[483] = 32'b11111111111111111111111010100010;
assign LUT_4[484] = 32'b00000000000000000100010100100010;
assign LUT_4[485] = 32'b11111111111111111101100000011010;
assign LUT_4[486] = 32'b00000000000000000011101111000110;
assign LUT_4[487] = 32'b11111111111111111100111010111110;
assign LUT_4[488] = 32'b00000000000000000000100000011011;
assign LUT_4[489] = 32'b11111111111111111001101100010011;
assign LUT_4[490] = 32'b11111111111111111111111010111111;
assign LUT_4[491] = 32'b11111111111111111001000110110111;
assign LUT_4[492] = 32'b11111111111111111101100000110111;
assign LUT_4[493] = 32'b11111111111111110110101100101111;
assign LUT_4[494] = 32'b11111111111111111100111011011011;
assign LUT_4[495] = 32'b11111111111111110110000111010011;
assign LUT_4[496] = 32'b00000000000000000101000101110100;
assign LUT_4[497] = 32'b11111111111111111110010001101100;
assign LUT_4[498] = 32'b00000000000000000100100000011000;
assign LUT_4[499] = 32'b11111111111111111101101100010000;
assign LUT_4[500] = 32'b00000000000000000010000110010000;
assign LUT_4[501] = 32'b11111111111111111011010010001000;
assign LUT_4[502] = 32'b00000000000000000001100000110100;
assign LUT_4[503] = 32'b11111111111111111010101100101100;
assign LUT_4[504] = 32'b11111111111111111110010010001001;
assign LUT_4[505] = 32'b11111111111111110111011110000001;
assign LUT_4[506] = 32'b11111111111111111101101100101101;
assign LUT_4[507] = 32'b11111111111111110110111000100101;
assign LUT_4[508] = 32'b11111111111111111011010010100101;
assign LUT_4[509] = 32'b11111111111111110100011110011101;
assign LUT_4[510] = 32'b11111111111111111010101101001001;
assign LUT_4[511] = 32'b11111111111111110011111001000001;
assign LUT_4[512] = 32'b11111111111111111111000100001000;
assign LUT_4[513] = 32'b11111111111111111000010000000000;
assign LUT_4[514] = 32'b11111111111111111110011110101100;
assign LUT_4[515] = 32'b11111111111111110111101010100100;
assign LUT_4[516] = 32'b11111111111111111100000100100100;
assign LUT_4[517] = 32'b11111111111111110101010000011100;
assign LUT_4[518] = 32'b11111111111111111011011111001000;
assign LUT_4[519] = 32'b11111111111111110100101011000000;
assign LUT_4[520] = 32'b11111111111111111000010000011101;
assign LUT_4[521] = 32'b11111111111111110001011100010101;
assign LUT_4[522] = 32'b11111111111111110111101011000001;
assign LUT_4[523] = 32'b11111111111111110000110110111001;
assign LUT_4[524] = 32'b11111111111111110101010000111001;
assign LUT_4[525] = 32'b11111111111111101110011100110001;
assign LUT_4[526] = 32'b11111111111111110100101011011101;
assign LUT_4[527] = 32'b11111111111111101101110111010101;
assign LUT_4[528] = 32'b11111111111111111100110101110110;
assign LUT_4[529] = 32'b11111111111111110110000001101110;
assign LUT_4[530] = 32'b11111111111111111100010000011010;
assign LUT_4[531] = 32'b11111111111111110101011100010010;
assign LUT_4[532] = 32'b11111111111111111001110110010010;
assign LUT_4[533] = 32'b11111111111111110011000010001010;
assign LUT_4[534] = 32'b11111111111111111001010000110110;
assign LUT_4[535] = 32'b11111111111111110010011100101110;
assign LUT_4[536] = 32'b11111111111111110110000010001011;
assign LUT_4[537] = 32'b11111111111111101111001110000011;
assign LUT_4[538] = 32'b11111111111111110101011100101111;
assign LUT_4[539] = 32'b11111111111111101110101000100111;
assign LUT_4[540] = 32'b11111111111111110011000010100111;
assign LUT_4[541] = 32'b11111111111111101100001110011111;
assign LUT_4[542] = 32'b11111111111111110010011101001011;
assign LUT_4[543] = 32'b11111111111111101011101001000011;
assign LUT_4[544] = 32'b11111111111111111101011111001111;
assign LUT_4[545] = 32'b11111111111111110110101011000111;
assign LUT_4[546] = 32'b11111111111111111100111001110011;
assign LUT_4[547] = 32'b11111111111111110110000101101011;
assign LUT_4[548] = 32'b11111111111111111010011111101011;
assign LUT_4[549] = 32'b11111111111111110011101011100011;
assign LUT_4[550] = 32'b11111111111111111001111010001111;
assign LUT_4[551] = 32'b11111111111111110011000110000111;
assign LUT_4[552] = 32'b11111111111111110110101011100100;
assign LUT_4[553] = 32'b11111111111111101111110111011100;
assign LUT_4[554] = 32'b11111111111111110110000110001000;
assign LUT_4[555] = 32'b11111111111111101111010010000000;
assign LUT_4[556] = 32'b11111111111111110011101100000000;
assign LUT_4[557] = 32'b11111111111111101100110111111000;
assign LUT_4[558] = 32'b11111111111111110011000110100100;
assign LUT_4[559] = 32'b11111111111111101100010010011100;
assign LUT_4[560] = 32'b11111111111111111011010000111101;
assign LUT_4[561] = 32'b11111111111111110100011100110101;
assign LUT_4[562] = 32'b11111111111111111010101011100001;
assign LUT_4[563] = 32'b11111111111111110011110111011001;
assign LUT_4[564] = 32'b11111111111111111000010001011001;
assign LUT_4[565] = 32'b11111111111111110001011101010001;
assign LUT_4[566] = 32'b11111111111111110111101011111101;
assign LUT_4[567] = 32'b11111111111111110000110111110101;
assign LUT_4[568] = 32'b11111111111111110100011101010010;
assign LUT_4[569] = 32'b11111111111111101101101001001010;
assign LUT_4[570] = 32'b11111111111111110011110111110110;
assign LUT_4[571] = 32'b11111111111111101101000011101110;
assign LUT_4[572] = 32'b11111111111111110001011101101110;
assign LUT_4[573] = 32'b11111111111111101010101001100110;
assign LUT_4[574] = 32'b11111111111111110000111000010010;
assign LUT_4[575] = 32'b11111111111111101010000100001010;
assign LUT_4[576] = 32'b00000000000000000000011011011100;
assign LUT_4[577] = 32'b11111111111111111001100111010100;
assign LUT_4[578] = 32'b11111111111111111111110110000000;
assign LUT_4[579] = 32'b11111111111111111001000001111000;
assign LUT_4[580] = 32'b11111111111111111101011011111000;
assign LUT_4[581] = 32'b11111111111111110110100111110000;
assign LUT_4[582] = 32'b11111111111111111100110110011100;
assign LUT_4[583] = 32'b11111111111111110110000010010100;
assign LUT_4[584] = 32'b11111111111111111001100111110001;
assign LUT_4[585] = 32'b11111111111111110010110011101001;
assign LUT_4[586] = 32'b11111111111111111001000010010101;
assign LUT_4[587] = 32'b11111111111111110010001110001101;
assign LUT_4[588] = 32'b11111111111111110110101000001101;
assign LUT_4[589] = 32'b11111111111111101111110100000101;
assign LUT_4[590] = 32'b11111111111111110110000010110001;
assign LUT_4[591] = 32'b11111111111111101111001110101001;
assign LUT_4[592] = 32'b11111111111111111110001101001010;
assign LUT_4[593] = 32'b11111111111111110111011001000010;
assign LUT_4[594] = 32'b11111111111111111101100111101110;
assign LUT_4[595] = 32'b11111111111111110110110011100110;
assign LUT_4[596] = 32'b11111111111111111011001101100110;
assign LUT_4[597] = 32'b11111111111111110100011001011110;
assign LUT_4[598] = 32'b11111111111111111010101000001010;
assign LUT_4[599] = 32'b11111111111111110011110100000010;
assign LUT_4[600] = 32'b11111111111111110111011001011111;
assign LUT_4[601] = 32'b11111111111111110000100101010111;
assign LUT_4[602] = 32'b11111111111111110110110100000011;
assign LUT_4[603] = 32'b11111111111111101111111111111011;
assign LUT_4[604] = 32'b11111111111111110100011001111011;
assign LUT_4[605] = 32'b11111111111111101101100101110011;
assign LUT_4[606] = 32'b11111111111111110011110100011111;
assign LUT_4[607] = 32'b11111111111111101101000000010111;
assign LUT_4[608] = 32'b11111111111111111110110110100011;
assign LUT_4[609] = 32'b11111111111111111000000010011011;
assign LUT_4[610] = 32'b11111111111111111110010001000111;
assign LUT_4[611] = 32'b11111111111111110111011100111111;
assign LUT_4[612] = 32'b11111111111111111011110110111111;
assign LUT_4[613] = 32'b11111111111111110101000010110111;
assign LUT_4[614] = 32'b11111111111111111011010001100011;
assign LUT_4[615] = 32'b11111111111111110100011101011011;
assign LUT_4[616] = 32'b11111111111111111000000010111000;
assign LUT_4[617] = 32'b11111111111111110001001110110000;
assign LUT_4[618] = 32'b11111111111111110111011101011100;
assign LUT_4[619] = 32'b11111111111111110000101001010100;
assign LUT_4[620] = 32'b11111111111111110101000011010100;
assign LUT_4[621] = 32'b11111111111111101110001111001100;
assign LUT_4[622] = 32'b11111111111111110100011101111000;
assign LUT_4[623] = 32'b11111111111111101101101001110000;
assign LUT_4[624] = 32'b11111111111111111100101000010001;
assign LUT_4[625] = 32'b11111111111111110101110100001001;
assign LUT_4[626] = 32'b11111111111111111100000010110101;
assign LUT_4[627] = 32'b11111111111111110101001110101101;
assign LUT_4[628] = 32'b11111111111111111001101000101101;
assign LUT_4[629] = 32'b11111111111111110010110100100101;
assign LUT_4[630] = 32'b11111111111111111001000011010001;
assign LUT_4[631] = 32'b11111111111111110010001111001001;
assign LUT_4[632] = 32'b11111111111111110101110100100110;
assign LUT_4[633] = 32'b11111111111111101111000000011110;
assign LUT_4[634] = 32'b11111111111111110101001111001010;
assign LUT_4[635] = 32'b11111111111111101110011011000010;
assign LUT_4[636] = 32'b11111111111111110010110101000010;
assign LUT_4[637] = 32'b11111111111111101100000000111010;
assign LUT_4[638] = 32'b11111111111111110010001111100110;
assign LUT_4[639] = 32'b11111111111111101011011011011110;
assign LUT_4[640] = 32'b00000000000000000001101010010000;
assign LUT_4[641] = 32'b11111111111111111010110110001000;
assign LUT_4[642] = 32'b00000000000000000001000100110100;
assign LUT_4[643] = 32'b11111111111111111010010000101100;
assign LUT_4[644] = 32'b11111111111111111110101010101100;
assign LUT_4[645] = 32'b11111111111111110111110110100100;
assign LUT_4[646] = 32'b11111111111111111110000101010000;
assign LUT_4[647] = 32'b11111111111111110111010001001000;
assign LUT_4[648] = 32'b11111111111111111010110110100101;
assign LUT_4[649] = 32'b11111111111111110100000010011101;
assign LUT_4[650] = 32'b11111111111111111010010001001001;
assign LUT_4[651] = 32'b11111111111111110011011101000001;
assign LUT_4[652] = 32'b11111111111111110111110111000001;
assign LUT_4[653] = 32'b11111111111111110001000010111001;
assign LUT_4[654] = 32'b11111111111111110111010001100101;
assign LUT_4[655] = 32'b11111111111111110000011101011101;
assign LUT_4[656] = 32'b11111111111111111111011011111110;
assign LUT_4[657] = 32'b11111111111111111000100111110110;
assign LUT_4[658] = 32'b11111111111111111110110110100010;
assign LUT_4[659] = 32'b11111111111111111000000010011010;
assign LUT_4[660] = 32'b11111111111111111100011100011010;
assign LUT_4[661] = 32'b11111111111111110101101000010010;
assign LUT_4[662] = 32'b11111111111111111011110110111110;
assign LUT_4[663] = 32'b11111111111111110101000010110110;
assign LUT_4[664] = 32'b11111111111111111000101000010011;
assign LUT_4[665] = 32'b11111111111111110001110100001011;
assign LUT_4[666] = 32'b11111111111111111000000010110111;
assign LUT_4[667] = 32'b11111111111111110001001110101111;
assign LUT_4[668] = 32'b11111111111111110101101000101111;
assign LUT_4[669] = 32'b11111111111111101110110100100111;
assign LUT_4[670] = 32'b11111111111111110101000011010011;
assign LUT_4[671] = 32'b11111111111111101110001111001011;
assign LUT_4[672] = 32'b00000000000000000000000101010111;
assign LUT_4[673] = 32'b11111111111111111001010001001111;
assign LUT_4[674] = 32'b11111111111111111111011111111011;
assign LUT_4[675] = 32'b11111111111111111000101011110011;
assign LUT_4[676] = 32'b11111111111111111101000101110011;
assign LUT_4[677] = 32'b11111111111111110110010001101011;
assign LUT_4[678] = 32'b11111111111111111100100000010111;
assign LUT_4[679] = 32'b11111111111111110101101100001111;
assign LUT_4[680] = 32'b11111111111111111001010001101100;
assign LUT_4[681] = 32'b11111111111111110010011101100100;
assign LUT_4[682] = 32'b11111111111111111000101100010000;
assign LUT_4[683] = 32'b11111111111111110001111000001000;
assign LUT_4[684] = 32'b11111111111111110110010010001000;
assign LUT_4[685] = 32'b11111111111111101111011110000000;
assign LUT_4[686] = 32'b11111111111111110101101100101100;
assign LUT_4[687] = 32'b11111111111111101110111000100100;
assign LUT_4[688] = 32'b11111111111111111101110111000101;
assign LUT_4[689] = 32'b11111111111111110111000010111101;
assign LUT_4[690] = 32'b11111111111111111101010001101001;
assign LUT_4[691] = 32'b11111111111111110110011101100001;
assign LUT_4[692] = 32'b11111111111111111010110111100001;
assign LUT_4[693] = 32'b11111111111111110100000011011001;
assign LUT_4[694] = 32'b11111111111111111010010010000101;
assign LUT_4[695] = 32'b11111111111111110011011101111101;
assign LUT_4[696] = 32'b11111111111111110111000011011010;
assign LUT_4[697] = 32'b11111111111111110000001111010010;
assign LUT_4[698] = 32'b11111111111111110110011101111110;
assign LUT_4[699] = 32'b11111111111111101111101001110110;
assign LUT_4[700] = 32'b11111111111111110100000011110110;
assign LUT_4[701] = 32'b11111111111111101101001111101110;
assign LUT_4[702] = 32'b11111111111111110011011110011010;
assign LUT_4[703] = 32'b11111111111111101100101010010010;
assign LUT_4[704] = 32'b00000000000000000011000001100100;
assign LUT_4[705] = 32'b11111111111111111100001101011100;
assign LUT_4[706] = 32'b00000000000000000010011100001000;
assign LUT_4[707] = 32'b11111111111111111011101000000000;
assign LUT_4[708] = 32'b00000000000000000000000010000000;
assign LUT_4[709] = 32'b11111111111111111001001101111000;
assign LUT_4[710] = 32'b11111111111111111111011100100100;
assign LUT_4[711] = 32'b11111111111111111000101000011100;
assign LUT_4[712] = 32'b11111111111111111100001101111001;
assign LUT_4[713] = 32'b11111111111111110101011001110001;
assign LUT_4[714] = 32'b11111111111111111011101000011101;
assign LUT_4[715] = 32'b11111111111111110100110100010101;
assign LUT_4[716] = 32'b11111111111111111001001110010101;
assign LUT_4[717] = 32'b11111111111111110010011010001101;
assign LUT_4[718] = 32'b11111111111111111000101000111001;
assign LUT_4[719] = 32'b11111111111111110001110100110001;
assign LUT_4[720] = 32'b00000000000000000000110011010010;
assign LUT_4[721] = 32'b11111111111111111001111111001010;
assign LUT_4[722] = 32'b00000000000000000000001101110110;
assign LUT_4[723] = 32'b11111111111111111001011001101110;
assign LUT_4[724] = 32'b11111111111111111101110011101110;
assign LUT_4[725] = 32'b11111111111111110110111111100110;
assign LUT_4[726] = 32'b11111111111111111101001110010010;
assign LUT_4[727] = 32'b11111111111111110110011010001010;
assign LUT_4[728] = 32'b11111111111111111001111111100111;
assign LUT_4[729] = 32'b11111111111111110011001011011111;
assign LUT_4[730] = 32'b11111111111111111001011010001011;
assign LUT_4[731] = 32'b11111111111111110010100110000011;
assign LUT_4[732] = 32'b11111111111111110111000000000011;
assign LUT_4[733] = 32'b11111111111111110000001011111011;
assign LUT_4[734] = 32'b11111111111111110110011010100111;
assign LUT_4[735] = 32'b11111111111111101111100110011111;
assign LUT_4[736] = 32'b00000000000000000001011100101011;
assign LUT_4[737] = 32'b11111111111111111010101000100011;
assign LUT_4[738] = 32'b00000000000000000000110111001111;
assign LUT_4[739] = 32'b11111111111111111010000011000111;
assign LUT_4[740] = 32'b11111111111111111110011101000111;
assign LUT_4[741] = 32'b11111111111111110111101000111111;
assign LUT_4[742] = 32'b11111111111111111101110111101011;
assign LUT_4[743] = 32'b11111111111111110111000011100011;
assign LUT_4[744] = 32'b11111111111111111010101001000000;
assign LUT_4[745] = 32'b11111111111111110011110100111000;
assign LUT_4[746] = 32'b11111111111111111010000011100100;
assign LUT_4[747] = 32'b11111111111111110011001111011100;
assign LUT_4[748] = 32'b11111111111111110111101001011100;
assign LUT_4[749] = 32'b11111111111111110000110101010100;
assign LUT_4[750] = 32'b11111111111111110111000100000000;
assign LUT_4[751] = 32'b11111111111111110000001111111000;
assign LUT_4[752] = 32'b11111111111111111111001110011001;
assign LUT_4[753] = 32'b11111111111111111000011010010001;
assign LUT_4[754] = 32'b11111111111111111110101000111101;
assign LUT_4[755] = 32'b11111111111111110111110100110101;
assign LUT_4[756] = 32'b11111111111111111100001110110101;
assign LUT_4[757] = 32'b11111111111111110101011010101101;
assign LUT_4[758] = 32'b11111111111111111011101001011001;
assign LUT_4[759] = 32'b11111111111111110100110101010001;
assign LUT_4[760] = 32'b11111111111111111000011010101110;
assign LUT_4[761] = 32'b11111111111111110001100110100110;
assign LUT_4[762] = 32'b11111111111111110111110101010010;
assign LUT_4[763] = 32'b11111111111111110001000001001010;
assign LUT_4[764] = 32'b11111111111111110101011011001010;
assign LUT_4[765] = 32'b11111111111111101110100111000010;
assign LUT_4[766] = 32'b11111111111111110100110101101110;
assign LUT_4[767] = 32'b11111111111111101110000001100110;
assign LUT_4[768] = 32'b00000000000000000011111111101011;
assign LUT_4[769] = 32'b11111111111111111101001011100011;
assign LUT_4[770] = 32'b00000000000000000011011010001111;
assign LUT_4[771] = 32'b11111111111111111100100110000111;
assign LUT_4[772] = 32'b00000000000000000001000000000111;
assign LUT_4[773] = 32'b11111111111111111010001011111111;
assign LUT_4[774] = 32'b00000000000000000000011010101011;
assign LUT_4[775] = 32'b11111111111111111001100110100011;
assign LUT_4[776] = 32'b11111111111111111101001100000000;
assign LUT_4[777] = 32'b11111111111111110110010111111000;
assign LUT_4[778] = 32'b11111111111111111100100110100100;
assign LUT_4[779] = 32'b11111111111111110101110010011100;
assign LUT_4[780] = 32'b11111111111111111010001100011100;
assign LUT_4[781] = 32'b11111111111111110011011000010100;
assign LUT_4[782] = 32'b11111111111111111001100111000000;
assign LUT_4[783] = 32'b11111111111111110010110010111000;
assign LUT_4[784] = 32'b00000000000000000001110001011001;
assign LUT_4[785] = 32'b11111111111111111010111101010001;
assign LUT_4[786] = 32'b00000000000000000001001011111101;
assign LUT_4[787] = 32'b11111111111111111010010111110101;
assign LUT_4[788] = 32'b11111111111111111110110001110101;
assign LUT_4[789] = 32'b11111111111111110111111101101101;
assign LUT_4[790] = 32'b11111111111111111110001100011001;
assign LUT_4[791] = 32'b11111111111111110111011000010001;
assign LUT_4[792] = 32'b11111111111111111010111101101110;
assign LUT_4[793] = 32'b11111111111111110100001001100110;
assign LUT_4[794] = 32'b11111111111111111010011000010010;
assign LUT_4[795] = 32'b11111111111111110011100100001010;
assign LUT_4[796] = 32'b11111111111111110111111110001010;
assign LUT_4[797] = 32'b11111111111111110001001010000010;
assign LUT_4[798] = 32'b11111111111111110111011000101110;
assign LUT_4[799] = 32'b11111111111111110000100100100110;
assign LUT_4[800] = 32'b00000000000000000010011010110010;
assign LUT_4[801] = 32'b11111111111111111011100110101010;
assign LUT_4[802] = 32'b00000000000000000001110101010110;
assign LUT_4[803] = 32'b11111111111111111011000001001110;
assign LUT_4[804] = 32'b11111111111111111111011011001110;
assign LUT_4[805] = 32'b11111111111111111000100111000110;
assign LUT_4[806] = 32'b11111111111111111110110101110010;
assign LUT_4[807] = 32'b11111111111111111000000001101010;
assign LUT_4[808] = 32'b11111111111111111011100111000111;
assign LUT_4[809] = 32'b11111111111111110100110010111111;
assign LUT_4[810] = 32'b11111111111111111011000001101011;
assign LUT_4[811] = 32'b11111111111111110100001101100011;
assign LUT_4[812] = 32'b11111111111111111000100111100011;
assign LUT_4[813] = 32'b11111111111111110001110011011011;
assign LUT_4[814] = 32'b11111111111111111000000010000111;
assign LUT_4[815] = 32'b11111111111111110001001101111111;
assign LUT_4[816] = 32'b00000000000000000000001100100000;
assign LUT_4[817] = 32'b11111111111111111001011000011000;
assign LUT_4[818] = 32'b11111111111111111111100111000100;
assign LUT_4[819] = 32'b11111111111111111000110010111100;
assign LUT_4[820] = 32'b11111111111111111101001100111100;
assign LUT_4[821] = 32'b11111111111111110110011000110100;
assign LUT_4[822] = 32'b11111111111111111100100111100000;
assign LUT_4[823] = 32'b11111111111111110101110011011000;
assign LUT_4[824] = 32'b11111111111111111001011000110101;
assign LUT_4[825] = 32'b11111111111111110010100100101101;
assign LUT_4[826] = 32'b11111111111111111000110011011001;
assign LUT_4[827] = 32'b11111111111111110001111111010001;
assign LUT_4[828] = 32'b11111111111111110110011001010001;
assign LUT_4[829] = 32'b11111111111111101111100101001001;
assign LUT_4[830] = 32'b11111111111111110101110011110101;
assign LUT_4[831] = 32'b11111111111111101110111111101101;
assign LUT_4[832] = 32'b00000000000000000101010110111111;
assign LUT_4[833] = 32'b11111111111111111110100010110111;
assign LUT_4[834] = 32'b00000000000000000100110001100011;
assign LUT_4[835] = 32'b11111111111111111101111101011011;
assign LUT_4[836] = 32'b00000000000000000010010111011011;
assign LUT_4[837] = 32'b11111111111111111011100011010011;
assign LUT_4[838] = 32'b00000000000000000001110001111111;
assign LUT_4[839] = 32'b11111111111111111010111101110111;
assign LUT_4[840] = 32'b11111111111111111110100011010100;
assign LUT_4[841] = 32'b11111111111111110111101111001100;
assign LUT_4[842] = 32'b11111111111111111101111101111000;
assign LUT_4[843] = 32'b11111111111111110111001001110000;
assign LUT_4[844] = 32'b11111111111111111011100011110000;
assign LUT_4[845] = 32'b11111111111111110100101111101000;
assign LUT_4[846] = 32'b11111111111111111010111110010100;
assign LUT_4[847] = 32'b11111111111111110100001010001100;
assign LUT_4[848] = 32'b00000000000000000011001000101101;
assign LUT_4[849] = 32'b11111111111111111100010100100101;
assign LUT_4[850] = 32'b00000000000000000010100011010001;
assign LUT_4[851] = 32'b11111111111111111011101111001001;
assign LUT_4[852] = 32'b00000000000000000000001001001001;
assign LUT_4[853] = 32'b11111111111111111001010101000001;
assign LUT_4[854] = 32'b11111111111111111111100011101101;
assign LUT_4[855] = 32'b11111111111111111000101111100101;
assign LUT_4[856] = 32'b11111111111111111100010101000010;
assign LUT_4[857] = 32'b11111111111111110101100000111010;
assign LUT_4[858] = 32'b11111111111111111011101111100110;
assign LUT_4[859] = 32'b11111111111111110100111011011110;
assign LUT_4[860] = 32'b11111111111111111001010101011110;
assign LUT_4[861] = 32'b11111111111111110010100001010110;
assign LUT_4[862] = 32'b11111111111111111000110000000010;
assign LUT_4[863] = 32'b11111111111111110001111011111010;
assign LUT_4[864] = 32'b00000000000000000011110010000110;
assign LUT_4[865] = 32'b11111111111111111100111101111110;
assign LUT_4[866] = 32'b00000000000000000011001100101010;
assign LUT_4[867] = 32'b11111111111111111100011000100010;
assign LUT_4[868] = 32'b00000000000000000000110010100010;
assign LUT_4[869] = 32'b11111111111111111001111110011010;
assign LUT_4[870] = 32'b00000000000000000000001101000110;
assign LUT_4[871] = 32'b11111111111111111001011000111110;
assign LUT_4[872] = 32'b11111111111111111100111110011011;
assign LUT_4[873] = 32'b11111111111111110110001010010011;
assign LUT_4[874] = 32'b11111111111111111100011000111111;
assign LUT_4[875] = 32'b11111111111111110101100100110111;
assign LUT_4[876] = 32'b11111111111111111001111110110111;
assign LUT_4[877] = 32'b11111111111111110011001010101111;
assign LUT_4[878] = 32'b11111111111111111001011001011011;
assign LUT_4[879] = 32'b11111111111111110010100101010011;
assign LUT_4[880] = 32'b00000000000000000001100011110100;
assign LUT_4[881] = 32'b11111111111111111010101111101100;
assign LUT_4[882] = 32'b00000000000000000000111110011000;
assign LUT_4[883] = 32'b11111111111111111010001010010000;
assign LUT_4[884] = 32'b11111111111111111110100100010000;
assign LUT_4[885] = 32'b11111111111111110111110000001000;
assign LUT_4[886] = 32'b11111111111111111101111110110100;
assign LUT_4[887] = 32'b11111111111111110111001010101100;
assign LUT_4[888] = 32'b11111111111111111010110000001001;
assign LUT_4[889] = 32'b11111111111111110011111100000001;
assign LUT_4[890] = 32'b11111111111111111010001010101101;
assign LUT_4[891] = 32'b11111111111111110011010110100101;
assign LUT_4[892] = 32'b11111111111111110111110000100101;
assign LUT_4[893] = 32'b11111111111111110000111100011101;
assign LUT_4[894] = 32'b11111111111111110111001011001001;
assign LUT_4[895] = 32'b11111111111111110000010111000001;
assign LUT_4[896] = 32'b00000000000000000110100101110011;
assign LUT_4[897] = 32'b11111111111111111111110001101011;
assign LUT_4[898] = 32'b00000000000000000110000000010111;
assign LUT_4[899] = 32'b11111111111111111111001100001111;
assign LUT_4[900] = 32'b00000000000000000011100110001111;
assign LUT_4[901] = 32'b11111111111111111100110010000111;
assign LUT_4[902] = 32'b00000000000000000011000000110011;
assign LUT_4[903] = 32'b11111111111111111100001100101011;
assign LUT_4[904] = 32'b11111111111111111111110010001000;
assign LUT_4[905] = 32'b11111111111111111000111110000000;
assign LUT_4[906] = 32'b11111111111111111111001100101100;
assign LUT_4[907] = 32'b11111111111111111000011000100100;
assign LUT_4[908] = 32'b11111111111111111100110010100100;
assign LUT_4[909] = 32'b11111111111111110101111110011100;
assign LUT_4[910] = 32'b11111111111111111100001101001000;
assign LUT_4[911] = 32'b11111111111111110101011001000000;
assign LUT_4[912] = 32'b00000000000000000100010111100001;
assign LUT_4[913] = 32'b11111111111111111101100011011001;
assign LUT_4[914] = 32'b00000000000000000011110010000101;
assign LUT_4[915] = 32'b11111111111111111100111101111101;
assign LUT_4[916] = 32'b00000000000000000001010111111101;
assign LUT_4[917] = 32'b11111111111111111010100011110101;
assign LUT_4[918] = 32'b00000000000000000000110010100001;
assign LUT_4[919] = 32'b11111111111111111001111110011001;
assign LUT_4[920] = 32'b11111111111111111101100011110110;
assign LUT_4[921] = 32'b11111111111111110110101111101110;
assign LUT_4[922] = 32'b11111111111111111100111110011010;
assign LUT_4[923] = 32'b11111111111111110110001010010010;
assign LUT_4[924] = 32'b11111111111111111010100100010010;
assign LUT_4[925] = 32'b11111111111111110011110000001010;
assign LUT_4[926] = 32'b11111111111111111001111110110110;
assign LUT_4[927] = 32'b11111111111111110011001010101110;
assign LUT_4[928] = 32'b00000000000000000101000000111010;
assign LUT_4[929] = 32'b11111111111111111110001100110010;
assign LUT_4[930] = 32'b00000000000000000100011011011110;
assign LUT_4[931] = 32'b11111111111111111101100111010110;
assign LUT_4[932] = 32'b00000000000000000010000001010110;
assign LUT_4[933] = 32'b11111111111111111011001101001110;
assign LUT_4[934] = 32'b00000000000000000001011011111010;
assign LUT_4[935] = 32'b11111111111111111010100111110010;
assign LUT_4[936] = 32'b11111111111111111110001101001111;
assign LUT_4[937] = 32'b11111111111111110111011001000111;
assign LUT_4[938] = 32'b11111111111111111101100111110011;
assign LUT_4[939] = 32'b11111111111111110110110011101011;
assign LUT_4[940] = 32'b11111111111111111011001101101011;
assign LUT_4[941] = 32'b11111111111111110100011001100011;
assign LUT_4[942] = 32'b11111111111111111010101000001111;
assign LUT_4[943] = 32'b11111111111111110011110100000111;
assign LUT_4[944] = 32'b00000000000000000010110010101000;
assign LUT_4[945] = 32'b11111111111111111011111110100000;
assign LUT_4[946] = 32'b00000000000000000010001101001100;
assign LUT_4[947] = 32'b11111111111111111011011001000100;
assign LUT_4[948] = 32'b11111111111111111111110011000100;
assign LUT_4[949] = 32'b11111111111111111000111110111100;
assign LUT_4[950] = 32'b11111111111111111111001101101000;
assign LUT_4[951] = 32'b11111111111111111000011001100000;
assign LUT_4[952] = 32'b11111111111111111011111110111101;
assign LUT_4[953] = 32'b11111111111111110101001010110101;
assign LUT_4[954] = 32'b11111111111111111011011001100001;
assign LUT_4[955] = 32'b11111111111111110100100101011001;
assign LUT_4[956] = 32'b11111111111111111000111111011001;
assign LUT_4[957] = 32'b11111111111111110010001011010001;
assign LUT_4[958] = 32'b11111111111111111000011001111101;
assign LUT_4[959] = 32'b11111111111111110001100101110101;
assign LUT_4[960] = 32'b00000000000000000111111101000111;
assign LUT_4[961] = 32'b00000000000000000001001000111111;
assign LUT_4[962] = 32'b00000000000000000111010111101011;
assign LUT_4[963] = 32'b00000000000000000000100011100011;
assign LUT_4[964] = 32'b00000000000000000100111101100011;
assign LUT_4[965] = 32'b11111111111111111110001001011011;
assign LUT_4[966] = 32'b00000000000000000100011000000111;
assign LUT_4[967] = 32'b11111111111111111101100011111111;
assign LUT_4[968] = 32'b00000000000000000001001001011100;
assign LUT_4[969] = 32'b11111111111111111010010101010100;
assign LUT_4[970] = 32'b00000000000000000000100100000000;
assign LUT_4[971] = 32'b11111111111111111001101111111000;
assign LUT_4[972] = 32'b11111111111111111110001001111000;
assign LUT_4[973] = 32'b11111111111111110111010101110000;
assign LUT_4[974] = 32'b11111111111111111101100100011100;
assign LUT_4[975] = 32'b11111111111111110110110000010100;
assign LUT_4[976] = 32'b00000000000000000101101110110101;
assign LUT_4[977] = 32'b11111111111111111110111010101101;
assign LUT_4[978] = 32'b00000000000000000101001001011001;
assign LUT_4[979] = 32'b11111111111111111110010101010001;
assign LUT_4[980] = 32'b00000000000000000010101111010001;
assign LUT_4[981] = 32'b11111111111111111011111011001001;
assign LUT_4[982] = 32'b00000000000000000010001001110101;
assign LUT_4[983] = 32'b11111111111111111011010101101101;
assign LUT_4[984] = 32'b11111111111111111110111011001010;
assign LUT_4[985] = 32'b11111111111111111000000111000010;
assign LUT_4[986] = 32'b11111111111111111110010101101110;
assign LUT_4[987] = 32'b11111111111111110111100001100110;
assign LUT_4[988] = 32'b11111111111111111011111011100110;
assign LUT_4[989] = 32'b11111111111111110101000111011110;
assign LUT_4[990] = 32'b11111111111111111011010110001010;
assign LUT_4[991] = 32'b11111111111111110100100010000010;
assign LUT_4[992] = 32'b00000000000000000110011000001110;
assign LUT_4[993] = 32'b11111111111111111111100100000110;
assign LUT_4[994] = 32'b00000000000000000101110010110010;
assign LUT_4[995] = 32'b11111111111111111110111110101010;
assign LUT_4[996] = 32'b00000000000000000011011000101010;
assign LUT_4[997] = 32'b11111111111111111100100100100010;
assign LUT_4[998] = 32'b00000000000000000010110011001110;
assign LUT_4[999] = 32'b11111111111111111011111111000110;
assign LUT_4[1000] = 32'b11111111111111111111100100100011;
assign LUT_4[1001] = 32'b11111111111111111000110000011011;
assign LUT_4[1002] = 32'b11111111111111111110111111000111;
assign LUT_4[1003] = 32'b11111111111111111000001010111111;
assign LUT_4[1004] = 32'b11111111111111111100100100111111;
assign LUT_4[1005] = 32'b11111111111111110101110000110111;
assign LUT_4[1006] = 32'b11111111111111111011111111100011;
assign LUT_4[1007] = 32'b11111111111111110101001011011011;
assign LUT_4[1008] = 32'b00000000000000000100001001111100;
assign LUT_4[1009] = 32'b11111111111111111101010101110100;
assign LUT_4[1010] = 32'b00000000000000000011100100100000;
assign LUT_4[1011] = 32'b11111111111111111100110000011000;
assign LUT_4[1012] = 32'b00000000000000000001001010011000;
assign LUT_4[1013] = 32'b11111111111111111010010110010000;
assign LUT_4[1014] = 32'b00000000000000000000100100111100;
assign LUT_4[1015] = 32'b11111111111111111001110000110100;
assign LUT_4[1016] = 32'b11111111111111111101010110010001;
assign LUT_4[1017] = 32'b11111111111111110110100010001001;
assign LUT_4[1018] = 32'b11111111111111111100110000110101;
assign LUT_4[1019] = 32'b11111111111111110101111100101101;
assign LUT_4[1020] = 32'b11111111111111111010010110101101;
assign LUT_4[1021] = 32'b11111111111111110011100010100101;
assign LUT_4[1022] = 32'b11111111111111111001110001010001;
assign LUT_4[1023] = 32'b11111111111111110010111101001001;
assign LUT_4[1024] = 32'b00000000000000000001101010011111;
assign LUT_4[1025] = 32'b11111111111111111010110110010111;
assign LUT_4[1026] = 32'b00000000000000000001000101000011;
assign LUT_4[1027] = 32'b11111111111111111010010000111011;
assign LUT_4[1028] = 32'b11111111111111111110101010111011;
assign LUT_4[1029] = 32'b11111111111111110111110110110011;
assign LUT_4[1030] = 32'b11111111111111111110000101011111;
assign LUT_4[1031] = 32'b11111111111111110111010001010111;
assign LUT_4[1032] = 32'b11111111111111111010110110110100;
assign LUT_4[1033] = 32'b11111111111111110100000010101100;
assign LUT_4[1034] = 32'b11111111111111111010010001011000;
assign LUT_4[1035] = 32'b11111111111111110011011101010000;
assign LUT_4[1036] = 32'b11111111111111110111110111010000;
assign LUT_4[1037] = 32'b11111111111111110001000011001000;
assign LUT_4[1038] = 32'b11111111111111110111010001110100;
assign LUT_4[1039] = 32'b11111111111111110000011101101100;
assign LUT_4[1040] = 32'b11111111111111111111011100001101;
assign LUT_4[1041] = 32'b11111111111111111000101000000101;
assign LUT_4[1042] = 32'b11111111111111111110110110110001;
assign LUT_4[1043] = 32'b11111111111111111000000010101001;
assign LUT_4[1044] = 32'b11111111111111111100011100101001;
assign LUT_4[1045] = 32'b11111111111111110101101000100001;
assign LUT_4[1046] = 32'b11111111111111111011110111001101;
assign LUT_4[1047] = 32'b11111111111111110101000011000101;
assign LUT_4[1048] = 32'b11111111111111111000101000100010;
assign LUT_4[1049] = 32'b11111111111111110001110100011010;
assign LUT_4[1050] = 32'b11111111111111111000000011000110;
assign LUT_4[1051] = 32'b11111111111111110001001110111110;
assign LUT_4[1052] = 32'b11111111111111110101101000111110;
assign LUT_4[1053] = 32'b11111111111111101110110100110110;
assign LUT_4[1054] = 32'b11111111111111110101000011100010;
assign LUT_4[1055] = 32'b11111111111111101110001111011010;
assign LUT_4[1056] = 32'b00000000000000000000000101100110;
assign LUT_4[1057] = 32'b11111111111111111001010001011110;
assign LUT_4[1058] = 32'b11111111111111111111100000001010;
assign LUT_4[1059] = 32'b11111111111111111000101100000010;
assign LUT_4[1060] = 32'b11111111111111111101000110000010;
assign LUT_4[1061] = 32'b11111111111111110110010001111010;
assign LUT_4[1062] = 32'b11111111111111111100100000100110;
assign LUT_4[1063] = 32'b11111111111111110101101100011110;
assign LUT_4[1064] = 32'b11111111111111111001010001111011;
assign LUT_4[1065] = 32'b11111111111111110010011101110011;
assign LUT_4[1066] = 32'b11111111111111111000101100011111;
assign LUT_4[1067] = 32'b11111111111111110001111000010111;
assign LUT_4[1068] = 32'b11111111111111110110010010010111;
assign LUT_4[1069] = 32'b11111111111111101111011110001111;
assign LUT_4[1070] = 32'b11111111111111110101101100111011;
assign LUT_4[1071] = 32'b11111111111111101110111000110011;
assign LUT_4[1072] = 32'b11111111111111111101110111010100;
assign LUT_4[1073] = 32'b11111111111111110111000011001100;
assign LUT_4[1074] = 32'b11111111111111111101010001111000;
assign LUT_4[1075] = 32'b11111111111111110110011101110000;
assign LUT_4[1076] = 32'b11111111111111111010110111110000;
assign LUT_4[1077] = 32'b11111111111111110100000011101000;
assign LUT_4[1078] = 32'b11111111111111111010010010010100;
assign LUT_4[1079] = 32'b11111111111111110011011110001100;
assign LUT_4[1080] = 32'b11111111111111110111000011101001;
assign LUT_4[1081] = 32'b11111111111111110000001111100001;
assign LUT_4[1082] = 32'b11111111111111110110011110001101;
assign LUT_4[1083] = 32'b11111111111111101111101010000101;
assign LUT_4[1084] = 32'b11111111111111110100000100000101;
assign LUT_4[1085] = 32'b11111111111111101101001111111101;
assign LUT_4[1086] = 32'b11111111111111110011011110101001;
assign LUT_4[1087] = 32'b11111111111111101100101010100001;
assign LUT_4[1088] = 32'b00000000000000000011000001110011;
assign LUT_4[1089] = 32'b11111111111111111100001101101011;
assign LUT_4[1090] = 32'b00000000000000000010011100010111;
assign LUT_4[1091] = 32'b11111111111111111011101000001111;
assign LUT_4[1092] = 32'b00000000000000000000000010001111;
assign LUT_4[1093] = 32'b11111111111111111001001110000111;
assign LUT_4[1094] = 32'b11111111111111111111011100110011;
assign LUT_4[1095] = 32'b11111111111111111000101000101011;
assign LUT_4[1096] = 32'b11111111111111111100001110001000;
assign LUT_4[1097] = 32'b11111111111111110101011010000000;
assign LUT_4[1098] = 32'b11111111111111111011101000101100;
assign LUT_4[1099] = 32'b11111111111111110100110100100100;
assign LUT_4[1100] = 32'b11111111111111111001001110100100;
assign LUT_4[1101] = 32'b11111111111111110010011010011100;
assign LUT_4[1102] = 32'b11111111111111111000101001001000;
assign LUT_4[1103] = 32'b11111111111111110001110101000000;
assign LUT_4[1104] = 32'b00000000000000000000110011100001;
assign LUT_4[1105] = 32'b11111111111111111001111111011001;
assign LUT_4[1106] = 32'b00000000000000000000001110000101;
assign LUT_4[1107] = 32'b11111111111111111001011001111101;
assign LUT_4[1108] = 32'b11111111111111111101110011111101;
assign LUT_4[1109] = 32'b11111111111111110110111111110101;
assign LUT_4[1110] = 32'b11111111111111111101001110100001;
assign LUT_4[1111] = 32'b11111111111111110110011010011001;
assign LUT_4[1112] = 32'b11111111111111111001111111110110;
assign LUT_4[1113] = 32'b11111111111111110011001011101110;
assign LUT_4[1114] = 32'b11111111111111111001011010011010;
assign LUT_4[1115] = 32'b11111111111111110010100110010010;
assign LUT_4[1116] = 32'b11111111111111110111000000010010;
assign LUT_4[1117] = 32'b11111111111111110000001100001010;
assign LUT_4[1118] = 32'b11111111111111110110011010110110;
assign LUT_4[1119] = 32'b11111111111111101111100110101110;
assign LUT_4[1120] = 32'b00000000000000000001011100111010;
assign LUT_4[1121] = 32'b11111111111111111010101000110010;
assign LUT_4[1122] = 32'b00000000000000000000110111011110;
assign LUT_4[1123] = 32'b11111111111111111010000011010110;
assign LUT_4[1124] = 32'b11111111111111111110011101010110;
assign LUT_4[1125] = 32'b11111111111111110111101001001110;
assign LUT_4[1126] = 32'b11111111111111111101110111111010;
assign LUT_4[1127] = 32'b11111111111111110111000011110010;
assign LUT_4[1128] = 32'b11111111111111111010101001001111;
assign LUT_4[1129] = 32'b11111111111111110011110101000111;
assign LUT_4[1130] = 32'b11111111111111111010000011110011;
assign LUT_4[1131] = 32'b11111111111111110011001111101011;
assign LUT_4[1132] = 32'b11111111111111110111101001101011;
assign LUT_4[1133] = 32'b11111111111111110000110101100011;
assign LUT_4[1134] = 32'b11111111111111110111000100001111;
assign LUT_4[1135] = 32'b11111111111111110000010000000111;
assign LUT_4[1136] = 32'b11111111111111111111001110101000;
assign LUT_4[1137] = 32'b11111111111111111000011010100000;
assign LUT_4[1138] = 32'b11111111111111111110101001001100;
assign LUT_4[1139] = 32'b11111111111111110111110101000100;
assign LUT_4[1140] = 32'b11111111111111111100001111000100;
assign LUT_4[1141] = 32'b11111111111111110101011010111100;
assign LUT_4[1142] = 32'b11111111111111111011101001101000;
assign LUT_4[1143] = 32'b11111111111111110100110101100000;
assign LUT_4[1144] = 32'b11111111111111111000011010111101;
assign LUT_4[1145] = 32'b11111111111111110001100110110101;
assign LUT_4[1146] = 32'b11111111111111110111110101100001;
assign LUT_4[1147] = 32'b11111111111111110001000001011001;
assign LUT_4[1148] = 32'b11111111111111110101011011011001;
assign LUT_4[1149] = 32'b11111111111111101110100111010001;
assign LUT_4[1150] = 32'b11111111111111110100110101111101;
assign LUT_4[1151] = 32'b11111111111111101110000001110101;
assign LUT_4[1152] = 32'b00000000000000000100010000100111;
assign LUT_4[1153] = 32'b11111111111111111101011100011111;
assign LUT_4[1154] = 32'b00000000000000000011101011001011;
assign LUT_4[1155] = 32'b11111111111111111100110111000011;
assign LUT_4[1156] = 32'b00000000000000000001010001000011;
assign LUT_4[1157] = 32'b11111111111111111010011100111011;
assign LUT_4[1158] = 32'b00000000000000000000101011100111;
assign LUT_4[1159] = 32'b11111111111111111001110111011111;
assign LUT_4[1160] = 32'b11111111111111111101011100111100;
assign LUT_4[1161] = 32'b11111111111111110110101000110100;
assign LUT_4[1162] = 32'b11111111111111111100110111100000;
assign LUT_4[1163] = 32'b11111111111111110110000011011000;
assign LUT_4[1164] = 32'b11111111111111111010011101011000;
assign LUT_4[1165] = 32'b11111111111111110011101001010000;
assign LUT_4[1166] = 32'b11111111111111111001110111111100;
assign LUT_4[1167] = 32'b11111111111111110011000011110100;
assign LUT_4[1168] = 32'b00000000000000000010000010010101;
assign LUT_4[1169] = 32'b11111111111111111011001110001101;
assign LUT_4[1170] = 32'b00000000000000000001011100111001;
assign LUT_4[1171] = 32'b11111111111111111010101000110001;
assign LUT_4[1172] = 32'b11111111111111111111000010110001;
assign LUT_4[1173] = 32'b11111111111111111000001110101001;
assign LUT_4[1174] = 32'b11111111111111111110011101010101;
assign LUT_4[1175] = 32'b11111111111111110111101001001101;
assign LUT_4[1176] = 32'b11111111111111111011001110101010;
assign LUT_4[1177] = 32'b11111111111111110100011010100010;
assign LUT_4[1178] = 32'b11111111111111111010101001001110;
assign LUT_4[1179] = 32'b11111111111111110011110101000110;
assign LUT_4[1180] = 32'b11111111111111111000001111000110;
assign LUT_4[1181] = 32'b11111111111111110001011010111110;
assign LUT_4[1182] = 32'b11111111111111110111101001101010;
assign LUT_4[1183] = 32'b11111111111111110000110101100010;
assign LUT_4[1184] = 32'b00000000000000000010101011101110;
assign LUT_4[1185] = 32'b11111111111111111011110111100110;
assign LUT_4[1186] = 32'b00000000000000000010000110010010;
assign LUT_4[1187] = 32'b11111111111111111011010010001010;
assign LUT_4[1188] = 32'b11111111111111111111101100001010;
assign LUT_4[1189] = 32'b11111111111111111000111000000010;
assign LUT_4[1190] = 32'b11111111111111111111000110101110;
assign LUT_4[1191] = 32'b11111111111111111000010010100110;
assign LUT_4[1192] = 32'b11111111111111111011111000000011;
assign LUT_4[1193] = 32'b11111111111111110101000011111011;
assign LUT_4[1194] = 32'b11111111111111111011010010100111;
assign LUT_4[1195] = 32'b11111111111111110100011110011111;
assign LUT_4[1196] = 32'b11111111111111111000111000011111;
assign LUT_4[1197] = 32'b11111111111111110010000100010111;
assign LUT_4[1198] = 32'b11111111111111111000010011000011;
assign LUT_4[1199] = 32'b11111111111111110001011110111011;
assign LUT_4[1200] = 32'b00000000000000000000011101011100;
assign LUT_4[1201] = 32'b11111111111111111001101001010100;
assign LUT_4[1202] = 32'b11111111111111111111111000000000;
assign LUT_4[1203] = 32'b11111111111111111001000011111000;
assign LUT_4[1204] = 32'b11111111111111111101011101111000;
assign LUT_4[1205] = 32'b11111111111111110110101001110000;
assign LUT_4[1206] = 32'b11111111111111111100111000011100;
assign LUT_4[1207] = 32'b11111111111111110110000100010100;
assign LUT_4[1208] = 32'b11111111111111111001101001110001;
assign LUT_4[1209] = 32'b11111111111111110010110101101001;
assign LUT_4[1210] = 32'b11111111111111111001000100010101;
assign LUT_4[1211] = 32'b11111111111111110010010000001101;
assign LUT_4[1212] = 32'b11111111111111110110101010001101;
assign LUT_4[1213] = 32'b11111111111111101111110110000101;
assign LUT_4[1214] = 32'b11111111111111110110000100110001;
assign LUT_4[1215] = 32'b11111111111111101111010000101001;
assign LUT_4[1216] = 32'b00000000000000000101100111111011;
assign LUT_4[1217] = 32'b11111111111111111110110011110011;
assign LUT_4[1218] = 32'b00000000000000000101000010011111;
assign LUT_4[1219] = 32'b11111111111111111110001110010111;
assign LUT_4[1220] = 32'b00000000000000000010101000010111;
assign LUT_4[1221] = 32'b11111111111111111011110100001111;
assign LUT_4[1222] = 32'b00000000000000000010000010111011;
assign LUT_4[1223] = 32'b11111111111111111011001110110011;
assign LUT_4[1224] = 32'b11111111111111111110110100010000;
assign LUT_4[1225] = 32'b11111111111111111000000000001000;
assign LUT_4[1226] = 32'b11111111111111111110001110110100;
assign LUT_4[1227] = 32'b11111111111111110111011010101100;
assign LUT_4[1228] = 32'b11111111111111111011110100101100;
assign LUT_4[1229] = 32'b11111111111111110101000000100100;
assign LUT_4[1230] = 32'b11111111111111111011001111010000;
assign LUT_4[1231] = 32'b11111111111111110100011011001000;
assign LUT_4[1232] = 32'b00000000000000000011011001101001;
assign LUT_4[1233] = 32'b11111111111111111100100101100001;
assign LUT_4[1234] = 32'b00000000000000000010110100001101;
assign LUT_4[1235] = 32'b11111111111111111100000000000101;
assign LUT_4[1236] = 32'b00000000000000000000011010000101;
assign LUT_4[1237] = 32'b11111111111111111001100101111101;
assign LUT_4[1238] = 32'b11111111111111111111110100101001;
assign LUT_4[1239] = 32'b11111111111111111001000000100001;
assign LUT_4[1240] = 32'b11111111111111111100100101111110;
assign LUT_4[1241] = 32'b11111111111111110101110001110110;
assign LUT_4[1242] = 32'b11111111111111111100000000100010;
assign LUT_4[1243] = 32'b11111111111111110101001100011010;
assign LUT_4[1244] = 32'b11111111111111111001100110011010;
assign LUT_4[1245] = 32'b11111111111111110010110010010010;
assign LUT_4[1246] = 32'b11111111111111111001000000111110;
assign LUT_4[1247] = 32'b11111111111111110010001100110110;
assign LUT_4[1248] = 32'b00000000000000000100000011000010;
assign LUT_4[1249] = 32'b11111111111111111101001110111010;
assign LUT_4[1250] = 32'b00000000000000000011011101100110;
assign LUT_4[1251] = 32'b11111111111111111100101001011110;
assign LUT_4[1252] = 32'b00000000000000000001000011011110;
assign LUT_4[1253] = 32'b11111111111111111010001111010110;
assign LUT_4[1254] = 32'b00000000000000000000011110000010;
assign LUT_4[1255] = 32'b11111111111111111001101001111010;
assign LUT_4[1256] = 32'b11111111111111111101001111010111;
assign LUT_4[1257] = 32'b11111111111111110110011011001111;
assign LUT_4[1258] = 32'b11111111111111111100101001111011;
assign LUT_4[1259] = 32'b11111111111111110101110101110011;
assign LUT_4[1260] = 32'b11111111111111111010001111110011;
assign LUT_4[1261] = 32'b11111111111111110011011011101011;
assign LUT_4[1262] = 32'b11111111111111111001101010010111;
assign LUT_4[1263] = 32'b11111111111111110010110110001111;
assign LUT_4[1264] = 32'b00000000000000000001110100110000;
assign LUT_4[1265] = 32'b11111111111111111011000000101000;
assign LUT_4[1266] = 32'b00000000000000000001001111010100;
assign LUT_4[1267] = 32'b11111111111111111010011011001100;
assign LUT_4[1268] = 32'b11111111111111111110110101001100;
assign LUT_4[1269] = 32'b11111111111111111000000001000100;
assign LUT_4[1270] = 32'b11111111111111111110001111110000;
assign LUT_4[1271] = 32'b11111111111111110111011011101000;
assign LUT_4[1272] = 32'b11111111111111111011000001000101;
assign LUT_4[1273] = 32'b11111111111111110100001100111101;
assign LUT_4[1274] = 32'b11111111111111111010011011101001;
assign LUT_4[1275] = 32'b11111111111111110011100111100001;
assign LUT_4[1276] = 32'b11111111111111111000000001100001;
assign LUT_4[1277] = 32'b11111111111111110001001101011001;
assign LUT_4[1278] = 32'b11111111111111110111011100000101;
assign LUT_4[1279] = 32'b11111111111111110000100111111101;
assign LUT_4[1280] = 32'b00000000000000000110100110000010;
assign LUT_4[1281] = 32'b11111111111111111111110001111010;
assign LUT_4[1282] = 32'b00000000000000000110000000100110;
assign LUT_4[1283] = 32'b11111111111111111111001100011110;
assign LUT_4[1284] = 32'b00000000000000000011100110011110;
assign LUT_4[1285] = 32'b11111111111111111100110010010110;
assign LUT_4[1286] = 32'b00000000000000000011000001000010;
assign LUT_4[1287] = 32'b11111111111111111100001100111010;
assign LUT_4[1288] = 32'b11111111111111111111110010010111;
assign LUT_4[1289] = 32'b11111111111111111000111110001111;
assign LUT_4[1290] = 32'b11111111111111111111001100111011;
assign LUT_4[1291] = 32'b11111111111111111000011000110011;
assign LUT_4[1292] = 32'b11111111111111111100110010110011;
assign LUT_4[1293] = 32'b11111111111111110101111110101011;
assign LUT_4[1294] = 32'b11111111111111111100001101010111;
assign LUT_4[1295] = 32'b11111111111111110101011001001111;
assign LUT_4[1296] = 32'b00000000000000000100010111110000;
assign LUT_4[1297] = 32'b11111111111111111101100011101000;
assign LUT_4[1298] = 32'b00000000000000000011110010010100;
assign LUT_4[1299] = 32'b11111111111111111100111110001100;
assign LUT_4[1300] = 32'b00000000000000000001011000001100;
assign LUT_4[1301] = 32'b11111111111111111010100100000100;
assign LUT_4[1302] = 32'b00000000000000000000110010110000;
assign LUT_4[1303] = 32'b11111111111111111001111110101000;
assign LUT_4[1304] = 32'b11111111111111111101100100000101;
assign LUT_4[1305] = 32'b11111111111111110110101111111101;
assign LUT_4[1306] = 32'b11111111111111111100111110101001;
assign LUT_4[1307] = 32'b11111111111111110110001010100001;
assign LUT_4[1308] = 32'b11111111111111111010100100100001;
assign LUT_4[1309] = 32'b11111111111111110011110000011001;
assign LUT_4[1310] = 32'b11111111111111111001111111000101;
assign LUT_4[1311] = 32'b11111111111111110011001010111101;
assign LUT_4[1312] = 32'b00000000000000000101000001001001;
assign LUT_4[1313] = 32'b11111111111111111110001101000001;
assign LUT_4[1314] = 32'b00000000000000000100011011101101;
assign LUT_4[1315] = 32'b11111111111111111101100111100101;
assign LUT_4[1316] = 32'b00000000000000000010000001100101;
assign LUT_4[1317] = 32'b11111111111111111011001101011101;
assign LUT_4[1318] = 32'b00000000000000000001011100001001;
assign LUT_4[1319] = 32'b11111111111111111010101000000001;
assign LUT_4[1320] = 32'b11111111111111111110001101011110;
assign LUT_4[1321] = 32'b11111111111111110111011001010110;
assign LUT_4[1322] = 32'b11111111111111111101101000000010;
assign LUT_4[1323] = 32'b11111111111111110110110011111010;
assign LUT_4[1324] = 32'b11111111111111111011001101111010;
assign LUT_4[1325] = 32'b11111111111111110100011001110010;
assign LUT_4[1326] = 32'b11111111111111111010101000011110;
assign LUT_4[1327] = 32'b11111111111111110011110100010110;
assign LUT_4[1328] = 32'b00000000000000000010110010110111;
assign LUT_4[1329] = 32'b11111111111111111011111110101111;
assign LUT_4[1330] = 32'b00000000000000000010001101011011;
assign LUT_4[1331] = 32'b11111111111111111011011001010011;
assign LUT_4[1332] = 32'b11111111111111111111110011010011;
assign LUT_4[1333] = 32'b11111111111111111000111111001011;
assign LUT_4[1334] = 32'b11111111111111111111001101110111;
assign LUT_4[1335] = 32'b11111111111111111000011001101111;
assign LUT_4[1336] = 32'b11111111111111111011111111001100;
assign LUT_4[1337] = 32'b11111111111111110101001011000100;
assign LUT_4[1338] = 32'b11111111111111111011011001110000;
assign LUT_4[1339] = 32'b11111111111111110100100101101000;
assign LUT_4[1340] = 32'b11111111111111111000111111101000;
assign LUT_4[1341] = 32'b11111111111111110010001011100000;
assign LUT_4[1342] = 32'b11111111111111111000011010001100;
assign LUT_4[1343] = 32'b11111111111111110001100110000100;
assign LUT_4[1344] = 32'b00000000000000000111111101010110;
assign LUT_4[1345] = 32'b00000000000000000001001001001110;
assign LUT_4[1346] = 32'b00000000000000000111010111111010;
assign LUT_4[1347] = 32'b00000000000000000000100011110010;
assign LUT_4[1348] = 32'b00000000000000000100111101110010;
assign LUT_4[1349] = 32'b11111111111111111110001001101010;
assign LUT_4[1350] = 32'b00000000000000000100011000010110;
assign LUT_4[1351] = 32'b11111111111111111101100100001110;
assign LUT_4[1352] = 32'b00000000000000000001001001101011;
assign LUT_4[1353] = 32'b11111111111111111010010101100011;
assign LUT_4[1354] = 32'b00000000000000000000100100001111;
assign LUT_4[1355] = 32'b11111111111111111001110000000111;
assign LUT_4[1356] = 32'b11111111111111111110001010000111;
assign LUT_4[1357] = 32'b11111111111111110111010101111111;
assign LUT_4[1358] = 32'b11111111111111111101100100101011;
assign LUT_4[1359] = 32'b11111111111111110110110000100011;
assign LUT_4[1360] = 32'b00000000000000000101101111000100;
assign LUT_4[1361] = 32'b11111111111111111110111010111100;
assign LUT_4[1362] = 32'b00000000000000000101001001101000;
assign LUT_4[1363] = 32'b11111111111111111110010101100000;
assign LUT_4[1364] = 32'b00000000000000000010101111100000;
assign LUT_4[1365] = 32'b11111111111111111011111011011000;
assign LUT_4[1366] = 32'b00000000000000000010001010000100;
assign LUT_4[1367] = 32'b11111111111111111011010101111100;
assign LUT_4[1368] = 32'b11111111111111111110111011011001;
assign LUT_4[1369] = 32'b11111111111111111000000111010001;
assign LUT_4[1370] = 32'b11111111111111111110010101111101;
assign LUT_4[1371] = 32'b11111111111111110111100001110101;
assign LUT_4[1372] = 32'b11111111111111111011111011110101;
assign LUT_4[1373] = 32'b11111111111111110101000111101101;
assign LUT_4[1374] = 32'b11111111111111111011010110011001;
assign LUT_4[1375] = 32'b11111111111111110100100010010001;
assign LUT_4[1376] = 32'b00000000000000000110011000011101;
assign LUT_4[1377] = 32'b11111111111111111111100100010101;
assign LUT_4[1378] = 32'b00000000000000000101110011000001;
assign LUT_4[1379] = 32'b11111111111111111110111110111001;
assign LUT_4[1380] = 32'b00000000000000000011011000111001;
assign LUT_4[1381] = 32'b11111111111111111100100100110001;
assign LUT_4[1382] = 32'b00000000000000000010110011011101;
assign LUT_4[1383] = 32'b11111111111111111011111111010101;
assign LUT_4[1384] = 32'b11111111111111111111100100110010;
assign LUT_4[1385] = 32'b11111111111111111000110000101010;
assign LUT_4[1386] = 32'b11111111111111111110111111010110;
assign LUT_4[1387] = 32'b11111111111111111000001011001110;
assign LUT_4[1388] = 32'b11111111111111111100100101001110;
assign LUT_4[1389] = 32'b11111111111111110101110001000110;
assign LUT_4[1390] = 32'b11111111111111111011111111110010;
assign LUT_4[1391] = 32'b11111111111111110101001011101010;
assign LUT_4[1392] = 32'b00000000000000000100001010001011;
assign LUT_4[1393] = 32'b11111111111111111101010110000011;
assign LUT_4[1394] = 32'b00000000000000000011100100101111;
assign LUT_4[1395] = 32'b11111111111111111100110000100111;
assign LUT_4[1396] = 32'b00000000000000000001001010100111;
assign LUT_4[1397] = 32'b11111111111111111010010110011111;
assign LUT_4[1398] = 32'b00000000000000000000100101001011;
assign LUT_4[1399] = 32'b11111111111111111001110001000011;
assign LUT_4[1400] = 32'b11111111111111111101010110100000;
assign LUT_4[1401] = 32'b11111111111111110110100010011000;
assign LUT_4[1402] = 32'b11111111111111111100110001000100;
assign LUT_4[1403] = 32'b11111111111111110101111100111100;
assign LUT_4[1404] = 32'b11111111111111111010010110111100;
assign LUT_4[1405] = 32'b11111111111111110011100010110100;
assign LUT_4[1406] = 32'b11111111111111111001110001100000;
assign LUT_4[1407] = 32'b11111111111111110010111101011000;
assign LUT_4[1408] = 32'b00000000000000001001001100001010;
assign LUT_4[1409] = 32'b00000000000000000010011000000010;
assign LUT_4[1410] = 32'b00000000000000001000100110101110;
assign LUT_4[1411] = 32'b00000000000000000001110010100110;
assign LUT_4[1412] = 32'b00000000000000000110001100100110;
assign LUT_4[1413] = 32'b11111111111111111111011000011110;
assign LUT_4[1414] = 32'b00000000000000000101100111001010;
assign LUT_4[1415] = 32'b11111111111111111110110011000010;
assign LUT_4[1416] = 32'b00000000000000000010011000011111;
assign LUT_4[1417] = 32'b11111111111111111011100100010111;
assign LUT_4[1418] = 32'b00000000000000000001110011000011;
assign LUT_4[1419] = 32'b11111111111111111010111110111011;
assign LUT_4[1420] = 32'b11111111111111111111011000111011;
assign LUT_4[1421] = 32'b11111111111111111000100100110011;
assign LUT_4[1422] = 32'b11111111111111111110110011011111;
assign LUT_4[1423] = 32'b11111111111111110111111111010111;
assign LUT_4[1424] = 32'b00000000000000000110111101111000;
assign LUT_4[1425] = 32'b00000000000000000000001001110000;
assign LUT_4[1426] = 32'b00000000000000000110011000011100;
assign LUT_4[1427] = 32'b11111111111111111111100100010100;
assign LUT_4[1428] = 32'b00000000000000000011111110010100;
assign LUT_4[1429] = 32'b11111111111111111101001010001100;
assign LUT_4[1430] = 32'b00000000000000000011011000111000;
assign LUT_4[1431] = 32'b11111111111111111100100100110000;
assign LUT_4[1432] = 32'b00000000000000000000001010001101;
assign LUT_4[1433] = 32'b11111111111111111001010110000101;
assign LUT_4[1434] = 32'b11111111111111111111100100110001;
assign LUT_4[1435] = 32'b11111111111111111000110000101001;
assign LUT_4[1436] = 32'b11111111111111111101001010101001;
assign LUT_4[1437] = 32'b11111111111111110110010110100001;
assign LUT_4[1438] = 32'b11111111111111111100100101001101;
assign LUT_4[1439] = 32'b11111111111111110101110001000101;
assign LUT_4[1440] = 32'b00000000000000000111100111010001;
assign LUT_4[1441] = 32'b00000000000000000000110011001001;
assign LUT_4[1442] = 32'b00000000000000000111000001110101;
assign LUT_4[1443] = 32'b00000000000000000000001101101101;
assign LUT_4[1444] = 32'b00000000000000000100100111101101;
assign LUT_4[1445] = 32'b11111111111111111101110011100101;
assign LUT_4[1446] = 32'b00000000000000000100000010010001;
assign LUT_4[1447] = 32'b11111111111111111101001110001001;
assign LUT_4[1448] = 32'b00000000000000000000110011100110;
assign LUT_4[1449] = 32'b11111111111111111001111111011110;
assign LUT_4[1450] = 32'b00000000000000000000001110001010;
assign LUT_4[1451] = 32'b11111111111111111001011010000010;
assign LUT_4[1452] = 32'b11111111111111111101110100000010;
assign LUT_4[1453] = 32'b11111111111111110110111111111010;
assign LUT_4[1454] = 32'b11111111111111111101001110100110;
assign LUT_4[1455] = 32'b11111111111111110110011010011110;
assign LUT_4[1456] = 32'b00000000000000000101011000111111;
assign LUT_4[1457] = 32'b11111111111111111110100100110111;
assign LUT_4[1458] = 32'b00000000000000000100110011100011;
assign LUT_4[1459] = 32'b11111111111111111101111111011011;
assign LUT_4[1460] = 32'b00000000000000000010011001011011;
assign LUT_4[1461] = 32'b11111111111111111011100101010011;
assign LUT_4[1462] = 32'b00000000000000000001110011111111;
assign LUT_4[1463] = 32'b11111111111111111010111111110111;
assign LUT_4[1464] = 32'b11111111111111111110100101010100;
assign LUT_4[1465] = 32'b11111111111111110111110001001100;
assign LUT_4[1466] = 32'b11111111111111111101111111111000;
assign LUT_4[1467] = 32'b11111111111111110111001011110000;
assign LUT_4[1468] = 32'b11111111111111111011100101110000;
assign LUT_4[1469] = 32'b11111111111111110100110001101000;
assign LUT_4[1470] = 32'b11111111111111111011000000010100;
assign LUT_4[1471] = 32'b11111111111111110100001100001100;
assign LUT_4[1472] = 32'b00000000000000001010100011011110;
assign LUT_4[1473] = 32'b00000000000000000011101111010110;
assign LUT_4[1474] = 32'b00000000000000001001111110000010;
assign LUT_4[1475] = 32'b00000000000000000011001001111010;
assign LUT_4[1476] = 32'b00000000000000000111100011111010;
assign LUT_4[1477] = 32'b00000000000000000000101111110010;
assign LUT_4[1478] = 32'b00000000000000000110111110011110;
assign LUT_4[1479] = 32'b00000000000000000000001010010110;
assign LUT_4[1480] = 32'b00000000000000000011101111110011;
assign LUT_4[1481] = 32'b11111111111111111100111011101011;
assign LUT_4[1482] = 32'b00000000000000000011001010010111;
assign LUT_4[1483] = 32'b11111111111111111100010110001111;
assign LUT_4[1484] = 32'b00000000000000000000110000001111;
assign LUT_4[1485] = 32'b11111111111111111001111100000111;
assign LUT_4[1486] = 32'b00000000000000000000001010110011;
assign LUT_4[1487] = 32'b11111111111111111001010110101011;
assign LUT_4[1488] = 32'b00000000000000001000010101001100;
assign LUT_4[1489] = 32'b00000000000000000001100001000100;
assign LUT_4[1490] = 32'b00000000000000000111101111110000;
assign LUT_4[1491] = 32'b00000000000000000000111011101000;
assign LUT_4[1492] = 32'b00000000000000000101010101101000;
assign LUT_4[1493] = 32'b11111111111111111110100001100000;
assign LUT_4[1494] = 32'b00000000000000000100110000001100;
assign LUT_4[1495] = 32'b11111111111111111101111100000100;
assign LUT_4[1496] = 32'b00000000000000000001100001100001;
assign LUT_4[1497] = 32'b11111111111111111010101101011001;
assign LUT_4[1498] = 32'b00000000000000000000111100000101;
assign LUT_4[1499] = 32'b11111111111111111010000111111101;
assign LUT_4[1500] = 32'b11111111111111111110100001111101;
assign LUT_4[1501] = 32'b11111111111111110111101101110101;
assign LUT_4[1502] = 32'b11111111111111111101111100100001;
assign LUT_4[1503] = 32'b11111111111111110111001000011001;
assign LUT_4[1504] = 32'b00000000000000001000111110100101;
assign LUT_4[1505] = 32'b00000000000000000010001010011101;
assign LUT_4[1506] = 32'b00000000000000001000011001001001;
assign LUT_4[1507] = 32'b00000000000000000001100101000001;
assign LUT_4[1508] = 32'b00000000000000000101111111000001;
assign LUT_4[1509] = 32'b11111111111111111111001010111001;
assign LUT_4[1510] = 32'b00000000000000000101011001100101;
assign LUT_4[1511] = 32'b11111111111111111110100101011101;
assign LUT_4[1512] = 32'b00000000000000000010001010111010;
assign LUT_4[1513] = 32'b11111111111111111011010110110010;
assign LUT_4[1514] = 32'b00000000000000000001100101011110;
assign LUT_4[1515] = 32'b11111111111111111010110001010110;
assign LUT_4[1516] = 32'b11111111111111111111001011010110;
assign LUT_4[1517] = 32'b11111111111111111000010111001110;
assign LUT_4[1518] = 32'b11111111111111111110100101111010;
assign LUT_4[1519] = 32'b11111111111111110111110001110010;
assign LUT_4[1520] = 32'b00000000000000000110110000010011;
assign LUT_4[1521] = 32'b11111111111111111111111100001011;
assign LUT_4[1522] = 32'b00000000000000000110001010110111;
assign LUT_4[1523] = 32'b11111111111111111111010110101111;
assign LUT_4[1524] = 32'b00000000000000000011110000101111;
assign LUT_4[1525] = 32'b11111111111111111100111100100111;
assign LUT_4[1526] = 32'b00000000000000000011001011010011;
assign LUT_4[1527] = 32'b11111111111111111100010111001011;
assign LUT_4[1528] = 32'b11111111111111111111111100101000;
assign LUT_4[1529] = 32'b11111111111111111001001000100000;
assign LUT_4[1530] = 32'b11111111111111111111010111001100;
assign LUT_4[1531] = 32'b11111111111111111000100011000100;
assign LUT_4[1532] = 32'b11111111111111111100111101000100;
assign LUT_4[1533] = 32'b11111111111111110110001000111100;
assign LUT_4[1534] = 32'b11111111111111111100010111101000;
assign LUT_4[1535] = 32'b11111111111111110101100011100000;
assign LUT_4[1536] = 32'b00000000000000000000101110100111;
assign LUT_4[1537] = 32'b11111111111111111001111010011111;
assign LUT_4[1538] = 32'b00000000000000000000001001001011;
assign LUT_4[1539] = 32'b11111111111111111001010101000011;
assign LUT_4[1540] = 32'b11111111111111111101101111000011;
assign LUT_4[1541] = 32'b11111111111111110110111010111011;
assign LUT_4[1542] = 32'b11111111111111111101001001100111;
assign LUT_4[1543] = 32'b11111111111111110110010101011111;
assign LUT_4[1544] = 32'b11111111111111111001111010111100;
assign LUT_4[1545] = 32'b11111111111111110011000110110100;
assign LUT_4[1546] = 32'b11111111111111111001010101100000;
assign LUT_4[1547] = 32'b11111111111111110010100001011000;
assign LUT_4[1548] = 32'b11111111111111110110111011011000;
assign LUT_4[1549] = 32'b11111111111111110000000111010000;
assign LUT_4[1550] = 32'b11111111111111110110010101111100;
assign LUT_4[1551] = 32'b11111111111111101111100001110100;
assign LUT_4[1552] = 32'b11111111111111111110100000010101;
assign LUT_4[1553] = 32'b11111111111111110111101100001101;
assign LUT_4[1554] = 32'b11111111111111111101111010111001;
assign LUT_4[1555] = 32'b11111111111111110111000110110001;
assign LUT_4[1556] = 32'b11111111111111111011100000110001;
assign LUT_4[1557] = 32'b11111111111111110100101100101001;
assign LUT_4[1558] = 32'b11111111111111111010111011010101;
assign LUT_4[1559] = 32'b11111111111111110100000111001101;
assign LUT_4[1560] = 32'b11111111111111110111101100101010;
assign LUT_4[1561] = 32'b11111111111111110000111000100010;
assign LUT_4[1562] = 32'b11111111111111110111000111001110;
assign LUT_4[1563] = 32'b11111111111111110000010011000110;
assign LUT_4[1564] = 32'b11111111111111110100101101000110;
assign LUT_4[1565] = 32'b11111111111111101101111000111110;
assign LUT_4[1566] = 32'b11111111111111110100000111101010;
assign LUT_4[1567] = 32'b11111111111111101101010011100010;
assign LUT_4[1568] = 32'b11111111111111111111001001101110;
assign LUT_4[1569] = 32'b11111111111111111000010101100110;
assign LUT_4[1570] = 32'b11111111111111111110100100010010;
assign LUT_4[1571] = 32'b11111111111111110111110000001010;
assign LUT_4[1572] = 32'b11111111111111111100001010001010;
assign LUT_4[1573] = 32'b11111111111111110101010110000010;
assign LUT_4[1574] = 32'b11111111111111111011100100101110;
assign LUT_4[1575] = 32'b11111111111111110100110000100110;
assign LUT_4[1576] = 32'b11111111111111111000010110000011;
assign LUT_4[1577] = 32'b11111111111111110001100001111011;
assign LUT_4[1578] = 32'b11111111111111110111110000100111;
assign LUT_4[1579] = 32'b11111111111111110000111100011111;
assign LUT_4[1580] = 32'b11111111111111110101010110011111;
assign LUT_4[1581] = 32'b11111111111111101110100010010111;
assign LUT_4[1582] = 32'b11111111111111110100110001000011;
assign LUT_4[1583] = 32'b11111111111111101101111100111011;
assign LUT_4[1584] = 32'b11111111111111111100111011011100;
assign LUT_4[1585] = 32'b11111111111111110110000111010100;
assign LUT_4[1586] = 32'b11111111111111111100010110000000;
assign LUT_4[1587] = 32'b11111111111111110101100001111000;
assign LUT_4[1588] = 32'b11111111111111111001111011111000;
assign LUT_4[1589] = 32'b11111111111111110011000111110000;
assign LUT_4[1590] = 32'b11111111111111111001010110011100;
assign LUT_4[1591] = 32'b11111111111111110010100010010100;
assign LUT_4[1592] = 32'b11111111111111110110000111110001;
assign LUT_4[1593] = 32'b11111111111111101111010011101001;
assign LUT_4[1594] = 32'b11111111111111110101100010010101;
assign LUT_4[1595] = 32'b11111111111111101110101110001101;
assign LUT_4[1596] = 32'b11111111111111110011001000001101;
assign LUT_4[1597] = 32'b11111111111111101100010100000101;
assign LUT_4[1598] = 32'b11111111111111110010100010110001;
assign LUT_4[1599] = 32'b11111111111111101011101110101001;
assign LUT_4[1600] = 32'b00000000000000000010000101111011;
assign LUT_4[1601] = 32'b11111111111111111011010001110011;
assign LUT_4[1602] = 32'b00000000000000000001100000011111;
assign LUT_4[1603] = 32'b11111111111111111010101100010111;
assign LUT_4[1604] = 32'b11111111111111111111000110010111;
assign LUT_4[1605] = 32'b11111111111111111000010010001111;
assign LUT_4[1606] = 32'b11111111111111111110100000111011;
assign LUT_4[1607] = 32'b11111111111111110111101100110011;
assign LUT_4[1608] = 32'b11111111111111111011010010010000;
assign LUT_4[1609] = 32'b11111111111111110100011110001000;
assign LUT_4[1610] = 32'b11111111111111111010101100110100;
assign LUT_4[1611] = 32'b11111111111111110011111000101100;
assign LUT_4[1612] = 32'b11111111111111111000010010101100;
assign LUT_4[1613] = 32'b11111111111111110001011110100100;
assign LUT_4[1614] = 32'b11111111111111110111101101010000;
assign LUT_4[1615] = 32'b11111111111111110000111001001000;
assign LUT_4[1616] = 32'b11111111111111111111110111101001;
assign LUT_4[1617] = 32'b11111111111111111001000011100001;
assign LUT_4[1618] = 32'b11111111111111111111010010001101;
assign LUT_4[1619] = 32'b11111111111111111000011110000101;
assign LUT_4[1620] = 32'b11111111111111111100111000000101;
assign LUT_4[1621] = 32'b11111111111111110110000011111101;
assign LUT_4[1622] = 32'b11111111111111111100010010101001;
assign LUT_4[1623] = 32'b11111111111111110101011110100001;
assign LUT_4[1624] = 32'b11111111111111111001000011111110;
assign LUT_4[1625] = 32'b11111111111111110010001111110110;
assign LUT_4[1626] = 32'b11111111111111111000011110100010;
assign LUT_4[1627] = 32'b11111111111111110001101010011010;
assign LUT_4[1628] = 32'b11111111111111110110000100011010;
assign LUT_4[1629] = 32'b11111111111111101111010000010010;
assign LUT_4[1630] = 32'b11111111111111110101011110111110;
assign LUT_4[1631] = 32'b11111111111111101110101010110110;
assign LUT_4[1632] = 32'b00000000000000000000100001000010;
assign LUT_4[1633] = 32'b11111111111111111001101100111010;
assign LUT_4[1634] = 32'b11111111111111111111111011100110;
assign LUT_4[1635] = 32'b11111111111111111001000111011110;
assign LUT_4[1636] = 32'b11111111111111111101100001011110;
assign LUT_4[1637] = 32'b11111111111111110110101101010110;
assign LUT_4[1638] = 32'b11111111111111111100111100000010;
assign LUT_4[1639] = 32'b11111111111111110110000111111010;
assign LUT_4[1640] = 32'b11111111111111111001101101010111;
assign LUT_4[1641] = 32'b11111111111111110010111001001111;
assign LUT_4[1642] = 32'b11111111111111111001000111111011;
assign LUT_4[1643] = 32'b11111111111111110010010011110011;
assign LUT_4[1644] = 32'b11111111111111110110101101110011;
assign LUT_4[1645] = 32'b11111111111111101111111001101011;
assign LUT_4[1646] = 32'b11111111111111110110001000010111;
assign LUT_4[1647] = 32'b11111111111111101111010100001111;
assign LUT_4[1648] = 32'b11111111111111111110010010110000;
assign LUT_4[1649] = 32'b11111111111111110111011110101000;
assign LUT_4[1650] = 32'b11111111111111111101101101010100;
assign LUT_4[1651] = 32'b11111111111111110110111001001100;
assign LUT_4[1652] = 32'b11111111111111111011010011001100;
assign LUT_4[1653] = 32'b11111111111111110100011111000100;
assign LUT_4[1654] = 32'b11111111111111111010101101110000;
assign LUT_4[1655] = 32'b11111111111111110011111001101000;
assign LUT_4[1656] = 32'b11111111111111110111011111000101;
assign LUT_4[1657] = 32'b11111111111111110000101010111101;
assign LUT_4[1658] = 32'b11111111111111110110111001101001;
assign LUT_4[1659] = 32'b11111111111111110000000101100001;
assign LUT_4[1660] = 32'b11111111111111110100011111100001;
assign LUT_4[1661] = 32'b11111111111111101101101011011001;
assign LUT_4[1662] = 32'b11111111111111110011111010000101;
assign LUT_4[1663] = 32'b11111111111111101101000101111101;
assign LUT_4[1664] = 32'b00000000000000000011010100101111;
assign LUT_4[1665] = 32'b11111111111111111100100000100111;
assign LUT_4[1666] = 32'b00000000000000000010101111010011;
assign LUT_4[1667] = 32'b11111111111111111011111011001011;
assign LUT_4[1668] = 32'b00000000000000000000010101001011;
assign LUT_4[1669] = 32'b11111111111111111001100001000011;
assign LUT_4[1670] = 32'b11111111111111111111101111101111;
assign LUT_4[1671] = 32'b11111111111111111000111011100111;
assign LUT_4[1672] = 32'b11111111111111111100100001000100;
assign LUT_4[1673] = 32'b11111111111111110101101100111100;
assign LUT_4[1674] = 32'b11111111111111111011111011101000;
assign LUT_4[1675] = 32'b11111111111111110101000111100000;
assign LUT_4[1676] = 32'b11111111111111111001100001100000;
assign LUT_4[1677] = 32'b11111111111111110010101101011000;
assign LUT_4[1678] = 32'b11111111111111111000111100000100;
assign LUT_4[1679] = 32'b11111111111111110010000111111100;
assign LUT_4[1680] = 32'b00000000000000000001000110011101;
assign LUT_4[1681] = 32'b11111111111111111010010010010101;
assign LUT_4[1682] = 32'b00000000000000000000100001000001;
assign LUT_4[1683] = 32'b11111111111111111001101100111001;
assign LUT_4[1684] = 32'b11111111111111111110000110111001;
assign LUT_4[1685] = 32'b11111111111111110111010010110001;
assign LUT_4[1686] = 32'b11111111111111111101100001011101;
assign LUT_4[1687] = 32'b11111111111111110110101101010101;
assign LUT_4[1688] = 32'b11111111111111111010010010110010;
assign LUT_4[1689] = 32'b11111111111111110011011110101010;
assign LUT_4[1690] = 32'b11111111111111111001101101010110;
assign LUT_4[1691] = 32'b11111111111111110010111001001110;
assign LUT_4[1692] = 32'b11111111111111110111010011001110;
assign LUT_4[1693] = 32'b11111111111111110000011111000110;
assign LUT_4[1694] = 32'b11111111111111110110101101110010;
assign LUT_4[1695] = 32'b11111111111111101111111001101010;
assign LUT_4[1696] = 32'b00000000000000000001101111110110;
assign LUT_4[1697] = 32'b11111111111111111010111011101110;
assign LUT_4[1698] = 32'b00000000000000000001001010011010;
assign LUT_4[1699] = 32'b11111111111111111010010110010010;
assign LUT_4[1700] = 32'b11111111111111111110110000010010;
assign LUT_4[1701] = 32'b11111111111111110111111100001010;
assign LUT_4[1702] = 32'b11111111111111111110001010110110;
assign LUT_4[1703] = 32'b11111111111111110111010110101110;
assign LUT_4[1704] = 32'b11111111111111111010111100001011;
assign LUT_4[1705] = 32'b11111111111111110100001000000011;
assign LUT_4[1706] = 32'b11111111111111111010010110101111;
assign LUT_4[1707] = 32'b11111111111111110011100010100111;
assign LUT_4[1708] = 32'b11111111111111110111111100100111;
assign LUT_4[1709] = 32'b11111111111111110001001000011111;
assign LUT_4[1710] = 32'b11111111111111110111010111001011;
assign LUT_4[1711] = 32'b11111111111111110000100011000011;
assign LUT_4[1712] = 32'b11111111111111111111100001100100;
assign LUT_4[1713] = 32'b11111111111111111000101101011100;
assign LUT_4[1714] = 32'b11111111111111111110111100001000;
assign LUT_4[1715] = 32'b11111111111111111000001000000000;
assign LUT_4[1716] = 32'b11111111111111111100100010000000;
assign LUT_4[1717] = 32'b11111111111111110101101101111000;
assign LUT_4[1718] = 32'b11111111111111111011111100100100;
assign LUT_4[1719] = 32'b11111111111111110101001000011100;
assign LUT_4[1720] = 32'b11111111111111111000101101111001;
assign LUT_4[1721] = 32'b11111111111111110001111001110001;
assign LUT_4[1722] = 32'b11111111111111111000001000011101;
assign LUT_4[1723] = 32'b11111111111111110001010100010101;
assign LUT_4[1724] = 32'b11111111111111110101101110010101;
assign LUT_4[1725] = 32'b11111111111111101110111010001101;
assign LUT_4[1726] = 32'b11111111111111110101001000111001;
assign LUT_4[1727] = 32'b11111111111111101110010100110001;
assign LUT_4[1728] = 32'b00000000000000000100101100000011;
assign LUT_4[1729] = 32'b11111111111111111101110111111011;
assign LUT_4[1730] = 32'b00000000000000000100000110100111;
assign LUT_4[1731] = 32'b11111111111111111101010010011111;
assign LUT_4[1732] = 32'b00000000000000000001101100011111;
assign LUT_4[1733] = 32'b11111111111111111010111000010111;
assign LUT_4[1734] = 32'b00000000000000000001000111000011;
assign LUT_4[1735] = 32'b11111111111111111010010010111011;
assign LUT_4[1736] = 32'b11111111111111111101111000011000;
assign LUT_4[1737] = 32'b11111111111111110111000100010000;
assign LUT_4[1738] = 32'b11111111111111111101010010111100;
assign LUT_4[1739] = 32'b11111111111111110110011110110100;
assign LUT_4[1740] = 32'b11111111111111111010111000110100;
assign LUT_4[1741] = 32'b11111111111111110100000100101100;
assign LUT_4[1742] = 32'b11111111111111111010010011011000;
assign LUT_4[1743] = 32'b11111111111111110011011111010000;
assign LUT_4[1744] = 32'b00000000000000000010011101110001;
assign LUT_4[1745] = 32'b11111111111111111011101001101001;
assign LUT_4[1746] = 32'b00000000000000000001111000010101;
assign LUT_4[1747] = 32'b11111111111111111011000100001101;
assign LUT_4[1748] = 32'b11111111111111111111011110001101;
assign LUT_4[1749] = 32'b11111111111111111000101010000101;
assign LUT_4[1750] = 32'b11111111111111111110111000110001;
assign LUT_4[1751] = 32'b11111111111111111000000100101001;
assign LUT_4[1752] = 32'b11111111111111111011101010000110;
assign LUT_4[1753] = 32'b11111111111111110100110101111110;
assign LUT_4[1754] = 32'b11111111111111111011000100101010;
assign LUT_4[1755] = 32'b11111111111111110100010000100010;
assign LUT_4[1756] = 32'b11111111111111111000101010100010;
assign LUT_4[1757] = 32'b11111111111111110001110110011010;
assign LUT_4[1758] = 32'b11111111111111111000000101000110;
assign LUT_4[1759] = 32'b11111111111111110001010000111110;
assign LUT_4[1760] = 32'b00000000000000000011000111001010;
assign LUT_4[1761] = 32'b11111111111111111100010011000010;
assign LUT_4[1762] = 32'b00000000000000000010100001101110;
assign LUT_4[1763] = 32'b11111111111111111011101101100110;
assign LUT_4[1764] = 32'b00000000000000000000000111100110;
assign LUT_4[1765] = 32'b11111111111111111001010011011110;
assign LUT_4[1766] = 32'b11111111111111111111100010001010;
assign LUT_4[1767] = 32'b11111111111111111000101110000010;
assign LUT_4[1768] = 32'b11111111111111111100010011011111;
assign LUT_4[1769] = 32'b11111111111111110101011111010111;
assign LUT_4[1770] = 32'b11111111111111111011101110000011;
assign LUT_4[1771] = 32'b11111111111111110100111001111011;
assign LUT_4[1772] = 32'b11111111111111111001010011111011;
assign LUT_4[1773] = 32'b11111111111111110010011111110011;
assign LUT_4[1774] = 32'b11111111111111111000101110011111;
assign LUT_4[1775] = 32'b11111111111111110001111010010111;
assign LUT_4[1776] = 32'b00000000000000000000111000111000;
assign LUT_4[1777] = 32'b11111111111111111010000100110000;
assign LUT_4[1778] = 32'b00000000000000000000010011011100;
assign LUT_4[1779] = 32'b11111111111111111001011111010100;
assign LUT_4[1780] = 32'b11111111111111111101111001010100;
assign LUT_4[1781] = 32'b11111111111111110111000101001100;
assign LUT_4[1782] = 32'b11111111111111111101010011111000;
assign LUT_4[1783] = 32'b11111111111111110110011111110000;
assign LUT_4[1784] = 32'b11111111111111111010000101001101;
assign LUT_4[1785] = 32'b11111111111111110011010001000101;
assign LUT_4[1786] = 32'b11111111111111111001011111110001;
assign LUT_4[1787] = 32'b11111111111111110010101011101001;
assign LUT_4[1788] = 32'b11111111111111110111000101101001;
assign LUT_4[1789] = 32'b11111111111111110000010001100001;
assign LUT_4[1790] = 32'b11111111111111110110100000001101;
assign LUT_4[1791] = 32'b11111111111111101111101100000101;
assign LUT_4[1792] = 32'b00000000000000000101101010001010;
assign LUT_4[1793] = 32'b11111111111111111110110110000010;
assign LUT_4[1794] = 32'b00000000000000000101000100101110;
assign LUT_4[1795] = 32'b11111111111111111110010000100110;
assign LUT_4[1796] = 32'b00000000000000000010101010100110;
assign LUT_4[1797] = 32'b11111111111111111011110110011110;
assign LUT_4[1798] = 32'b00000000000000000010000101001010;
assign LUT_4[1799] = 32'b11111111111111111011010001000010;
assign LUT_4[1800] = 32'b11111111111111111110110110011111;
assign LUT_4[1801] = 32'b11111111111111111000000010010111;
assign LUT_4[1802] = 32'b11111111111111111110010001000011;
assign LUT_4[1803] = 32'b11111111111111110111011100111011;
assign LUT_4[1804] = 32'b11111111111111111011110110111011;
assign LUT_4[1805] = 32'b11111111111111110101000010110011;
assign LUT_4[1806] = 32'b11111111111111111011010001011111;
assign LUT_4[1807] = 32'b11111111111111110100011101010111;
assign LUT_4[1808] = 32'b00000000000000000011011011111000;
assign LUT_4[1809] = 32'b11111111111111111100100111110000;
assign LUT_4[1810] = 32'b00000000000000000010110110011100;
assign LUT_4[1811] = 32'b11111111111111111100000010010100;
assign LUT_4[1812] = 32'b00000000000000000000011100010100;
assign LUT_4[1813] = 32'b11111111111111111001101000001100;
assign LUT_4[1814] = 32'b11111111111111111111110110111000;
assign LUT_4[1815] = 32'b11111111111111111001000010110000;
assign LUT_4[1816] = 32'b11111111111111111100101000001101;
assign LUT_4[1817] = 32'b11111111111111110101110100000101;
assign LUT_4[1818] = 32'b11111111111111111100000010110001;
assign LUT_4[1819] = 32'b11111111111111110101001110101001;
assign LUT_4[1820] = 32'b11111111111111111001101000101001;
assign LUT_4[1821] = 32'b11111111111111110010110100100001;
assign LUT_4[1822] = 32'b11111111111111111001000011001101;
assign LUT_4[1823] = 32'b11111111111111110010001111000101;
assign LUT_4[1824] = 32'b00000000000000000100000101010001;
assign LUT_4[1825] = 32'b11111111111111111101010001001001;
assign LUT_4[1826] = 32'b00000000000000000011011111110101;
assign LUT_4[1827] = 32'b11111111111111111100101011101101;
assign LUT_4[1828] = 32'b00000000000000000001000101101101;
assign LUT_4[1829] = 32'b11111111111111111010010001100101;
assign LUT_4[1830] = 32'b00000000000000000000100000010001;
assign LUT_4[1831] = 32'b11111111111111111001101100001001;
assign LUT_4[1832] = 32'b11111111111111111101010001100110;
assign LUT_4[1833] = 32'b11111111111111110110011101011110;
assign LUT_4[1834] = 32'b11111111111111111100101100001010;
assign LUT_4[1835] = 32'b11111111111111110101111000000010;
assign LUT_4[1836] = 32'b11111111111111111010010010000010;
assign LUT_4[1837] = 32'b11111111111111110011011101111010;
assign LUT_4[1838] = 32'b11111111111111111001101100100110;
assign LUT_4[1839] = 32'b11111111111111110010111000011110;
assign LUT_4[1840] = 32'b00000000000000000001110110111111;
assign LUT_4[1841] = 32'b11111111111111111011000010110111;
assign LUT_4[1842] = 32'b00000000000000000001010001100011;
assign LUT_4[1843] = 32'b11111111111111111010011101011011;
assign LUT_4[1844] = 32'b11111111111111111110110111011011;
assign LUT_4[1845] = 32'b11111111111111111000000011010011;
assign LUT_4[1846] = 32'b11111111111111111110010001111111;
assign LUT_4[1847] = 32'b11111111111111110111011101110111;
assign LUT_4[1848] = 32'b11111111111111111011000011010100;
assign LUT_4[1849] = 32'b11111111111111110100001111001100;
assign LUT_4[1850] = 32'b11111111111111111010011101111000;
assign LUT_4[1851] = 32'b11111111111111110011101001110000;
assign LUT_4[1852] = 32'b11111111111111111000000011110000;
assign LUT_4[1853] = 32'b11111111111111110001001111101000;
assign LUT_4[1854] = 32'b11111111111111110111011110010100;
assign LUT_4[1855] = 32'b11111111111111110000101010001100;
assign LUT_4[1856] = 32'b00000000000000000111000001011110;
assign LUT_4[1857] = 32'b00000000000000000000001101010110;
assign LUT_4[1858] = 32'b00000000000000000110011100000010;
assign LUT_4[1859] = 32'b11111111111111111111100111111010;
assign LUT_4[1860] = 32'b00000000000000000100000001111010;
assign LUT_4[1861] = 32'b11111111111111111101001101110010;
assign LUT_4[1862] = 32'b00000000000000000011011100011110;
assign LUT_4[1863] = 32'b11111111111111111100101000010110;
assign LUT_4[1864] = 32'b00000000000000000000001101110011;
assign LUT_4[1865] = 32'b11111111111111111001011001101011;
assign LUT_4[1866] = 32'b11111111111111111111101000010111;
assign LUT_4[1867] = 32'b11111111111111111000110100001111;
assign LUT_4[1868] = 32'b11111111111111111101001110001111;
assign LUT_4[1869] = 32'b11111111111111110110011010000111;
assign LUT_4[1870] = 32'b11111111111111111100101000110011;
assign LUT_4[1871] = 32'b11111111111111110101110100101011;
assign LUT_4[1872] = 32'b00000000000000000100110011001100;
assign LUT_4[1873] = 32'b11111111111111111101111111000100;
assign LUT_4[1874] = 32'b00000000000000000100001101110000;
assign LUT_4[1875] = 32'b11111111111111111101011001101000;
assign LUT_4[1876] = 32'b00000000000000000001110011101000;
assign LUT_4[1877] = 32'b11111111111111111010111111100000;
assign LUT_4[1878] = 32'b00000000000000000001001110001100;
assign LUT_4[1879] = 32'b11111111111111111010011010000100;
assign LUT_4[1880] = 32'b11111111111111111101111111100001;
assign LUT_4[1881] = 32'b11111111111111110111001011011001;
assign LUT_4[1882] = 32'b11111111111111111101011010000101;
assign LUT_4[1883] = 32'b11111111111111110110100101111101;
assign LUT_4[1884] = 32'b11111111111111111010111111111101;
assign LUT_4[1885] = 32'b11111111111111110100001011110101;
assign LUT_4[1886] = 32'b11111111111111111010011010100001;
assign LUT_4[1887] = 32'b11111111111111110011100110011001;
assign LUT_4[1888] = 32'b00000000000000000101011100100101;
assign LUT_4[1889] = 32'b11111111111111111110101000011101;
assign LUT_4[1890] = 32'b00000000000000000100110111001001;
assign LUT_4[1891] = 32'b11111111111111111110000011000001;
assign LUT_4[1892] = 32'b00000000000000000010011101000001;
assign LUT_4[1893] = 32'b11111111111111111011101000111001;
assign LUT_4[1894] = 32'b00000000000000000001110111100101;
assign LUT_4[1895] = 32'b11111111111111111011000011011101;
assign LUT_4[1896] = 32'b11111111111111111110101000111010;
assign LUT_4[1897] = 32'b11111111111111110111110100110010;
assign LUT_4[1898] = 32'b11111111111111111110000011011110;
assign LUT_4[1899] = 32'b11111111111111110111001111010110;
assign LUT_4[1900] = 32'b11111111111111111011101001010110;
assign LUT_4[1901] = 32'b11111111111111110100110101001110;
assign LUT_4[1902] = 32'b11111111111111111011000011111010;
assign LUT_4[1903] = 32'b11111111111111110100001111110010;
assign LUT_4[1904] = 32'b00000000000000000011001110010011;
assign LUT_4[1905] = 32'b11111111111111111100011010001011;
assign LUT_4[1906] = 32'b00000000000000000010101000110111;
assign LUT_4[1907] = 32'b11111111111111111011110100101111;
assign LUT_4[1908] = 32'b00000000000000000000001110101111;
assign LUT_4[1909] = 32'b11111111111111111001011010100111;
assign LUT_4[1910] = 32'b11111111111111111111101001010011;
assign LUT_4[1911] = 32'b11111111111111111000110101001011;
assign LUT_4[1912] = 32'b11111111111111111100011010101000;
assign LUT_4[1913] = 32'b11111111111111110101100110100000;
assign LUT_4[1914] = 32'b11111111111111111011110101001100;
assign LUT_4[1915] = 32'b11111111111111110101000001000100;
assign LUT_4[1916] = 32'b11111111111111111001011011000100;
assign LUT_4[1917] = 32'b11111111111111110010100110111100;
assign LUT_4[1918] = 32'b11111111111111111000110101101000;
assign LUT_4[1919] = 32'b11111111111111110010000001100000;
assign LUT_4[1920] = 32'b00000000000000001000010000010010;
assign LUT_4[1921] = 32'b00000000000000000001011100001010;
assign LUT_4[1922] = 32'b00000000000000000111101010110110;
assign LUT_4[1923] = 32'b00000000000000000000110110101110;
assign LUT_4[1924] = 32'b00000000000000000101010000101110;
assign LUT_4[1925] = 32'b11111111111111111110011100100110;
assign LUT_4[1926] = 32'b00000000000000000100101011010010;
assign LUT_4[1927] = 32'b11111111111111111101110111001010;
assign LUT_4[1928] = 32'b00000000000000000001011100100111;
assign LUT_4[1929] = 32'b11111111111111111010101000011111;
assign LUT_4[1930] = 32'b00000000000000000000110111001011;
assign LUT_4[1931] = 32'b11111111111111111010000011000011;
assign LUT_4[1932] = 32'b11111111111111111110011101000011;
assign LUT_4[1933] = 32'b11111111111111110111101000111011;
assign LUT_4[1934] = 32'b11111111111111111101110111100111;
assign LUT_4[1935] = 32'b11111111111111110111000011011111;
assign LUT_4[1936] = 32'b00000000000000000110000010000000;
assign LUT_4[1937] = 32'b11111111111111111111001101111000;
assign LUT_4[1938] = 32'b00000000000000000101011100100100;
assign LUT_4[1939] = 32'b11111111111111111110101000011100;
assign LUT_4[1940] = 32'b00000000000000000011000010011100;
assign LUT_4[1941] = 32'b11111111111111111100001110010100;
assign LUT_4[1942] = 32'b00000000000000000010011101000000;
assign LUT_4[1943] = 32'b11111111111111111011101000111000;
assign LUT_4[1944] = 32'b11111111111111111111001110010101;
assign LUT_4[1945] = 32'b11111111111111111000011010001101;
assign LUT_4[1946] = 32'b11111111111111111110101000111001;
assign LUT_4[1947] = 32'b11111111111111110111110100110001;
assign LUT_4[1948] = 32'b11111111111111111100001110110001;
assign LUT_4[1949] = 32'b11111111111111110101011010101001;
assign LUT_4[1950] = 32'b11111111111111111011101001010101;
assign LUT_4[1951] = 32'b11111111111111110100110101001101;
assign LUT_4[1952] = 32'b00000000000000000110101011011001;
assign LUT_4[1953] = 32'b11111111111111111111110111010001;
assign LUT_4[1954] = 32'b00000000000000000110000101111101;
assign LUT_4[1955] = 32'b11111111111111111111010001110101;
assign LUT_4[1956] = 32'b00000000000000000011101011110101;
assign LUT_4[1957] = 32'b11111111111111111100110111101101;
assign LUT_4[1958] = 32'b00000000000000000011000110011001;
assign LUT_4[1959] = 32'b11111111111111111100010010010001;
assign LUT_4[1960] = 32'b11111111111111111111110111101110;
assign LUT_4[1961] = 32'b11111111111111111001000011100110;
assign LUT_4[1962] = 32'b11111111111111111111010010010010;
assign LUT_4[1963] = 32'b11111111111111111000011110001010;
assign LUT_4[1964] = 32'b11111111111111111100111000001010;
assign LUT_4[1965] = 32'b11111111111111110110000100000010;
assign LUT_4[1966] = 32'b11111111111111111100010010101110;
assign LUT_4[1967] = 32'b11111111111111110101011110100110;
assign LUT_4[1968] = 32'b00000000000000000100011101000111;
assign LUT_4[1969] = 32'b11111111111111111101101000111111;
assign LUT_4[1970] = 32'b00000000000000000011110111101011;
assign LUT_4[1971] = 32'b11111111111111111101000011100011;
assign LUT_4[1972] = 32'b00000000000000000001011101100011;
assign LUT_4[1973] = 32'b11111111111111111010101001011011;
assign LUT_4[1974] = 32'b00000000000000000000111000000111;
assign LUT_4[1975] = 32'b11111111111111111010000011111111;
assign LUT_4[1976] = 32'b11111111111111111101101001011100;
assign LUT_4[1977] = 32'b11111111111111110110110101010100;
assign LUT_4[1978] = 32'b11111111111111111101000100000000;
assign LUT_4[1979] = 32'b11111111111111110110001111111000;
assign LUT_4[1980] = 32'b11111111111111111010101001111000;
assign LUT_4[1981] = 32'b11111111111111110011110101110000;
assign LUT_4[1982] = 32'b11111111111111111010000100011100;
assign LUT_4[1983] = 32'b11111111111111110011010000010100;
assign LUT_4[1984] = 32'b00000000000000001001100111100110;
assign LUT_4[1985] = 32'b00000000000000000010110011011110;
assign LUT_4[1986] = 32'b00000000000000001001000010001010;
assign LUT_4[1987] = 32'b00000000000000000010001110000010;
assign LUT_4[1988] = 32'b00000000000000000110101000000010;
assign LUT_4[1989] = 32'b11111111111111111111110011111010;
assign LUT_4[1990] = 32'b00000000000000000110000010100110;
assign LUT_4[1991] = 32'b11111111111111111111001110011110;
assign LUT_4[1992] = 32'b00000000000000000010110011111011;
assign LUT_4[1993] = 32'b11111111111111111011111111110011;
assign LUT_4[1994] = 32'b00000000000000000010001110011111;
assign LUT_4[1995] = 32'b11111111111111111011011010010111;
assign LUT_4[1996] = 32'b11111111111111111111110100010111;
assign LUT_4[1997] = 32'b11111111111111111001000000001111;
assign LUT_4[1998] = 32'b11111111111111111111001110111011;
assign LUT_4[1999] = 32'b11111111111111111000011010110011;
assign LUT_4[2000] = 32'b00000000000000000111011001010100;
assign LUT_4[2001] = 32'b00000000000000000000100101001100;
assign LUT_4[2002] = 32'b00000000000000000110110011111000;
assign LUT_4[2003] = 32'b11111111111111111111111111110000;
assign LUT_4[2004] = 32'b00000000000000000100011001110000;
assign LUT_4[2005] = 32'b11111111111111111101100101101000;
assign LUT_4[2006] = 32'b00000000000000000011110100010100;
assign LUT_4[2007] = 32'b11111111111111111101000000001100;
assign LUT_4[2008] = 32'b00000000000000000000100101101001;
assign LUT_4[2009] = 32'b11111111111111111001110001100001;
assign LUT_4[2010] = 32'b00000000000000000000000000001101;
assign LUT_4[2011] = 32'b11111111111111111001001100000101;
assign LUT_4[2012] = 32'b11111111111111111101100110000101;
assign LUT_4[2013] = 32'b11111111111111110110110001111101;
assign LUT_4[2014] = 32'b11111111111111111101000000101001;
assign LUT_4[2015] = 32'b11111111111111110110001100100001;
assign LUT_4[2016] = 32'b00000000000000001000000010101101;
assign LUT_4[2017] = 32'b00000000000000000001001110100101;
assign LUT_4[2018] = 32'b00000000000000000111011101010001;
assign LUT_4[2019] = 32'b00000000000000000000101001001001;
assign LUT_4[2020] = 32'b00000000000000000101000011001001;
assign LUT_4[2021] = 32'b11111111111111111110001111000001;
assign LUT_4[2022] = 32'b00000000000000000100011101101101;
assign LUT_4[2023] = 32'b11111111111111111101101001100101;
assign LUT_4[2024] = 32'b00000000000000000001001111000010;
assign LUT_4[2025] = 32'b11111111111111111010011010111010;
assign LUT_4[2026] = 32'b00000000000000000000101001100110;
assign LUT_4[2027] = 32'b11111111111111111001110101011110;
assign LUT_4[2028] = 32'b11111111111111111110001111011110;
assign LUT_4[2029] = 32'b11111111111111110111011011010110;
assign LUT_4[2030] = 32'b11111111111111111101101010000010;
assign LUT_4[2031] = 32'b11111111111111110110110101111010;
assign LUT_4[2032] = 32'b00000000000000000101110100011011;
assign LUT_4[2033] = 32'b11111111111111111111000000010011;
assign LUT_4[2034] = 32'b00000000000000000101001110111111;
assign LUT_4[2035] = 32'b11111111111111111110011010110111;
assign LUT_4[2036] = 32'b00000000000000000010110100110111;
assign LUT_4[2037] = 32'b11111111111111111100000000101111;
assign LUT_4[2038] = 32'b00000000000000000010001111011011;
assign LUT_4[2039] = 32'b11111111111111111011011011010011;
assign LUT_4[2040] = 32'b11111111111111111111000000110000;
assign LUT_4[2041] = 32'b11111111111111111000001100101000;
assign LUT_4[2042] = 32'b11111111111111111110011011010100;
assign LUT_4[2043] = 32'b11111111111111110111100111001100;
assign LUT_4[2044] = 32'b11111111111111111100000001001100;
assign LUT_4[2045] = 32'b11111111111111110101001101000100;
assign LUT_4[2046] = 32'b11111111111111111011011011110000;
assign LUT_4[2047] = 32'b11111111111111110100100111101000;
assign LUT_4[2048] = 32'b11111111111111111011011111001010;
assign LUT_4[2049] = 32'b11111111111111110100101011000010;
assign LUT_4[2050] = 32'b11111111111111111010111001101110;
assign LUT_4[2051] = 32'b11111111111111110100000101100110;
assign LUT_4[2052] = 32'b11111111111111111000011111100110;
assign LUT_4[2053] = 32'b11111111111111110001101011011110;
assign LUT_4[2054] = 32'b11111111111111110111111010001010;
assign LUT_4[2055] = 32'b11111111111111110001000110000010;
assign LUT_4[2056] = 32'b11111111111111110100101011011111;
assign LUT_4[2057] = 32'b11111111111111101101110111010111;
assign LUT_4[2058] = 32'b11111111111111110100000110000011;
assign LUT_4[2059] = 32'b11111111111111101101010001111011;
assign LUT_4[2060] = 32'b11111111111111110001101011111011;
assign LUT_4[2061] = 32'b11111111111111101010110111110011;
assign LUT_4[2062] = 32'b11111111111111110001000110011111;
assign LUT_4[2063] = 32'b11111111111111101010010010010111;
assign LUT_4[2064] = 32'b11111111111111111001010000111000;
assign LUT_4[2065] = 32'b11111111111111110010011100110000;
assign LUT_4[2066] = 32'b11111111111111111000101011011100;
assign LUT_4[2067] = 32'b11111111111111110001110111010100;
assign LUT_4[2068] = 32'b11111111111111110110010001010100;
assign LUT_4[2069] = 32'b11111111111111101111011101001100;
assign LUT_4[2070] = 32'b11111111111111110101101011111000;
assign LUT_4[2071] = 32'b11111111111111101110110111110000;
assign LUT_4[2072] = 32'b11111111111111110010011101001101;
assign LUT_4[2073] = 32'b11111111111111101011101001000101;
assign LUT_4[2074] = 32'b11111111111111110001110111110001;
assign LUT_4[2075] = 32'b11111111111111101011000011101001;
assign LUT_4[2076] = 32'b11111111111111101111011101101001;
assign LUT_4[2077] = 32'b11111111111111101000101001100001;
assign LUT_4[2078] = 32'b11111111111111101110111000001101;
assign LUT_4[2079] = 32'b11111111111111101000000100000101;
assign LUT_4[2080] = 32'b11111111111111111001111010010001;
assign LUT_4[2081] = 32'b11111111111111110011000110001001;
assign LUT_4[2082] = 32'b11111111111111111001010100110101;
assign LUT_4[2083] = 32'b11111111111111110010100000101101;
assign LUT_4[2084] = 32'b11111111111111110110111010101101;
assign LUT_4[2085] = 32'b11111111111111110000000110100101;
assign LUT_4[2086] = 32'b11111111111111110110010101010001;
assign LUT_4[2087] = 32'b11111111111111101111100001001001;
assign LUT_4[2088] = 32'b11111111111111110011000110100110;
assign LUT_4[2089] = 32'b11111111111111101100010010011110;
assign LUT_4[2090] = 32'b11111111111111110010100001001010;
assign LUT_4[2091] = 32'b11111111111111101011101101000010;
assign LUT_4[2092] = 32'b11111111111111110000000111000010;
assign LUT_4[2093] = 32'b11111111111111101001010010111010;
assign LUT_4[2094] = 32'b11111111111111101111100001100110;
assign LUT_4[2095] = 32'b11111111111111101000101101011110;
assign LUT_4[2096] = 32'b11111111111111110111101011111111;
assign LUT_4[2097] = 32'b11111111111111110000110111110111;
assign LUT_4[2098] = 32'b11111111111111110111000110100011;
assign LUT_4[2099] = 32'b11111111111111110000010010011011;
assign LUT_4[2100] = 32'b11111111111111110100101100011011;
assign LUT_4[2101] = 32'b11111111111111101101111000010011;
assign LUT_4[2102] = 32'b11111111111111110100000110111111;
assign LUT_4[2103] = 32'b11111111111111101101010010110111;
assign LUT_4[2104] = 32'b11111111111111110000111000010100;
assign LUT_4[2105] = 32'b11111111111111101010000100001100;
assign LUT_4[2106] = 32'b11111111111111110000010010111000;
assign LUT_4[2107] = 32'b11111111111111101001011110110000;
assign LUT_4[2108] = 32'b11111111111111101101111000110000;
assign LUT_4[2109] = 32'b11111111111111100111000100101000;
assign LUT_4[2110] = 32'b11111111111111101101010011010100;
assign LUT_4[2111] = 32'b11111111111111100110011111001100;
assign LUT_4[2112] = 32'b11111111111111111100110110011110;
assign LUT_4[2113] = 32'b11111111111111110110000010010110;
assign LUT_4[2114] = 32'b11111111111111111100010001000010;
assign LUT_4[2115] = 32'b11111111111111110101011100111010;
assign LUT_4[2116] = 32'b11111111111111111001110110111010;
assign LUT_4[2117] = 32'b11111111111111110011000010110010;
assign LUT_4[2118] = 32'b11111111111111111001010001011110;
assign LUT_4[2119] = 32'b11111111111111110010011101010110;
assign LUT_4[2120] = 32'b11111111111111110110000010110011;
assign LUT_4[2121] = 32'b11111111111111101111001110101011;
assign LUT_4[2122] = 32'b11111111111111110101011101010111;
assign LUT_4[2123] = 32'b11111111111111101110101001001111;
assign LUT_4[2124] = 32'b11111111111111110011000011001111;
assign LUT_4[2125] = 32'b11111111111111101100001111000111;
assign LUT_4[2126] = 32'b11111111111111110010011101110011;
assign LUT_4[2127] = 32'b11111111111111101011101001101011;
assign LUT_4[2128] = 32'b11111111111111111010101000001100;
assign LUT_4[2129] = 32'b11111111111111110011110100000100;
assign LUT_4[2130] = 32'b11111111111111111010000010110000;
assign LUT_4[2131] = 32'b11111111111111110011001110101000;
assign LUT_4[2132] = 32'b11111111111111110111101000101000;
assign LUT_4[2133] = 32'b11111111111111110000110100100000;
assign LUT_4[2134] = 32'b11111111111111110111000011001100;
assign LUT_4[2135] = 32'b11111111111111110000001111000100;
assign LUT_4[2136] = 32'b11111111111111110011110100100001;
assign LUT_4[2137] = 32'b11111111111111101101000000011001;
assign LUT_4[2138] = 32'b11111111111111110011001111000101;
assign LUT_4[2139] = 32'b11111111111111101100011010111101;
assign LUT_4[2140] = 32'b11111111111111110000110100111101;
assign LUT_4[2141] = 32'b11111111111111101010000000110101;
assign LUT_4[2142] = 32'b11111111111111110000001111100001;
assign LUT_4[2143] = 32'b11111111111111101001011011011001;
assign LUT_4[2144] = 32'b11111111111111111011010001100101;
assign LUT_4[2145] = 32'b11111111111111110100011101011101;
assign LUT_4[2146] = 32'b11111111111111111010101100001001;
assign LUT_4[2147] = 32'b11111111111111110011111000000001;
assign LUT_4[2148] = 32'b11111111111111111000010010000001;
assign LUT_4[2149] = 32'b11111111111111110001011101111001;
assign LUT_4[2150] = 32'b11111111111111110111101100100101;
assign LUT_4[2151] = 32'b11111111111111110000111000011101;
assign LUT_4[2152] = 32'b11111111111111110100011101111010;
assign LUT_4[2153] = 32'b11111111111111101101101001110010;
assign LUT_4[2154] = 32'b11111111111111110011111000011110;
assign LUT_4[2155] = 32'b11111111111111101101000100010110;
assign LUT_4[2156] = 32'b11111111111111110001011110010110;
assign LUT_4[2157] = 32'b11111111111111101010101010001110;
assign LUT_4[2158] = 32'b11111111111111110000111000111010;
assign LUT_4[2159] = 32'b11111111111111101010000100110010;
assign LUT_4[2160] = 32'b11111111111111111001000011010011;
assign LUT_4[2161] = 32'b11111111111111110010001111001011;
assign LUT_4[2162] = 32'b11111111111111111000011101110111;
assign LUT_4[2163] = 32'b11111111111111110001101001101111;
assign LUT_4[2164] = 32'b11111111111111110110000011101111;
assign LUT_4[2165] = 32'b11111111111111101111001111100111;
assign LUT_4[2166] = 32'b11111111111111110101011110010011;
assign LUT_4[2167] = 32'b11111111111111101110101010001011;
assign LUT_4[2168] = 32'b11111111111111110010001111101000;
assign LUT_4[2169] = 32'b11111111111111101011011011100000;
assign LUT_4[2170] = 32'b11111111111111110001101010001100;
assign LUT_4[2171] = 32'b11111111111111101010110110000100;
assign LUT_4[2172] = 32'b11111111111111101111010000000100;
assign LUT_4[2173] = 32'b11111111111111101000011011111100;
assign LUT_4[2174] = 32'b11111111111111101110101010101000;
assign LUT_4[2175] = 32'b11111111111111100111110110100000;
assign LUT_4[2176] = 32'b11111111111111111110000101010010;
assign LUT_4[2177] = 32'b11111111111111110111010001001010;
assign LUT_4[2178] = 32'b11111111111111111101011111110110;
assign LUT_4[2179] = 32'b11111111111111110110101011101110;
assign LUT_4[2180] = 32'b11111111111111111011000101101110;
assign LUT_4[2181] = 32'b11111111111111110100010001100110;
assign LUT_4[2182] = 32'b11111111111111111010100000010010;
assign LUT_4[2183] = 32'b11111111111111110011101100001010;
assign LUT_4[2184] = 32'b11111111111111110111010001100111;
assign LUT_4[2185] = 32'b11111111111111110000011101011111;
assign LUT_4[2186] = 32'b11111111111111110110101100001011;
assign LUT_4[2187] = 32'b11111111111111101111111000000011;
assign LUT_4[2188] = 32'b11111111111111110100010010000011;
assign LUT_4[2189] = 32'b11111111111111101101011101111011;
assign LUT_4[2190] = 32'b11111111111111110011101100100111;
assign LUT_4[2191] = 32'b11111111111111101100111000011111;
assign LUT_4[2192] = 32'b11111111111111111011110111000000;
assign LUT_4[2193] = 32'b11111111111111110101000010111000;
assign LUT_4[2194] = 32'b11111111111111111011010001100100;
assign LUT_4[2195] = 32'b11111111111111110100011101011100;
assign LUT_4[2196] = 32'b11111111111111111000110111011100;
assign LUT_4[2197] = 32'b11111111111111110010000011010100;
assign LUT_4[2198] = 32'b11111111111111111000010010000000;
assign LUT_4[2199] = 32'b11111111111111110001011101111000;
assign LUT_4[2200] = 32'b11111111111111110101000011010101;
assign LUT_4[2201] = 32'b11111111111111101110001111001101;
assign LUT_4[2202] = 32'b11111111111111110100011101111001;
assign LUT_4[2203] = 32'b11111111111111101101101001110001;
assign LUT_4[2204] = 32'b11111111111111110010000011110001;
assign LUT_4[2205] = 32'b11111111111111101011001111101001;
assign LUT_4[2206] = 32'b11111111111111110001011110010101;
assign LUT_4[2207] = 32'b11111111111111101010101010001101;
assign LUT_4[2208] = 32'b11111111111111111100100000011001;
assign LUT_4[2209] = 32'b11111111111111110101101100010001;
assign LUT_4[2210] = 32'b11111111111111111011111010111101;
assign LUT_4[2211] = 32'b11111111111111110101000110110101;
assign LUT_4[2212] = 32'b11111111111111111001100000110101;
assign LUT_4[2213] = 32'b11111111111111110010101100101101;
assign LUT_4[2214] = 32'b11111111111111111000111011011001;
assign LUT_4[2215] = 32'b11111111111111110010000111010001;
assign LUT_4[2216] = 32'b11111111111111110101101100101110;
assign LUT_4[2217] = 32'b11111111111111101110111000100110;
assign LUT_4[2218] = 32'b11111111111111110101000111010010;
assign LUT_4[2219] = 32'b11111111111111101110010011001010;
assign LUT_4[2220] = 32'b11111111111111110010101101001010;
assign LUT_4[2221] = 32'b11111111111111101011111001000010;
assign LUT_4[2222] = 32'b11111111111111110010000111101110;
assign LUT_4[2223] = 32'b11111111111111101011010011100110;
assign LUT_4[2224] = 32'b11111111111111111010010010000111;
assign LUT_4[2225] = 32'b11111111111111110011011101111111;
assign LUT_4[2226] = 32'b11111111111111111001101100101011;
assign LUT_4[2227] = 32'b11111111111111110010111000100011;
assign LUT_4[2228] = 32'b11111111111111110111010010100011;
assign LUT_4[2229] = 32'b11111111111111110000011110011011;
assign LUT_4[2230] = 32'b11111111111111110110101101000111;
assign LUT_4[2231] = 32'b11111111111111101111111000111111;
assign LUT_4[2232] = 32'b11111111111111110011011110011100;
assign LUT_4[2233] = 32'b11111111111111101100101010010100;
assign LUT_4[2234] = 32'b11111111111111110010111001000000;
assign LUT_4[2235] = 32'b11111111111111101100000100111000;
assign LUT_4[2236] = 32'b11111111111111110000011110111000;
assign LUT_4[2237] = 32'b11111111111111101001101010110000;
assign LUT_4[2238] = 32'b11111111111111101111111001011100;
assign LUT_4[2239] = 32'b11111111111111101001000101010100;
assign LUT_4[2240] = 32'b11111111111111111111011100100110;
assign LUT_4[2241] = 32'b11111111111111111000101000011110;
assign LUT_4[2242] = 32'b11111111111111111110110111001010;
assign LUT_4[2243] = 32'b11111111111111111000000011000010;
assign LUT_4[2244] = 32'b11111111111111111100011101000010;
assign LUT_4[2245] = 32'b11111111111111110101101000111010;
assign LUT_4[2246] = 32'b11111111111111111011110111100110;
assign LUT_4[2247] = 32'b11111111111111110101000011011110;
assign LUT_4[2248] = 32'b11111111111111111000101000111011;
assign LUT_4[2249] = 32'b11111111111111110001110100110011;
assign LUT_4[2250] = 32'b11111111111111111000000011011111;
assign LUT_4[2251] = 32'b11111111111111110001001111010111;
assign LUT_4[2252] = 32'b11111111111111110101101001010111;
assign LUT_4[2253] = 32'b11111111111111101110110101001111;
assign LUT_4[2254] = 32'b11111111111111110101000011111011;
assign LUT_4[2255] = 32'b11111111111111101110001111110011;
assign LUT_4[2256] = 32'b11111111111111111101001110010100;
assign LUT_4[2257] = 32'b11111111111111110110011010001100;
assign LUT_4[2258] = 32'b11111111111111111100101000111000;
assign LUT_4[2259] = 32'b11111111111111110101110100110000;
assign LUT_4[2260] = 32'b11111111111111111010001110110000;
assign LUT_4[2261] = 32'b11111111111111110011011010101000;
assign LUT_4[2262] = 32'b11111111111111111001101001010100;
assign LUT_4[2263] = 32'b11111111111111110010110101001100;
assign LUT_4[2264] = 32'b11111111111111110110011010101001;
assign LUT_4[2265] = 32'b11111111111111101111100110100001;
assign LUT_4[2266] = 32'b11111111111111110101110101001101;
assign LUT_4[2267] = 32'b11111111111111101111000001000101;
assign LUT_4[2268] = 32'b11111111111111110011011011000101;
assign LUT_4[2269] = 32'b11111111111111101100100110111101;
assign LUT_4[2270] = 32'b11111111111111110010110101101001;
assign LUT_4[2271] = 32'b11111111111111101100000001100001;
assign LUT_4[2272] = 32'b11111111111111111101110111101101;
assign LUT_4[2273] = 32'b11111111111111110111000011100101;
assign LUT_4[2274] = 32'b11111111111111111101010010010001;
assign LUT_4[2275] = 32'b11111111111111110110011110001001;
assign LUT_4[2276] = 32'b11111111111111111010111000001001;
assign LUT_4[2277] = 32'b11111111111111110100000100000001;
assign LUT_4[2278] = 32'b11111111111111111010010010101101;
assign LUT_4[2279] = 32'b11111111111111110011011110100101;
assign LUT_4[2280] = 32'b11111111111111110111000100000010;
assign LUT_4[2281] = 32'b11111111111111110000001111111010;
assign LUT_4[2282] = 32'b11111111111111110110011110100110;
assign LUT_4[2283] = 32'b11111111111111101111101010011110;
assign LUT_4[2284] = 32'b11111111111111110100000100011110;
assign LUT_4[2285] = 32'b11111111111111101101010000010110;
assign LUT_4[2286] = 32'b11111111111111110011011111000010;
assign LUT_4[2287] = 32'b11111111111111101100101010111010;
assign LUT_4[2288] = 32'b11111111111111111011101001011011;
assign LUT_4[2289] = 32'b11111111111111110100110101010011;
assign LUT_4[2290] = 32'b11111111111111111011000011111111;
assign LUT_4[2291] = 32'b11111111111111110100001111110111;
assign LUT_4[2292] = 32'b11111111111111111000101001110111;
assign LUT_4[2293] = 32'b11111111111111110001110101101111;
assign LUT_4[2294] = 32'b11111111111111111000000100011011;
assign LUT_4[2295] = 32'b11111111111111110001010000010011;
assign LUT_4[2296] = 32'b11111111111111110100110101110000;
assign LUT_4[2297] = 32'b11111111111111101110000001101000;
assign LUT_4[2298] = 32'b11111111111111110100010000010100;
assign LUT_4[2299] = 32'b11111111111111101101011100001100;
assign LUT_4[2300] = 32'b11111111111111110001110110001100;
assign LUT_4[2301] = 32'b11111111111111101011000010000100;
assign LUT_4[2302] = 32'b11111111111111110001010000110000;
assign LUT_4[2303] = 32'b11111111111111101010011100101000;
assign LUT_4[2304] = 32'b00000000000000000000011010101101;
assign LUT_4[2305] = 32'b11111111111111111001100110100101;
assign LUT_4[2306] = 32'b11111111111111111111110101010001;
assign LUT_4[2307] = 32'b11111111111111111001000001001001;
assign LUT_4[2308] = 32'b11111111111111111101011011001001;
assign LUT_4[2309] = 32'b11111111111111110110100111000001;
assign LUT_4[2310] = 32'b11111111111111111100110101101101;
assign LUT_4[2311] = 32'b11111111111111110110000001100101;
assign LUT_4[2312] = 32'b11111111111111111001100111000010;
assign LUT_4[2313] = 32'b11111111111111110010110010111010;
assign LUT_4[2314] = 32'b11111111111111111001000001100110;
assign LUT_4[2315] = 32'b11111111111111110010001101011110;
assign LUT_4[2316] = 32'b11111111111111110110100111011110;
assign LUT_4[2317] = 32'b11111111111111101111110011010110;
assign LUT_4[2318] = 32'b11111111111111110110000010000010;
assign LUT_4[2319] = 32'b11111111111111101111001101111010;
assign LUT_4[2320] = 32'b11111111111111111110001100011011;
assign LUT_4[2321] = 32'b11111111111111110111011000010011;
assign LUT_4[2322] = 32'b11111111111111111101100110111111;
assign LUT_4[2323] = 32'b11111111111111110110110010110111;
assign LUT_4[2324] = 32'b11111111111111111011001100110111;
assign LUT_4[2325] = 32'b11111111111111110100011000101111;
assign LUT_4[2326] = 32'b11111111111111111010100111011011;
assign LUT_4[2327] = 32'b11111111111111110011110011010011;
assign LUT_4[2328] = 32'b11111111111111110111011000110000;
assign LUT_4[2329] = 32'b11111111111111110000100100101000;
assign LUT_4[2330] = 32'b11111111111111110110110011010100;
assign LUT_4[2331] = 32'b11111111111111101111111111001100;
assign LUT_4[2332] = 32'b11111111111111110100011001001100;
assign LUT_4[2333] = 32'b11111111111111101101100101000100;
assign LUT_4[2334] = 32'b11111111111111110011110011110000;
assign LUT_4[2335] = 32'b11111111111111101100111111101000;
assign LUT_4[2336] = 32'b11111111111111111110110101110100;
assign LUT_4[2337] = 32'b11111111111111111000000001101100;
assign LUT_4[2338] = 32'b11111111111111111110010000011000;
assign LUT_4[2339] = 32'b11111111111111110111011100010000;
assign LUT_4[2340] = 32'b11111111111111111011110110010000;
assign LUT_4[2341] = 32'b11111111111111110101000010001000;
assign LUT_4[2342] = 32'b11111111111111111011010000110100;
assign LUT_4[2343] = 32'b11111111111111110100011100101100;
assign LUT_4[2344] = 32'b11111111111111111000000010001001;
assign LUT_4[2345] = 32'b11111111111111110001001110000001;
assign LUT_4[2346] = 32'b11111111111111110111011100101101;
assign LUT_4[2347] = 32'b11111111111111110000101000100101;
assign LUT_4[2348] = 32'b11111111111111110101000010100101;
assign LUT_4[2349] = 32'b11111111111111101110001110011101;
assign LUT_4[2350] = 32'b11111111111111110100011101001001;
assign LUT_4[2351] = 32'b11111111111111101101101001000001;
assign LUT_4[2352] = 32'b11111111111111111100100111100010;
assign LUT_4[2353] = 32'b11111111111111110101110011011010;
assign LUT_4[2354] = 32'b11111111111111111100000010000110;
assign LUT_4[2355] = 32'b11111111111111110101001101111110;
assign LUT_4[2356] = 32'b11111111111111111001100111111110;
assign LUT_4[2357] = 32'b11111111111111110010110011110110;
assign LUT_4[2358] = 32'b11111111111111111001000010100010;
assign LUT_4[2359] = 32'b11111111111111110010001110011010;
assign LUT_4[2360] = 32'b11111111111111110101110011110111;
assign LUT_4[2361] = 32'b11111111111111101110111111101111;
assign LUT_4[2362] = 32'b11111111111111110101001110011011;
assign LUT_4[2363] = 32'b11111111111111101110011010010011;
assign LUT_4[2364] = 32'b11111111111111110010110100010011;
assign LUT_4[2365] = 32'b11111111111111101100000000001011;
assign LUT_4[2366] = 32'b11111111111111110010001110110111;
assign LUT_4[2367] = 32'b11111111111111101011011010101111;
assign LUT_4[2368] = 32'b00000000000000000001110010000001;
assign LUT_4[2369] = 32'b11111111111111111010111101111001;
assign LUT_4[2370] = 32'b00000000000000000001001100100101;
assign LUT_4[2371] = 32'b11111111111111111010011000011101;
assign LUT_4[2372] = 32'b11111111111111111110110010011101;
assign LUT_4[2373] = 32'b11111111111111110111111110010101;
assign LUT_4[2374] = 32'b11111111111111111110001101000001;
assign LUT_4[2375] = 32'b11111111111111110111011000111001;
assign LUT_4[2376] = 32'b11111111111111111010111110010110;
assign LUT_4[2377] = 32'b11111111111111110100001010001110;
assign LUT_4[2378] = 32'b11111111111111111010011000111010;
assign LUT_4[2379] = 32'b11111111111111110011100100110010;
assign LUT_4[2380] = 32'b11111111111111110111111110110010;
assign LUT_4[2381] = 32'b11111111111111110001001010101010;
assign LUT_4[2382] = 32'b11111111111111110111011001010110;
assign LUT_4[2383] = 32'b11111111111111110000100101001110;
assign LUT_4[2384] = 32'b11111111111111111111100011101111;
assign LUT_4[2385] = 32'b11111111111111111000101111100111;
assign LUT_4[2386] = 32'b11111111111111111110111110010011;
assign LUT_4[2387] = 32'b11111111111111111000001010001011;
assign LUT_4[2388] = 32'b11111111111111111100100100001011;
assign LUT_4[2389] = 32'b11111111111111110101110000000011;
assign LUT_4[2390] = 32'b11111111111111111011111110101111;
assign LUT_4[2391] = 32'b11111111111111110101001010100111;
assign LUT_4[2392] = 32'b11111111111111111000110000000100;
assign LUT_4[2393] = 32'b11111111111111110001111011111100;
assign LUT_4[2394] = 32'b11111111111111111000001010101000;
assign LUT_4[2395] = 32'b11111111111111110001010110100000;
assign LUT_4[2396] = 32'b11111111111111110101110000100000;
assign LUT_4[2397] = 32'b11111111111111101110111100011000;
assign LUT_4[2398] = 32'b11111111111111110101001011000100;
assign LUT_4[2399] = 32'b11111111111111101110010110111100;
assign LUT_4[2400] = 32'b00000000000000000000001101001000;
assign LUT_4[2401] = 32'b11111111111111111001011001000000;
assign LUT_4[2402] = 32'b11111111111111111111100111101100;
assign LUT_4[2403] = 32'b11111111111111111000110011100100;
assign LUT_4[2404] = 32'b11111111111111111101001101100100;
assign LUT_4[2405] = 32'b11111111111111110110011001011100;
assign LUT_4[2406] = 32'b11111111111111111100101000001000;
assign LUT_4[2407] = 32'b11111111111111110101110100000000;
assign LUT_4[2408] = 32'b11111111111111111001011001011101;
assign LUT_4[2409] = 32'b11111111111111110010100101010101;
assign LUT_4[2410] = 32'b11111111111111111000110100000001;
assign LUT_4[2411] = 32'b11111111111111110001111111111001;
assign LUT_4[2412] = 32'b11111111111111110110011001111001;
assign LUT_4[2413] = 32'b11111111111111101111100101110001;
assign LUT_4[2414] = 32'b11111111111111110101110100011101;
assign LUT_4[2415] = 32'b11111111111111101111000000010101;
assign LUT_4[2416] = 32'b11111111111111111101111110110110;
assign LUT_4[2417] = 32'b11111111111111110111001010101110;
assign LUT_4[2418] = 32'b11111111111111111101011001011010;
assign LUT_4[2419] = 32'b11111111111111110110100101010010;
assign LUT_4[2420] = 32'b11111111111111111010111111010010;
assign LUT_4[2421] = 32'b11111111111111110100001011001010;
assign LUT_4[2422] = 32'b11111111111111111010011001110110;
assign LUT_4[2423] = 32'b11111111111111110011100101101110;
assign LUT_4[2424] = 32'b11111111111111110111001011001011;
assign LUT_4[2425] = 32'b11111111111111110000010111000011;
assign LUT_4[2426] = 32'b11111111111111110110100101101111;
assign LUT_4[2427] = 32'b11111111111111101111110001100111;
assign LUT_4[2428] = 32'b11111111111111110100001011100111;
assign LUT_4[2429] = 32'b11111111111111101101010111011111;
assign LUT_4[2430] = 32'b11111111111111110011100110001011;
assign LUT_4[2431] = 32'b11111111111111101100110010000011;
assign LUT_4[2432] = 32'b00000000000000000011000000110101;
assign LUT_4[2433] = 32'b11111111111111111100001100101101;
assign LUT_4[2434] = 32'b00000000000000000010011011011001;
assign LUT_4[2435] = 32'b11111111111111111011100111010001;
assign LUT_4[2436] = 32'b00000000000000000000000001010001;
assign LUT_4[2437] = 32'b11111111111111111001001101001001;
assign LUT_4[2438] = 32'b11111111111111111111011011110101;
assign LUT_4[2439] = 32'b11111111111111111000100111101101;
assign LUT_4[2440] = 32'b11111111111111111100001101001010;
assign LUT_4[2441] = 32'b11111111111111110101011001000010;
assign LUT_4[2442] = 32'b11111111111111111011100111101110;
assign LUT_4[2443] = 32'b11111111111111110100110011100110;
assign LUT_4[2444] = 32'b11111111111111111001001101100110;
assign LUT_4[2445] = 32'b11111111111111110010011001011110;
assign LUT_4[2446] = 32'b11111111111111111000101000001010;
assign LUT_4[2447] = 32'b11111111111111110001110100000010;
assign LUT_4[2448] = 32'b00000000000000000000110010100011;
assign LUT_4[2449] = 32'b11111111111111111001111110011011;
assign LUT_4[2450] = 32'b00000000000000000000001101000111;
assign LUT_4[2451] = 32'b11111111111111111001011000111111;
assign LUT_4[2452] = 32'b11111111111111111101110010111111;
assign LUT_4[2453] = 32'b11111111111111110110111110110111;
assign LUT_4[2454] = 32'b11111111111111111101001101100011;
assign LUT_4[2455] = 32'b11111111111111110110011001011011;
assign LUT_4[2456] = 32'b11111111111111111001111110111000;
assign LUT_4[2457] = 32'b11111111111111110011001010110000;
assign LUT_4[2458] = 32'b11111111111111111001011001011100;
assign LUT_4[2459] = 32'b11111111111111110010100101010100;
assign LUT_4[2460] = 32'b11111111111111110110111111010100;
assign LUT_4[2461] = 32'b11111111111111110000001011001100;
assign LUT_4[2462] = 32'b11111111111111110110011001111000;
assign LUT_4[2463] = 32'b11111111111111101111100101110000;
assign LUT_4[2464] = 32'b00000000000000000001011011111100;
assign LUT_4[2465] = 32'b11111111111111111010100111110100;
assign LUT_4[2466] = 32'b00000000000000000000110110100000;
assign LUT_4[2467] = 32'b11111111111111111010000010011000;
assign LUT_4[2468] = 32'b11111111111111111110011100011000;
assign LUT_4[2469] = 32'b11111111111111110111101000010000;
assign LUT_4[2470] = 32'b11111111111111111101110110111100;
assign LUT_4[2471] = 32'b11111111111111110111000010110100;
assign LUT_4[2472] = 32'b11111111111111111010101000010001;
assign LUT_4[2473] = 32'b11111111111111110011110100001001;
assign LUT_4[2474] = 32'b11111111111111111010000010110101;
assign LUT_4[2475] = 32'b11111111111111110011001110101101;
assign LUT_4[2476] = 32'b11111111111111110111101000101101;
assign LUT_4[2477] = 32'b11111111111111110000110100100101;
assign LUT_4[2478] = 32'b11111111111111110111000011010001;
assign LUT_4[2479] = 32'b11111111111111110000001111001001;
assign LUT_4[2480] = 32'b11111111111111111111001101101010;
assign LUT_4[2481] = 32'b11111111111111111000011001100010;
assign LUT_4[2482] = 32'b11111111111111111110101000001110;
assign LUT_4[2483] = 32'b11111111111111110111110100000110;
assign LUT_4[2484] = 32'b11111111111111111100001110000110;
assign LUT_4[2485] = 32'b11111111111111110101011001111110;
assign LUT_4[2486] = 32'b11111111111111111011101000101010;
assign LUT_4[2487] = 32'b11111111111111110100110100100010;
assign LUT_4[2488] = 32'b11111111111111111000011001111111;
assign LUT_4[2489] = 32'b11111111111111110001100101110111;
assign LUT_4[2490] = 32'b11111111111111110111110100100011;
assign LUT_4[2491] = 32'b11111111111111110001000000011011;
assign LUT_4[2492] = 32'b11111111111111110101011010011011;
assign LUT_4[2493] = 32'b11111111111111101110100110010011;
assign LUT_4[2494] = 32'b11111111111111110100110100111111;
assign LUT_4[2495] = 32'b11111111111111101110000000110111;
assign LUT_4[2496] = 32'b00000000000000000100011000001001;
assign LUT_4[2497] = 32'b11111111111111111101100100000001;
assign LUT_4[2498] = 32'b00000000000000000011110010101101;
assign LUT_4[2499] = 32'b11111111111111111100111110100101;
assign LUT_4[2500] = 32'b00000000000000000001011000100101;
assign LUT_4[2501] = 32'b11111111111111111010100100011101;
assign LUT_4[2502] = 32'b00000000000000000000110011001001;
assign LUT_4[2503] = 32'b11111111111111111001111111000001;
assign LUT_4[2504] = 32'b11111111111111111101100100011110;
assign LUT_4[2505] = 32'b11111111111111110110110000010110;
assign LUT_4[2506] = 32'b11111111111111111100111111000010;
assign LUT_4[2507] = 32'b11111111111111110110001010111010;
assign LUT_4[2508] = 32'b11111111111111111010100100111010;
assign LUT_4[2509] = 32'b11111111111111110011110000110010;
assign LUT_4[2510] = 32'b11111111111111111001111111011110;
assign LUT_4[2511] = 32'b11111111111111110011001011010110;
assign LUT_4[2512] = 32'b00000000000000000010001001110111;
assign LUT_4[2513] = 32'b11111111111111111011010101101111;
assign LUT_4[2514] = 32'b00000000000000000001100100011011;
assign LUT_4[2515] = 32'b11111111111111111010110000010011;
assign LUT_4[2516] = 32'b11111111111111111111001010010011;
assign LUT_4[2517] = 32'b11111111111111111000010110001011;
assign LUT_4[2518] = 32'b11111111111111111110100100110111;
assign LUT_4[2519] = 32'b11111111111111110111110000101111;
assign LUT_4[2520] = 32'b11111111111111111011010110001100;
assign LUT_4[2521] = 32'b11111111111111110100100010000100;
assign LUT_4[2522] = 32'b11111111111111111010110000110000;
assign LUT_4[2523] = 32'b11111111111111110011111100101000;
assign LUT_4[2524] = 32'b11111111111111111000010110101000;
assign LUT_4[2525] = 32'b11111111111111110001100010100000;
assign LUT_4[2526] = 32'b11111111111111110111110001001100;
assign LUT_4[2527] = 32'b11111111111111110000111101000100;
assign LUT_4[2528] = 32'b00000000000000000010110011010000;
assign LUT_4[2529] = 32'b11111111111111111011111111001000;
assign LUT_4[2530] = 32'b00000000000000000010001101110100;
assign LUT_4[2531] = 32'b11111111111111111011011001101100;
assign LUT_4[2532] = 32'b11111111111111111111110011101100;
assign LUT_4[2533] = 32'b11111111111111111000111111100100;
assign LUT_4[2534] = 32'b11111111111111111111001110010000;
assign LUT_4[2535] = 32'b11111111111111111000011010001000;
assign LUT_4[2536] = 32'b11111111111111111011111111100101;
assign LUT_4[2537] = 32'b11111111111111110101001011011101;
assign LUT_4[2538] = 32'b11111111111111111011011010001001;
assign LUT_4[2539] = 32'b11111111111111110100100110000001;
assign LUT_4[2540] = 32'b11111111111111111001000000000001;
assign LUT_4[2541] = 32'b11111111111111110010001011111001;
assign LUT_4[2542] = 32'b11111111111111111000011010100101;
assign LUT_4[2543] = 32'b11111111111111110001100110011101;
assign LUT_4[2544] = 32'b00000000000000000000100100111110;
assign LUT_4[2545] = 32'b11111111111111111001110000110110;
assign LUT_4[2546] = 32'b11111111111111111111111111100010;
assign LUT_4[2547] = 32'b11111111111111111001001011011010;
assign LUT_4[2548] = 32'b11111111111111111101100101011010;
assign LUT_4[2549] = 32'b11111111111111110110110001010010;
assign LUT_4[2550] = 32'b11111111111111111100111111111110;
assign LUT_4[2551] = 32'b11111111111111110110001011110110;
assign LUT_4[2552] = 32'b11111111111111111001110001010011;
assign LUT_4[2553] = 32'b11111111111111110010111101001011;
assign LUT_4[2554] = 32'b11111111111111111001001011110111;
assign LUT_4[2555] = 32'b11111111111111110010010111101111;
assign LUT_4[2556] = 32'b11111111111111110110110001101111;
assign LUT_4[2557] = 32'b11111111111111101111111101100111;
assign LUT_4[2558] = 32'b11111111111111110110001100010011;
assign LUT_4[2559] = 32'b11111111111111101111011000001011;
assign LUT_4[2560] = 32'b11111111111111111010100011010010;
assign LUT_4[2561] = 32'b11111111111111110011101111001010;
assign LUT_4[2562] = 32'b11111111111111111001111101110110;
assign LUT_4[2563] = 32'b11111111111111110011001001101110;
assign LUT_4[2564] = 32'b11111111111111110111100011101110;
assign LUT_4[2565] = 32'b11111111111111110000101111100110;
assign LUT_4[2566] = 32'b11111111111111110110111110010010;
assign LUT_4[2567] = 32'b11111111111111110000001010001010;
assign LUT_4[2568] = 32'b11111111111111110011101111100111;
assign LUT_4[2569] = 32'b11111111111111101100111011011111;
assign LUT_4[2570] = 32'b11111111111111110011001010001011;
assign LUT_4[2571] = 32'b11111111111111101100010110000011;
assign LUT_4[2572] = 32'b11111111111111110000110000000011;
assign LUT_4[2573] = 32'b11111111111111101001111011111011;
assign LUT_4[2574] = 32'b11111111111111110000001010100111;
assign LUT_4[2575] = 32'b11111111111111101001010110011111;
assign LUT_4[2576] = 32'b11111111111111111000010101000000;
assign LUT_4[2577] = 32'b11111111111111110001100000111000;
assign LUT_4[2578] = 32'b11111111111111110111101111100100;
assign LUT_4[2579] = 32'b11111111111111110000111011011100;
assign LUT_4[2580] = 32'b11111111111111110101010101011100;
assign LUT_4[2581] = 32'b11111111111111101110100001010100;
assign LUT_4[2582] = 32'b11111111111111110100110000000000;
assign LUT_4[2583] = 32'b11111111111111101101111011111000;
assign LUT_4[2584] = 32'b11111111111111110001100001010101;
assign LUT_4[2585] = 32'b11111111111111101010101101001101;
assign LUT_4[2586] = 32'b11111111111111110000111011111001;
assign LUT_4[2587] = 32'b11111111111111101010000111110001;
assign LUT_4[2588] = 32'b11111111111111101110100001110001;
assign LUT_4[2589] = 32'b11111111111111100111101101101001;
assign LUT_4[2590] = 32'b11111111111111101101111100010101;
assign LUT_4[2591] = 32'b11111111111111100111001000001101;
assign LUT_4[2592] = 32'b11111111111111111000111110011001;
assign LUT_4[2593] = 32'b11111111111111110010001010010001;
assign LUT_4[2594] = 32'b11111111111111111000011000111101;
assign LUT_4[2595] = 32'b11111111111111110001100100110101;
assign LUT_4[2596] = 32'b11111111111111110101111110110101;
assign LUT_4[2597] = 32'b11111111111111101111001010101101;
assign LUT_4[2598] = 32'b11111111111111110101011001011001;
assign LUT_4[2599] = 32'b11111111111111101110100101010001;
assign LUT_4[2600] = 32'b11111111111111110010001010101110;
assign LUT_4[2601] = 32'b11111111111111101011010110100110;
assign LUT_4[2602] = 32'b11111111111111110001100101010010;
assign LUT_4[2603] = 32'b11111111111111101010110001001010;
assign LUT_4[2604] = 32'b11111111111111101111001011001010;
assign LUT_4[2605] = 32'b11111111111111101000010111000010;
assign LUT_4[2606] = 32'b11111111111111101110100101101110;
assign LUT_4[2607] = 32'b11111111111111100111110001100110;
assign LUT_4[2608] = 32'b11111111111111110110110000000111;
assign LUT_4[2609] = 32'b11111111111111101111111011111111;
assign LUT_4[2610] = 32'b11111111111111110110001010101011;
assign LUT_4[2611] = 32'b11111111111111101111010110100011;
assign LUT_4[2612] = 32'b11111111111111110011110000100011;
assign LUT_4[2613] = 32'b11111111111111101100111100011011;
assign LUT_4[2614] = 32'b11111111111111110011001011000111;
assign LUT_4[2615] = 32'b11111111111111101100010110111111;
assign LUT_4[2616] = 32'b11111111111111101111111100011100;
assign LUT_4[2617] = 32'b11111111111111101001001000010100;
assign LUT_4[2618] = 32'b11111111111111101111010111000000;
assign LUT_4[2619] = 32'b11111111111111101000100010111000;
assign LUT_4[2620] = 32'b11111111111111101100111100111000;
assign LUT_4[2621] = 32'b11111111111111100110001000110000;
assign LUT_4[2622] = 32'b11111111111111101100010111011100;
assign LUT_4[2623] = 32'b11111111111111100101100011010100;
assign LUT_4[2624] = 32'b11111111111111111011111010100110;
assign LUT_4[2625] = 32'b11111111111111110101000110011110;
assign LUT_4[2626] = 32'b11111111111111111011010101001010;
assign LUT_4[2627] = 32'b11111111111111110100100001000010;
assign LUT_4[2628] = 32'b11111111111111111000111011000010;
assign LUT_4[2629] = 32'b11111111111111110010000110111010;
assign LUT_4[2630] = 32'b11111111111111111000010101100110;
assign LUT_4[2631] = 32'b11111111111111110001100001011110;
assign LUT_4[2632] = 32'b11111111111111110101000110111011;
assign LUT_4[2633] = 32'b11111111111111101110010010110011;
assign LUT_4[2634] = 32'b11111111111111110100100001011111;
assign LUT_4[2635] = 32'b11111111111111101101101101010111;
assign LUT_4[2636] = 32'b11111111111111110010000111010111;
assign LUT_4[2637] = 32'b11111111111111101011010011001111;
assign LUT_4[2638] = 32'b11111111111111110001100001111011;
assign LUT_4[2639] = 32'b11111111111111101010101101110011;
assign LUT_4[2640] = 32'b11111111111111111001101100010100;
assign LUT_4[2641] = 32'b11111111111111110010111000001100;
assign LUT_4[2642] = 32'b11111111111111111001000110111000;
assign LUT_4[2643] = 32'b11111111111111110010010010110000;
assign LUT_4[2644] = 32'b11111111111111110110101100110000;
assign LUT_4[2645] = 32'b11111111111111101111111000101000;
assign LUT_4[2646] = 32'b11111111111111110110000111010100;
assign LUT_4[2647] = 32'b11111111111111101111010011001100;
assign LUT_4[2648] = 32'b11111111111111110010111000101001;
assign LUT_4[2649] = 32'b11111111111111101100000100100001;
assign LUT_4[2650] = 32'b11111111111111110010010011001101;
assign LUT_4[2651] = 32'b11111111111111101011011111000101;
assign LUT_4[2652] = 32'b11111111111111101111111001000101;
assign LUT_4[2653] = 32'b11111111111111101001000100111101;
assign LUT_4[2654] = 32'b11111111111111101111010011101001;
assign LUT_4[2655] = 32'b11111111111111101000011111100001;
assign LUT_4[2656] = 32'b11111111111111111010010101101101;
assign LUT_4[2657] = 32'b11111111111111110011100001100101;
assign LUT_4[2658] = 32'b11111111111111111001110000010001;
assign LUT_4[2659] = 32'b11111111111111110010111100001001;
assign LUT_4[2660] = 32'b11111111111111110111010110001001;
assign LUT_4[2661] = 32'b11111111111111110000100010000001;
assign LUT_4[2662] = 32'b11111111111111110110110000101101;
assign LUT_4[2663] = 32'b11111111111111101111111100100101;
assign LUT_4[2664] = 32'b11111111111111110011100010000010;
assign LUT_4[2665] = 32'b11111111111111101100101101111010;
assign LUT_4[2666] = 32'b11111111111111110010111100100110;
assign LUT_4[2667] = 32'b11111111111111101100001000011110;
assign LUT_4[2668] = 32'b11111111111111110000100010011110;
assign LUT_4[2669] = 32'b11111111111111101001101110010110;
assign LUT_4[2670] = 32'b11111111111111101111111101000010;
assign LUT_4[2671] = 32'b11111111111111101001001000111010;
assign LUT_4[2672] = 32'b11111111111111111000000111011011;
assign LUT_4[2673] = 32'b11111111111111110001010011010011;
assign LUT_4[2674] = 32'b11111111111111110111100001111111;
assign LUT_4[2675] = 32'b11111111111111110000101101110111;
assign LUT_4[2676] = 32'b11111111111111110101000111110111;
assign LUT_4[2677] = 32'b11111111111111101110010011101111;
assign LUT_4[2678] = 32'b11111111111111110100100010011011;
assign LUT_4[2679] = 32'b11111111111111101101101110010011;
assign LUT_4[2680] = 32'b11111111111111110001010011110000;
assign LUT_4[2681] = 32'b11111111111111101010011111101000;
assign LUT_4[2682] = 32'b11111111111111110000101110010100;
assign LUT_4[2683] = 32'b11111111111111101001111010001100;
assign LUT_4[2684] = 32'b11111111111111101110010100001100;
assign LUT_4[2685] = 32'b11111111111111100111100000000100;
assign LUT_4[2686] = 32'b11111111111111101101101110110000;
assign LUT_4[2687] = 32'b11111111111111100110111010101000;
assign LUT_4[2688] = 32'b11111111111111111101001001011010;
assign LUT_4[2689] = 32'b11111111111111110110010101010010;
assign LUT_4[2690] = 32'b11111111111111111100100011111110;
assign LUT_4[2691] = 32'b11111111111111110101101111110110;
assign LUT_4[2692] = 32'b11111111111111111010001001110110;
assign LUT_4[2693] = 32'b11111111111111110011010101101110;
assign LUT_4[2694] = 32'b11111111111111111001100100011010;
assign LUT_4[2695] = 32'b11111111111111110010110000010010;
assign LUT_4[2696] = 32'b11111111111111110110010101101111;
assign LUT_4[2697] = 32'b11111111111111101111100001100111;
assign LUT_4[2698] = 32'b11111111111111110101110000010011;
assign LUT_4[2699] = 32'b11111111111111101110111100001011;
assign LUT_4[2700] = 32'b11111111111111110011010110001011;
assign LUT_4[2701] = 32'b11111111111111101100100010000011;
assign LUT_4[2702] = 32'b11111111111111110010110000101111;
assign LUT_4[2703] = 32'b11111111111111101011111100100111;
assign LUT_4[2704] = 32'b11111111111111111010111011001000;
assign LUT_4[2705] = 32'b11111111111111110100000111000000;
assign LUT_4[2706] = 32'b11111111111111111010010101101100;
assign LUT_4[2707] = 32'b11111111111111110011100001100100;
assign LUT_4[2708] = 32'b11111111111111110111111011100100;
assign LUT_4[2709] = 32'b11111111111111110001000111011100;
assign LUT_4[2710] = 32'b11111111111111110111010110001000;
assign LUT_4[2711] = 32'b11111111111111110000100010000000;
assign LUT_4[2712] = 32'b11111111111111110100000111011101;
assign LUT_4[2713] = 32'b11111111111111101101010011010101;
assign LUT_4[2714] = 32'b11111111111111110011100010000001;
assign LUT_4[2715] = 32'b11111111111111101100101101111001;
assign LUT_4[2716] = 32'b11111111111111110001000111111001;
assign LUT_4[2717] = 32'b11111111111111101010010011110001;
assign LUT_4[2718] = 32'b11111111111111110000100010011101;
assign LUT_4[2719] = 32'b11111111111111101001101110010101;
assign LUT_4[2720] = 32'b11111111111111111011100100100001;
assign LUT_4[2721] = 32'b11111111111111110100110000011001;
assign LUT_4[2722] = 32'b11111111111111111010111111000101;
assign LUT_4[2723] = 32'b11111111111111110100001010111101;
assign LUT_4[2724] = 32'b11111111111111111000100100111101;
assign LUT_4[2725] = 32'b11111111111111110001110000110101;
assign LUT_4[2726] = 32'b11111111111111110111111111100001;
assign LUT_4[2727] = 32'b11111111111111110001001011011001;
assign LUT_4[2728] = 32'b11111111111111110100110000110110;
assign LUT_4[2729] = 32'b11111111111111101101111100101110;
assign LUT_4[2730] = 32'b11111111111111110100001011011010;
assign LUT_4[2731] = 32'b11111111111111101101010111010010;
assign LUT_4[2732] = 32'b11111111111111110001110001010010;
assign LUT_4[2733] = 32'b11111111111111101010111101001010;
assign LUT_4[2734] = 32'b11111111111111110001001011110110;
assign LUT_4[2735] = 32'b11111111111111101010010111101110;
assign LUT_4[2736] = 32'b11111111111111111001010110001111;
assign LUT_4[2737] = 32'b11111111111111110010100010000111;
assign LUT_4[2738] = 32'b11111111111111111000110000110011;
assign LUT_4[2739] = 32'b11111111111111110001111100101011;
assign LUT_4[2740] = 32'b11111111111111110110010110101011;
assign LUT_4[2741] = 32'b11111111111111101111100010100011;
assign LUT_4[2742] = 32'b11111111111111110101110001001111;
assign LUT_4[2743] = 32'b11111111111111101110111101000111;
assign LUT_4[2744] = 32'b11111111111111110010100010100100;
assign LUT_4[2745] = 32'b11111111111111101011101110011100;
assign LUT_4[2746] = 32'b11111111111111110001111101001000;
assign LUT_4[2747] = 32'b11111111111111101011001001000000;
assign LUT_4[2748] = 32'b11111111111111101111100011000000;
assign LUT_4[2749] = 32'b11111111111111101000101110111000;
assign LUT_4[2750] = 32'b11111111111111101110111101100100;
assign LUT_4[2751] = 32'b11111111111111101000001001011100;
assign LUT_4[2752] = 32'b11111111111111111110100000101110;
assign LUT_4[2753] = 32'b11111111111111110111101100100110;
assign LUT_4[2754] = 32'b11111111111111111101111011010010;
assign LUT_4[2755] = 32'b11111111111111110111000111001010;
assign LUT_4[2756] = 32'b11111111111111111011100001001010;
assign LUT_4[2757] = 32'b11111111111111110100101101000010;
assign LUT_4[2758] = 32'b11111111111111111010111011101110;
assign LUT_4[2759] = 32'b11111111111111110100000111100110;
assign LUT_4[2760] = 32'b11111111111111110111101101000011;
assign LUT_4[2761] = 32'b11111111111111110000111000111011;
assign LUT_4[2762] = 32'b11111111111111110111000111100111;
assign LUT_4[2763] = 32'b11111111111111110000010011011111;
assign LUT_4[2764] = 32'b11111111111111110100101101011111;
assign LUT_4[2765] = 32'b11111111111111101101111001010111;
assign LUT_4[2766] = 32'b11111111111111110100001000000011;
assign LUT_4[2767] = 32'b11111111111111101101010011111011;
assign LUT_4[2768] = 32'b11111111111111111100010010011100;
assign LUT_4[2769] = 32'b11111111111111110101011110010100;
assign LUT_4[2770] = 32'b11111111111111111011101101000000;
assign LUT_4[2771] = 32'b11111111111111110100111000111000;
assign LUT_4[2772] = 32'b11111111111111111001010010111000;
assign LUT_4[2773] = 32'b11111111111111110010011110110000;
assign LUT_4[2774] = 32'b11111111111111111000101101011100;
assign LUT_4[2775] = 32'b11111111111111110001111001010100;
assign LUT_4[2776] = 32'b11111111111111110101011110110001;
assign LUT_4[2777] = 32'b11111111111111101110101010101001;
assign LUT_4[2778] = 32'b11111111111111110100111001010101;
assign LUT_4[2779] = 32'b11111111111111101110000101001101;
assign LUT_4[2780] = 32'b11111111111111110010011111001101;
assign LUT_4[2781] = 32'b11111111111111101011101011000101;
assign LUT_4[2782] = 32'b11111111111111110001111001110001;
assign LUT_4[2783] = 32'b11111111111111101011000101101001;
assign LUT_4[2784] = 32'b11111111111111111100111011110101;
assign LUT_4[2785] = 32'b11111111111111110110000111101101;
assign LUT_4[2786] = 32'b11111111111111111100010110011001;
assign LUT_4[2787] = 32'b11111111111111110101100010010001;
assign LUT_4[2788] = 32'b11111111111111111001111100010001;
assign LUT_4[2789] = 32'b11111111111111110011001000001001;
assign LUT_4[2790] = 32'b11111111111111111001010110110101;
assign LUT_4[2791] = 32'b11111111111111110010100010101101;
assign LUT_4[2792] = 32'b11111111111111110110001000001010;
assign LUT_4[2793] = 32'b11111111111111101111010100000010;
assign LUT_4[2794] = 32'b11111111111111110101100010101110;
assign LUT_4[2795] = 32'b11111111111111101110101110100110;
assign LUT_4[2796] = 32'b11111111111111110011001000100110;
assign LUT_4[2797] = 32'b11111111111111101100010100011110;
assign LUT_4[2798] = 32'b11111111111111110010100011001010;
assign LUT_4[2799] = 32'b11111111111111101011101111000010;
assign LUT_4[2800] = 32'b11111111111111111010101101100011;
assign LUT_4[2801] = 32'b11111111111111110011111001011011;
assign LUT_4[2802] = 32'b11111111111111111010001000000111;
assign LUT_4[2803] = 32'b11111111111111110011010011111111;
assign LUT_4[2804] = 32'b11111111111111110111101101111111;
assign LUT_4[2805] = 32'b11111111111111110000111001110111;
assign LUT_4[2806] = 32'b11111111111111110111001000100011;
assign LUT_4[2807] = 32'b11111111111111110000010100011011;
assign LUT_4[2808] = 32'b11111111111111110011111001111000;
assign LUT_4[2809] = 32'b11111111111111101101000101110000;
assign LUT_4[2810] = 32'b11111111111111110011010100011100;
assign LUT_4[2811] = 32'b11111111111111101100100000010100;
assign LUT_4[2812] = 32'b11111111111111110000111010010100;
assign LUT_4[2813] = 32'b11111111111111101010000110001100;
assign LUT_4[2814] = 32'b11111111111111110000010100111000;
assign LUT_4[2815] = 32'b11111111111111101001100000110000;
assign LUT_4[2816] = 32'b11111111111111111111011110110101;
assign LUT_4[2817] = 32'b11111111111111111000101010101101;
assign LUT_4[2818] = 32'b11111111111111111110111001011001;
assign LUT_4[2819] = 32'b11111111111111111000000101010001;
assign LUT_4[2820] = 32'b11111111111111111100011111010001;
assign LUT_4[2821] = 32'b11111111111111110101101011001001;
assign LUT_4[2822] = 32'b11111111111111111011111001110101;
assign LUT_4[2823] = 32'b11111111111111110101000101101101;
assign LUT_4[2824] = 32'b11111111111111111000101011001010;
assign LUT_4[2825] = 32'b11111111111111110001110111000010;
assign LUT_4[2826] = 32'b11111111111111111000000101101110;
assign LUT_4[2827] = 32'b11111111111111110001010001100110;
assign LUT_4[2828] = 32'b11111111111111110101101011100110;
assign LUT_4[2829] = 32'b11111111111111101110110111011110;
assign LUT_4[2830] = 32'b11111111111111110101000110001010;
assign LUT_4[2831] = 32'b11111111111111101110010010000010;
assign LUT_4[2832] = 32'b11111111111111111101010000100011;
assign LUT_4[2833] = 32'b11111111111111110110011100011011;
assign LUT_4[2834] = 32'b11111111111111111100101011000111;
assign LUT_4[2835] = 32'b11111111111111110101110110111111;
assign LUT_4[2836] = 32'b11111111111111111010010000111111;
assign LUT_4[2837] = 32'b11111111111111110011011100110111;
assign LUT_4[2838] = 32'b11111111111111111001101011100011;
assign LUT_4[2839] = 32'b11111111111111110010110111011011;
assign LUT_4[2840] = 32'b11111111111111110110011100111000;
assign LUT_4[2841] = 32'b11111111111111101111101000110000;
assign LUT_4[2842] = 32'b11111111111111110101110111011100;
assign LUT_4[2843] = 32'b11111111111111101111000011010100;
assign LUT_4[2844] = 32'b11111111111111110011011101010100;
assign LUT_4[2845] = 32'b11111111111111101100101001001100;
assign LUT_4[2846] = 32'b11111111111111110010110111111000;
assign LUT_4[2847] = 32'b11111111111111101100000011110000;
assign LUT_4[2848] = 32'b11111111111111111101111001111100;
assign LUT_4[2849] = 32'b11111111111111110111000101110100;
assign LUT_4[2850] = 32'b11111111111111111101010100100000;
assign LUT_4[2851] = 32'b11111111111111110110100000011000;
assign LUT_4[2852] = 32'b11111111111111111010111010011000;
assign LUT_4[2853] = 32'b11111111111111110100000110010000;
assign LUT_4[2854] = 32'b11111111111111111010010100111100;
assign LUT_4[2855] = 32'b11111111111111110011100000110100;
assign LUT_4[2856] = 32'b11111111111111110111000110010001;
assign LUT_4[2857] = 32'b11111111111111110000010010001001;
assign LUT_4[2858] = 32'b11111111111111110110100000110101;
assign LUT_4[2859] = 32'b11111111111111101111101100101101;
assign LUT_4[2860] = 32'b11111111111111110100000110101101;
assign LUT_4[2861] = 32'b11111111111111101101010010100101;
assign LUT_4[2862] = 32'b11111111111111110011100001010001;
assign LUT_4[2863] = 32'b11111111111111101100101101001001;
assign LUT_4[2864] = 32'b11111111111111111011101011101010;
assign LUT_4[2865] = 32'b11111111111111110100110111100010;
assign LUT_4[2866] = 32'b11111111111111111011000110001110;
assign LUT_4[2867] = 32'b11111111111111110100010010000110;
assign LUT_4[2868] = 32'b11111111111111111000101100000110;
assign LUT_4[2869] = 32'b11111111111111110001110111111110;
assign LUT_4[2870] = 32'b11111111111111111000000110101010;
assign LUT_4[2871] = 32'b11111111111111110001010010100010;
assign LUT_4[2872] = 32'b11111111111111110100110111111111;
assign LUT_4[2873] = 32'b11111111111111101110000011110111;
assign LUT_4[2874] = 32'b11111111111111110100010010100011;
assign LUT_4[2875] = 32'b11111111111111101101011110011011;
assign LUT_4[2876] = 32'b11111111111111110001111000011011;
assign LUT_4[2877] = 32'b11111111111111101011000100010011;
assign LUT_4[2878] = 32'b11111111111111110001010010111111;
assign LUT_4[2879] = 32'b11111111111111101010011110110111;
assign LUT_4[2880] = 32'b00000000000000000000110110001001;
assign LUT_4[2881] = 32'b11111111111111111010000010000001;
assign LUT_4[2882] = 32'b00000000000000000000010000101101;
assign LUT_4[2883] = 32'b11111111111111111001011100100101;
assign LUT_4[2884] = 32'b11111111111111111101110110100101;
assign LUT_4[2885] = 32'b11111111111111110111000010011101;
assign LUT_4[2886] = 32'b11111111111111111101010001001001;
assign LUT_4[2887] = 32'b11111111111111110110011101000001;
assign LUT_4[2888] = 32'b11111111111111111010000010011110;
assign LUT_4[2889] = 32'b11111111111111110011001110010110;
assign LUT_4[2890] = 32'b11111111111111111001011101000010;
assign LUT_4[2891] = 32'b11111111111111110010101000111010;
assign LUT_4[2892] = 32'b11111111111111110111000010111010;
assign LUT_4[2893] = 32'b11111111111111110000001110110010;
assign LUT_4[2894] = 32'b11111111111111110110011101011110;
assign LUT_4[2895] = 32'b11111111111111101111101001010110;
assign LUT_4[2896] = 32'b11111111111111111110100111110111;
assign LUT_4[2897] = 32'b11111111111111110111110011101111;
assign LUT_4[2898] = 32'b11111111111111111110000010011011;
assign LUT_4[2899] = 32'b11111111111111110111001110010011;
assign LUT_4[2900] = 32'b11111111111111111011101000010011;
assign LUT_4[2901] = 32'b11111111111111110100110100001011;
assign LUT_4[2902] = 32'b11111111111111111011000010110111;
assign LUT_4[2903] = 32'b11111111111111110100001110101111;
assign LUT_4[2904] = 32'b11111111111111110111110100001100;
assign LUT_4[2905] = 32'b11111111111111110001000000000100;
assign LUT_4[2906] = 32'b11111111111111110111001110110000;
assign LUT_4[2907] = 32'b11111111111111110000011010101000;
assign LUT_4[2908] = 32'b11111111111111110100110100101000;
assign LUT_4[2909] = 32'b11111111111111101110000000100000;
assign LUT_4[2910] = 32'b11111111111111110100001111001100;
assign LUT_4[2911] = 32'b11111111111111101101011011000100;
assign LUT_4[2912] = 32'b11111111111111111111010001010000;
assign LUT_4[2913] = 32'b11111111111111111000011101001000;
assign LUT_4[2914] = 32'b11111111111111111110101011110100;
assign LUT_4[2915] = 32'b11111111111111110111110111101100;
assign LUT_4[2916] = 32'b11111111111111111100010001101100;
assign LUT_4[2917] = 32'b11111111111111110101011101100100;
assign LUT_4[2918] = 32'b11111111111111111011101100010000;
assign LUT_4[2919] = 32'b11111111111111110100111000001000;
assign LUT_4[2920] = 32'b11111111111111111000011101100101;
assign LUT_4[2921] = 32'b11111111111111110001101001011101;
assign LUT_4[2922] = 32'b11111111111111110111111000001001;
assign LUT_4[2923] = 32'b11111111111111110001000100000001;
assign LUT_4[2924] = 32'b11111111111111110101011110000001;
assign LUT_4[2925] = 32'b11111111111111101110101001111001;
assign LUT_4[2926] = 32'b11111111111111110100111000100101;
assign LUT_4[2927] = 32'b11111111111111101110000100011101;
assign LUT_4[2928] = 32'b11111111111111111101000010111110;
assign LUT_4[2929] = 32'b11111111111111110110001110110110;
assign LUT_4[2930] = 32'b11111111111111111100011101100010;
assign LUT_4[2931] = 32'b11111111111111110101101001011010;
assign LUT_4[2932] = 32'b11111111111111111010000011011010;
assign LUT_4[2933] = 32'b11111111111111110011001111010010;
assign LUT_4[2934] = 32'b11111111111111111001011101111110;
assign LUT_4[2935] = 32'b11111111111111110010101001110110;
assign LUT_4[2936] = 32'b11111111111111110110001111010011;
assign LUT_4[2937] = 32'b11111111111111101111011011001011;
assign LUT_4[2938] = 32'b11111111111111110101101001110111;
assign LUT_4[2939] = 32'b11111111111111101110110101101111;
assign LUT_4[2940] = 32'b11111111111111110011001111101111;
assign LUT_4[2941] = 32'b11111111111111101100011011100111;
assign LUT_4[2942] = 32'b11111111111111110010101010010011;
assign LUT_4[2943] = 32'b11111111111111101011110110001011;
assign LUT_4[2944] = 32'b00000000000000000010000100111101;
assign LUT_4[2945] = 32'b11111111111111111011010000110101;
assign LUT_4[2946] = 32'b00000000000000000001011111100001;
assign LUT_4[2947] = 32'b11111111111111111010101011011001;
assign LUT_4[2948] = 32'b11111111111111111111000101011001;
assign LUT_4[2949] = 32'b11111111111111111000010001010001;
assign LUT_4[2950] = 32'b11111111111111111110011111111101;
assign LUT_4[2951] = 32'b11111111111111110111101011110101;
assign LUT_4[2952] = 32'b11111111111111111011010001010010;
assign LUT_4[2953] = 32'b11111111111111110100011101001010;
assign LUT_4[2954] = 32'b11111111111111111010101011110110;
assign LUT_4[2955] = 32'b11111111111111110011110111101110;
assign LUT_4[2956] = 32'b11111111111111111000010001101110;
assign LUT_4[2957] = 32'b11111111111111110001011101100110;
assign LUT_4[2958] = 32'b11111111111111110111101100010010;
assign LUT_4[2959] = 32'b11111111111111110000111000001010;
assign LUT_4[2960] = 32'b11111111111111111111110110101011;
assign LUT_4[2961] = 32'b11111111111111111001000010100011;
assign LUT_4[2962] = 32'b11111111111111111111010001001111;
assign LUT_4[2963] = 32'b11111111111111111000011101000111;
assign LUT_4[2964] = 32'b11111111111111111100110111000111;
assign LUT_4[2965] = 32'b11111111111111110110000010111111;
assign LUT_4[2966] = 32'b11111111111111111100010001101011;
assign LUT_4[2967] = 32'b11111111111111110101011101100011;
assign LUT_4[2968] = 32'b11111111111111111001000011000000;
assign LUT_4[2969] = 32'b11111111111111110010001110111000;
assign LUT_4[2970] = 32'b11111111111111111000011101100100;
assign LUT_4[2971] = 32'b11111111111111110001101001011100;
assign LUT_4[2972] = 32'b11111111111111110110000011011100;
assign LUT_4[2973] = 32'b11111111111111101111001111010100;
assign LUT_4[2974] = 32'b11111111111111110101011110000000;
assign LUT_4[2975] = 32'b11111111111111101110101001111000;
assign LUT_4[2976] = 32'b00000000000000000000100000000100;
assign LUT_4[2977] = 32'b11111111111111111001101011111100;
assign LUT_4[2978] = 32'b11111111111111111111111010101000;
assign LUT_4[2979] = 32'b11111111111111111001000110100000;
assign LUT_4[2980] = 32'b11111111111111111101100000100000;
assign LUT_4[2981] = 32'b11111111111111110110101100011000;
assign LUT_4[2982] = 32'b11111111111111111100111011000100;
assign LUT_4[2983] = 32'b11111111111111110110000110111100;
assign LUT_4[2984] = 32'b11111111111111111001101100011001;
assign LUT_4[2985] = 32'b11111111111111110010111000010001;
assign LUT_4[2986] = 32'b11111111111111111001000110111101;
assign LUT_4[2987] = 32'b11111111111111110010010010110101;
assign LUT_4[2988] = 32'b11111111111111110110101100110101;
assign LUT_4[2989] = 32'b11111111111111101111111000101101;
assign LUT_4[2990] = 32'b11111111111111110110000111011001;
assign LUT_4[2991] = 32'b11111111111111101111010011010001;
assign LUT_4[2992] = 32'b11111111111111111110010001110010;
assign LUT_4[2993] = 32'b11111111111111110111011101101010;
assign LUT_4[2994] = 32'b11111111111111111101101100010110;
assign LUT_4[2995] = 32'b11111111111111110110111000001110;
assign LUT_4[2996] = 32'b11111111111111111011010010001110;
assign LUT_4[2997] = 32'b11111111111111110100011110000110;
assign LUT_4[2998] = 32'b11111111111111111010101100110010;
assign LUT_4[2999] = 32'b11111111111111110011111000101010;
assign LUT_4[3000] = 32'b11111111111111110111011110000111;
assign LUT_4[3001] = 32'b11111111111111110000101001111111;
assign LUT_4[3002] = 32'b11111111111111110110111000101011;
assign LUT_4[3003] = 32'b11111111111111110000000100100011;
assign LUT_4[3004] = 32'b11111111111111110100011110100011;
assign LUT_4[3005] = 32'b11111111111111101101101010011011;
assign LUT_4[3006] = 32'b11111111111111110011111001000111;
assign LUT_4[3007] = 32'b11111111111111101101000100111111;
assign LUT_4[3008] = 32'b00000000000000000011011100010001;
assign LUT_4[3009] = 32'b11111111111111111100101000001001;
assign LUT_4[3010] = 32'b00000000000000000010110110110101;
assign LUT_4[3011] = 32'b11111111111111111100000010101101;
assign LUT_4[3012] = 32'b00000000000000000000011100101101;
assign LUT_4[3013] = 32'b11111111111111111001101000100101;
assign LUT_4[3014] = 32'b11111111111111111111110111010001;
assign LUT_4[3015] = 32'b11111111111111111001000011001001;
assign LUT_4[3016] = 32'b11111111111111111100101000100110;
assign LUT_4[3017] = 32'b11111111111111110101110100011110;
assign LUT_4[3018] = 32'b11111111111111111100000011001010;
assign LUT_4[3019] = 32'b11111111111111110101001111000010;
assign LUT_4[3020] = 32'b11111111111111111001101001000010;
assign LUT_4[3021] = 32'b11111111111111110010110100111010;
assign LUT_4[3022] = 32'b11111111111111111001000011100110;
assign LUT_4[3023] = 32'b11111111111111110010001111011110;
assign LUT_4[3024] = 32'b00000000000000000001001101111111;
assign LUT_4[3025] = 32'b11111111111111111010011001110111;
assign LUT_4[3026] = 32'b00000000000000000000101000100011;
assign LUT_4[3027] = 32'b11111111111111111001110100011011;
assign LUT_4[3028] = 32'b11111111111111111110001110011011;
assign LUT_4[3029] = 32'b11111111111111110111011010010011;
assign LUT_4[3030] = 32'b11111111111111111101101000111111;
assign LUT_4[3031] = 32'b11111111111111110110110100110111;
assign LUT_4[3032] = 32'b11111111111111111010011010010100;
assign LUT_4[3033] = 32'b11111111111111110011100110001100;
assign LUT_4[3034] = 32'b11111111111111111001110100111000;
assign LUT_4[3035] = 32'b11111111111111110011000000110000;
assign LUT_4[3036] = 32'b11111111111111110111011010110000;
assign LUT_4[3037] = 32'b11111111111111110000100110101000;
assign LUT_4[3038] = 32'b11111111111111110110110101010100;
assign LUT_4[3039] = 32'b11111111111111110000000001001100;
assign LUT_4[3040] = 32'b00000000000000000001110111011000;
assign LUT_4[3041] = 32'b11111111111111111011000011010000;
assign LUT_4[3042] = 32'b00000000000000000001010001111100;
assign LUT_4[3043] = 32'b11111111111111111010011101110100;
assign LUT_4[3044] = 32'b11111111111111111110110111110100;
assign LUT_4[3045] = 32'b11111111111111111000000011101100;
assign LUT_4[3046] = 32'b11111111111111111110010010011000;
assign LUT_4[3047] = 32'b11111111111111110111011110010000;
assign LUT_4[3048] = 32'b11111111111111111011000011101101;
assign LUT_4[3049] = 32'b11111111111111110100001111100101;
assign LUT_4[3050] = 32'b11111111111111111010011110010001;
assign LUT_4[3051] = 32'b11111111111111110011101010001001;
assign LUT_4[3052] = 32'b11111111111111111000000100001001;
assign LUT_4[3053] = 32'b11111111111111110001010000000001;
assign LUT_4[3054] = 32'b11111111111111110111011110101101;
assign LUT_4[3055] = 32'b11111111111111110000101010100101;
assign LUT_4[3056] = 32'b11111111111111111111101001000110;
assign LUT_4[3057] = 32'b11111111111111111000110100111110;
assign LUT_4[3058] = 32'b11111111111111111111000011101010;
assign LUT_4[3059] = 32'b11111111111111111000001111100010;
assign LUT_4[3060] = 32'b11111111111111111100101001100010;
assign LUT_4[3061] = 32'b11111111111111110101110101011010;
assign LUT_4[3062] = 32'b11111111111111111100000100000110;
assign LUT_4[3063] = 32'b11111111111111110101001111111110;
assign LUT_4[3064] = 32'b11111111111111111000110101011011;
assign LUT_4[3065] = 32'b11111111111111110010000001010011;
assign LUT_4[3066] = 32'b11111111111111111000001111111111;
assign LUT_4[3067] = 32'b11111111111111110001011011110111;
assign LUT_4[3068] = 32'b11111111111111110101110101110111;
assign LUT_4[3069] = 32'b11111111111111101111000001101111;
assign LUT_4[3070] = 32'b11111111111111110101010000011011;
assign LUT_4[3071] = 32'b11111111111111101110011100010011;
assign LUT_4[3072] = 32'b11111111111111111101001001101001;
assign LUT_4[3073] = 32'b11111111111111110110010101100001;
assign LUT_4[3074] = 32'b11111111111111111100100100001101;
assign LUT_4[3075] = 32'b11111111111111110101110000000101;
assign LUT_4[3076] = 32'b11111111111111111010001010000101;
assign LUT_4[3077] = 32'b11111111111111110011010101111101;
assign LUT_4[3078] = 32'b11111111111111111001100100101001;
assign LUT_4[3079] = 32'b11111111111111110010110000100001;
assign LUT_4[3080] = 32'b11111111111111110110010101111110;
assign LUT_4[3081] = 32'b11111111111111101111100001110110;
assign LUT_4[3082] = 32'b11111111111111110101110000100010;
assign LUT_4[3083] = 32'b11111111111111101110111100011010;
assign LUT_4[3084] = 32'b11111111111111110011010110011010;
assign LUT_4[3085] = 32'b11111111111111101100100010010010;
assign LUT_4[3086] = 32'b11111111111111110010110000111110;
assign LUT_4[3087] = 32'b11111111111111101011111100110110;
assign LUT_4[3088] = 32'b11111111111111111010111011010111;
assign LUT_4[3089] = 32'b11111111111111110100000111001111;
assign LUT_4[3090] = 32'b11111111111111111010010101111011;
assign LUT_4[3091] = 32'b11111111111111110011100001110011;
assign LUT_4[3092] = 32'b11111111111111110111111011110011;
assign LUT_4[3093] = 32'b11111111111111110001000111101011;
assign LUT_4[3094] = 32'b11111111111111110111010110010111;
assign LUT_4[3095] = 32'b11111111111111110000100010001111;
assign LUT_4[3096] = 32'b11111111111111110100000111101100;
assign LUT_4[3097] = 32'b11111111111111101101010011100100;
assign LUT_4[3098] = 32'b11111111111111110011100010010000;
assign LUT_4[3099] = 32'b11111111111111101100101110001000;
assign LUT_4[3100] = 32'b11111111111111110001001000001000;
assign LUT_4[3101] = 32'b11111111111111101010010100000000;
assign LUT_4[3102] = 32'b11111111111111110000100010101100;
assign LUT_4[3103] = 32'b11111111111111101001101110100100;
assign LUT_4[3104] = 32'b11111111111111111011100100110000;
assign LUT_4[3105] = 32'b11111111111111110100110000101000;
assign LUT_4[3106] = 32'b11111111111111111010111111010100;
assign LUT_4[3107] = 32'b11111111111111110100001011001100;
assign LUT_4[3108] = 32'b11111111111111111000100101001100;
assign LUT_4[3109] = 32'b11111111111111110001110001000100;
assign LUT_4[3110] = 32'b11111111111111110111111111110000;
assign LUT_4[3111] = 32'b11111111111111110001001011101000;
assign LUT_4[3112] = 32'b11111111111111110100110001000101;
assign LUT_4[3113] = 32'b11111111111111101101111100111101;
assign LUT_4[3114] = 32'b11111111111111110100001011101001;
assign LUT_4[3115] = 32'b11111111111111101101010111100001;
assign LUT_4[3116] = 32'b11111111111111110001110001100001;
assign LUT_4[3117] = 32'b11111111111111101010111101011001;
assign LUT_4[3118] = 32'b11111111111111110001001100000101;
assign LUT_4[3119] = 32'b11111111111111101010010111111101;
assign LUT_4[3120] = 32'b11111111111111111001010110011110;
assign LUT_4[3121] = 32'b11111111111111110010100010010110;
assign LUT_4[3122] = 32'b11111111111111111000110001000010;
assign LUT_4[3123] = 32'b11111111111111110001111100111010;
assign LUT_4[3124] = 32'b11111111111111110110010110111010;
assign LUT_4[3125] = 32'b11111111111111101111100010110010;
assign LUT_4[3126] = 32'b11111111111111110101110001011110;
assign LUT_4[3127] = 32'b11111111111111101110111101010110;
assign LUT_4[3128] = 32'b11111111111111110010100010110011;
assign LUT_4[3129] = 32'b11111111111111101011101110101011;
assign LUT_4[3130] = 32'b11111111111111110001111101010111;
assign LUT_4[3131] = 32'b11111111111111101011001001001111;
assign LUT_4[3132] = 32'b11111111111111101111100011001111;
assign LUT_4[3133] = 32'b11111111111111101000101111000111;
assign LUT_4[3134] = 32'b11111111111111101110111101110011;
assign LUT_4[3135] = 32'b11111111111111101000001001101011;
assign LUT_4[3136] = 32'b11111111111111111110100000111101;
assign LUT_4[3137] = 32'b11111111111111110111101100110101;
assign LUT_4[3138] = 32'b11111111111111111101111011100001;
assign LUT_4[3139] = 32'b11111111111111110111000111011001;
assign LUT_4[3140] = 32'b11111111111111111011100001011001;
assign LUT_4[3141] = 32'b11111111111111110100101101010001;
assign LUT_4[3142] = 32'b11111111111111111010111011111101;
assign LUT_4[3143] = 32'b11111111111111110100000111110101;
assign LUT_4[3144] = 32'b11111111111111110111101101010010;
assign LUT_4[3145] = 32'b11111111111111110000111001001010;
assign LUT_4[3146] = 32'b11111111111111110111000111110110;
assign LUT_4[3147] = 32'b11111111111111110000010011101110;
assign LUT_4[3148] = 32'b11111111111111110100101101101110;
assign LUT_4[3149] = 32'b11111111111111101101111001100110;
assign LUT_4[3150] = 32'b11111111111111110100001000010010;
assign LUT_4[3151] = 32'b11111111111111101101010100001010;
assign LUT_4[3152] = 32'b11111111111111111100010010101011;
assign LUT_4[3153] = 32'b11111111111111110101011110100011;
assign LUT_4[3154] = 32'b11111111111111111011101101001111;
assign LUT_4[3155] = 32'b11111111111111110100111001000111;
assign LUT_4[3156] = 32'b11111111111111111001010011000111;
assign LUT_4[3157] = 32'b11111111111111110010011110111111;
assign LUT_4[3158] = 32'b11111111111111111000101101101011;
assign LUT_4[3159] = 32'b11111111111111110001111001100011;
assign LUT_4[3160] = 32'b11111111111111110101011111000000;
assign LUT_4[3161] = 32'b11111111111111101110101010111000;
assign LUT_4[3162] = 32'b11111111111111110100111001100100;
assign LUT_4[3163] = 32'b11111111111111101110000101011100;
assign LUT_4[3164] = 32'b11111111111111110010011111011100;
assign LUT_4[3165] = 32'b11111111111111101011101011010100;
assign LUT_4[3166] = 32'b11111111111111110001111010000000;
assign LUT_4[3167] = 32'b11111111111111101011000101111000;
assign LUT_4[3168] = 32'b11111111111111111100111100000100;
assign LUT_4[3169] = 32'b11111111111111110110000111111100;
assign LUT_4[3170] = 32'b11111111111111111100010110101000;
assign LUT_4[3171] = 32'b11111111111111110101100010100000;
assign LUT_4[3172] = 32'b11111111111111111001111100100000;
assign LUT_4[3173] = 32'b11111111111111110011001000011000;
assign LUT_4[3174] = 32'b11111111111111111001010111000100;
assign LUT_4[3175] = 32'b11111111111111110010100010111100;
assign LUT_4[3176] = 32'b11111111111111110110001000011001;
assign LUT_4[3177] = 32'b11111111111111101111010100010001;
assign LUT_4[3178] = 32'b11111111111111110101100010111101;
assign LUT_4[3179] = 32'b11111111111111101110101110110101;
assign LUT_4[3180] = 32'b11111111111111110011001000110101;
assign LUT_4[3181] = 32'b11111111111111101100010100101101;
assign LUT_4[3182] = 32'b11111111111111110010100011011001;
assign LUT_4[3183] = 32'b11111111111111101011101111010001;
assign LUT_4[3184] = 32'b11111111111111111010101101110010;
assign LUT_4[3185] = 32'b11111111111111110011111001101010;
assign LUT_4[3186] = 32'b11111111111111111010001000010110;
assign LUT_4[3187] = 32'b11111111111111110011010100001110;
assign LUT_4[3188] = 32'b11111111111111110111101110001110;
assign LUT_4[3189] = 32'b11111111111111110000111010000110;
assign LUT_4[3190] = 32'b11111111111111110111001000110010;
assign LUT_4[3191] = 32'b11111111111111110000010100101010;
assign LUT_4[3192] = 32'b11111111111111110011111010000111;
assign LUT_4[3193] = 32'b11111111111111101101000101111111;
assign LUT_4[3194] = 32'b11111111111111110011010100101011;
assign LUT_4[3195] = 32'b11111111111111101100100000100011;
assign LUT_4[3196] = 32'b11111111111111110000111010100011;
assign LUT_4[3197] = 32'b11111111111111101010000110011011;
assign LUT_4[3198] = 32'b11111111111111110000010101000111;
assign LUT_4[3199] = 32'b11111111111111101001100000111111;
assign LUT_4[3200] = 32'b11111111111111111111101111110001;
assign LUT_4[3201] = 32'b11111111111111111000111011101001;
assign LUT_4[3202] = 32'b11111111111111111111001010010101;
assign LUT_4[3203] = 32'b11111111111111111000010110001101;
assign LUT_4[3204] = 32'b11111111111111111100110000001101;
assign LUT_4[3205] = 32'b11111111111111110101111100000101;
assign LUT_4[3206] = 32'b11111111111111111100001010110001;
assign LUT_4[3207] = 32'b11111111111111110101010110101001;
assign LUT_4[3208] = 32'b11111111111111111000111100000110;
assign LUT_4[3209] = 32'b11111111111111110010000111111110;
assign LUT_4[3210] = 32'b11111111111111111000010110101010;
assign LUT_4[3211] = 32'b11111111111111110001100010100010;
assign LUT_4[3212] = 32'b11111111111111110101111100100010;
assign LUT_4[3213] = 32'b11111111111111101111001000011010;
assign LUT_4[3214] = 32'b11111111111111110101010111000110;
assign LUT_4[3215] = 32'b11111111111111101110100010111110;
assign LUT_4[3216] = 32'b11111111111111111101100001011111;
assign LUT_4[3217] = 32'b11111111111111110110101101010111;
assign LUT_4[3218] = 32'b11111111111111111100111100000011;
assign LUT_4[3219] = 32'b11111111111111110110000111111011;
assign LUT_4[3220] = 32'b11111111111111111010100001111011;
assign LUT_4[3221] = 32'b11111111111111110011101101110011;
assign LUT_4[3222] = 32'b11111111111111111001111100011111;
assign LUT_4[3223] = 32'b11111111111111110011001000010111;
assign LUT_4[3224] = 32'b11111111111111110110101101110100;
assign LUT_4[3225] = 32'b11111111111111101111111001101100;
assign LUT_4[3226] = 32'b11111111111111110110001000011000;
assign LUT_4[3227] = 32'b11111111111111101111010100010000;
assign LUT_4[3228] = 32'b11111111111111110011101110010000;
assign LUT_4[3229] = 32'b11111111111111101100111010001000;
assign LUT_4[3230] = 32'b11111111111111110011001000110100;
assign LUT_4[3231] = 32'b11111111111111101100010100101100;
assign LUT_4[3232] = 32'b11111111111111111110001010111000;
assign LUT_4[3233] = 32'b11111111111111110111010110110000;
assign LUT_4[3234] = 32'b11111111111111111101100101011100;
assign LUT_4[3235] = 32'b11111111111111110110110001010100;
assign LUT_4[3236] = 32'b11111111111111111011001011010100;
assign LUT_4[3237] = 32'b11111111111111110100010111001100;
assign LUT_4[3238] = 32'b11111111111111111010100101111000;
assign LUT_4[3239] = 32'b11111111111111110011110001110000;
assign LUT_4[3240] = 32'b11111111111111110111010111001101;
assign LUT_4[3241] = 32'b11111111111111110000100011000101;
assign LUT_4[3242] = 32'b11111111111111110110110001110001;
assign LUT_4[3243] = 32'b11111111111111101111111101101001;
assign LUT_4[3244] = 32'b11111111111111110100010111101001;
assign LUT_4[3245] = 32'b11111111111111101101100011100001;
assign LUT_4[3246] = 32'b11111111111111110011110010001101;
assign LUT_4[3247] = 32'b11111111111111101100111110000101;
assign LUT_4[3248] = 32'b11111111111111111011111100100110;
assign LUT_4[3249] = 32'b11111111111111110101001000011110;
assign LUT_4[3250] = 32'b11111111111111111011010111001010;
assign LUT_4[3251] = 32'b11111111111111110100100011000010;
assign LUT_4[3252] = 32'b11111111111111111000111101000010;
assign LUT_4[3253] = 32'b11111111111111110010001000111010;
assign LUT_4[3254] = 32'b11111111111111111000010111100110;
assign LUT_4[3255] = 32'b11111111111111110001100011011110;
assign LUT_4[3256] = 32'b11111111111111110101001000111011;
assign LUT_4[3257] = 32'b11111111111111101110010100110011;
assign LUT_4[3258] = 32'b11111111111111110100100011011111;
assign LUT_4[3259] = 32'b11111111111111101101101111010111;
assign LUT_4[3260] = 32'b11111111111111110010001001010111;
assign LUT_4[3261] = 32'b11111111111111101011010101001111;
assign LUT_4[3262] = 32'b11111111111111110001100011111011;
assign LUT_4[3263] = 32'b11111111111111101010101111110011;
assign LUT_4[3264] = 32'b00000000000000000001000111000101;
assign LUT_4[3265] = 32'b11111111111111111010010010111101;
assign LUT_4[3266] = 32'b00000000000000000000100001101001;
assign LUT_4[3267] = 32'b11111111111111111001101101100001;
assign LUT_4[3268] = 32'b11111111111111111110000111100001;
assign LUT_4[3269] = 32'b11111111111111110111010011011001;
assign LUT_4[3270] = 32'b11111111111111111101100010000101;
assign LUT_4[3271] = 32'b11111111111111110110101101111101;
assign LUT_4[3272] = 32'b11111111111111111010010011011010;
assign LUT_4[3273] = 32'b11111111111111110011011111010010;
assign LUT_4[3274] = 32'b11111111111111111001101101111110;
assign LUT_4[3275] = 32'b11111111111111110010111001110110;
assign LUT_4[3276] = 32'b11111111111111110111010011110110;
assign LUT_4[3277] = 32'b11111111111111110000011111101110;
assign LUT_4[3278] = 32'b11111111111111110110101110011010;
assign LUT_4[3279] = 32'b11111111111111101111111010010010;
assign LUT_4[3280] = 32'b11111111111111111110111000110011;
assign LUT_4[3281] = 32'b11111111111111111000000100101011;
assign LUT_4[3282] = 32'b11111111111111111110010011010111;
assign LUT_4[3283] = 32'b11111111111111110111011111001111;
assign LUT_4[3284] = 32'b11111111111111111011111001001111;
assign LUT_4[3285] = 32'b11111111111111110101000101000111;
assign LUT_4[3286] = 32'b11111111111111111011010011110011;
assign LUT_4[3287] = 32'b11111111111111110100011111101011;
assign LUT_4[3288] = 32'b11111111111111111000000101001000;
assign LUT_4[3289] = 32'b11111111111111110001010001000000;
assign LUT_4[3290] = 32'b11111111111111110111011111101100;
assign LUT_4[3291] = 32'b11111111111111110000101011100100;
assign LUT_4[3292] = 32'b11111111111111110101000101100100;
assign LUT_4[3293] = 32'b11111111111111101110010001011100;
assign LUT_4[3294] = 32'b11111111111111110100100000001000;
assign LUT_4[3295] = 32'b11111111111111101101101100000000;
assign LUT_4[3296] = 32'b11111111111111111111100010001100;
assign LUT_4[3297] = 32'b11111111111111111000101110000100;
assign LUT_4[3298] = 32'b11111111111111111110111100110000;
assign LUT_4[3299] = 32'b11111111111111111000001000101000;
assign LUT_4[3300] = 32'b11111111111111111100100010101000;
assign LUT_4[3301] = 32'b11111111111111110101101110100000;
assign LUT_4[3302] = 32'b11111111111111111011111101001100;
assign LUT_4[3303] = 32'b11111111111111110101001001000100;
assign LUT_4[3304] = 32'b11111111111111111000101110100001;
assign LUT_4[3305] = 32'b11111111111111110001111010011001;
assign LUT_4[3306] = 32'b11111111111111111000001001000101;
assign LUT_4[3307] = 32'b11111111111111110001010100111101;
assign LUT_4[3308] = 32'b11111111111111110101101110111101;
assign LUT_4[3309] = 32'b11111111111111101110111010110101;
assign LUT_4[3310] = 32'b11111111111111110101001001100001;
assign LUT_4[3311] = 32'b11111111111111101110010101011001;
assign LUT_4[3312] = 32'b11111111111111111101010011111010;
assign LUT_4[3313] = 32'b11111111111111110110011111110010;
assign LUT_4[3314] = 32'b11111111111111111100101110011110;
assign LUT_4[3315] = 32'b11111111111111110101111010010110;
assign LUT_4[3316] = 32'b11111111111111111010010100010110;
assign LUT_4[3317] = 32'b11111111111111110011100000001110;
assign LUT_4[3318] = 32'b11111111111111111001101110111010;
assign LUT_4[3319] = 32'b11111111111111110010111010110010;
assign LUT_4[3320] = 32'b11111111111111110110100000001111;
assign LUT_4[3321] = 32'b11111111111111101111101100000111;
assign LUT_4[3322] = 32'b11111111111111110101111010110011;
assign LUT_4[3323] = 32'b11111111111111101111000110101011;
assign LUT_4[3324] = 32'b11111111111111110011100000101011;
assign LUT_4[3325] = 32'b11111111111111101100101100100011;
assign LUT_4[3326] = 32'b11111111111111110010111011001111;
assign LUT_4[3327] = 32'b11111111111111101100000111000111;
assign LUT_4[3328] = 32'b00000000000000000010000101001100;
assign LUT_4[3329] = 32'b11111111111111111011010001000100;
assign LUT_4[3330] = 32'b00000000000000000001011111110000;
assign LUT_4[3331] = 32'b11111111111111111010101011101000;
assign LUT_4[3332] = 32'b11111111111111111111000101101000;
assign LUT_4[3333] = 32'b11111111111111111000010001100000;
assign LUT_4[3334] = 32'b11111111111111111110100000001100;
assign LUT_4[3335] = 32'b11111111111111110111101100000100;
assign LUT_4[3336] = 32'b11111111111111111011010001100001;
assign LUT_4[3337] = 32'b11111111111111110100011101011001;
assign LUT_4[3338] = 32'b11111111111111111010101100000101;
assign LUT_4[3339] = 32'b11111111111111110011110111111101;
assign LUT_4[3340] = 32'b11111111111111111000010001111101;
assign LUT_4[3341] = 32'b11111111111111110001011101110101;
assign LUT_4[3342] = 32'b11111111111111110111101100100001;
assign LUT_4[3343] = 32'b11111111111111110000111000011001;
assign LUT_4[3344] = 32'b11111111111111111111110110111010;
assign LUT_4[3345] = 32'b11111111111111111001000010110010;
assign LUT_4[3346] = 32'b11111111111111111111010001011110;
assign LUT_4[3347] = 32'b11111111111111111000011101010110;
assign LUT_4[3348] = 32'b11111111111111111100110111010110;
assign LUT_4[3349] = 32'b11111111111111110110000011001110;
assign LUT_4[3350] = 32'b11111111111111111100010001111010;
assign LUT_4[3351] = 32'b11111111111111110101011101110010;
assign LUT_4[3352] = 32'b11111111111111111001000011001111;
assign LUT_4[3353] = 32'b11111111111111110010001111000111;
assign LUT_4[3354] = 32'b11111111111111111000011101110011;
assign LUT_4[3355] = 32'b11111111111111110001101001101011;
assign LUT_4[3356] = 32'b11111111111111110110000011101011;
assign LUT_4[3357] = 32'b11111111111111101111001111100011;
assign LUT_4[3358] = 32'b11111111111111110101011110001111;
assign LUT_4[3359] = 32'b11111111111111101110101010000111;
assign LUT_4[3360] = 32'b00000000000000000000100000010011;
assign LUT_4[3361] = 32'b11111111111111111001101100001011;
assign LUT_4[3362] = 32'b11111111111111111111111010110111;
assign LUT_4[3363] = 32'b11111111111111111001000110101111;
assign LUT_4[3364] = 32'b11111111111111111101100000101111;
assign LUT_4[3365] = 32'b11111111111111110110101100100111;
assign LUT_4[3366] = 32'b11111111111111111100111011010011;
assign LUT_4[3367] = 32'b11111111111111110110000111001011;
assign LUT_4[3368] = 32'b11111111111111111001101100101000;
assign LUT_4[3369] = 32'b11111111111111110010111000100000;
assign LUT_4[3370] = 32'b11111111111111111001000111001100;
assign LUT_4[3371] = 32'b11111111111111110010010011000100;
assign LUT_4[3372] = 32'b11111111111111110110101101000100;
assign LUT_4[3373] = 32'b11111111111111101111111000111100;
assign LUT_4[3374] = 32'b11111111111111110110000111101000;
assign LUT_4[3375] = 32'b11111111111111101111010011100000;
assign LUT_4[3376] = 32'b11111111111111111110010010000001;
assign LUT_4[3377] = 32'b11111111111111110111011101111001;
assign LUT_4[3378] = 32'b11111111111111111101101100100101;
assign LUT_4[3379] = 32'b11111111111111110110111000011101;
assign LUT_4[3380] = 32'b11111111111111111011010010011101;
assign LUT_4[3381] = 32'b11111111111111110100011110010101;
assign LUT_4[3382] = 32'b11111111111111111010101101000001;
assign LUT_4[3383] = 32'b11111111111111110011111000111001;
assign LUT_4[3384] = 32'b11111111111111110111011110010110;
assign LUT_4[3385] = 32'b11111111111111110000101010001110;
assign LUT_4[3386] = 32'b11111111111111110110111000111010;
assign LUT_4[3387] = 32'b11111111111111110000000100110010;
assign LUT_4[3388] = 32'b11111111111111110100011110110010;
assign LUT_4[3389] = 32'b11111111111111101101101010101010;
assign LUT_4[3390] = 32'b11111111111111110011111001010110;
assign LUT_4[3391] = 32'b11111111111111101101000101001110;
assign LUT_4[3392] = 32'b00000000000000000011011100100000;
assign LUT_4[3393] = 32'b11111111111111111100101000011000;
assign LUT_4[3394] = 32'b00000000000000000010110111000100;
assign LUT_4[3395] = 32'b11111111111111111100000010111100;
assign LUT_4[3396] = 32'b00000000000000000000011100111100;
assign LUT_4[3397] = 32'b11111111111111111001101000110100;
assign LUT_4[3398] = 32'b11111111111111111111110111100000;
assign LUT_4[3399] = 32'b11111111111111111001000011011000;
assign LUT_4[3400] = 32'b11111111111111111100101000110101;
assign LUT_4[3401] = 32'b11111111111111110101110100101101;
assign LUT_4[3402] = 32'b11111111111111111100000011011001;
assign LUT_4[3403] = 32'b11111111111111110101001111010001;
assign LUT_4[3404] = 32'b11111111111111111001101001010001;
assign LUT_4[3405] = 32'b11111111111111110010110101001001;
assign LUT_4[3406] = 32'b11111111111111111001000011110101;
assign LUT_4[3407] = 32'b11111111111111110010001111101101;
assign LUT_4[3408] = 32'b00000000000000000001001110001110;
assign LUT_4[3409] = 32'b11111111111111111010011010000110;
assign LUT_4[3410] = 32'b00000000000000000000101000110010;
assign LUT_4[3411] = 32'b11111111111111111001110100101010;
assign LUT_4[3412] = 32'b11111111111111111110001110101010;
assign LUT_4[3413] = 32'b11111111111111110111011010100010;
assign LUT_4[3414] = 32'b11111111111111111101101001001110;
assign LUT_4[3415] = 32'b11111111111111110110110101000110;
assign LUT_4[3416] = 32'b11111111111111111010011010100011;
assign LUT_4[3417] = 32'b11111111111111110011100110011011;
assign LUT_4[3418] = 32'b11111111111111111001110101000111;
assign LUT_4[3419] = 32'b11111111111111110011000000111111;
assign LUT_4[3420] = 32'b11111111111111110111011010111111;
assign LUT_4[3421] = 32'b11111111111111110000100110110111;
assign LUT_4[3422] = 32'b11111111111111110110110101100011;
assign LUT_4[3423] = 32'b11111111111111110000000001011011;
assign LUT_4[3424] = 32'b00000000000000000001110111100111;
assign LUT_4[3425] = 32'b11111111111111111011000011011111;
assign LUT_4[3426] = 32'b00000000000000000001010010001011;
assign LUT_4[3427] = 32'b11111111111111111010011110000011;
assign LUT_4[3428] = 32'b11111111111111111110111000000011;
assign LUT_4[3429] = 32'b11111111111111111000000011111011;
assign LUT_4[3430] = 32'b11111111111111111110010010100111;
assign LUT_4[3431] = 32'b11111111111111110111011110011111;
assign LUT_4[3432] = 32'b11111111111111111011000011111100;
assign LUT_4[3433] = 32'b11111111111111110100001111110100;
assign LUT_4[3434] = 32'b11111111111111111010011110100000;
assign LUT_4[3435] = 32'b11111111111111110011101010011000;
assign LUT_4[3436] = 32'b11111111111111111000000100011000;
assign LUT_4[3437] = 32'b11111111111111110001010000010000;
assign LUT_4[3438] = 32'b11111111111111110111011110111100;
assign LUT_4[3439] = 32'b11111111111111110000101010110100;
assign LUT_4[3440] = 32'b11111111111111111111101001010101;
assign LUT_4[3441] = 32'b11111111111111111000110101001101;
assign LUT_4[3442] = 32'b11111111111111111111000011111001;
assign LUT_4[3443] = 32'b11111111111111111000001111110001;
assign LUT_4[3444] = 32'b11111111111111111100101001110001;
assign LUT_4[3445] = 32'b11111111111111110101110101101001;
assign LUT_4[3446] = 32'b11111111111111111100000100010101;
assign LUT_4[3447] = 32'b11111111111111110101010000001101;
assign LUT_4[3448] = 32'b11111111111111111000110101101010;
assign LUT_4[3449] = 32'b11111111111111110010000001100010;
assign LUT_4[3450] = 32'b11111111111111111000010000001110;
assign LUT_4[3451] = 32'b11111111111111110001011100000110;
assign LUT_4[3452] = 32'b11111111111111110101110110000110;
assign LUT_4[3453] = 32'b11111111111111101111000001111110;
assign LUT_4[3454] = 32'b11111111111111110101010000101010;
assign LUT_4[3455] = 32'b11111111111111101110011100100010;
assign LUT_4[3456] = 32'b00000000000000000100101011010100;
assign LUT_4[3457] = 32'b11111111111111111101110111001100;
assign LUT_4[3458] = 32'b00000000000000000100000101111000;
assign LUT_4[3459] = 32'b11111111111111111101010001110000;
assign LUT_4[3460] = 32'b00000000000000000001101011110000;
assign LUT_4[3461] = 32'b11111111111111111010110111101000;
assign LUT_4[3462] = 32'b00000000000000000001000110010100;
assign LUT_4[3463] = 32'b11111111111111111010010010001100;
assign LUT_4[3464] = 32'b11111111111111111101110111101001;
assign LUT_4[3465] = 32'b11111111111111110111000011100001;
assign LUT_4[3466] = 32'b11111111111111111101010010001101;
assign LUT_4[3467] = 32'b11111111111111110110011110000101;
assign LUT_4[3468] = 32'b11111111111111111010111000000101;
assign LUT_4[3469] = 32'b11111111111111110100000011111101;
assign LUT_4[3470] = 32'b11111111111111111010010010101001;
assign LUT_4[3471] = 32'b11111111111111110011011110100001;
assign LUT_4[3472] = 32'b00000000000000000010011101000010;
assign LUT_4[3473] = 32'b11111111111111111011101000111010;
assign LUT_4[3474] = 32'b00000000000000000001110111100110;
assign LUT_4[3475] = 32'b11111111111111111011000011011110;
assign LUT_4[3476] = 32'b11111111111111111111011101011110;
assign LUT_4[3477] = 32'b11111111111111111000101001010110;
assign LUT_4[3478] = 32'b11111111111111111110111000000010;
assign LUT_4[3479] = 32'b11111111111111111000000011111010;
assign LUT_4[3480] = 32'b11111111111111111011101001010111;
assign LUT_4[3481] = 32'b11111111111111110100110101001111;
assign LUT_4[3482] = 32'b11111111111111111011000011111011;
assign LUT_4[3483] = 32'b11111111111111110100001111110011;
assign LUT_4[3484] = 32'b11111111111111111000101001110011;
assign LUT_4[3485] = 32'b11111111111111110001110101101011;
assign LUT_4[3486] = 32'b11111111111111111000000100010111;
assign LUT_4[3487] = 32'b11111111111111110001010000001111;
assign LUT_4[3488] = 32'b00000000000000000011000110011011;
assign LUT_4[3489] = 32'b11111111111111111100010010010011;
assign LUT_4[3490] = 32'b00000000000000000010100000111111;
assign LUT_4[3491] = 32'b11111111111111111011101100110111;
assign LUT_4[3492] = 32'b00000000000000000000000110110111;
assign LUT_4[3493] = 32'b11111111111111111001010010101111;
assign LUT_4[3494] = 32'b11111111111111111111100001011011;
assign LUT_4[3495] = 32'b11111111111111111000101101010011;
assign LUT_4[3496] = 32'b11111111111111111100010010110000;
assign LUT_4[3497] = 32'b11111111111111110101011110101000;
assign LUT_4[3498] = 32'b11111111111111111011101101010100;
assign LUT_4[3499] = 32'b11111111111111110100111001001100;
assign LUT_4[3500] = 32'b11111111111111111001010011001100;
assign LUT_4[3501] = 32'b11111111111111110010011111000100;
assign LUT_4[3502] = 32'b11111111111111111000101101110000;
assign LUT_4[3503] = 32'b11111111111111110001111001101000;
assign LUT_4[3504] = 32'b00000000000000000000111000001001;
assign LUT_4[3505] = 32'b11111111111111111010000100000001;
assign LUT_4[3506] = 32'b00000000000000000000010010101101;
assign LUT_4[3507] = 32'b11111111111111111001011110100101;
assign LUT_4[3508] = 32'b11111111111111111101111000100101;
assign LUT_4[3509] = 32'b11111111111111110111000100011101;
assign LUT_4[3510] = 32'b11111111111111111101010011001001;
assign LUT_4[3511] = 32'b11111111111111110110011111000001;
assign LUT_4[3512] = 32'b11111111111111111010000100011110;
assign LUT_4[3513] = 32'b11111111111111110011010000010110;
assign LUT_4[3514] = 32'b11111111111111111001011111000010;
assign LUT_4[3515] = 32'b11111111111111110010101010111010;
assign LUT_4[3516] = 32'b11111111111111110111000100111010;
assign LUT_4[3517] = 32'b11111111111111110000010000110010;
assign LUT_4[3518] = 32'b11111111111111110110011111011110;
assign LUT_4[3519] = 32'b11111111111111101111101011010110;
assign LUT_4[3520] = 32'b00000000000000000110000010101000;
assign LUT_4[3521] = 32'b11111111111111111111001110100000;
assign LUT_4[3522] = 32'b00000000000000000101011101001100;
assign LUT_4[3523] = 32'b11111111111111111110101001000100;
assign LUT_4[3524] = 32'b00000000000000000011000011000100;
assign LUT_4[3525] = 32'b11111111111111111100001110111100;
assign LUT_4[3526] = 32'b00000000000000000010011101101000;
assign LUT_4[3527] = 32'b11111111111111111011101001100000;
assign LUT_4[3528] = 32'b11111111111111111111001110111101;
assign LUT_4[3529] = 32'b11111111111111111000011010110101;
assign LUT_4[3530] = 32'b11111111111111111110101001100001;
assign LUT_4[3531] = 32'b11111111111111110111110101011001;
assign LUT_4[3532] = 32'b11111111111111111100001111011001;
assign LUT_4[3533] = 32'b11111111111111110101011011010001;
assign LUT_4[3534] = 32'b11111111111111111011101001111101;
assign LUT_4[3535] = 32'b11111111111111110100110101110101;
assign LUT_4[3536] = 32'b00000000000000000011110100010110;
assign LUT_4[3537] = 32'b11111111111111111101000000001110;
assign LUT_4[3538] = 32'b00000000000000000011001110111010;
assign LUT_4[3539] = 32'b11111111111111111100011010110010;
assign LUT_4[3540] = 32'b00000000000000000000110100110010;
assign LUT_4[3541] = 32'b11111111111111111010000000101010;
assign LUT_4[3542] = 32'b00000000000000000000001111010110;
assign LUT_4[3543] = 32'b11111111111111111001011011001110;
assign LUT_4[3544] = 32'b11111111111111111101000000101011;
assign LUT_4[3545] = 32'b11111111111111110110001100100011;
assign LUT_4[3546] = 32'b11111111111111111100011011001111;
assign LUT_4[3547] = 32'b11111111111111110101100111000111;
assign LUT_4[3548] = 32'b11111111111111111010000001000111;
assign LUT_4[3549] = 32'b11111111111111110011001100111111;
assign LUT_4[3550] = 32'b11111111111111111001011011101011;
assign LUT_4[3551] = 32'b11111111111111110010100111100011;
assign LUT_4[3552] = 32'b00000000000000000100011101101111;
assign LUT_4[3553] = 32'b11111111111111111101101001100111;
assign LUT_4[3554] = 32'b00000000000000000011111000010011;
assign LUT_4[3555] = 32'b11111111111111111101000100001011;
assign LUT_4[3556] = 32'b00000000000000000001011110001011;
assign LUT_4[3557] = 32'b11111111111111111010101010000011;
assign LUT_4[3558] = 32'b00000000000000000000111000101111;
assign LUT_4[3559] = 32'b11111111111111111010000100100111;
assign LUT_4[3560] = 32'b11111111111111111101101010000100;
assign LUT_4[3561] = 32'b11111111111111110110110101111100;
assign LUT_4[3562] = 32'b11111111111111111101000100101000;
assign LUT_4[3563] = 32'b11111111111111110110010000100000;
assign LUT_4[3564] = 32'b11111111111111111010101010100000;
assign LUT_4[3565] = 32'b11111111111111110011110110011000;
assign LUT_4[3566] = 32'b11111111111111111010000101000100;
assign LUT_4[3567] = 32'b11111111111111110011010000111100;
assign LUT_4[3568] = 32'b00000000000000000010001111011101;
assign LUT_4[3569] = 32'b11111111111111111011011011010101;
assign LUT_4[3570] = 32'b00000000000000000001101010000001;
assign LUT_4[3571] = 32'b11111111111111111010110101111001;
assign LUT_4[3572] = 32'b11111111111111111111001111111001;
assign LUT_4[3573] = 32'b11111111111111111000011011110001;
assign LUT_4[3574] = 32'b11111111111111111110101010011101;
assign LUT_4[3575] = 32'b11111111111111110111110110010101;
assign LUT_4[3576] = 32'b11111111111111111011011011110010;
assign LUT_4[3577] = 32'b11111111111111110100100111101010;
assign LUT_4[3578] = 32'b11111111111111111010110110010110;
assign LUT_4[3579] = 32'b11111111111111110100000010001110;
assign LUT_4[3580] = 32'b11111111111111111000011100001110;
assign LUT_4[3581] = 32'b11111111111111110001101000000110;
assign LUT_4[3582] = 32'b11111111111111110111110110110010;
assign LUT_4[3583] = 32'b11111111111111110001000010101010;
assign LUT_4[3584] = 32'b11111111111111111100001101110001;
assign LUT_4[3585] = 32'b11111111111111110101011001101001;
assign LUT_4[3586] = 32'b11111111111111111011101000010101;
assign LUT_4[3587] = 32'b11111111111111110100110100001101;
assign LUT_4[3588] = 32'b11111111111111111001001110001101;
assign LUT_4[3589] = 32'b11111111111111110010011010000101;
assign LUT_4[3590] = 32'b11111111111111111000101000110001;
assign LUT_4[3591] = 32'b11111111111111110001110100101001;
assign LUT_4[3592] = 32'b11111111111111110101011010000110;
assign LUT_4[3593] = 32'b11111111111111101110100101111110;
assign LUT_4[3594] = 32'b11111111111111110100110100101010;
assign LUT_4[3595] = 32'b11111111111111101110000000100010;
assign LUT_4[3596] = 32'b11111111111111110010011010100010;
assign LUT_4[3597] = 32'b11111111111111101011100110011010;
assign LUT_4[3598] = 32'b11111111111111110001110101000110;
assign LUT_4[3599] = 32'b11111111111111101011000000111110;
assign LUT_4[3600] = 32'b11111111111111111001111111011111;
assign LUT_4[3601] = 32'b11111111111111110011001011010111;
assign LUT_4[3602] = 32'b11111111111111111001011010000011;
assign LUT_4[3603] = 32'b11111111111111110010100101111011;
assign LUT_4[3604] = 32'b11111111111111110110111111111011;
assign LUT_4[3605] = 32'b11111111111111110000001011110011;
assign LUT_4[3606] = 32'b11111111111111110110011010011111;
assign LUT_4[3607] = 32'b11111111111111101111100110010111;
assign LUT_4[3608] = 32'b11111111111111110011001011110100;
assign LUT_4[3609] = 32'b11111111111111101100010111101100;
assign LUT_4[3610] = 32'b11111111111111110010100110011000;
assign LUT_4[3611] = 32'b11111111111111101011110010010000;
assign LUT_4[3612] = 32'b11111111111111110000001100010000;
assign LUT_4[3613] = 32'b11111111111111101001011000001000;
assign LUT_4[3614] = 32'b11111111111111101111100110110100;
assign LUT_4[3615] = 32'b11111111111111101000110010101100;
assign LUT_4[3616] = 32'b11111111111111111010101000111000;
assign LUT_4[3617] = 32'b11111111111111110011110100110000;
assign LUT_4[3618] = 32'b11111111111111111010000011011100;
assign LUT_4[3619] = 32'b11111111111111110011001111010100;
assign LUT_4[3620] = 32'b11111111111111110111101001010100;
assign LUT_4[3621] = 32'b11111111111111110000110101001100;
assign LUT_4[3622] = 32'b11111111111111110111000011111000;
assign LUT_4[3623] = 32'b11111111111111110000001111110000;
assign LUT_4[3624] = 32'b11111111111111110011110101001101;
assign LUT_4[3625] = 32'b11111111111111101101000001000101;
assign LUT_4[3626] = 32'b11111111111111110011001111110001;
assign LUT_4[3627] = 32'b11111111111111101100011011101001;
assign LUT_4[3628] = 32'b11111111111111110000110101101001;
assign LUT_4[3629] = 32'b11111111111111101010000001100001;
assign LUT_4[3630] = 32'b11111111111111110000010000001101;
assign LUT_4[3631] = 32'b11111111111111101001011100000101;
assign LUT_4[3632] = 32'b11111111111111111000011010100110;
assign LUT_4[3633] = 32'b11111111111111110001100110011110;
assign LUT_4[3634] = 32'b11111111111111110111110101001010;
assign LUT_4[3635] = 32'b11111111111111110001000001000010;
assign LUT_4[3636] = 32'b11111111111111110101011011000010;
assign LUT_4[3637] = 32'b11111111111111101110100110111010;
assign LUT_4[3638] = 32'b11111111111111110100110101100110;
assign LUT_4[3639] = 32'b11111111111111101110000001011110;
assign LUT_4[3640] = 32'b11111111111111110001100110111011;
assign LUT_4[3641] = 32'b11111111111111101010110010110011;
assign LUT_4[3642] = 32'b11111111111111110001000001011111;
assign LUT_4[3643] = 32'b11111111111111101010001101010111;
assign LUT_4[3644] = 32'b11111111111111101110100111010111;
assign LUT_4[3645] = 32'b11111111111111100111110011001111;
assign LUT_4[3646] = 32'b11111111111111101110000001111011;
assign LUT_4[3647] = 32'b11111111111111100111001101110011;
assign LUT_4[3648] = 32'b11111111111111111101100101000101;
assign LUT_4[3649] = 32'b11111111111111110110110000111101;
assign LUT_4[3650] = 32'b11111111111111111100111111101001;
assign LUT_4[3651] = 32'b11111111111111110110001011100001;
assign LUT_4[3652] = 32'b11111111111111111010100101100001;
assign LUT_4[3653] = 32'b11111111111111110011110001011001;
assign LUT_4[3654] = 32'b11111111111111111010000000000101;
assign LUT_4[3655] = 32'b11111111111111110011001011111101;
assign LUT_4[3656] = 32'b11111111111111110110110001011010;
assign LUT_4[3657] = 32'b11111111111111101111111101010010;
assign LUT_4[3658] = 32'b11111111111111110110001011111110;
assign LUT_4[3659] = 32'b11111111111111101111010111110110;
assign LUT_4[3660] = 32'b11111111111111110011110001110110;
assign LUT_4[3661] = 32'b11111111111111101100111101101110;
assign LUT_4[3662] = 32'b11111111111111110011001100011010;
assign LUT_4[3663] = 32'b11111111111111101100011000010010;
assign LUT_4[3664] = 32'b11111111111111111011010110110011;
assign LUT_4[3665] = 32'b11111111111111110100100010101011;
assign LUT_4[3666] = 32'b11111111111111111010110001010111;
assign LUT_4[3667] = 32'b11111111111111110011111101001111;
assign LUT_4[3668] = 32'b11111111111111111000010111001111;
assign LUT_4[3669] = 32'b11111111111111110001100011000111;
assign LUT_4[3670] = 32'b11111111111111110111110001110011;
assign LUT_4[3671] = 32'b11111111111111110000111101101011;
assign LUT_4[3672] = 32'b11111111111111110100100011001000;
assign LUT_4[3673] = 32'b11111111111111101101101111000000;
assign LUT_4[3674] = 32'b11111111111111110011111101101100;
assign LUT_4[3675] = 32'b11111111111111101101001001100100;
assign LUT_4[3676] = 32'b11111111111111110001100011100100;
assign LUT_4[3677] = 32'b11111111111111101010101111011100;
assign LUT_4[3678] = 32'b11111111111111110000111110001000;
assign LUT_4[3679] = 32'b11111111111111101010001010000000;
assign LUT_4[3680] = 32'b11111111111111111100000000001100;
assign LUT_4[3681] = 32'b11111111111111110101001100000100;
assign LUT_4[3682] = 32'b11111111111111111011011010110000;
assign LUT_4[3683] = 32'b11111111111111110100100110101000;
assign LUT_4[3684] = 32'b11111111111111111001000000101000;
assign LUT_4[3685] = 32'b11111111111111110010001100100000;
assign LUT_4[3686] = 32'b11111111111111111000011011001100;
assign LUT_4[3687] = 32'b11111111111111110001100111000100;
assign LUT_4[3688] = 32'b11111111111111110101001100100001;
assign LUT_4[3689] = 32'b11111111111111101110011000011001;
assign LUT_4[3690] = 32'b11111111111111110100100111000101;
assign LUT_4[3691] = 32'b11111111111111101101110010111101;
assign LUT_4[3692] = 32'b11111111111111110010001100111101;
assign LUT_4[3693] = 32'b11111111111111101011011000110101;
assign LUT_4[3694] = 32'b11111111111111110001100111100001;
assign LUT_4[3695] = 32'b11111111111111101010110011011001;
assign LUT_4[3696] = 32'b11111111111111111001110001111010;
assign LUT_4[3697] = 32'b11111111111111110010111101110010;
assign LUT_4[3698] = 32'b11111111111111111001001100011110;
assign LUT_4[3699] = 32'b11111111111111110010011000010110;
assign LUT_4[3700] = 32'b11111111111111110110110010010110;
assign LUT_4[3701] = 32'b11111111111111101111111110001110;
assign LUT_4[3702] = 32'b11111111111111110110001100111010;
assign LUT_4[3703] = 32'b11111111111111101111011000110010;
assign LUT_4[3704] = 32'b11111111111111110010111110001111;
assign LUT_4[3705] = 32'b11111111111111101100001010000111;
assign LUT_4[3706] = 32'b11111111111111110010011000110011;
assign LUT_4[3707] = 32'b11111111111111101011100100101011;
assign LUT_4[3708] = 32'b11111111111111101111111110101011;
assign LUT_4[3709] = 32'b11111111111111101001001010100011;
assign LUT_4[3710] = 32'b11111111111111101111011001001111;
assign LUT_4[3711] = 32'b11111111111111101000100101000111;
assign LUT_4[3712] = 32'b11111111111111111110110011111001;
assign LUT_4[3713] = 32'b11111111111111110111111111110001;
assign LUT_4[3714] = 32'b11111111111111111110001110011101;
assign LUT_4[3715] = 32'b11111111111111110111011010010101;
assign LUT_4[3716] = 32'b11111111111111111011110100010101;
assign LUT_4[3717] = 32'b11111111111111110101000000001101;
assign LUT_4[3718] = 32'b11111111111111111011001110111001;
assign LUT_4[3719] = 32'b11111111111111110100011010110001;
assign LUT_4[3720] = 32'b11111111111111111000000000001110;
assign LUT_4[3721] = 32'b11111111111111110001001100000110;
assign LUT_4[3722] = 32'b11111111111111110111011010110010;
assign LUT_4[3723] = 32'b11111111111111110000100110101010;
assign LUT_4[3724] = 32'b11111111111111110101000000101010;
assign LUT_4[3725] = 32'b11111111111111101110001100100010;
assign LUT_4[3726] = 32'b11111111111111110100011011001110;
assign LUT_4[3727] = 32'b11111111111111101101100111000110;
assign LUT_4[3728] = 32'b11111111111111111100100101100111;
assign LUT_4[3729] = 32'b11111111111111110101110001011111;
assign LUT_4[3730] = 32'b11111111111111111100000000001011;
assign LUT_4[3731] = 32'b11111111111111110101001100000011;
assign LUT_4[3732] = 32'b11111111111111111001100110000011;
assign LUT_4[3733] = 32'b11111111111111110010110001111011;
assign LUT_4[3734] = 32'b11111111111111111001000000100111;
assign LUT_4[3735] = 32'b11111111111111110010001100011111;
assign LUT_4[3736] = 32'b11111111111111110101110001111100;
assign LUT_4[3737] = 32'b11111111111111101110111101110100;
assign LUT_4[3738] = 32'b11111111111111110101001100100000;
assign LUT_4[3739] = 32'b11111111111111101110011000011000;
assign LUT_4[3740] = 32'b11111111111111110010110010011000;
assign LUT_4[3741] = 32'b11111111111111101011111110010000;
assign LUT_4[3742] = 32'b11111111111111110010001100111100;
assign LUT_4[3743] = 32'b11111111111111101011011000110100;
assign LUT_4[3744] = 32'b11111111111111111101001111000000;
assign LUT_4[3745] = 32'b11111111111111110110011010111000;
assign LUT_4[3746] = 32'b11111111111111111100101001100100;
assign LUT_4[3747] = 32'b11111111111111110101110101011100;
assign LUT_4[3748] = 32'b11111111111111111010001111011100;
assign LUT_4[3749] = 32'b11111111111111110011011011010100;
assign LUT_4[3750] = 32'b11111111111111111001101010000000;
assign LUT_4[3751] = 32'b11111111111111110010110101111000;
assign LUT_4[3752] = 32'b11111111111111110110011011010101;
assign LUT_4[3753] = 32'b11111111111111101111100111001101;
assign LUT_4[3754] = 32'b11111111111111110101110101111001;
assign LUT_4[3755] = 32'b11111111111111101111000001110001;
assign LUT_4[3756] = 32'b11111111111111110011011011110001;
assign LUT_4[3757] = 32'b11111111111111101100100111101001;
assign LUT_4[3758] = 32'b11111111111111110010110110010101;
assign LUT_4[3759] = 32'b11111111111111101100000010001101;
assign LUT_4[3760] = 32'b11111111111111111011000000101110;
assign LUT_4[3761] = 32'b11111111111111110100001100100110;
assign LUT_4[3762] = 32'b11111111111111111010011011010010;
assign LUT_4[3763] = 32'b11111111111111110011100111001010;
assign LUT_4[3764] = 32'b11111111111111111000000001001010;
assign LUT_4[3765] = 32'b11111111111111110001001101000010;
assign LUT_4[3766] = 32'b11111111111111110111011011101110;
assign LUT_4[3767] = 32'b11111111111111110000100111100110;
assign LUT_4[3768] = 32'b11111111111111110100001101000011;
assign LUT_4[3769] = 32'b11111111111111101101011000111011;
assign LUT_4[3770] = 32'b11111111111111110011100111100111;
assign LUT_4[3771] = 32'b11111111111111101100110011011111;
assign LUT_4[3772] = 32'b11111111111111110001001101011111;
assign LUT_4[3773] = 32'b11111111111111101010011001010111;
assign LUT_4[3774] = 32'b11111111111111110000101000000011;
assign LUT_4[3775] = 32'b11111111111111101001110011111011;
assign LUT_4[3776] = 32'b00000000000000000000001011001101;
assign LUT_4[3777] = 32'b11111111111111111001010111000101;
assign LUT_4[3778] = 32'b11111111111111111111100101110001;
assign LUT_4[3779] = 32'b11111111111111111000110001101001;
assign LUT_4[3780] = 32'b11111111111111111101001011101001;
assign LUT_4[3781] = 32'b11111111111111110110010111100001;
assign LUT_4[3782] = 32'b11111111111111111100100110001101;
assign LUT_4[3783] = 32'b11111111111111110101110010000101;
assign LUT_4[3784] = 32'b11111111111111111001010111100010;
assign LUT_4[3785] = 32'b11111111111111110010100011011010;
assign LUT_4[3786] = 32'b11111111111111111000110010000110;
assign LUT_4[3787] = 32'b11111111111111110001111101111110;
assign LUT_4[3788] = 32'b11111111111111110110010111111110;
assign LUT_4[3789] = 32'b11111111111111101111100011110110;
assign LUT_4[3790] = 32'b11111111111111110101110010100010;
assign LUT_4[3791] = 32'b11111111111111101110111110011010;
assign LUT_4[3792] = 32'b11111111111111111101111100111011;
assign LUT_4[3793] = 32'b11111111111111110111001000110011;
assign LUT_4[3794] = 32'b11111111111111111101010111011111;
assign LUT_4[3795] = 32'b11111111111111110110100011010111;
assign LUT_4[3796] = 32'b11111111111111111010111101010111;
assign LUT_4[3797] = 32'b11111111111111110100001001001111;
assign LUT_4[3798] = 32'b11111111111111111010010111111011;
assign LUT_4[3799] = 32'b11111111111111110011100011110011;
assign LUT_4[3800] = 32'b11111111111111110111001001010000;
assign LUT_4[3801] = 32'b11111111111111110000010101001000;
assign LUT_4[3802] = 32'b11111111111111110110100011110100;
assign LUT_4[3803] = 32'b11111111111111101111101111101100;
assign LUT_4[3804] = 32'b11111111111111110100001001101100;
assign LUT_4[3805] = 32'b11111111111111101101010101100100;
assign LUT_4[3806] = 32'b11111111111111110011100100010000;
assign LUT_4[3807] = 32'b11111111111111101100110000001000;
assign LUT_4[3808] = 32'b11111111111111111110100110010100;
assign LUT_4[3809] = 32'b11111111111111110111110010001100;
assign LUT_4[3810] = 32'b11111111111111111110000000111000;
assign LUT_4[3811] = 32'b11111111111111110111001100110000;
assign LUT_4[3812] = 32'b11111111111111111011100110110000;
assign LUT_4[3813] = 32'b11111111111111110100110010101000;
assign LUT_4[3814] = 32'b11111111111111111011000001010100;
assign LUT_4[3815] = 32'b11111111111111110100001101001100;
assign LUT_4[3816] = 32'b11111111111111110111110010101001;
assign LUT_4[3817] = 32'b11111111111111110000111110100001;
assign LUT_4[3818] = 32'b11111111111111110111001101001101;
assign LUT_4[3819] = 32'b11111111111111110000011001000101;
assign LUT_4[3820] = 32'b11111111111111110100110011000101;
assign LUT_4[3821] = 32'b11111111111111101101111110111101;
assign LUT_4[3822] = 32'b11111111111111110100001101101001;
assign LUT_4[3823] = 32'b11111111111111101101011001100001;
assign LUT_4[3824] = 32'b11111111111111111100011000000010;
assign LUT_4[3825] = 32'b11111111111111110101100011111010;
assign LUT_4[3826] = 32'b11111111111111111011110010100110;
assign LUT_4[3827] = 32'b11111111111111110100111110011110;
assign LUT_4[3828] = 32'b11111111111111111001011000011110;
assign LUT_4[3829] = 32'b11111111111111110010100100010110;
assign LUT_4[3830] = 32'b11111111111111111000110011000010;
assign LUT_4[3831] = 32'b11111111111111110001111110111010;
assign LUT_4[3832] = 32'b11111111111111110101100100010111;
assign LUT_4[3833] = 32'b11111111111111101110110000001111;
assign LUT_4[3834] = 32'b11111111111111110100111110111011;
assign LUT_4[3835] = 32'b11111111111111101110001010110011;
assign LUT_4[3836] = 32'b11111111111111110010100100110011;
assign LUT_4[3837] = 32'b11111111111111101011110000101011;
assign LUT_4[3838] = 32'b11111111111111110001111111010111;
assign LUT_4[3839] = 32'b11111111111111101011001011001111;
assign LUT_4[3840] = 32'b00000000000000000001001001010100;
assign LUT_4[3841] = 32'b11111111111111111010010101001100;
assign LUT_4[3842] = 32'b00000000000000000000100011111000;
assign LUT_4[3843] = 32'b11111111111111111001101111110000;
assign LUT_4[3844] = 32'b11111111111111111110001001110000;
assign LUT_4[3845] = 32'b11111111111111110111010101101000;
assign LUT_4[3846] = 32'b11111111111111111101100100010100;
assign LUT_4[3847] = 32'b11111111111111110110110000001100;
assign LUT_4[3848] = 32'b11111111111111111010010101101001;
assign LUT_4[3849] = 32'b11111111111111110011100001100001;
assign LUT_4[3850] = 32'b11111111111111111001110000001101;
assign LUT_4[3851] = 32'b11111111111111110010111100000101;
assign LUT_4[3852] = 32'b11111111111111110111010110000101;
assign LUT_4[3853] = 32'b11111111111111110000100001111101;
assign LUT_4[3854] = 32'b11111111111111110110110000101001;
assign LUT_4[3855] = 32'b11111111111111101111111100100001;
assign LUT_4[3856] = 32'b11111111111111111110111011000010;
assign LUT_4[3857] = 32'b11111111111111111000000110111010;
assign LUT_4[3858] = 32'b11111111111111111110010101100110;
assign LUT_4[3859] = 32'b11111111111111110111100001011110;
assign LUT_4[3860] = 32'b11111111111111111011111011011110;
assign LUT_4[3861] = 32'b11111111111111110101000111010110;
assign LUT_4[3862] = 32'b11111111111111111011010110000010;
assign LUT_4[3863] = 32'b11111111111111110100100001111010;
assign LUT_4[3864] = 32'b11111111111111111000000111010111;
assign LUT_4[3865] = 32'b11111111111111110001010011001111;
assign LUT_4[3866] = 32'b11111111111111110111100001111011;
assign LUT_4[3867] = 32'b11111111111111110000101101110011;
assign LUT_4[3868] = 32'b11111111111111110101000111110011;
assign LUT_4[3869] = 32'b11111111111111101110010011101011;
assign LUT_4[3870] = 32'b11111111111111110100100010010111;
assign LUT_4[3871] = 32'b11111111111111101101101110001111;
assign LUT_4[3872] = 32'b11111111111111111111100100011011;
assign LUT_4[3873] = 32'b11111111111111111000110000010011;
assign LUT_4[3874] = 32'b11111111111111111110111110111111;
assign LUT_4[3875] = 32'b11111111111111111000001010110111;
assign LUT_4[3876] = 32'b11111111111111111100100100110111;
assign LUT_4[3877] = 32'b11111111111111110101110000101111;
assign LUT_4[3878] = 32'b11111111111111111011111111011011;
assign LUT_4[3879] = 32'b11111111111111110101001011010011;
assign LUT_4[3880] = 32'b11111111111111111000110000110000;
assign LUT_4[3881] = 32'b11111111111111110001111100101000;
assign LUT_4[3882] = 32'b11111111111111111000001011010100;
assign LUT_4[3883] = 32'b11111111111111110001010111001100;
assign LUT_4[3884] = 32'b11111111111111110101110001001100;
assign LUT_4[3885] = 32'b11111111111111101110111101000100;
assign LUT_4[3886] = 32'b11111111111111110101001011110000;
assign LUT_4[3887] = 32'b11111111111111101110010111101000;
assign LUT_4[3888] = 32'b11111111111111111101010110001001;
assign LUT_4[3889] = 32'b11111111111111110110100010000001;
assign LUT_4[3890] = 32'b11111111111111111100110000101101;
assign LUT_4[3891] = 32'b11111111111111110101111100100101;
assign LUT_4[3892] = 32'b11111111111111111010010110100101;
assign LUT_4[3893] = 32'b11111111111111110011100010011101;
assign LUT_4[3894] = 32'b11111111111111111001110001001001;
assign LUT_4[3895] = 32'b11111111111111110010111101000001;
assign LUT_4[3896] = 32'b11111111111111110110100010011110;
assign LUT_4[3897] = 32'b11111111111111101111101110010110;
assign LUT_4[3898] = 32'b11111111111111110101111101000010;
assign LUT_4[3899] = 32'b11111111111111101111001000111010;
assign LUT_4[3900] = 32'b11111111111111110011100010111010;
assign LUT_4[3901] = 32'b11111111111111101100101110110010;
assign LUT_4[3902] = 32'b11111111111111110010111101011110;
assign LUT_4[3903] = 32'b11111111111111101100001001010110;
assign LUT_4[3904] = 32'b00000000000000000010100000101000;
assign LUT_4[3905] = 32'b11111111111111111011101100100000;
assign LUT_4[3906] = 32'b00000000000000000001111011001100;
assign LUT_4[3907] = 32'b11111111111111111011000111000100;
assign LUT_4[3908] = 32'b11111111111111111111100001000100;
assign LUT_4[3909] = 32'b11111111111111111000101100111100;
assign LUT_4[3910] = 32'b11111111111111111110111011101000;
assign LUT_4[3911] = 32'b11111111111111111000000111100000;
assign LUT_4[3912] = 32'b11111111111111111011101100111101;
assign LUT_4[3913] = 32'b11111111111111110100111000110101;
assign LUT_4[3914] = 32'b11111111111111111011000111100001;
assign LUT_4[3915] = 32'b11111111111111110100010011011001;
assign LUT_4[3916] = 32'b11111111111111111000101101011001;
assign LUT_4[3917] = 32'b11111111111111110001111001010001;
assign LUT_4[3918] = 32'b11111111111111111000000111111101;
assign LUT_4[3919] = 32'b11111111111111110001010011110101;
assign LUT_4[3920] = 32'b00000000000000000000010010010110;
assign LUT_4[3921] = 32'b11111111111111111001011110001110;
assign LUT_4[3922] = 32'b11111111111111111111101100111010;
assign LUT_4[3923] = 32'b11111111111111111000111000110010;
assign LUT_4[3924] = 32'b11111111111111111101010010110010;
assign LUT_4[3925] = 32'b11111111111111110110011110101010;
assign LUT_4[3926] = 32'b11111111111111111100101101010110;
assign LUT_4[3927] = 32'b11111111111111110101111001001110;
assign LUT_4[3928] = 32'b11111111111111111001011110101011;
assign LUT_4[3929] = 32'b11111111111111110010101010100011;
assign LUT_4[3930] = 32'b11111111111111111000111001001111;
assign LUT_4[3931] = 32'b11111111111111110010000101000111;
assign LUT_4[3932] = 32'b11111111111111110110011111000111;
assign LUT_4[3933] = 32'b11111111111111101111101010111111;
assign LUT_4[3934] = 32'b11111111111111110101111001101011;
assign LUT_4[3935] = 32'b11111111111111101111000101100011;
assign LUT_4[3936] = 32'b00000000000000000000111011101111;
assign LUT_4[3937] = 32'b11111111111111111010000111100111;
assign LUT_4[3938] = 32'b00000000000000000000010110010011;
assign LUT_4[3939] = 32'b11111111111111111001100010001011;
assign LUT_4[3940] = 32'b11111111111111111101111100001011;
assign LUT_4[3941] = 32'b11111111111111110111001000000011;
assign LUT_4[3942] = 32'b11111111111111111101010110101111;
assign LUT_4[3943] = 32'b11111111111111110110100010100111;
assign LUT_4[3944] = 32'b11111111111111111010001000000100;
assign LUT_4[3945] = 32'b11111111111111110011010011111100;
assign LUT_4[3946] = 32'b11111111111111111001100010101000;
assign LUT_4[3947] = 32'b11111111111111110010101110100000;
assign LUT_4[3948] = 32'b11111111111111110111001000100000;
assign LUT_4[3949] = 32'b11111111111111110000010100011000;
assign LUT_4[3950] = 32'b11111111111111110110100011000100;
assign LUT_4[3951] = 32'b11111111111111101111101110111100;
assign LUT_4[3952] = 32'b11111111111111111110101101011101;
assign LUT_4[3953] = 32'b11111111111111110111111001010101;
assign LUT_4[3954] = 32'b11111111111111111110001000000001;
assign LUT_4[3955] = 32'b11111111111111110111010011111001;
assign LUT_4[3956] = 32'b11111111111111111011101101111001;
assign LUT_4[3957] = 32'b11111111111111110100111001110001;
assign LUT_4[3958] = 32'b11111111111111111011001000011101;
assign LUT_4[3959] = 32'b11111111111111110100010100010101;
assign LUT_4[3960] = 32'b11111111111111110111111001110010;
assign LUT_4[3961] = 32'b11111111111111110001000101101010;
assign LUT_4[3962] = 32'b11111111111111110111010100010110;
assign LUT_4[3963] = 32'b11111111111111110000100000001110;
assign LUT_4[3964] = 32'b11111111111111110100111010001110;
assign LUT_4[3965] = 32'b11111111111111101110000110000110;
assign LUT_4[3966] = 32'b11111111111111110100010100110010;
assign LUT_4[3967] = 32'b11111111111111101101100000101010;
assign LUT_4[3968] = 32'b00000000000000000011101111011100;
assign LUT_4[3969] = 32'b11111111111111111100111011010100;
assign LUT_4[3970] = 32'b00000000000000000011001010000000;
assign LUT_4[3971] = 32'b11111111111111111100010101111000;
assign LUT_4[3972] = 32'b00000000000000000000101111111000;
assign LUT_4[3973] = 32'b11111111111111111001111011110000;
assign LUT_4[3974] = 32'b00000000000000000000001010011100;
assign LUT_4[3975] = 32'b11111111111111111001010110010100;
assign LUT_4[3976] = 32'b11111111111111111100111011110001;
assign LUT_4[3977] = 32'b11111111111111110110000111101001;
assign LUT_4[3978] = 32'b11111111111111111100010110010101;
assign LUT_4[3979] = 32'b11111111111111110101100010001101;
assign LUT_4[3980] = 32'b11111111111111111001111100001101;
assign LUT_4[3981] = 32'b11111111111111110011001000000101;
assign LUT_4[3982] = 32'b11111111111111111001010110110001;
assign LUT_4[3983] = 32'b11111111111111110010100010101001;
assign LUT_4[3984] = 32'b00000000000000000001100001001010;
assign LUT_4[3985] = 32'b11111111111111111010101101000010;
assign LUT_4[3986] = 32'b00000000000000000000111011101110;
assign LUT_4[3987] = 32'b11111111111111111010000111100110;
assign LUT_4[3988] = 32'b11111111111111111110100001100110;
assign LUT_4[3989] = 32'b11111111111111110111101101011110;
assign LUT_4[3990] = 32'b11111111111111111101111100001010;
assign LUT_4[3991] = 32'b11111111111111110111001000000010;
assign LUT_4[3992] = 32'b11111111111111111010101101011111;
assign LUT_4[3993] = 32'b11111111111111110011111001010111;
assign LUT_4[3994] = 32'b11111111111111111010001000000011;
assign LUT_4[3995] = 32'b11111111111111110011010011111011;
assign LUT_4[3996] = 32'b11111111111111110111101101111011;
assign LUT_4[3997] = 32'b11111111111111110000111001110011;
assign LUT_4[3998] = 32'b11111111111111110111001000011111;
assign LUT_4[3999] = 32'b11111111111111110000010100010111;
assign LUT_4[4000] = 32'b00000000000000000010001010100011;
assign LUT_4[4001] = 32'b11111111111111111011010110011011;
assign LUT_4[4002] = 32'b00000000000000000001100101000111;
assign LUT_4[4003] = 32'b11111111111111111010110000111111;
assign LUT_4[4004] = 32'b11111111111111111111001010111111;
assign LUT_4[4005] = 32'b11111111111111111000010110110111;
assign LUT_4[4006] = 32'b11111111111111111110100101100011;
assign LUT_4[4007] = 32'b11111111111111110111110001011011;
assign LUT_4[4008] = 32'b11111111111111111011010110111000;
assign LUT_4[4009] = 32'b11111111111111110100100010110000;
assign LUT_4[4010] = 32'b11111111111111111010110001011100;
assign LUT_4[4011] = 32'b11111111111111110011111101010100;
assign LUT_4[4012] = 32'b11111111111111111000010111010100;
assign LUT_4[4013] = 32'b11111111111111110001100011001100;
assign LUT_4[4014] = 32'b11111111111111110111110001111000;
assign LUT_4[4015] = 32'b11111111111111110000111101110000;
assign LUT_4[4016] = 32'b11111111111111111111111100010001;
assign LUT_4[4017] = 32'b11111111111111111001001000001001;
assign LUT_4[4018] = 32'b11111111111111111111010110110101;
assign LUT_4[4019] = 32'b11111111111111111000100010101101;
assign LUT_4[4020] = 32'b11111111111111111100111100101101;
assign LUT_4[4021] = 32'b11111111111111110110001000100101;
assign LUT_4[4022] = 32'b11111111111111111100010111010001;
assign LUT_4[4023] = 32'b11111111111111110101100011001001;
assign LUT_4[4024] = 32'b11111111111111111001001000100110;
assign LUT_4[4025] = 32'b11111111111111110010010100011110;
assign LUT_4[4026] = 32'b11111111111111111000100011001010;
assign LUT_4[4027] = 32'b11111111111111110001101111000010;
assign LUT_4[4028] = 32'b11111111111111110110001001000010;
assign LUT_4[4029] = 32'b11111111111111101111010100111010;
assign LUT_4[4030] = 32'b11111111111111110101100011100110;
assign LUT_4[4031] = 32'b11111111111111101110101111011110;
assign LUT_4[4032] = 32'b00000000000000000101000110110000;
assign LUT_4[4033] = 32'b11111111111111111110010010101000;
assign LUT_4[4034] = 32'b00000000000000000100100001010100;
assign LUT_4[4035] = 32'b11111111111111111101101101001100;
assign LUT_4[4036] = 32'b00000000000000000010000111001100;
assign LUT_4[4037] = 32'b11111111111111111011010011000100;
assign LUT_4[4038] = 32'b00000000000000000001100001110000;
assign LUT_4[4039] = 32'b11111111111111111010101101101000;
assign LUT_4[4040] = 32'b11111111111111111110010011000101;
assign LUT_4[4041] = 32'b11111111111111110111011110111101;
assign LUT_4[4042] = 32'b11111111111111111101101101101001;
assign LUT_4[4043] = 32'b11111111111111110110111001100001;
assign LUT_4[4044] = 32'b11111111111111111011010011100001;
assign LUT_4[4045] = 32'b11111111111111110100011111011001;
assign LUT_4[4046] = 32'b11111111111111111010101110000101;
assign LUT_4[4047] = 32'b11111111111111110011111001111101;
assign LUT_4[4048] = 32'b00000000000000000010111000011110;
assign LUT_4[4049] = 32'b11111111111111111100000100010110;
assign LUT_4[4050] = 32'b00000000000000000010010011000010;
assign LUT_4[4051] = 32'b11111111111111111011011110111010;
assign LUT_4[4052] = 32'b11111111111111111111111000111010;
assign LUT_4[4053] = 32'b11111111111111111001000100110010;
assign LUT_4[4054] = 32'b11111111111111111111010011011110;
assign LUT_4[4055] = 32'b11111111111111111000011111010110;
assign LUT_4[4056] = 32'b11111111111111111100000100110011;
assign LUT_4[4057] = 32'b11111111111111110101010000101011;
assign LUT_4[4058] = 32'b11111111111111111011011111010111;
assign LUT_4[4059] = 32'b11111111111111110100101011001111;
assign LUT_4[4060] = 32'b11111111111111111001000101001111;
assign LUT_4[4061] = 32'b11111111111111110010010001000111;
assign LUT_4[4062] = 32'b11111111111111111000011111110011;
assign LUT_4[4063] = 32'b11111111111111110001101011101011;
assign LUT_4[4064] = 32'b00000000000000000011100001110111;
assign LUT_4[4065] = 32'b11111111111111111100101101101111;
assign LUT_4[4066] = 32'b00000000000000000010111100011011;
assign LUT_4[4067] = 32'b11111111111111111100001000010011;
assign LUT_4[4068] = 32'b00000000000000000000100010010011;
assign LUT_4[4069] = 32'b11111111111111111001101110001011;
assign LUT_4[4070] = 32'b11111111111111111111111100110111;
assign LUT_4[4071] = 32'b11111111111111111001001000101111;
assign LUT_4[4072] = 32'b11111111111111111100101110001100;
assign LUT_4[4073] = 32'b11111111111111110101111010000100;
assign LUT_4[4074] = 32'b11111111111111111100001000110000;
assign LUT_4[4075] = 32'b11111111111111110101010100101000;
assign LUT_4[4076] = 32'b11111111111111111001101110101000;
assign LUT_4[4077] = 32'b11111111111111110010111010100000;
assign LUT_4[4078] = 32'b11111111111111111001001001001100;
assign LUT_4[4079] = 32'b11111111111111110010010101000100;
assign LUT_4[4080] = 32'b00000000000000000001010011100101;
assign LUT_4[4081] = 32'b11111111111111111010011111011101;
assign LUT_4[4082] = 32'b00000000000000000000101110001001;
assign LUT_4[4083] = 32'b11111111111111111001111010000001;
assign LUT_4[4084] = 32'b11111111111111111110010100000001;
assign LUT_4[4085] = 32'b11111111111111110111011111111001;
assign LUT_4[4086] = 32'b11111111111111111101101110100101;
assign LUT_4[4087] = 32'b11111111111111110110111010011101;
assign LUT_4[4088] = 32'b11111111111111111010011111111010;
assign LUT_4[4089] = 32'b11111111111111110011101011110010;
assign LUT_4[4090] = 32'b11111111111111111001111010011110;
assign LUT_4[4091] = 32'b11111111111111110011000110010110;
assign LUT_4[4092] = 32'b11111111111111110111100000010110;
assign LUT_4[4093] = 32'b11111111111111110000101100001110;
assign LUT_4[4094] = 32'b11111111111111110110111010111010;
assign LUT_4[4095] = 32'b11111111111111110000000110110010;
assign LUT_4[4096] = 32'b11111111111111111100001111110001;
assign LUT_4[4097] = 32'b11111111111111110101011011101001;
assign LUT_4[4098] = 32'b11111111111111111011101010010101;
assign LUT_4[4099] = 32'b11111111111111110100110110001101;
assign LUT_4[4100] = 32'b11111111111111111001010000001101;
assign LUT_4[4101] = 32'b11111111111111110010011100000101;
assign LUT_4[4102] = 32'b11111111111111111000101010110001;
assign LUT_4[4103] = 32'b11111111111111110001110110101001;
assign LUT_4[4104] = 32'b11111111111111110101011100000110;
assign LUT_4[4105] = 32'b11111111111111101110100111111110;
assign LUT_4[4106] = 32'b11111111111111110100110110101010;
assign LUT_4[4107] = 32'b11111111111111101110000010100010;
assign LUT_4[4108] = 32'b11111111111111110010011100100010;
assign LUT_4[4109] = 32'b11111111111111101011101000011010;
assign LUT_4[4110] = 32'b11111111111111110001110111000110;
assign LUT_4[4111] = 32'b11111111111111101011000010111110;
assign LUT_4[4112] = 32'b11111111111111111010000001011111;
assign LUT_4[4113] = 32'b11111111111111110011001101010111;
assign LUT_4[4114] = 32'b11111111111111111001011100000011;
assign LUT_4[4115] = 32'b11111111111111110010100111111011;
assign LUT_4[4116] = 32'b11111111111111110111000001111011;
assign LUT_4[4117] = 32'b11111111111111110000001101110011;
assign LUT_4[4118] = 32'b11111111111111110110011100011111;
assign LUT_4[4119] = 32'b11111111111111101111101000010111;
assign LUT_4[4120] = 32'b11111111111111110011001101110100;
assign LUT_4[4121] = 32'b11111111111111101100011001101100;
assign LUT_4[4122] = 32'b11111111111111110010101000011000;
assign LUT_4[4123] = 32'b11111111111111101011110100010000;
assign LUT_4[4124] = 32'b11111111111111110000001110010000;
assign LUT_4[4125] = 32'b11111111111111101001011010001000;
assign LUT_4[4126] = 32'b11111111111111101111101000110100;
assign LUT_4[4127] = 32'b11111111111111101000110100101100;
assign LUT_4[4128] = 32'b11111111111111111010101010111000;
assign LUT_4[4129] = 32'b11111111111111110011110110110000;
assign LUT_4[4130] = 32'b11111111111111111010000101011100;
assign LUT_4[4131] = 32'b11111111111111110011010001010100;
assign LUT_4[4132] = 32'b11111111111111110111101011010100;
assign LUT_4[4133] = 32'b11111111111111110000110111001100;
assign LUT_4[4134] = 32'b11111111111111110111000101111000;
assign LUT_4[4135] = 32'b11111111111111110000010001110000;
assign LUT_4[4136] = 32'b11111111111111110011110111001101;
assign LUT_4[4137] = 32'b11111111111111101101000011000101;
assign LUT_4[4138] = 32'b11111111111111110011010001110001;
assign LUT_4[4139] = 32'b11111111111111101100011101101001;
assign LUT_4[4140] = 32'b11111111111111110000110111101001;
assign LUT_4[4141] = 32'b11111111111111101010000011100001;
assign LUT_4[4142] = 32'b11111111111111110000010010001101;
assign LUT_4[4143] = 32'b11111111111111101001011110000101;
assign LUT_4[4144] = 32'b11111111111111111000011100100110;
assign LUT_4[4145] = 32'b11111111111111110001101000011110;
assign LUT_4[4146] = 32'b11111111111111110111110111001010;
assign LUT_4[4147] = 32'b11111111111111110001000011000010;
assign LUT_4[4148] = 32'b11111111111111110101011101000010;
assign LUT_4[4149] = 32'b11111111111111101110101000111010;
assign LUT_4[4150] = 32'b11111111111111110100110111100110;
assign LUT_4[4151] = 32'b11111111111111101110000011011110;
assign LUT_4[4152] = 32'b11111111111111110001101000111011;
assign LUT_4[4153] = 32'b11111111111111101010110100110011;
assign LUT_4[4154] = 32'b11111111111111110001000011011111;
assign LUT_4[4155] = 32'b11111111111111101010001111010111;
assign LUT_4[4156] = 32'b11111111111111101110101001010111;
assign LUT_4[4157] = 32'b11111111111111100111110101001111;
assign LUT_4[4158] = 32'b11111111111111101110000011111011;
assign LUT_4[4159] = 32'b11111111111111100111001111110011;
assign LUT_4[4160] = 32'b11111111111111111101100111000101;
assign LUT_4[4161] = 32'b11111111111111110110110010111101;
assign LUT_4[4162] = 32'b11111111111111111101000001101001;
assign LUT_4[4163] = 32'b11111111111111110110001101100001;
assign LUT_4[4164] = 32'b11111111111111111010100111100001;
assign LUT_4[4165] = 32'b11111111111111110011110011011001;
assign LUT_4[4166] = 32'b11111111111111111010000010000101;
assign LUT_4[4167] = 32'b11111111111111110011001101111101;
assign LUT_4[4168] = 32'b11111111111111110110110011011010;
assign LUT_4[4169] = 32'b11111111111111101111111111010010;
assign LUT_4[4170] = 32'b11111111111111110110001101111110;
assign LUT_4[4171] = 32'b11111111111111101111011001110110;
assign LUT_4[4172] = 32'b11111111111111110011110011110110;
assign LUT_4[4173] = 32'b11111111111111101100111111101110;
assign LUT_4[4174] = 32'b11111111111111110011001110011010;
assign LUT_4[4175] = 32'b11111111111111101100011010010010;
assign LUT_4[4176] = 32'b11111111111111111011011000110011;
assign LUT_4[4177] = 32'b11111111111111110100100100101011;
assign LUT_4[4178] = 32'b11111111111111111010110011010111;
assign LUT_4[4179] = 32'b11111111111111110011111111001111;
assign LUT_4[4180] = 32'b11111111111111111000011001001111;
assign LUT_4[4181] = 32'b11111111111111110001100101000111;
assign LUT_4[4182] = 32'b11111111111111110111110011110011;
assign LUT_4[4183] = 32'b11111111111111110000111111101011;
assign LUT_4[4184] = 32'b11111111111111110100100101001000;
assign LUT_4[4185] = 32'b11111111111111101101110001000000;
assign LUT_4[4186] = 32'b11111111111111110011111111101100;
assign LUT_4[4187] = 32'b11111111111111101101001011100100;
assign LUT_4[4188] = 32'b11111111111111110001100101100100;
assign LUT_4[4189] = 32'b11111111111111101010110001011100;
assign LUT_4[4190] = 32'b11111111111111110001000000001000;
assign LUT_4[4191] = 32'b11111111111111101010001100000000;
assign LUT_4[4192] = 32'b11111111111111111100000010001100;
assign LUT_4[4193] = 32'b11111111111111110101001110000100;
assign LUT_4[4194] = 32'b11111111111111111011011100110000;
assign LUT_4[4195] = 32'b11111111111111110100101000101000;
assign LUT_4[4196] = 32'b11111111111111111001000010101000;
assign LUT_4[4197] = 32'b11111111111111110010001110100000;
assign LUT_4[4198] = 32'b11111111111111111000011101001100;
assign LUT_4[4199] = 32'b11111111111111110001101001000100;
assign LUT_4[4200] = 32'b11111111111111110101001110100001;
assign LUT_4[4201] = 32'b11111111111111101110011010011001;
assign LUT_4[4202] = 32'b11111111111111110100101001000101;
assign LUT_4[4203] = 32'b11111111111111101101110100111101;
assign LUT_4[4204] = 32'b11111111111111110010001110111101;
assign LUT_4[4205] = 32'b11111111111111101011011010110101;
assign LUT_4[4206] = 32'b11111111111111110001101001100001;
assign LUT_4[4207] = 32'b11111111111111101010110101011001;
assign LUT_4[4208] = 32'b11111111111111111001110011111010;
assign LUT_4[4209] = 32'b11111111111111110010111111110010;
assign LUT_4[4210] = 32'b11111111111111111001001110011110;
assign LUT_4[4211] = 32'b11111111111111110010011010010110;
assign LUT_4[4212] = 32'b11111111111111110110110100010110;
assign LUT_4[4213] = 32'b11111111111111110000000000001110;
assign LUT_4[4214] = 32'b11111111111111110110001110111010;
assign LUT_4[4215] = 32'b11111111111111101111011010110010;
assign LUT_4[4216] = 32'b11111111111111110011000000001111;
assign LUT_4[4217] = 32'b11111111111111101100001100000111;
assign LUT_4[4218] = 32'b11111111111111110010011010110011;
assign LUT_4[4219] = 32'b11111111111111101011100110101011;
assign LUT_4[4220] = 32'b11111111111111110000000000101011;
assign LUT_4[4221] = 32'b11111111111111101001001100100011;
assign LUT_4[4222] = 32'b11111111111111101111011011001111;
assign LUT_4[4223] = 32'b11111111111111101000100111000111;
assign LUT_4[4224] = 32'b11111111111111111110110101111001;
assign LUT_4[4225] = 32'b11111111111111111000000001110001;
assign LUT_4[4226] = 32'b11111111111111111110010000011101;
assign LUT_4[4227] = 32'b11111111111111110111011100010101;
assign LUT_4[4228] = 32'b11111111111111111011110110010101;
assign LUT_4[4229] = 32'b11111111111111110101000010001101;
assign LUT_4[4230] = 32'b11111111111111111011010000111001;
assign LUT_4[4231] = 32'b11111111111111110100011100110001;
assign LUT_4[4232] = 32'b11111111111111111000000010001110;
assign LUT_4[4233] = 32'b11111111111111110001001110000110;
assign LUT_4[4234] = 32'b11111111111111110111011100110010;
assign LUT_4[4235] = 32'b11111111111111110000101000101010;
assign LUT_4[4236] = 32'b11111111111111110101000010101010;
assign LUT_4[4237] = 32'b11111111111111101110001110100010;
assign LUT_4[4238] = 32'b11111111111111110100011101001110;
assign LUT_4[4239] = 32'b11111111111111101101101001000110;
assign LUT_4[4240] = 32'b11111111111111111100100111100111;
assign LUT_4[4241] = 32'b11111111111111110101110011011111;
assign LUT_4[4242] = 32'b11111111111111111100000010001011;
assign LUT_4[4243] = 32'b11111111111111110101001110000011;
assign LUT_4[4244] = 32'b11111111111111111001101000000011;
assign LUT_4[4245] = 32'b11111111111111110010110011111011;
assign LUT_4[4246] = 32'b11111111111111111001000010100111;
assign LUT_4[4247] = 32'b11111111111111110010001110011111;
assign LUT_4[4248] = 32'b11111111111111110101110011111100;
assign LUT_4[4249] = 32'b11111111111111101110111111110100;
assign LUT_4[4250] = 32'b11111111111111110101001110100000;
assign LUT_4[4251] = 32'b11111111111111101110011010011000;
assign LUT_4[4252] = 32'b11111111111111110010110100011000;
assign LUT_4[4253] = 32'b11111111111111101100000000010000;
assign LUT_4[4254] = 32'b11111111111111110010001110111100;
assign LUT_4[4255] = 32'b11111111111111101011011010110100;
assign LUT_4[4256] = 32'b11111111111111111101010001000000;
assign LUT_4[4257] = 32'b11111111111111110110011100111000;
assign LUT_4[4258] = 32'b11111111111111111100101011100100;
assign LUT_4[4259] = 32'b11111111111111110101110111011100;
assign LUT_4[4260] = 32'b11111111111111111010010001011100;
assign LUT_4[4261] = 32'b11111111111111110011011101010100;
assign LUT_4[4262] = 32'b11111111111111111001101100000000;
assign LUT_4[4263] = 32'b11111111111111110010110111111000;
assign LUT_4[4264] = 32'b11111111111111110110011101010101;
assign LUT_4[4265] = 32'b11111111111111101111101001001101;
assign LUT_4[4266] = 32'b11111111111111110101110111111001;
assign LUT_4[4267] = 32'b11111111111111101111000011110001;
assign LUT_4[4268] = 32'b11111111111111110011011101110001;
assign LUT_4[4269] = 32'b11111111111111101100101001101001;
assign LUT_4[4270] = 32'b11111111111111110010111000010101;
assign LUT_4[4271] = 32'b11111111111111101100000100001101;
assign LUT_4[4272] = 32'b11111111111111111011000010101110;
assign LUT_4[4273] = 32'b11111111111111110100001110100110;
assign LUT_4[4274] = 32'b11111111111111111010011101010010;
assign LUT_4[4275] = 32'b11111111111111110011101001001010;
assign LUT_4[4276] = 32'b11111111111111111000000011001010;
assign LUT_4[4277] = 32'b11111111111111110001001111000010;
assign LUT_4[4278] = 32'b11111111111111110111011101101110;
assign LUT_4[4279] = 32'b11111111111111110000101001100110;
assign LUT_4[4280] = 32'b11111111111111110100001111000011;
assign LUT_4[4281] = 32'b11111111111111101101011010111011;
assign LUT_4[4282] = 32'b11111111111111110011101001100111;
assign LUT_4[4283] = 32'b11111111111111101100110101011111;
assign LUT_4[4284] = 32'b11111111111111110001001111011111;
assign LUT_4[4285] = 32'b11111111111111101010011011010111;
assign LUT_4[4286] = 32'b11111111111111110000101010000011;
assign LUT_4[4287] = 32'b11111111111111101001110101111011;
assign LUT_4[4288] = 32'b00000000000000000000001101001101;
assign LUT_4[4289] = 32'b11111111111111111001011001000101;
assign LUT_4[4290] = 32'b11111111111111111111100111110001;
assign LUT_4[4291] = 32'b11111111111111111000110011101001;
assign LUT_4[4292] = 32'b11111111111111111101001101101001;
assign LUT_4[4293] = 32'b11111111111111110110011001100001;
assign LUT_4[4294] = 32'b11111111111111111100101000001101;
assign LUT_4[4295] = 32'b11111111111111110101110100000101;
assign LUT_4[4296] = 32'b11111111111111111001011001100010;
assign LUT_4[4297] = 32'b11111111111111110010100101011010;
assign LUT_4[4298] = 32'b11111111111111111000110100000110;
assign LUT_4[4299] = 32'b11111111111111110001111111111110;
assign LUT_4[4300] = 32'b11111111111111110110011001111110;
assign LUT_4[4301] = 32'b11111111111111101111100101110110;
assign LUT_4[4302] = 32'b11111111111111110101110100100010;
assign LUT_4[4303] = 32'b11111111111111101111000000011010;
assign LUT_4[4304] = 32'b11111111111111111101111110111011;
assign LUT_4[4305] = 32'b11111111111111110111001010110011;
assign LUT_4[4306] = 32'b11111111111111111101011001011111;
assign LUT_4[4307] = 32'b11111111111111110110100101010111;
assign LUT_4[4308] = 32'b11111111111111111010111111010111;
assign LUT_4[4309] = 32'b11111111111111110100001011001111;
assign LUT_4[4310] = 32'b11111111111111111010011001111011;
assign LUT_4[4311] = 32'b11111111111111110011100101110011;
assign LUT_4[4312] = 32'b11111111111111110111001011010000;
assign LUT_4[4313] = 32'b11111111111111110000010111001000;
assign LUT_4[4314] = 32'b11111111111111110110100101110100;
assign LUT_4[4315] = 32'b11111111111111101111110001101100;
assign LUT_4[4316] = 32'b11111111111111110100001011101100;
assign LUT_4[4317] = 32'b11111111111111101101010111100100;
assign LUT_4[4318] = 32'b11111111111111110011100110010000;
assign LUT_4[4319] = 32'b11111111111111101100110010001000;
assign LUT_4[4320] = 32'b11111111111111111110101000010100;
assign LUT_4[4321] = 32'b11111111111111110111110100001100;
assign LUT_4[4322] = 32'b11111111111111111110000010111000;
assign LUT_4[4323] = 32'b11111111111111110111001110110000;
assign LUT_4[4324] = 32'b11111111111111111011101000110000;
assign LUT_4[4325] = 32'b11111111111111110100110100101000;
assign LUT_4[4326] = 32'b11111111111111111011000011010100;
assign LUT_4[4327] = 32'b11111111111111110100001111001100;
assign LUT_4[4328] = 32'b11111111111111110111110100101001;
assign LUT_4[4329] = 32'b11111111111111110001000000100001;
assign LUT_4[4330] = 32'b11111111111111110111001111001101;
assign LUT_4[4331] = 32'b11111111111111110000011011000101;
assign LUT_4[4332] = 32'b11111111111111110100110101000101;
assign LUT_4[4333] = 32'b11111111111111101110000000111101;
assign LUT_4[4334] = 32'b11111111111111110100001111101001;
assign LUT_4[4335] = 32'b11111111111111101101011011100001;
assign LUT_4[4336] = 32'b11111111111111111100011010000010;
assign LUT_4[4337] = 32'b11111111111111110101100101111010;
assign LUT_4[4338] = 32'b11111111111111111011110100100110;
assign LUT_4[4339] = 32'b11111111111111110101000000011110;
assign LUT_4[4340] = 32'b11111111111111111001011010011110;
assign LUT_4[4341] = 32'b11111111111111110010100110010110;
assign LUT_4[4342] = 32'b11111111111111111000110101000010;
assign LUT_4[4343] = 32'b11111111111111110010000000111010;
assign LUT_4[4344] = 32'b11111111111111110101100110010111;
assign LUT_4[4345] = 32'b11111111111111101110110010001111;
assign LUT_4[4346] = 32'b11111111111111110101000000111011;
assign LUT_4[4347] = 32'b11111111111111101110001100110011;
assign LUT_4[4348] = 32'b11111111111111110010100110110011;
assign LUT_4[4349] = 32'b11111111111111101011110010101011;
assign LUT_4[4350] = 32'b11111111111111110010000001010111;
assign LUT_4[4351] = 32'b11111111111111101011001101001111;
assign LUT_4[4352] = 32'b00000000000000000001001011010100;
assign LUT_4[4353] = 32'b11111111111111111010010111001100;
assign LUT_4[4354] = 32'b00000000000000000000100101111000;
assign LUT_4[4355] = 32'b11111111111111111001110001110000;
assign LUT_4[4356] = 32'b11111111111111111110001011110000;
assign LUT_4[4357] = 32'b11111111111111110111010111101000;
assign LUT_4[4358] = 32'b11111111111111111101100110010100;
assign LUT_4[4359] = 32'b11111111111111110110110010001100;
assign LUT_4[4360] = 32'b11111111111111111010010111101001;
assign LUT_4[4361] = 32'b11111111111111110011100011100001;
assign LUT_4[4362] = 32'b11111111111111111001110010001101;
assign LUT_4[4363] = 32'b11111111111111110010111110000101;
assign LUT_4[4364] = 32'b11111111111111110111011000000101;
assign LUT_4[4365] = 32'b11111111111111110000100011111101;
assign LUT_4[4366] = 32'b11111111111111110110110010101001;
assign LUT_4[4367] = 32'b11111111111111101111111110100001;
assign LUT_4[4368] = 32'b11111111111111111110111101000010;
assign LUT_4[4369] = 32'b11111111111111111000001000111010;
assign LUT_4[4370] = 32'b11111111111111111110010111100110;
assign LUT_4[4371] = 32'b11111111111111110111100011011110;
assign LUT_4[4372] = 32'b11111111111111111011111101011110;
assign LUT_4[4373] = 32'b11111111111111110101001001010110;
assign LUT_4[4374] = 32'b11111111111111111011011000000010;
assign LUT_4[4375] = 32'b11111111111111110100100011111010;
assign LUT_4[4376] = 32'b11111111111111111000001001010111;
assign LUT_4[4377] = 32'b11111111111111110001010101001111;
assign LUT_4[4378] = 32'b11111111111111110111100011111011;
assign LUT_4[4379] = 32'b11111111111111110000101111110011;
assign LUT_4[4380] = 32'b11111111111111110101001001110011;
assign LUT_4[4381] = 32'b11111111111111101110010101101011;
assign LUT_4[4382] = 32'b11111111111111110100100100010111;
assign LUT_4[4383] = 32'b11111111111111101101110000001111;
assign LUT_4[4384] = 32'b11111111111111111111100110011011;
assign LUT_4[4385] = 32'b11111111111111111000110010010011;
assign LUT_4[4386] = 32'b11111111111111111111000000111111;
assign LUT_4[4387] = 32'b11111111111111111000001100110111;
assign LUT_4[4388] = 32'b11111111111111111100100110110111;
assign LUT_4[4389] = 32'b11111111111111110101110010101111;
assign LUT_4[4390] = 32'b11111111111111111100000001011011;
assign LUT_4[4391] = 32'b11111111111111110101001101010011;
assign LUT_4[4392] = 32'b11111111111111111000110010110000;
assign LUT_4[4393] = 32'b11111111111111110001111110101000;
assign LUT_4[4394] = 32'b11111111111111111000001101010100;
assign LUT_4[4395] = 32'b11111111111111110001011001001100;
assign LUT_4[4396] = 32'b11111111111111110101110011001100;
assign LUT_4[4397] = 32'b11111111111111101110111111000100;
assign LUT_4[4398] = 32'b11111111111111110101001101110000;
assign LUT_4[4399] = 32'b11111111111111101110011001101000;
assign LUT_4[4400] = 32'b11111111111111111101011000001001;
assign LUT_4[4401] = 32'b11111111111111110110100100000001;
assign LUT_4[4402] = 32'b11111111111111111100110010101101;
assign LUT_4[4403] = 32'b11111111111111110101111110100101;
assign LUT_4[4404] = 32'b11111111111111111010011000100101;
assign LUT_4[4405] = 32'b11111111111111110011100100011101;
assign LUT_4[4406] = 32'b11111111111111111001110011001001;
assign LUT_4[4407] = 32'b11111111111111110010111111000001;
assign LUT_4[4408] = 32'b11111111111111110110100100011110;
assign LUT_4[4409] = 32'b11111111111111101111110000010110;
assign LUT_4[4410] = 32'b11111111111111110101111111000010;
assign LUT_4[4411] = 32'b11111111111111101111001010111010;
assign LUT_4[4412] = 32'b11111111111111110011100100111010;
assign LUT_4[4413] = 32'b11111111111111101100110000110010;
assign LUT_4[4414] = 32'b11111111111111110010111111011110;
assign LUT_4[4415] = 32'b11111111111111101100001011010110;
assign LUT_4[4416] = 32'b00000000000000000010100010101000;
assign LUT_4[4417] = 32'b11111111111111111011101110100000;
assign LUT_4[4418] = 32'b00000000000000000001111101001100;
assign LUT_4[4419] = 32'b11111111111111111011001001000100;
assign LUT_4[4420] = 32'b11111111111111111111100011000100;
assign LUT_4[4421] = 32'b11111111111111111000101110111100;
assign LUT_4[4422] = 32'b11111111111111111110111101101000;
assign LUT_4[4423] = 32'b11111111111111111000001001100000;
assign LUT_4[4424] = 32'b11111111111111111011101110111101;
assign LUT_4[4425] = 32'b11111111111111110100111010110101;
assign LUT_4[4426] = 32'b11111111111111111011001001100001;
assign LUT_4[4427] = 32'b11111111111111110100010101011001;
assign LUT_4[4428] = 32'b11111111111111111000101111011001;
assign LUT_4[4429] = 32'b11111111111111110001111011010001;
assign LUT_4[4430] = 32'b11111111111111111000001001111101;
assign LUT_4[4431] = 32'b11111111111111110001010101110101;
assign LUT_4[4432] = 32'b00000000000000000000010100010110;
assign LUT_4[4433] = 32'b11111111111111111001100000001110;
assign LUT_4[4434] = 32'b11111111111111111111101110111010;
assign LUT_4[4435] = 32'b11111111111111111000111010110010;
assign LUT_4[4436] = 32'b11111111111111111101010100110010;
assign LUT_4[4437] = 32'b11111111111111110110100000101010;
assign LUT_4[4438] = 32'b11111111111111111100101111010110;
assign LUT_4[4439] = 32'b11111111111111110101111011001110;
assign LUT_4[4440] = 32'b11111111111111111001100000101011;
assign LUT_4[4441] = 32'b11111111111111110010101100100011;
assign LUT_4[4442] = 32'b11111111111111111000111011001111;
assign LUT_4[4443] = 32'b11111111111111110010000111000111;
assign LUT_4[4444] = 32'b11111111111111110110100001000111;
assign LUT_4[4445] = 32'b11111111111111101111101100111111;
assign LUT_4[4446] = 32'b11111111111111110101111011101011;
assign LUT_4[4447] = 32'b11111111111111101111000111100011;
assign LUT_4[4448] = 32'b00000000000000000000111101101111;
assign LUT_4[4449] = 32'b11111111111111111010001001100111;
assign LUT_4[4450] = 32'b00000000000000000000011000010011;
assign LUT_4[4451] = 32'b11111111111111111001100100001011;
assign LUT_4[4452] = 32'b11111111111111111101111110001011;
assign LUT_4[4453] = 32'b11111111111111110111001010000011;
assign LUT_4[4454] = 32'b11111111111111111101011000101111;
assign LUT_4[4455] = 32'b11111111111111110110100100100111;
assign LUT_4[4456] = 32'b11111111111111111010001010000100;
assign LUT_4[4457] = 32'b11111111111111110011010101111100;
assign LUT_4[4458] = 32'b11111111111111111001100100101000;
assign LUT_4[4459] = 32'b11111111111111110010110000100000;
assign LUT_4[4460] = 32'b11111111111111110111001010100000;
assign LUT_4[4461] = 32'b11111111111111110000010110011000;
assign LUT_4[4462] = 32'b11111111111111110110100101000100;
assign LUT_4[4463] = 32'b11111111111111101111110000111100;
assign LUT_4[4464] = 32'b11111111111111111110101111011101;
assign LUT_4[4465] = 32'b11111111111111110111111011010101;
assign LUT_4[4466] = 32'b11111111111111111110001010000001;
assign LUT_4[4467] = 32'b11111111111111110111010101111001;
assign LUT_4[4468] = 32'b11111111111111111011101111111001;
assign LUT_4[4469] = 32'b11111111111111110100111011110001;
assign LUT_4[4470] = 32'b11111111111111111011001010011101;
assign LUT_4[4471] = 32'b11111111111111110100010110010101;
assign LUT_4[4472] = 32'b11111111111111110111111011110010;
assign LUT_4[4473] = 32'b11111111111111110001000111101010;
assign LUT_4[4474] = 32'b11111111111111110111010110010110;
assign LUT_4[4475] = 32'b11111111111111110000100010001110;
assign LUT_4[4476] = 32'b11111111111111110100111100001110;
assign LUT_4[4477] = 32'b11111111111111101110001000000110;
assign LUT_4[4478] = 32'b11111111111111110100010110110010;
assign LUT_4[4479] = 32'b11111111111111101101100010101010;
assign LUT_4[4480] = 32'b00000000000000000011110001011100;
assign LUT_4[4481] = 32'b11111111111111111100111101010100;
assign LUT_4[4482] = 32'b00000000000000000011001100000000;
assign LUT_4[4483] = 32'b11111111111111111100010111111000;
assign LUT_4[4484] = 32'b00000000000000000000110001111000;
assign LUT_4[4485] = 32'b11111111111111111001111101110000;
assign LUT_4[4486] = 32'b00000000000000000000001100011100;
assign LUT_4[4487] = 32'b11111111111111111001011000010100;
assign LUT_4[4488] = 32'b11111111111111111100111101110001;
assign LUT_4[4489] = 32'b11111111111111110110001001101001;
assign LUT_4[4490] = 32'b11111111111111111100011000010101;
assign LUT_4[4491] = 32'b11111111111111110101100100001101;
assign LUT_4[4492] = 32'b11111111111111111001111110001101;
assign LUT_4[4493] = 32'b11111111111111110011001010000101;
assign LUT_4[4494] = 32'b11111111111111111001011000110001;
assign LUT_4[4495] = 32'b11111111111111110010100100101001;
assign LUT_4[4496] = 32'b00000000000000000001100011001010;
assign LUT_4[4497] = 32'b11111111111111111010101111000010;
assign LUT_4[4498] = 32'b00000000000000000000111101101110;
assign LUT_4[4499] = 32'b11111111111111111010001001100110;
assign LUT_4[4500] = 32'b11111111111111111110100011100110;
assign LUT_4[4501] = 32'b11111111111111110111101111011110;
assign LUT_4[4502] = 32'b11111111111111111101111110001010;
assign LUT_4[4503] = 32'b11111111111111110111001010000010;
assign LUT_4[4504] = 32'b11111111111111111010101111011111;
assign LUT_4[4505] = 32'b11111111111111110011111011010111;
assign LUT_4[4506] = 32'b11111111111111111010001010000011;
assign LUT_4[4507] = 32'b11111111111111110011010101111011;
assign LUT_4[4508] = 32'b11111111111111110111101111111011;
assign LUT_4[4509] = 32'b11111111111111110000111011110011;
assign LUT_4[4510] = 32'b11111111111111110111001010011111;
assign LUT_4[4511] = 32'b11111111111111110000010110010111;
assign LUT_4[4512] = 32'b00000000000000000010001100100011;
assign LUT_4[4513] = 32'b11111111111111111011011000011011;
assign LUT_4[4514] = 32'b00000000000000000001100111000111;
assign LUT_4[4515] = 32'b11111111111111111010110010111111;
assign LUT_4[4516] = 32'b11111111111111111111001100111111;
assign LUT_4[4517] = 32'b11111111111111111000011000110111;
assign LUT_4[4518] = 32'b11111111111111111110100111100011;
assign LUT_4[4519] = 32'b11111111111111110111110011011011;
assign LUT_4[4520] = 32'b11111111111111111011011000111000;
assign LUT_4[4521] = 32'b11111111111111110100100100110000;
assign LUT_4[4522] = 32'b11111111111111111010110011011100;
assign LUT_4[4523] = 32'b11111111111111110011111111010100;
assign LUT_4[4524] = 32'b11111111111111111000011001010100;
assign LUT_4[4525] = 32'b11111111111111110001100101001100;
assign LUT_4[4526] = 32'b11111111111111110111110011111000;
assign LUT_4[4527] = 32'b11111111111111110000111111110000;
assign LUT_4[4528] = 32'b11111111111111111111111110010001;
assign LUT_4[4529] = 32'b11111111111111111001001010001001;
assign LUT_4[4530] = 32'b11111111111111111111011000110101;
assign LUT_4[4531] = 32'b11111111111111111000100100101101;
assign LUT_4[4532] = 32'b11111111111111111100111110101101;
assign LUT_4[4533] = 32'b11111111111111110110001010100101;
assign LUT_4[4534] = 32'b11111111111111111100011001010001;
assign LUT_4[4535] = 32'b11111111111111110101100101001001;
assign LUT_4[4536] = 32'b11111111111111111001001010100110;
assign LUT_4[4537] = 32'b11111111111111110010010110011110;
assign LUT_4[4538] = 32'b11111111111111111000100101001010;
assign LUT_4[4539] = 32'b11111111111111110001110001000010;
assign LUT_4[4540] = 32'b11111111111111110110001011000010;
assign LUT_4[4541] = 32'b11111111111111101111010110111010;
assign LUT_4[4542] = 32'b11111111111111110101100101100110;
assign LUT_4[4543] = 32'b11111111111111101110110001011110;
assign LUT_4[4544] = 32'b00000000000000000101001000110000;
assign LUT_4[4545] = 32'b11111111111111111110010100101000;
assign LUT_4[4546] = 32'b00000000000000000100100011010100;
assign LUT_4[4547] = 32'b11111111111111111101101111001100;
assign LUT_4[4548] = 32'b00000000000000000010001001001100;
assign LUT_4[4549] = 32'b11111111111111111011010101000100;
assign LUT_4[4550] = 32'b00000000000000000001100011110000;
assign LUT_4[4551] = 32'b11111111111111111010101111101000;
assign LUT_4[4552] = 32'b11111111111111111110010101000101;
assign LUT_4[4553] = 32'b11111111111111110111100000111101;
assign LUT_4[4554] = 32'b11111111111111111101101111101001;
assign LUT_4[4555] = 32'b11111111111111110110111011100001;
assign LUT_4[4556] = 32'b11111111111111111011010101100001;
assign LUT_4[4557] = 32'b11111111111111110100100001011001;
assign LUT_4[4558] = 32'b11111111111111111010110000000101;
assign LUT_4[4559] = 32'b11111111111111110011111011111101;
assign LUT_4[4560] = 32'b00000000000000000010111010011110;
assign LUT_4[4561] = 32'b11111111111111111100000110010110;
assign LUT_4[4562] = 32'b00000000000000000010010101000010;
assign LUT_4[4563] = 32'b11111111111111111011100000111010;
assign LUT_4[4564] = 32'b11111111111111111111111010111010;
assign LUT_4[4565] = 32'b11111111111111111001000110110010;
assign LUT_4[4566] = 32'b11111111111111111111010101011110;
assign LUT_4[4567] = 32'b11111111111111111000100001010110;
assign LUT_4[4568] = 32'b11111111111111111100000110110011;
assign LUT_4[4569] = 32'b11111111111111110101010010101011;
assign LUT_4[4570] = 32'b11111111111111111011100001010111;
assign LUT_4[4571] = 32'b11111111111111110100101101001111;
assign LUT_4[4572] = 32'b11111111111111111001000111001111;
assign LUT_4[4573] = 32'b11111111111111110010010011000111;
assign LUT_4[4574] = 32'b11111111111111111000100001110011;
assign LUT_4[4575] = 32'b11111111111111110001101101101011;
assign LUT_4[4576] = 32'b00000000000000000011100011110111;
assign LUT_4[4577] = 32'b11111111111111111100101111101111;
assign LUT_4[4578] = 32'b00000000000000000010111110011011;
assign LUT_4[4579] = 32'b11111111111111111100001010010011;
assign LUT_4[4580] = 32'b00000000000000000000100100010011;
assign LUT_4[4581] = 32'b11111111111111111001110000001011;
assign LUT_4[4582] = 32'b11111111111111111111111110110111;
assign LUT_4[4583] = 32'b11111111111111111001001010101111;
assign LUT_4[4584] = 32'b11111111111111111100110000001100;
assign LUT_4[4585] = 32'b11111111111111110101111100000100;
assign LUT_4[4586] = 32'b11111111111111111100001010110000;
assign LUT_4[4587] = 32'b11111111111111110101010110101000;
assign LUT_4[4588] = 32'b11111111111111111001110000101000;
assign LUT_4[4589] = 32'b11111111111111110010111100100000;
assign LUT_4[4590] = 32'b11111111111111111001001011001100;
assign LUT_4[4591] = 32'b11111111111111110010010111000100;
assign LUT_4[4592] = 32'b00000000000000000001010101100101;
assign LUT_4[4593] = 32'b11111111111111111010100001011101;
assign LUT_4[4594] = 32'b00000000000000000000110000001001;
assign LUT_4[4595] = 32'b11111111111111111001111100000001;
assign LUT_4[4596] = 32'b11111111111111111110010110000001;
assign LUT_4[4597] = 32'b11111111111111110111100001111001;
assign LUT_4[4598] = 32'b11111111111111111101110000100101;
assign LUT_4[4599] = 32'b11111111111111110110111100011101;
assign LUT_4[4600] = 32'b11111111111111111010100001111010;
assign LUT_4[4601] = 32'b11111111111111110011101101110010;
assign LUT_4[4602] = 32'b11111111111111111001111100011110;
assign LUT_4[4603] = 32'b11111111111111110011001000010110;
assign LUT_4[4604] = 32'b11111111111111110111100010010110;
assign LUT_4[4605] = 32'b11111111111111110000101110001110;
assign LUT_4[4606] = 32'b11111111111111110110111100111010;
assign LUT_4[4607] = 32'b11111111111111110000001000110010;
assign LUT_4[4608] = 32'b11111111111111111011010011111001;
assign LUT_4[4609] = 32'b11111111111111110100011111110001;
assign LUT_4[4610] = 32'b11111111111111111010101110011101;
assign LUT_4[4611] = 32'b11111111111111110011111010010101;
assign LUT_4[4612] = 32'b11111111111111111000010100010101;
assign LUT_4[4613] = 32'b11111111111111110001100000001101;
assign LUT_4[4614] = 32'b11111111111111110111101110111001;
assign LUT_4[4615] = 32'b11111111111111110000111010110001;
assign LUT_4[4616] = 32'b11111111111111110100100000001110;
assign LUT_4[4617] = 32'b11111111111111101101101100000110;
assign LUT_4[4618] = 32'b11111111111111110011111010110010;
assign LUT_4[4619] = 32'b11111111111111101101000110101010;
assign LUT_4[4620] = 32'b11111111111111110001100000101010;
assign LUT_4[4621] = 32'b11111111111111101010101100100010;
assign LUT_4[4622] = 32'b11111111111111110000111011001110;
assign LUT_4[4623] = 32'b11111111111111101010000111000110;
assign LUT_4[4624] = 32'b11111111111111111001000101100111;
assign LUT_4[4625] = 32'b11111111111111110010010001011111;
assign LUT_4[4626] = 32'b11111111111111111000100000001011;
assign LUT_4[4627] = 32'b11111111111111110001101100000011;
assign LUT_4[4628] = 32'b11111111111111110110000110000011;
assign LUT_4[4629] = 32'b11111111111111101111010001111011;
assign LUT_4[4630] = 32'b11111111111111110101100000100111;
assign LUT_4[4631] = 32'b11111111111111101110101100011111;
assign LUT_4[4632] = 32'b11111111111111110010010001111100;
assign LUT_4[4633] = 32'b11111111111111101011011101110100;
assign LUT_4[4634] = 32'b11111111111111110001101100100000;
assign LUT_4[4635] = 32'b11111111111111101010111000011000;
assign LUT_4[4636] = 32'b11111111111111101111010010011000;
assign LUT_4[4637] = 32'b11111111111111101000011110010000;
assign LUT_4[4638] = 32'b11111111111111101110101100111100;
assign LUT_4[4639] = 32'b11111111111111100111111000110100;
assign LUT_4[4640] = 32'b11111111111111111001101111000000;
assign LUT_4[4641] = 32'b11111111111111110010111010111000;
assign LUT_4[4642] = 32'b11111111111111111001001001100100;
assign LUT_4[4643] = 32'b11111111111111110010010101011100;
assign LUT_4[4644] = 32'b11111111111111110110101111011100;
assign LUT_4[4645] = 32'b11111111111111101111111011010100;
assign LUT_4[4646] = 32'b11111111111111110110001010000000;
assign LUT_4[4647] = 32'b11111111111111101111010101111000;
assign LUT_4[4648] = 32'b11111111111111110010111011010101;
assign LUT_4[4649] = 32'b11111111111111101100000111001101;
assign LUT_4[4650] = 32'b11111111111111110010010101111001;
assign LUT_4[4651] = 32'b11111111111111101011100001110001;
assign LUT_4[4652] = 32'b11111111111111101111111011110001;
assign LUT_4[4653] = 32'b11111111111111101001000111101001;
assign LUT_4[4654] = 32'b11111111111111101111010110010101;
assign LUT_4[4655] = 32'b11111111111111101000100010001101;
assign LUT_4[4656] = 32'b11111111111111110111100000101110;
assign LUT_4[4657] = 32'b11111111111111110000101100100110;
assign LUT_4[4658] = 32'b11111111111111110110111011010010;
assign LUT_4[4659] = 32'b11111111111111110000000111001010;
assign LUT_4[4660] = 32'b11111111111111110100100001001010;
assign LUT_4[4661] = 32'b11111111111111101101101101000010;
assign LUT_4[4662] = 32'b11111111111111110011111011101110;
assign LUT_4[4663] = 32'b11111111111111101101000111100110;
assign LUT_4[4664] = 32'b11111111111111110000101101000011;
assign LUT_4[4665] = 32'b11111111111111101001111000111011;
assign LUT_4[4666] = 32'b11111111111111110000000111100111;
assign LUT_4[4667] = 32'b11111111111111101001010011011111;
assign LUT_4[4668] = 32'b11111111111111101101101101011111;
assign LUT_4[4669] = 32'b11111111111111100110111001010111;
assign LUT_4[4670] = 32'b11111111111111101101001000000011;
assign LUT_4[4671] = 32'b11111111111111100110010011111011;
assign LUT_4[4672] = 32'b11111111111111111100101011001101;
assign LUT_4[4673] = 32'b11111111111111110101110111000101;
assign LUT_4[4674] = 32'b11111111111111111100000101110001;
assign LUT_4[4675] = 32'b11111111111111110101010001101001;
assign LUT_4[4676] = 32'b11111111111111111001101011101001;
assign LUT_4[4677] = 32'b11111111111111110010110111100001;
assign LUT_4[4678] = 32'b11111111111111111001000110001101;
assign LUT_4[4679] = 32'b11111111111111110010010010000101;
assign LUT_4[4680] = 32'b11111111111111110101110111100010;
assign LUT_4[4681] = 32'b11111111111111101111000011011010;
assign LUT_4[4682] = 32'b11111111111111110101010010000110;
assign LUT_4[4683] = 32'b11111111111111101110011101111110;
assign LUT_4[4684] = 32'b11111111111111110010110111111110;
assign LUT_4[4685] = 32'b11111111111111101100000011110110;
assign LUT_4[4686] = 32'b11111111111111110010010010100010;
assign LUT_4[4687] = 32'b11111111111111101011011110011010;
assign LUT_4[4688] = 32'b11111111111111111010011100111011;
assign LUT_4[4689] = 32'b11111111111111110011101000110011;
assign LUT_4[4690] = 32'b11111111111111111001110111011111;
assign LUT_4[4691] = 32'b11111111111111110011000011010111;
assign LUT_4[4692] = 32'b11111111111111110111011101010111;
assign LUT_4[4693] = 32'b11111111111111110000101001001111;
assign LUT_4[4694] = 32'b11111111111111110110110111111011;
assign LUT_4[4695] = 32'b11111111111111110000000011110011;
assign LUT_4[4696] = 32'b11111111111111110011101001010000;
assign LUT_4[4697] = 32'b11111111111111101100110101001000;
assign LUT_4[4698] = 32'b11111111111111110011000011110100;
assign LUT_4[4699] = 32'b11111111111111101100001111101100;
assign LUT_4[4700] = 32'b11111111111111110000101001101100;
assign LUT_4[4701] = 32'b11111111111111101001110101100100;
assign LUT_4[4702] = 32'b11111111111111110000000100010000;
assign LUT_4[4703] = 32'b11111111111111101001010000001000;
assign LUT_4[4704] = 32'b11111111111111111011000110010100;
assign LUT_4[4705] = 32'b11111111111111110100010010001100;
assign LUT_4[4706] = 32'b11111111111111111010100000111000;
assign LUT_4[4707] = 32'b11111111111111110011101100110000;
assign LUT_4[4708] = 32'b11111111111111111000000110110000;
assign LUT_4[4709] = 32'b11111111111111110001010010101000;
assign LUT_4[4710] = 32'b11111111111111110111100001010100;
assign LUT_4[4711] = 32'b11111111111111110000101101001100;
assign LUT_4[4712] = 32'b11111111111111110100010010101001;
assign LUT_4[4713] = 32'b11111111111111101101011110100001;
assign LUT_4[4714] = 32'b11111111111111110011101101001101;
assign LUT_4[4715] = 32'b11111111111111101100111001000101;
assign LUT_4[4716] = 32'b11111111111111110001010011000101;
assign LUT_4[4717] = 32'b11111111111111101010011110111101;
assign LUT_4[4718] = 32'b11111111111111110000101101101001;
assign LUT_4[4719] = 32'b11111111111111101001111001100001;
assign LUT_4[4720] = 32'b11111111111111111000111000000010;
assign LUT_4[4721] = 32'b11111111111111110010000011111010;
assign LUT_4[4722] = 32'b11111111111111111000010010100110;
assign LUT_4[4723] = 32'b11111111111111110001011110011110;
assign LUT_4[4724] = 32'b11111111111111110101111000011110;
assign LUT_4[4725] = 32'b11111111111111101111000100010110;
assign LUT_4[4726] = 32'b11111111111111110101010011000010;
assign LUT_4[4727] = 32'b11111111111111101110011110111010;
assign LUT_4[4728] = 32'b11111111111111110010000100010111;
assign LUT_4[4729] = 32'b11111111111111101011010000001111;
assign LUT_4[4730] = 32'b11111111111111110001011110111011;
assign LUT_4[4731] = 32'b11111111111111101010101010110011;
assign LUT_4[4732] = 32'b11111111111111101111000100110011;
assign LUT_4[4733] = 32'b11111111111111101000010000101011;
assign LUT_4[4734] = 32'b11111111111111101110011111010111;
assign LUT_4[4735] = 32'b11111111111111100111101011001111;
assign LUT_4[4736] = 32'b11111111111111111101111010000001;
assign LUT_4[4737] = 32'b11111111111111110111000101111001;
assign LUT_4[4738] = 32'b11111111111111111101010100100101;
assign LUT_4[4739] = 32'b11111111111111110110100000011101;
assign LUT_4[4740] = 32'b11111111111111111010111010011101;
assign LUT_4[4741] = 32'b11111111111111110100000110010101;
assign LUT_4[4742] = 32'b11111111111111111010010101000001;
assign LUT_4[4743] = 32'b11111111111111110011100000111001;
assign LUT_4[4744] = 32'b11111111111111110111000110010110;
assign LUT_4[4745] = 32'b11111111111111110000010010001110;
assign LUT_4[4746] = 32'b11111111111111110110100000111010;
assign LUT_4[4747] = 32'b11111111111111101111101100110010;
assign LUT_4[4748] = 32'b11111111111111110100000110110010;
assign LUT_4[4749] = 32'b11111111111111101101010010101010;
assign LUT_4[4750] = 32'b11111111111111110011100001010110;
assign LUT_4[4751] = 32'b11111111111111101100101101001110;
assign LUT_4[4752] = 32'b11111111111111111011101011101111;
assign LUT_4[4753] = 32'b11111111111111110100110111100111;
assign LUT_4[4754] = 32'b11111111111111111011000110010011;
assign LUT_4[4755] = 32'b11111111111111110100010010001011;
assign LUT_4[4756] = 32'b11111111111111111000101100001011;
assign LUT_4[4757] = 32'b11111111111111110001111000000011;
assign LUT_4[4758] = 32'b11111111111111111000000110101111;
assign LUT_4[4759] = 32'b11111111111111110001010010100111;
assign LUT_4[4760] = 32'b11111111111111110100111000000100;
assign LUT_4[4761] = 32'b11111111111111101110000011111100;
assign LUT_4[4762] = 32'b11111111111111110100010010101000;
assign LUT_4[4763] = 32'b11111111111111101101011110100000;
assign LUT_4[4764] = 32'b11111111111111110001111000100000;
assign LUT_4[4765] = 32'b11111111111111101011000100011000;
assign LUT_4[4766] = 32'b11111111111111110001010011000100;
assign LUT_4[4767] = 32'b11111111111111101010011110111100;
assign LUT_4[4768] = 32'b11111111111111111100010101001000;
assign LUT_4[4769] = 32'b11111111111111110101100001000000;
assign LUT_4[4770] = 32'b11111111111111111011101111101100;
assign LUT_4[4771] = 32'b11111111111111110100111011100100;
assign LUT_4[4772] = 32'b11111111111111111001010101100100;
assign LUT_4[4773] = 32'b11111111111111110010100001011100;
assign LUT_4[4774] = 32'b11111111111111111000110000001000;
assign LUT_4[4775] = 32'b11111111111111110001111100000000;
assign LUT_4[4776] = 32'b11111111111111110101100001011101;
assign LUT_4[4777] = 32'b11111111111111101110101101010101;
assign LUT_4[4778] = 32'b11111111111111110100111100000001;
assign LUT_4[4779] = 32'b11111111111111101110000111111001;
assign LUT_4[4780] = 32'b11111111111111110010100001111001;
assign LUT_4[4781] = 32'b11111111111111101011101101110001;
assign LUT_4[4782] = 32'b11111111111111110001111100011101;
assign LUT_4[4783] = 32'b11111111111111101011001000010101;
assign LUT_4[4784] = 32'b11111111111111111010000110110110;
assign LUT_4[4785] = 32'b11111111111111110011010010101110;
assign LUT_4[4786] = 32'b11111111111111111001100001011010;
assign LUT_4[4787] = 32'b11111111111111110010101101010010;
assign LUT_4[4788] = 32'b11111111111111110111000111010010;
assign LUT_4[4789] = 32'b11111111111111110000010011001010;
assign LUT_4[4790] = 32'b11111111111111110110100001110110;
assign LUT_4[4791] = 32'b11111111111111101111101101101110;
assign LUT_4[4792] = 32'b11111111111111110011010011001011;
assign LUT_4[4793] = 32'b11111111111111101100011111000011;
assign LUT_4[4794] = 32'b11111111111111110010101101101111;
assign LUT_4[4795] = 32'b11111111111111101011111001100111;
assign LUT_4[4796] = 32'b11111111111111110000010011100111;
assign LUT_4[4797] = 32'b11111111111111101001011111011111;
assign LUT_4[4798] = 32'b11111111111111101111101110001011;
assign LUT_4[4799] = 32'b11111111111111101000111010000011;
assign LUT_4[4800] = 32'b11111111111111111111010001010101;
assign LUT_4[4801] = 32'b11111111111111111000011101001101;
assign LUT_4[4802] = 32'b11111111111111111110101011111001;
assign LUT_4[4803] = 32'b11111111111111110111110111110001;
assign LUT_4[4804] = 32'b11111111111111111100010001110001;
assign LUT_4[4805] = 32'b11111111111111110101011101101001;
assign LUT_4[4806] = 32'b11111111111111111011101100010101;
assign LUT_4[4807] = 32'b11111111111111110100111000001101;
assign LUT_4[4808] = 32'b11111111111111111000011101101010;
assign LUT_4[4809] = 32'b11111111111111110001101001100010;
assign LUT_4[4810] = 32'b11111111111111110111111000001110;
assign LUT_4[4811] = 32'b11111111111111110001000100000110;
assign LUT_4[4812] = 32'b11111111111111110101011110000110;
assign LUT_4[4813] = 32'b11111111111111101110101001111110;
assign LUT_4[4814] = 32'b11111111111111110100111000101010;
assign LUT_4[4815] = 32'b11111111111111101110000100100010;
assign LUT_4[4816] = 32'b11111111111111111101000011000011;
assign LUT_4[4817] = 32'b11111111111111110110001110111011;
assign LUT_4[4818] = 32'b11111111111111111100011101100111;
assign LUT_4[4819] = 32'b11111111111111110101101001011111;
assign LUT_4[4820] = 32'b11111111111111111010000011011111;
assign LUT_4[4821] = 32'b11111111111111110011001111010111;
assign LUT_4[4822] = 32'b11111111111111111001011110000011;
assign LUT_4[4823] = 32'b11111111111111110010101001111011;
assign LUT_4[4824] = 32'b11111111111111110110001111011000;
assign LUT_4[4825] = 32'b11111111111111101111011011010000;
assign LUT_4[4826] = 32'b11111111111111110101101001111100;
assign LUT_4[4827] = 32'b11111111111111101110110101110100;
assign LUT_4[4828] = 32'b11111111111111110011001111110100;
assign LUT_4[4829] = 32'b11111111111111101100011011101100;
assign LUT_4[4830] = 32'b11111111111111110010101010011000;
assign LUT_4[4831] = 32'b11111111111111101011110110010000;
assign LUT_4[4832] = 32'b11111111111111111101101100011100;
assign LUT_4[4833] = 32'b11111111111111110110111000010100;
assign LUT_4[4834] = 32'b11111111111111111101000111000000;
assign LUT_4[4835] = 32'b11111111111111110110010010111000;
assign LUT_4[4836] = 32'b11111111111111111010101100111000;
assign LUT_4[4837] = 32'b11111111111111110011111000110000;
assign LUT_4[4838] = 32'b11111111111111111010000111011100;
assign LUT_4[4839] = 32'b11111111111111110011010011010100;
assign LUT_4[4840] = 32'b11111111111111110110111000110001;
assign LUT_4[4841] = 32'b11111111111111110000000100101001;
assign LUT_4[4842] = 32'b11111111111111110110010011010101;
assign LUT_4[4843] = 32'b11111111111111101111011111001101;
assign LUT_4[4844] = 32'b11111111111111110011111001001101;
assign LUT_4[4845] = 32'b11111111111111101101000101000101;
assign LUT_4[4846] = 32'b11111111111111110011010011110001;
assign LUT_4[4847] = 32'b11111111111111101100011111101001;
assign LUT_4[4848] = 32'b11111111111111111011011110001010;
assign LUT_4[4849] = 32'b11111111111111110100101010000010;
assign LUT_4[4850] = 32'b11111111111111111010111000101110;
assign LUT_4[4851] = 32'b11111111111111110100000100100110;
assign LUT_4[4852] = 32'b11111111111111111000011110100110;
assign LUT_4[4853] = 32'b11111111111111110001101010011110;
assign LUT_4[4854] = 32'b11111111111111110111111001001010;
assign LUT_4[4855] = 32'b11111111111111110001000101000010;
assign LUT_4[4856] = 32'b11111111111111110100101010011111;
assign LUT_4[4857] = 32'b11111111111111101101110110010111;
assign LUT_4[4858] = 32'b11111111111111110100000101000011;
assign LUT_4[4859] = 32'b11111111111111101101010000111011;
assign LUT_4[4860] = 32'b11111111111111110001101010111011;
assign LUT_4[4861] = 32'b11111111111111101010110110110011;
assign LUT_4[4862] = 32'b11111111111111110001000101011111;
assign LUT_4[4863] = 32'b11111111111111101010010001010111;
assign LUT_4[4864] = 32'b00000000000000000000001111011100;
assign LUT_4[4865] = 32'b11111111111111111001011011010100;
assign LUT_4[4866] = 32'b11111111111111111111101010000000;
assign LUT_4[4867] = 32'b11111111111111111000110101111000;
assign LUT_4[4868] = 32'b11111111111111111101001111111000;
assign LUT_4[4869] = 32'b11111111111111110110011011110000;
assign LUT_4[4870] = 32'b11111111111111111100101010011100;
assign LUT_4[4871] = 32'b11111111111111110101110110010100;
assign LUT_4[4872] = 32'b11111111111111111001011011110001;
assign LUT_4[4873] = 32'b11111111111111110010100111101001;
assign LUT_4[4874] = 32'b11111111111111111000110110010101;
assign LUT_4[4875] = 32'b11111111111111110010000010001101;
assign LUT_4[4876] = 32'b11111111111111110110011100001101;
assign LUT_4[4877] = 32'b11111111111111101111101000000101;
assign LUT_4[4878] = 32'b11111111111111110101110110110001;
assign LUT_4[4879] = 32'b11111111111111101111000010101001;
assign LUT_4[4880] = 32'b11111111111111111110000001001010;
assign LUT_4[4881] = 32'b11111111111111110111001101000010;
assign LUT_4[4882] = 32'b11111111111111111101011011101110;
assign LUT_4[4883] = 32'b11111111111111110110100111100110;
assign LUT_4[4884] = 32'b11111111111111111011000001100110;
assign LUT_4[4885] = 32'b11111111111111110100001101011110;
assign LUT_4[4886] = 32'b11111111111111111010011100001010;
assign LUT_4[4887] = 32'b11111111111111110011101000000010;
assign LUT_4[4888] = 32'b11111111111111110111001101011111;
assign LUT_4[4889] = 32'b11111111111111110000011001010111;
assign LUT_4[4890] = 32'b11111111111111110110101000000011;
assign LUT_4[4891] = 32'b11111111111111101111110011111011;
assign LUT_4[4892] = 32'b11111111111111110100001101111011;
assign LUT_4[4893] = 32'b11111111111111101101011001110011;
assign LUT_4[4894] = 32'b11111111111111110011101000011111;
assign LUT_4[4895] = 32'b11111111111111101100110100010111;
assign LUT_4[4896] = 32'b11111111111111111110101010100011;
assign LUT_4[4897] = 32'b11111111111111110111110110011011;
assign LUT_4[4898] = 32'b11111111111111111110000101000111;
assign LUT_4[4899] = 32'b11111111111111110111010000111111;
assign LUT_4[4900] = 32'b11111111111111111011101010111111;
assign LUT_4[4901] = 32'b11111111111111110100110110110111;
assign LUT_4[4902] = 32'b11111111111111111011000101100011;
assign LUT_4[4903] = 32'b11111111111111110100010001011011;
assign LUT_4[4904] = 32'b11111111111111110111110110111000;
assign LUT_4[4905] = 32'b11111111111111110001000010110000;
assign LUT_4[4906] = 32'b11111111111111110111010001011100;
assign LUT_4[4907] = 32'b11111111111111110000011101010100;
assign LUT_4[4908] = 32'b11111111111111110100110111010100;
assign LUT_4[4909] = 32'b11111111111111101110000011001100;
assign LUT_4[4910] = 32'b11111111111111110100010001111000;
assign LUT_4[4911] = 32'b11111111111111101101011101110000;
assign LUT_4[4912] = 32'b11111111111111111100011100010001;
assign LUT_4[4913] = 32'b11111111111111110101101000001001;
assign LUT_4[4914] = 32'b11111111111111111011110110110101;
assign LUT_4[4915] = 32'b11111111111111110101000010101101;
assign LUT_4[4916] = 32'b11111111111111111001011100101101;
assign LUT_4[4917] = 32'b11111111111111110010101000100101;
assign LUT_4[4918] = 32'b11111111111111111000110111010001;
assign LUT_4[4919] = 32'b11111111111111110010000011001001;
assign LUT_4[4920] = 32'b11111111111111110101101000100110;
assign LUT_4[4921] = 32'b11111111111111101110110100011110;
assign LUT_4[4922] = 32'b11111111111111110101000011001010;
assign LUT_4[4923] = 32'b11111111111111101110001111000010;
assign LUT_4[4924] = 32'b11111111111111110010101001000010;
assign LUT_4[4925] = 32'b11111111111111101011110100111010;
assign LUT_4[4926] = 32'b11111111111111110010000011100110;
assign LUT_4[4927] = 32'b11111111111111101011001111011110;
assign LUT_4[4928] = 32'b00000000000000000001100110110000;
assign LUT_4[4929] = 32'b11111111111111111010110010101000;
assign LUT_4[4930] = 32'b00000000000000000001000001010100;
assign LUT_4[4931] = 32'b11111111111111111010001101001100;
assign LUT_4[4932] = 32'b11111111111111111110100111001100;
assign LUT_4[4933] = 32'b11111111111111110111110011000100;
assign LUT_4[4934] = 32'b11111111111111111110000001110000;
assign LUT_4[4935] = 32'b11111111111111110111001101101000;
assign LUT_4[4936] = 32'b11111111111111111010110011000101;
assign LUT_4[4937] = 32'b11111111111111110011111110111101;
assign LUT_4[4938] = 32'b11111111111111111010001101101001;
assign LUT_4[4939] = 32'b11111111111111110011011001100001;
assign LUT_4[4940] = 32'b11111111111111110111110011100001;
assign LUT_4[4941] = 32'b11111111111111110000111111011001;
assign LUT_4[4942] = 32'b11111111111111110111001110000101;
assign LUT_4[4943] = 32'b11111111111111110000011001111101;
assign LUT_4[4944] = 32'b11111111111111111111011000011110;
assign LUT_4[4945] = 32'b11111111111111111000100100010110;
assign LUT_4[4946] = 32'b11111111111111111110110011000010;
assign LUT_4[4947] = 32'b11111111111111110111111110111010;
assign LUT_4[4948] = 32'b11111111111111111100011000111010;
assign LUT_4[4949] = 32'b11111111111111110101100100110010;
assign LUT_4[4950] = 32'b11111111111111111011110011011110;
assign LUT_4[4951] = 32'b11111111111111110100111111010110;
assign LUT_4[4952] = 32'b11111111111111111000100100110011;
assign LUT_4[4953] = 32'b11111111111111110001110000101011;
assign LUT_4[4954] = 32'b11111111111111110111111111010111;
assign LUT_4[4955] = 32'b11111111111111110001001011001111;
assign LUT_4[4956] = 32'b11111111111111110101100101001111;
assign LUT_4[4957] = 32'b11111111111111101110110001000111;
assign LUT_4[4958] = 32'b11111111111111110100111111110011;
assign LUT_4[4959] = 32'b11111111111111101110001011101011;
assign LUT_4[4960] = 32'b00000000000000000000000001110111;
assign LUT_4[4961] = 32'b11111111111111111001001101101111;
assign LUT_4[4962] = 32'b11111111111111111111011100011011;
assign LUT_4[4963] = 32'b11111111111111111000101000010011;
assign LUT_4[4964] = 32'b11111111111111111101000010010011;
assign LUT_4[4965] = 32'b11111111111111110110001110001011;
assign LUT_4[4966] = 32'b11111111111111111100011100110111;
assign LUT_4[4967] = 32'b11111111111111110101101000101111;
assign LUT_4[4968] = 32'b11111111111111111001001110001100;
assign LUT_4[4969] = 32'b11111111111111110010011010000100;
assign LUT_4[4970] = 32'b11111111111111111000101000110000;
assign LUT_4[4971] = 32'b11111111111111110001110100101000;
assign LUT_4[4972] = 32'b11111111111111110110001110101000;
assign LUT_4[4973] = 32'b11111111111111101111011010100000;
assign LUT_4[4974] = 32'b11111111111111110101101001001100;
assign LUT_4[4975] = 32'b11111111111111101110110101000100;
assign LUT_4[4976] = 32'b11111111111111111101110011100101;
assign LUT_4[4977] = 32'b11111111111111110110111111011101;
assign LUT_4[4978] = 32'b11111111111111111101001110001001;
assign LUT_4[4979] = 32'b11111111111111110110011010000001;
assign LUT_4[4980] = 32'b11111111111111111010110100000001;
assign LUT_4[4981] = 32'b11111111111111110011111111111001;
assign LUT_4[4982] = 32'b11111111111111111010001110100101;
assign LUT_4[4983] = 32'b11111111111111110011011010011101;
assign LUT_4[4984] = 32'b11111111111111110110111111111010;
assign LUT_4[4985] = 32'b11111111111111110000001011110010;
assign LUT_4[4986] = 32'b11111111111111110110011010011110;
assign LUT_4[4987] = 32'b11111111111111101111100110010110;
assign LUT_4[4988] = 32'b11111111111111110100000000010110;
assign LUT_4[4989] = 32'b11111111111111101101001100001110;
assign LUT_4[4990] = 32'b11111111111111110011011010111010;
assign LUT_4[4991] = 32'b11111111111111101100100110110010;
assign LUT_4[4992] = 32'b00000000000000000010110101100100;
assign LUT_4[4993] = 32'b11111111111111111100000001011100;
assign LUT_4[4994] = 32'b00000000000000000010010000001000;
assign LUT_4[4995] = 32'b11111111111111111011011100000000;
assign LUT_4[4996] = 32'b11111111111111111111110110000000;
assign LUT_4[4997] = 32'b11111111111111111001000001111000;
assign LUT_4[4998] = 32'b11111111111111111111010000100100;
assign LUT_4[4999] = 32'b11111111111111111000011100011100;
assign LUT_4[5000] = 32'b11111111111111111100000001111001;
assign LUT_4[5001] = 32'b11111111111111110101001101110001;
assign LUT_4[5002] = 32'b11111111111111111011011100011101;
assign LUT_4[5003] = 32'b11111111111111110100101000010101;
assign LUT_4[5004] = 32'b11111111111111111001000010010101;
assign LUT_4[5005] = 32'b11111111111111110010001110001101;
assign LUT_4[5006] = 32'b11111111111111111000011100111001;
assign LUT_4[5007] = 32'b11111111111111110001101000110001;
assign LUT_4[5008] = 32'b00000000000000000000100111010010;
assign LUT_4[5009] = 32'b11111111111111111001110011001010;
assign LUT_4[5010] = 32'b00000000000000000000000001110110;
assign LUT_4[5011] = 32'b11111111111111111001001101101110;
assign LUT_4[5012] = 32'b11111111111111111101100111101110;
assign LUT_4[5013] = 32'b11111111111111110110110011100110;
assign LUT_4[5014] = 32'b11111111111111111101000010010010;
assign LUT_4[5015] = 32'b11111111111111110110001110001010;
assign LUT_4[5016] = 32'b11111111111111111001110011100111;
assign LUT_4[5017] = 32'b11111111111111110010111111011111;
assign LUT_4[5018] = 32'b11111111111111111001001110001011;
assign LUT_4[5019] = 32'b11111111111111110010011010000011;
assign LUT_4[5020] = 32'b11111111111111110110110100000011;
assign LUT_4[5021] = 32'b11111111111111101111111111111011;
assign LUT_4[5022] = 32'b11111111111111110110001110100111;
assign LUT_4[5023] = 32'b11111111111111101111011010011111;
assign LUT_4[5024] = 32'b00000000000000000001010000101011;
assign LUT_4[5025] = 32'b11111111111111111010011100100011;
assign LUT_4[5026] = 32'b00000000000000000000101011001111;
assign LUT_4[5027] = 32'b11111111111111111001110111000111;
assign LUT_4[5028] = 32'b11111111111111111110010001000111;
assign LUT_4[5029] = 32'b11111111111111110111011100111111;
assign LUT_4[5030] = 32'b11111111111111111101101011101011;
assign LUT_4[5031] = 32'b11111111111111110110110111100011;
assign LUT_4[5032] = 32'b11111111111111111010011101000000;
assign LUT_4[5033] = 32'b11111111111111110011101000111000;
assign LUT_4[5034] = 32'b11111111111111111001110111100100;
assign LUT_4[5035] = 32'b11111111111111110011000011011100;
assign LUT_4[5036] = 32'b11111111111111110111011101011100;
assign LUT_4[5037] = 32'b11111111111111110000101001010100;
assign LUT_4[5038] = 32'b11111111111111110110111000000000;
assign LUT_4[5039] = 32'b11111111111111110000000011111000;
assign LUT_4[5040] = 32'b11111111111111111111000010011001;
assign LUT_4[5041] = 32'b11111111111111111000001110010001;
assign LUT_4[5042] = 32'b11111111111111111110011100111101;
assign LUT_4[5043] = 32'b11111111111111110111101000110101;
assign LUT_4[5044] = 32'b11111111111111111100000010110101;
assign LUT_4[5045] = 32'b11111111111111110101001110101101;
assign LUT_4[5046] = 32'b11111111111111111011011101011001;
assign LUT_4[5047] = 32'b11111111111111110100101001010001;
assign LUT_4[5048] = 32'b11111111111111111000001110101110;
assign LUT_4[5049] = 32'b11111111111111110001011010100110;
assign LUT_4[5050] = 32'b11111111111111110111101001010010;
assign LUT_4[5051] = 32'b11111111111111110000110101001010;
assign LUT_4[5052] = 32'b11111111111111110101001111001010;
assign LUT_4[5053] = 32'b11111111111111101110011011000010;
assign LUT_4[5054] = 32'b11111111111111110100101001101110;
assign LUT_4[5055] = 32'b11111111111111101101110101100110;
assign LUT_4[5056] = 32'b00000000000000000100001100111000;
assign LUT_4[5057] = 32'b11111111111111111101011000110000;
assign LUT_4[5058] = 32'b00000000000000000011100111011100;
assign LUT_4[5059] = 32'b11111111111111111100110011010100;
assign LUT_4[5060] = 32'b00000000000000000001001101010100;
assign LUT_4[5061] = 32'b11111111111111111010011001001100;
assign LUT_4[5062] = 32'b00000000000000000000100111111000;
assign LUT_4[5063] = 32'b11111111111111111001110011110000;
assign LUT_4[5064] = 32'b11111111111111111101011001001101;
assign LUT_4[5065] = 32'b11111111111111110110100101000101;
assign LUT_4[5066] = 32'b11111111111111111100110011110001;
assign LUT_4[5067] = 32'b11111111111111110101111111101001;
assign LUT_4[5068] = 32'b11111111111111111010011001101001;
assign LUT_4[5069] = 32'b11111111111111110011100101100001;
assign LUT_4[5070] = 32'b11111111111111111001110100001101;
assign LUT_4[5071] = 32'b11111111111111110011000000000101;
assign LUT_4[5072] = 32'b00000000000000000001111110100110;
assign LUT_4[5073] = 32'b11111111111111111011001010011110;
assign LUT_4[5074] = 32'b00000000000000000001011001001010;
assign LUT_4[5075] = 32'b11111111111111111010100101000010;
assign LUT_4[5076] = 32'b11111111111111111110111111000010;
assign LUT_4[5077] = 32'b11111111111111111000001010111010;
assign LUT_4[5078] = 32'b11111111111111111110011001100110;
assign LUT_4[5079] = 32'b11111111111111110111100101011110;
assign LUT_4[5080] = 32'b11111111111111111011001010111011;
assign LUT_4[5081] = 32'b11111111111111110100010110110011;
assign LUT_4[5082] = 32'b11111111111111111010100101011111;
assign LUT_4[5083] = 32'b11111111111111110011110001010111;
assign LUT_4[5084] = 32'b11111111111111111000001011010111;
assign LUT_4[5085] = 32'b11111111111111110001010111001111;
assign LUT_4[5086] = 32'b11111111111111110111100101111011;
assign LUT_4[5087] = 32'b11111111111111110000110001110011;
assign LUT_4[5088] = 32'b00000000000000000010100111111111;
assign LUT_4[5089] = 32'b11111111111111111011110011110111;
assign LUT_4[5090] = 32'b00000000000000000010000010100011;
assign LUT_4[5091] = 32'b11111111111111111011001110011011;
assign LUT_4[5092] = 32'b11111111111111111111101000011011;
assign LUT_4[5093] = 32'b11111111111111111000110100010011;
assign LUT_4[5094] = 32'b11111111111111111111000010111111;
assign LUT_4[5095] = 32'b11111111111111111000001110110111;
assign LUT_4[5096] = 32'b11111111111111111011110100010100;
assign LUT_4[5097] = 32'b11111111111111110101000000001100;
assign LUT_4[5098] = 32'b11111111111111111011001110111000;
assign LUT_4[5099] = 32'b11111111111111110100011010110000;
assign LUT_4[5100] = 32'b11111111111111111000110100110000;
assign LUT_4[5101] = 32'b11111111111111110010000000101000;
assign LUT_4[5102] = 32'b11111111111111111000001111010100;
assign LUT_4[5103] = 32'b11111111111111110001011011001100;
assign LUT_4[5104] = 32'b00000000000000000000011001101101;
assign LUT_4[5105] = 32'b11111111111111111001100101100101;
assign LUT_4[5106] = 32'b11111111111111111111110100010001;
assign LUT_4[5107] = 32'b11111111111111111001000000001001;
assign LUT_4[5108] = 32'b11111111111111111101011010001001;
assign LUT_4[5109] = 32'b11111111111111110110100110000001;
assign LUT_4[5110] = 32'b11111111111111111100110100101101;
assign LUT_4[5111] = 32'b11111111111111110110000000100101;
assign LUT_4[5112] = 32'b11111111111111111001100110000010;
assign LUT_4[5113] = 32'b11111111111111110010110001111010;
assign LUT_4[5114] = 32'b11111111111111111001000000100110;
assign LUT_4[5115] = 32'b11111111111111110010001100011110;
assign LUT_4[5116] = 32'b11111111111111110110100110011110;
assign LUT_4[5117] = 32'b11111111111111101111110010010110;
assign LUT_4[5118] = 32'b11111111111111110110000001000010;
assign LUT_4[5119] = 32'b11111111111111101111001100111010;
assign LUT_4[5120] = 32'b11111111111111111101111010010000;
assign LUT_4[5121] = 32'b11111111111111110111000110001000;
assign LUT_4[5122] = 32'b11111111111111111101010100110100;
assign LUT_4[5123] = 32'b11111111111111110110100000101100;
assign LUT_4[5124] = 32'b11111111111111111010111010101100;
assign LUT_4[5125] = 32'b11111111111111110100000110100100;
assign LUT_4[5126] = 32'b11111111111111111010010101010000;
assign LUT_4[5127] = 32'b11111111111111110011100001001000;
assign LUT_4[5128] = 32'b11111111111111110111000110100101;
assign LUT_4[5129] = 32'b11111111111111110000010010011101;
assign LUT_4[5130] = 32'b11111111111111110110100001001001;
assign LUT_4[5131] = 32'b11111111111111101111101101000001;
assign LUT_4[5132] = 32'b11111111111111110100000111000001;
assign LUT_4[5133] = 32'b11111111111111101101010010111001;
assign LUT_4[5134] = 32'b11111111111111110011100001100101;
assign LUT_4[5135] = 32'b11111111111111101100101101011101;
assign LUT_4[5136] = 32'b11111111111111111011101011111110;
assign LUT_4[5137] = 32'b11111111111111110100110111110110;
assign LUT_4[5138] = 32'b11111111111111111011000110100010;
assign LUT_4[5139] = 32'b11111111111111110100010010011010;
assign LUT_4[5140] = 32'b11111111111111111000101100011010;
assign LUT_4[5141] = 32'b11111111111111110001111000010010;
assign LUT_4[5142] = 32'b11111111111111111000000110111110;
assign LUT_4[5143] = 32'b11111111111111110001010010110110;
assign LUT_4[5144] = 32'b11111111111111110100111000010011;
assign LUT_4[5145] = 32'b11111111111111101110000100001011;
assign LUT_4[5146] = 32'b11111111111111110100010010110111;
assign LUT_4[5147] = 32'b11111111111111101101011110101111;
assign LUT_4[5148] = 32'b11111111111111110001111000101111;
assign LUT_4[5149] = 32'b11111111111111101011000100100111;
assign LUT_4[5150] = 32'b11111111111111110001010011010011;
assign LUT_4[5151] = 32'b11111111111111101010011111001011;
assign LUT_4[5152] = 32'b11111111111111111100010101010111;
assign LUT_4[5153] = 32'b11111111111111110101100001001111;
assign LUT_4[5154] = 32'b11111111111111111011101111111011;
assign LUT_4[5155] = 32'b11111111111111110100111011110011;
assign LUT_4[5156] = 32'b11111111111111111001010101110011;
assign LUT_4[5157] = 32'b11111111111111110010100001101011;
assign LUT_4[5158] = 32'b11111111111111111000110000010111;
assign LUT_4[5159] = 32'b11111111111111110001111100001111;
assign LUT_4[5160] = 32'b11111111111111110101100001101100;
assign LUT_4[5161] = 32'b11111111111111101110101101100100;
assign LUT_4[5162] = 32'b11111111111111110100111100010000;
assign LUT_4[5163] = 32'b11111111111111101110001000001000;
assign LUT_4[5164] = 32'b11111111111111110010100010001000;
assign LUT_4[5165] = 32'b11111111111111101011101110000000;
assign LUT_4[5166] = 32'b11111111111111110001111100101100;
assign LUT_4[5167] = 32'b11111111111111101011001000100100;
assign LUT_4[5168] = 32'b11111111111111111010000111000101;
assign LUT_4[5169] = 32'b11111111111111110011010010111101;
assign LUT_4[5170] = 32'b11111111111111111001100001101001;
assign LUT_4[5171] = 32'b11111111111111110010101101100001;
assign LUT_4[5172] = 32'b11111111111111110111000111100001;
assign LUT_4[5173] = 32'b11111111111111110000010011011001;
assign LUT_4[5174] = 32'b11111111111111110110100010000101;
assign LUT_4[5175] = 32'b11111111111111101111101101111101;
assign LUT_4[5176] = 32'b11111111111111110011010011011010;
assign LUT_4[5177] = 32'b11111111111111101100011111010010;
assign LUT_4[5178] = 32'b11111111111111110010101101111110;
assign LUT_4[5179] = 32'b11111111111111101011111001110110;
assign LUT_4[5180] = 32'b11111111111111110000010011110110;
assign LUT_4[5181] = 32'b11111111111111101001011111101110;
assign LUT_4[5182] = 32'b11111111111111101111101110011010;
assign LUT_4[5183] = 32'b11111111111111101000111010010010;
assign LUT_4[5184] = 32'b11111111111111111111010001100100;
assign LUT_4[5185] = 32'b11111111111111111000011101011100;
assign LUT_4[5186] = 32'b11111111111111111110101100001000;
assign LUT_4[5187] = 32'b11111111111111110111111000000000;
assign LUT_4[5188] = 32'b11111111111111111100010010000000;
assign LUT_4[5189] = 32'b11111111111111110101011101111000;
assign LUT_4[5190] = 32'b11111111111111111011101100100100;
assign LUT_4[5191] = 32'b11111111111111110100111000011100;
assign LUT_4[5192] = 32'b11111111111111111000011101111001;
assign LUT_4[5193] = 32'b11111111111111110001101001110001;
assign LUT_4[5194] = 32'b11111111111111110111111000011101;
assign LUT_4[5195] = 32'b11111111111111110001000100010101;
assign LUT_4[5196] = 32'b11111111111111110101011110010101;
assign LUT_4[5197] = 32'b11111111111111101110101010001101;
assign LUT_4[5198] = 32'b11111111111111110100111000111001;
assign LUT_4[5199] = 32'b11111111111111101110000100110001;
assign LUT_4[5200] = 32'b11111111111111111101000011010010;
assign LUT_4[5201] = 32'b11111111111111110110001111001010;
assign LUT_4[5202] = 32'b11111111111111111100011101110110;
assign LUT_4[5203] = 32'b11111111111111110101101001101110;
assign LUT_4[5204] = 32'b11111111111111111010000011101110;
assign LUT_4[5205] = 32'b11111111111111110011001111100110;
assign LUT_4[5206] = 32'b11111111111111111001011110010010;
assign LUT_4[5207] = 32'b11111111111111110010101010001010;
assign LUT_4[5208] = 32'b11111111111111110110001111100111;
assign LUT_4[5209] = 32'b11111111111111101111011011011111;
assign LUT_4[5210] = 32'b11111111111111110101101010001011;
assign LUT_4[5211] = 32'b11111111111111101110110110000011;
assign LUT_4[5212] = 32'b11111111111111110011010000000011;
assign LUT_4[5213] = 32'b11111111111111101100011011111011;
assign LUT_4[5214] = 32'b11111111111111110010101010100111;
assign LUT_4[5215] = 32'b11111111111111101011110110011111;
assign LUT_4[5216] = 32'b11111111111111111101101100101011;
assign LUT_4[5217] = 32'b11111111111111110110111000100011;
assign LUT_4[5218] = 32'b11111111111111111101000111001111;
assign LUT_4[5219] = 32'b11111111111111110110010011000111;
assign LUT_4[5220] = 32'b11111111111111111010101101000111;
assign LUT_4[5221] = 32'b11111111111111110011111000111111;
assign LUT_4[5222] = 32'b11111111111111111010000111101011;
assign LUT_4[5223] = 32'b11111111111111110011010011100011;
assign LUT_4[5224] = 32'b11111111111111110110111001000000;
assign LUT_4[5225] = 32'b11111111111111110000000100111000;
assign LUT_4[5226] = 32'b11111111111111110110010011100100;
assign LUT_4[5227] = 32'b11111111111111101111011111011100;
assign LUT_4[5228] = 32'b11111111111111110011111001011100;
assign LUT_4[5229] = 32'b11111111111111101101000101010100;
assign LUT_4[5230] = 32'b11111111111111110011010100000000;
assign LUT_4[5231] = 32'b11111111111111101100011111111000;
assign LUT_4[5232] = 32'b11111111111111111011011110011001;
assign LUT_4[5233] = 32'b11111111111111110100101010010001;
assign LUT_4[5234] = 32'b11111111111111111010111000111101;
assign LUT_4[5235] = 32'b11111111111111110100000100110101;
assign LUT_4[5236] = 32'b11111111111111111000011110110101;
assign LUT_4[5237] = 32'b11111111111111110001101010101101;
assign LUT_4[5238] = 32'b11111111111111110111111001011001;
assign LUT_4[5239] = 32'b11111111111111110001000101010001;
assign LUT_4[5240] = 32'b11111111111111110100101010101110;
assign LUT_4[5241] = 32'b11111111111111101101110110100110;
assign LUT_4[5242] = 32'b11111111111111110100000101010010;
assign LUT_4[5243] = 32'b11111111111111101101010001001010;
assign LUT_4[5244] = 32'b11111111111111110001101011001010;
assign LUT_4[5245] = 32'b11111111111111101010110111000010;
assign LUT_4[5246] = 32'b11111111111111110001000101101110;
assign LUT_4[5247] = 32'b11111111111111101010010001100110;
assign LUT_4[5248] = 32'b00000000000000000000100000011000;
assign LUT_4[5249] = 32'b11111111111111111001101100010000;
assign LUT_4[5250] = 32'b11111111111111111111111010111100;
assign LUT_4[5251] = 32'b11111111111111111001000110110100;
assign LUT_4[5252] = 32'b11111111111111111101100000110100;
assign LUT_4[5253] = 32'b11111111111111110110101100101100;
assign LUT_4[5254] = 32'b11111111111111111100111011011000;
assign LUT_4[5255] = 32'b11111111111111110110000111010000;
assign LUT_4[5256] = 32'b11111111111111111001101100101101;
assign LUT_4[5257] = 32'b11111111111111110010111000100101;
assign LUT_4[5258] = 32'b11111111111111111001000111010001;
assign LUT_4[5259] = 32'b11111111111111110010010011001001;
assign LUT_4[5260] = 32'b11111111111111110110101101001001;
assign LUT_4[5261] = 32'b11111111111111101111111001000001;
assign LUT_4[5262] = 32'b11111111111111110110000111101101;
assign LUT_4[5263] = 32'b11111111111111101111010011100101;
assign LUT_4[5264] = 32'b11111111111111111110010010000110;
assign LUT_4[5265] = 32'b11111111111111110111011101111110;
assign LUT_4[5266] = 32'b11111111111111111101101100101010;
assign LUT_4[5267] = 32'b11111111111111110110111000100010;
assign LUT_4[5268] = 32'b11111111111111111011010010100010;
assign LUT_4[5269] = 32'b11111111111111110100011110011010;
assign LUT_4[5270] = 32'b11111111111111111010101101000110;
assign LUT_4[5271] = 32'b11111111111111110011111000111110;
assign LUT_4[5272] = 32'b11111111111111110111011110011011;
assign LUT_4[5273] = 32'b11111111111111110000101010010011;
assign LUT_4[5274] = 32'b11111111111111110110111000111111;
assign LUT_4[5275] = 32'b11111111111111110000000100110111;
assign LUT_4[5276] = 32'b11111111111111110100011110110111;
assign LUT_4[5277] = 32'b11111111111111101101101010101111;
assign LUT_4[5278] = 32'b11111111111111110011111001011011;
assign LUT_4[5279] = 32'b11111111111111101101000101010011;
assign LUT_4[5280] = 32'b11111111111111111110111011011111;
assign LUT_4[5281] = 32'b11111111111111111000000111010111;
assign LUT_4[5282] = 32'b11111111111111111110010110000011;
assign LUT_4[5283] = 32'b11111111111111110111100001111011;
assign LUT_4[5284] = 32'b11111111111111111011111011111011;
assign LUT_4[5285] = 32'b11111111111111110101000111110011;
assign LUT_4[5286] = 32'b11111111111111111011010110011111;
assign LUT_4[5287] = 32'b11111111111111110100100010010111;
assign LUT_4[5288] = 32'b11111111111111111000000111110100;
assign LUT_4[5289] = 32'b11111111111111110001010011101100;
assign LUT_4[5290] = 32'b11111111111111110111100010011000;
assign LUT_4[5291] = 32'b11111111111111110000101110010000;
assign LUT_4[5292] = 32'b11111111111111110101001000010000;
assign LUT_4[5293] = 32'b11111111111111101110010100001000;
assign LUT_4[5294] = 32'b11111111111111110100100010110100;
assign LUT_4[5295] = 32'b11111111111111101101101110101100;
assign LUT_4[5296] = 32'b11111111111111111100101101001101;
assign LUT_4[5297] = 32'b11111111111111110101111001000101;
assign LUT_4[5298] = 32'b11111111111111111100000111110001;
assign LUT_4[5299] = 32'b11111111111111110101010011101001;
assign LUT_4[5300] = 32'b11111111111111111001101101101001;
assign LUT_4[5301] = 32'b11111111111111110010111001100001;
assign LUT_4[5302] = 32'b11111111111111111001001000001101;
assign LUT_4[5303] = 32'b11111111111111110010010100000101;
assign LUT_4[5304] = 32'b11111111111111110101111001100010;
assign LUT_4[5305] = 32'b11111111111111101111000101011010;
assign LUT_4[5306] = 32'b11111111111111110101010100000110;
assign LUT_4[5307] = 32'b11111111111111101110011111111110;
assign LUT_4[5308] = 32'b11111111111111110010111001111110;
assign LUT_4[5309] = 32'b11111111111111101100000101110110;
assign LUT_4[5310] = 32'b11111111111111110010010100100010;
assign LUT_4[5311] = 32'b11111111111111101011100000011010;
assign LUT_4[5312] = 32'b00000000000000000001110111101100;
assign LUT_4[5313] = 32'b11111111111111111011000011100100;
assign LUT_4[5314] = 32'b00000000000000000001010010010000;
assign LUT_4[5315] = 32'b11111111111111111010011110001000;
assign LUT_4[5316] = 32'b11111111111111111110111000001000;
assign LUT_4[5317] = 32'b11111111111111111000000100000000;
assign LUT_4[5318] = 32'b11111111111111111110010010101100;
assign LUT_4[5319] = 32'b11111111111111110111011110100100;
assign LUT_4[5320] = 32'b11111111111111111011000100000001;
assign LUT_4[5321] = 32'b11111111111111110100001111111001;
assign LUT_4[5322] = 32'b11111111111111111010011110100101;
assign LUT_4[5323] = 32'b11111111111111110011101010011101;
assign LUT_4[5324] = 32'b11111111111111111000000100011101;
assign LUT_4[5325] = 32'b11111111111111110001010000010101;
assign LUT_4[5326] = 32'b11111111111111110111011111000001;
assign LUT_4[5327] = 32'b11111111111111110000101010111001;
assign LUT_4[5328] = 32'b11111111111111111111101001011010;
assign LUT_4[5329] = 32'b11111111111111111000110101010010;
assign LUT_4[5330] = 32'b11111111111111111111000011111110;
assign LUT_4[5331] = 32'b11111111111111111000001111110110;
assign LUT_4[5332] = 32'b11111111111111111100101001110110;
assign LUT_4[5333] = 32'b11111111111111110101110101101110;
assign LUT_4[5334] = 32'b11111111111111111100000100011010;
assign LUT_4[5335] = 32'b11111111111111110101010000010010;
assign LUT_4[5336] = 32'b11111111111111111000110101101111;
assign LUT_4[5337] = 32'b11111111111111110010000001100111;
assign LUT_4[5338] = 32'b11111111111111111000010000010011;
assign LUT_4[5339] = 32'b11111111111111110001011100001011;
assign LUT_4[5340] = 32'b11111111111111110101110110001011;
assign LUT_4[5341] = 32'b11111111111111101111000010000011;
assign LUT_4[5342] = 32'b11111111111111110101010000101111;
assign LUT_4[5343] = 32'b11111111111111101110011100100111;
assign LUT_4[5344] = 32'b00000000000000000000010010110011;
assign LUT_4[5345] = 32'b11111111111111111001011110101011;
assign LUT_4[5346] = 32'b11111111111111111111101101010111;
assign LUT_4[5347] = 32'b11111111111111111000111001001111;
assign LUT_4[5348] = 32'b11111111111111111101010011001111;
assign LUT_4[5349] = 32'b11111111111111110110011111000111;
assign LUT_4[5350] = 32'b11111111111111111100101101110011;
assign LUT_4[5351] = 32'b11111111111111110101111001101011;
assign LUT_4[5352] = 32'b11111111111111111001011111001000;
assign LUT_4[5353] = 32'b11111111111111110010101011000000;
assign LUT_4[5354] = 32'b11111111111111111000111001101100;
assign LUT_4[5355] = 32'b11111111111111110010000101100100;
assign LUT_4[5356] = 32'b11111111111111110110011111100100;
assign LUT_4[5357] = 32'b11111111111111101111101011011100;
assign LUT_4[5358] = 32'b11111111111111110101111010001000;
assign LUT_4[5359] = 32'b11111111111111101111000110000000;
assign LUT_4[5360] = 32'b11111111111111111110000100100001;
assign LUT_4[5361] = 32'b11111111111111110111010000011001;
assign LUT_4[5362] = 32'b11111111111111111101011111000101;
assign LUT_4[5363] = 32'b11111111111111110110101010111101;
assign LUT_4[5364] = 32'b11111111111111111011000100111101;
assign LUT_4[5365] = 32'b11111111111111110100010000110101;
assign LUT_4[5366] = 32'b11111111111111111010011111100001;
assign LUT_4[5367] = 32'b11111111111111110011101011011001;
assign LUT_4[5368] = 32'b11111111111111110111010000110110;
assign LUT_4[5369] = 32'b11111111111111110000011100101110;
assign LUT_4[5370] = 32'b11111111111111110110101011011010;
assign LUT_4[5371] = 32'b11111111111111101111110111010010;
assign LUT_4[5372] = 32'b11111111111111110100010001010010;
assign LUT_4[5373] = 32'b11111111111111101101011101001010;
assign LUT_4[5374] = 32'b11111111111111110011101011110110;
assign LUT_4[5375] = 32'b11111111111111101100110111101110;
assign LUT_4[5376] = 32'b00000000000000000010110101110011;
assign LUT_4[5377] = 32'b11111111111111111100000001101011;
assign LUT_4[5378] = 32'b00000000000000000010010000010111;
assign LUT_4[5379] = 32'b11111111111111111011011100001111;
assign LUT_4[5380] = 32'b11111111111111111111110110001111;
assign LUT_4[5381] = 32'b11111111111111111001000010000111;
assign LUT_4[5382] = 32'b11111111111111111111010000110011;
assign LUT_4[5383] = 32'b11111111111111111000011100101011;
assign LUT_4[5384] = 32'b11111111111111111100000010001000;
assign LUT_4[5385] = 32'b11111111111111110101001110000000;
assign LUT_4[5386] = 32'b11111111111111111011011100101100;
assign LUT_4[5387] = 32'b11111111111111110100101000100100;
assign LUT_4[5388] = 32'b11111111111111111001000010100100;
assign LUT_4[5389] = 32'b11111111111111110010001110011100;
assign LUT_4[5390] = 32'b11111111111111111000011101001000;
assign LUT_4[5391] = 32'b11111111111111110001101001000000;
assign LUT_4[5392] = 32'b00000000000000000000100111100001;
assign LUT_4[5393] = 32'b11111111111111111001110011011001;
assign LUT_4[5394] = 32'b00000000000000000000000010000101;
assign LUT_4[5395] = 32'b11111111111111111001001101111101;
assign LUT_4[5396] = 32'b11111111111111111101100111111101;
assign LUT_4[5397] = 32'b11111111111111110110110011110101;
assign LUT_4[5398] = 32'b11111111111111111101000010100001;
assign LUT_4[5399] = 32'b11111111111111110110001110011001;
assign LUT_4[5400] = 32'b11111111111111111001110011110110;
assign LUT_4[5401] = 32'b11111111111111110010111111101110;
assign LUT_4[5402] = 32'b11111111111111111001001110011010;
assign LUT_4[5403] = 32'b11111111111111110010011010010010;
assign LUT_4[5404] = 32'b11111111111111110110110100010010;
assign LUT_4[5405] = 32'b11111111111111110000000000001010;
assign LUT_4[5406] = 32'b11111111111111110110001110110110;
assign LUT_4[5407] = 32'b11111111111111101111011010101110;
assign LUT_4[5408] = 32'b00000000000000000001010000111010;
assign LUT_4[5409] = 32'b11111111111111111010011100110010;
assign LUT_4[5410] = 32'b00000000000000000000101011011110;
assign LUT_4[5411] = 32'b11111111111111111001110111010110;
assign LUT_4[5412] = 32'b11111111111111111110010001010110;
assign LUT_4[5413] = 32'b11111111111111110111011101001110;
assign LUT_4[5414] = 32'b11111111111111111101101011111010;
assign LUT_4[5415] = 32'b11111111111111110110110111110010;
assign LUT_4[5416] = 32'b11111111111111111010011101001111;
assign LUT_4[5417] = 32'b11111111111111110011101001000111;
assign LUT_4[5418] = 32'b11111111111111111001110111110011;
assign LUT_4[5419] = 32'b11111111111111110011000011101011;
assign LUT_4[5420] = 32'b11111111111111110111011101101011;
assign LUT_4[5421] = 32'b11111111111111110000101001100011;
assign LUT_4[5422] = 32'b11111111111111110110111000001111;
assign LUT_4[5423] = 32'b11111111111111110000000100000111;
assign LUT_4[5424] = 32'b11111111111111111111000010101000;
assign LUT_4[5425] = 32'b11111111111111111000001110100000;
assign LUT_4[5426] = 32'b11111111111111111110011101001100;
assign LUT_4[5427] = 32'b11111111111111110111101001000100;
assign LUT_4[5428] = 32'b11111111111111111100000011000100;
assign LUT_4[5429] = 32'b11111111111111110101001110111100;
assign LUT_4[5430] = 32'b11111111111111111011011101101000;
assign LUT_4[5431] = 32'b11111111111111110100101001100000;
assign LUT_4[5432] = 32'b11111111111111111000001110111101;
assign LUT_4[5433] = 32'b11111111111111110001011010110101;
assign LUT_4[5434] = 32'b11111111111111110111101001100001;
assign LUT_4[5435] = 32'b11111111111111110000110101011001;
assign LUT_4[5436] = 32'b11111111111111110101001111011001;
assign LUT_4[5437] = 32'b11111111111111101110011011010001;
assign LUT_4[5438] = 32'b11111111111111110100101001111101;
assign LUT_4[5439] = 32'b11111111111111101101110101110101;
assign LUT_4[5440] = 32'b00000000000000000100001101000111;
assign LUT_4[5441] = 32'b11111111111111111101011000111111;
assign LUT_4[5442] = 32'b00000000000000000011100111101011;
assign LUT_4[5443] = 32'b11111111111111111100110011100011;
assign LUT_4[5444] = 32'b00000000000000000001001101100011;
assign LUT_4[5445] = 32'b11111111111111111010011001011011;
assign LUT_4[5446] = 32'b00000000000000000000101000000111;
assign LUT_4[5447] = 32'b11111111111111111001110011111111;
assign LUT_4[5448] = 32'b11111111111111111101011001011100;
assign LUT_4[5449] = 32'b11111111111111110110100101010100;
assign LUT_4[5450] = 32'b11111111111111111100110100000000;
assign LUT_4[5451] = 32'b11111111111111110101111111111000;
assign LUT_4[5452] = 32'b11111111111111111010011001111000;
assign LUT_4[5453] = 32'b11111111111111110011100101110000;
assign LUT_4[5454] = 32'b11111111111111111001110100011100;
assign LUT_4[5455] = 32'b11111111111111110011000000010100;
assign LUT_4[5456] = 32'b00000000000000000001111110110101;
assign LUT_4[5457] = 32'b11111111111111111011001010101101;
assign LUT_4[5458] = 32'b00000000000000000001011001011001;
assign LUT_4[5459] = 32'b11111111111111111010100101010001;
assign LUT_4[5460] = 32'b11111111111111111110111111010001;
assign LUT_4[5461] = 32'b11111111111111111000001011001001;
assign LUT_4[5462] = 32'b11111111111111111110011001110101;
assign LUT_4[5463] = 32'b11111111111111110111100101101101;
assign LUT_4[5464] = 32'b11111111111111111011001011001010;
assign LUT_4[5465] = 32'b11111111111111110100010111000010;
assign LUT_4[5466] = 32'b11111111111111111010100101101110;
assign LUT_4[5467] = 32'b11111111111111110011110001100110;
assign LUT_4[5468] = 32'b11111111111111111000001011100110;
assign LUT_4[5469] = 32'b11111111111111110001010111011110;
assign LUT_4[5470] = 32'b11111111111111110111100110001010;
assign LUT_4[5471] = 32'b11111111111111110000110010000010;
assign LUT_4[5472] = 32'b00000000000000000010101000001110;
assign LUT_4[5473] = 32'b11111111111111111011110100000110;
assign LUT_4[5474] = 32'b00000000000000000010000010110010;
assign LUT_4[5475] = 32'b11111111111111111011001110101010;
assign LUT_4[5476] = 32'b11111111111111111111101000101010;
assign LUT_4[5477] = 32'b11111111111111111000110100100010;
assign LUT_4[5478] = 32'b11111111111111111111000011001110;
assign LUT_4[5479] = 32'b11111111111111111000001111000110;
assign LUT_4[5480] = 32'b11111111111111111011110100100011;
assign LUT_4[5481] = 32'b11111111111111110101000000011011;
assign LUT_4[5482] = 32'b11111111111111111011001111000111;
assign LUT_4[5483] = 32'b11111111111111110100011010111111;
assign LUT_4[5484] = 32'b11111111111111111000110100111111;
assign LUT_4[5485] = 32'b11111111111111110010000000110111;
assign LUT_4[5486] = 32'b11111111111111111000001111100011;
assign LUT_4[5487] = 32'b11111111111111110001011011011011;
assign LUT_4[5488] = 32'b00000000000000000000011001111100;
assign LUT_4[5489] = 32'b11111111111111111001100101110100;
assign LUT_4[5490] = 32'b11111111111111111111110100100000;
assign LUT_4[5491] = 32'b11111111111111111001000000011000;
assign LUT_4[5492] = 32'b11111111111111111101011010011000;
assign LUT_4[5493] = 32'b11111111111111110110100110010000;
assign LUT_4[5494] = 32'b11111111111111111100110100111100;
assign LUT_4[5495] = 32'b11111111111111110110000000110100;
assign LUT_4[5496] = 32'b11111111111111111001100110010001;
assign LUT_4[5497] = 32'b11111111111111110010110010001001;
assign LUT_4[5498] = 32'b11111111111111111001000000110101;
assign LUT_4[5499] = 32'b11111111111111110010001100101101;
assign LUT_4[5500] = 32'b11111111111111110110100110101101;
assign LUT_4[5501] = 32'b11111111111111101111110010100101;
assign LUT_4[5502] = 32'b11111111111111110110000001010001;
assign LUT_4[5503] = 32'b11111111111111101111001101001001;
assign LUT_4[5504] = 32'b00000000000000000101011011111011;
assign LUT_4[5505] = 32'b11111111111111111110100111110011;
assign LUT_4[5506] = 32'b00000000000000000100110110011111;
assign LUT_4[5507] = 32'b11111111111111111110000010010111;
assign LUT_4[5508] = 32'b00000000000000000010011100010111;
assign LUT_4[5509] = 32'b11111111111111111011101000001111;
assign LUT_4[5510] = 32'b00000000000000000001110110111011;
assign LUT_4[5511] = 32'b11111111111111111011000010110011;
assign LUT_4[5512] = 32'b11111111111111111110101000010000;
assign LUT_4[5513] = 32'b11111111111111110111110100001000;
assign LUT_4[5514] = 32'b11111111111111111110000010110100;
assign LUT_4[5515] = 32'b11111111111111110111001110101100;
assign LUT_4[5516] = 32'b11111111111111111011101000101100;
assign LUT_4[5517] = 32'b11111111111111110100110100100100;
assign LUT_4[5518] = 32'b11111111111111111011000011010000;
assign LUT_4[5519] = 32'b11111111111111110100001111001000;
assign LUT_4[5520] = 32'b00000000000000000011001101101001;
assign LUT_4[5521] = 32'b11111111111111111100011001100001;
assign LUT_4[5522] = 32'b00000000000000000010101000001101;
assign LUT_4[5523] = 32'b11111111111111111011110100000101;
assign LUT_4[5524] = 32'b00000000000000000000001110000101;
assign LUT_4[5525] = 32'b11111111111111111001011001111101;
assign LUT_4[5526] = 32'b11111111111111111111101000101001;
assign LUT_4[5527] = 32'b11111111111111111000110100100001;
assign LUT_4[5528] = 32'b11111111111111111100011001111110;
assign LUT_4[5529] = 32'b11111111111111110101100101110110;
assign LUT_4[5530] = 32'b11111111111111111011110100100010;
assign LUT_4[5531] = 32'b11111111111111110101000000011010;
assign LUT_4[5532] = 32'b11111111111111111001011010011010;
assign LUT_4[5533] = 32'b11111111111111110010100110010010;
assign LUT_4[5534] = 32'b11111111111111111000110100111110;
assign LUT_4[5535] = 32'b11111111111111110010000000110110;
assign LUT_4[5536] = 32'b00000000000000000011110111000010;
assign LUT_4[5537] = 32'b11111111111111111101000010111010;
assign LUT_4[5538] = 32'b00000000000000000011010001100110;
assign LUT_4[5539] = 32'b11111111111111111100011101011110;
assign LUT_4[5540] = 32'b00000000000000000000110111011110;
assign LUT_4[5541] = 32'b11111111111111111010000011010110;
assign LUT_4[5542] = 32'b00000000000000000000010010000010;
assign LUT_4[5543] = 32'b11111111111111111001011101111010;
assign LUT_4[5544] = 32'b11111111111111111101000011010111;
assign LUT_4[5545] = 32'b11111111111111110110001111001111;
assign LUT_4[5546] = 32'b11111111111111111100011101111011;
assign LUT_4[5547] = 32'b11111111111111110101101001110011;
assign LUT_4[5548] = 32'b11111111111111111010000011110011;
assign LUT_4[5549] = 32'b11111111111111110011001111101011;
assign LUT_4[5550] = 32'b11111111111111111001011110010111;
assign LUT_4[5551] = 32'b11111111111111110010101010001111;
assign LUT_4[5552] = 32'b00000000000000000001101000110000;
assign LUT_4[5553] = 32'b11111111111111111010110100101000;
assign LUT_4[5554] = 32'b00000000000000000001000011010100;
assign LUT_4[5555] = 32'b11111111111111111010001111001100;
assign LUT_4[5556] = 32'b11111111111111111110101001001100;
assign LUT_4[5557] = 32'b11111111111111110111110101000100;
assign LUT_4[5558] = 32'b11111111111111111110000011110000;
assign LUT_4[5559] = 32'b11111111111111110111001111101000;
assign LUT_4[5560] = 32'b11111111111111111010110101000101;
assign LUT_4[5561] = 32'b11111111111111110100000000111101;
assign LUT_4[5562] = 32'b11111111111111111010001111101001;
assign LUT_4[5563] = 32'b11111111111111110011011011100001;
assign LUT_4[5564] = 32'b11111111111111110111110101100001;
assign LUT_4[5565] = 32'b11111111111111110001000001011001;
assign LUT_4[5566] = 32'b11111111111111110111010000000101;
assign LUT_4[5567] = 32'b11111111111111110000011011111101;
assign LUT_4[5568] = 32'b00000000000000000110110011001111;
assign LUT_4[5569] = 32'b11111111111111111111111111000111;
assign LUT_4[5570] = 32'b00000000000000000110001101110011;
assign LUT_4[5571] = 32'b11111111111111111111011001101011;
assign LUT_4[5572] = 32'b00000000000000000011110011101011;
assign LUT_4[5573] = 32'b11111111111111111100111111100011;
assign LUT_4[5574] = 32'b00000000000000000011001110001111;
assign LUT_4[5575] = 32'b11111111111111111100011010000111;
assign LUT_4[5576] = 32'b11111111111111111111111111100100;
assign LUT_4[5577] = 32'b11111111111111111001001011011100;
assign LUT_4[5578] = 32'b11111111111111111111011010001000;
assign LUT_4[5579] = 32'b11111111111111111000100110000000;
assign LUT_4[5580] = 32'b11111111111111111101000000000000;
assign LUT_4[5581] = 32'b11111111111111110110001011111000;
assign LUT_4[5582] = 32'b11111111111111111100011010100100;
assign LUT_4[5583] = 32'b11111111111111110101100110011100;
assign LUT_4[5584] = 32'b00000000000000000100100100111101;
assign LUT_4[5585] = 32'b11111111111111111101110000110101;
assign LUT_4[5586] = 32'b00000000000000000011111111100001;
assign LUT_4[5587] = 32'b11111111111111111101001011011001;
assign LUT_4[5588] = 32'b00000000000000000001100101011001;
assign LUT_4[5589] = 32'b11111111111111111010110001010001;
assign LUT_4[5590] = 32'b00000000000000000000111111111101;
assign LUT_4[5591] = 32'b11111111111111111010001011110101;
assign LUT_4[5592] = 32'b11111111111111111101110001010010;
assign LUT_4[5593] = 32'b11111111111111110110111101001010;
assign LUT_4[5594] = 32'b11111111111111111101001011110110;
assign LUT_4[5595] = 32'b11111111111111110110010111101110;
assign LUT_4[5596] = 32'b11111111111111111010110001101110;
assign LUT_4[5597] = 32'b11111111111111110011111101100110;
assign LUT_4[5598] = 32'b11111111111111111010001100010010;
assign LUT_4[5599] = 32'b11111111111111110011011000001010;
assign LUT_4[5600] = 32'b00000000000000000101001110010110;
assign LUT_4[5601] = 32'b11111111111111111110011010001110;
assign LUT_4[5602] = 32'b00000000000000000100101000111010;
assign LUT_4[5603] = 32'b11111111111111111101110100110010;
assign LUT_4[5604] = 32'b00000000000000000010001110110010;
assign LUT_4[5605] = 32'b11111111111111111011011010101010;
assign LUT_4[5606] = 32'b00000000000000000001101001010110;
assign LUT_4[5607] = 32'b11111111111111111010110101001110;
assign LUT_4[5608] = 32'b11111111111111111110011010101011;
assign LUT_4[5609] = 32'b11111111111111110111100110100011;
assign LUT_4[5610] = 32'b11111111111111111101110101001111;
assign LUT_4[5611] = 32'b11111111111111110111000001000111;
assign LUT_4[5612] = 32'b11111111111111111011011011000111;
assign LUT_4[5613] = 32'b11111111111111110100100110111111;
assign LUT_4[5614] = 32'b11111111111111111010110101101011;
assign LUT_4[5615] = 32'b11111111111111110100000001100011;
assign LUT_4[5616] = 32'b00000000000000000011000000000100;
assign LUT_4[5617] = 32'b11111111111111111100001011111100;
assign LUT_4[5618] = 32'b00000000000000000010011010101000;
assign LUT_4[5619] = 32'b11111111111111111011100110100000;
assign LUT_4[5620] = 32'b00000000000000000000000000100000;
assign LUT_4[5621] = 32'b11111111111111111001001100011000;
assign LUT_4[5622] = 32'b11111111111111111111011011000100;
assign LUT_4[5623] = 32'b11111111111111111000100110111100;
assign LUT_4[5624] = 32'b11111111111111111100001100011001;
assign LUT_4[5625] = 32'b11111111111111110101011000010001;
assign LUT_4[5626] = 32'b11111111111111111011100110111101;
assign LUT_4[5627] = 32'b11111111111111110100110010110101;
assign LUT_4[5628] = 32'b11111111111111111001001100110101;
assign LUT_4[5629] = 32'b11111111111111110010011000101101;
assign LUT_4[5630] = 32'b11111111111111111000100111011001;
assign LUT_4[5631] = 32'b11111111111111110001110011010001;
assign LUT_4[5632] = 32'b11111111111111111100111110011000;
assign LUT_4[5633] = 32'b11111111111111110110001010010000;
assign LUT_4[5634] = 32'b11111111111111111100011000111100;
assign LUT_4[5635] = 32'b11111111111111110101100100110100;
assign LUT_4[5636] = 32'b11111111111111111001111110110100;
assign LUT_4[5637] = 32'b11111111111111110011001010101100;
assign LUT_4[5638] = 32'b11111111111111111001011001011000;
assign LUT_4[5639] = 32'b11111111111111110010100101010000;
assign LUT_4[5640] = 32'b11111111111111110110001010101101;
assign LUT_4[5641] = 32'b11111111111111101111010110100101;
assign LUT_4[5642] = 32'b11111111111111110101100101010001;
assign LUT_4[5643] = 32'b11111111111111101110110001001001;
assign LUT_4[5644] = 32'b11111111111111110011001011001001;
assign LUT_4[5645] = 32'b11111111111111101100010111000001;
assign LUT_4[5646] = 32'b11111111111111110010100101101101;
assign LUT_4[5647] = 32'b11111111111111101011110001100101;
assign LUT_4[5648] = 32'b11111111111111111010110000000110;
assign LUT_4[5649] = 32'b11111111111111110011111011111110;
assign LUT_4[5650] = 32'b11111111111111111010001010101010;
assign LUT_4[5651] = 32'b11111111111111110011010110100010;
assign LUT_4[5652] = 32'b11111111111111110111110000100010;
assign LUT_4[5653] = 32'b11111111111111110000111100011010;
assign LUT_4[5654] = 32'b11111111111111110111001011000110;
assign LUT_4[5655] = 32'b11111111111111110000010110111110;
assign LUT_4[5656] = 32'b11111111111111110011111100011011;
assign LUT_4[5657] = 32'b11111111111111101101001000010011;
assign LUT_4[5658] = 32'b11111111111111110011010110111111;
assign LUT_4[5659] = 32'b11111111111111101100100010110111;
assign LUT_4[5660] = 32'b11111111111111110000111100110111;
assign LUT_4[5661] = 32'b11111111111111101010001000101111;
assign LUT_4[5662] = 32'b11111111111111110000010111011011;
assign LUT_4[5663] = 32'b11111111111111101001100011010011;
assign LUT_4[5664] = 32'b11111111111111111011011001011111;
assign LUT_4[5665] = 32'b11111111111111110100100101010111;
assign LUT_4[5666] = 32'b11111111111111111010110100000011;
assign LUT_4[5667] = 32'b11111111111111110011111111111011;
assign LUT_4[5668] = 32'b11111111111111111000011001111011;
assign LUT_4[5669] = 32'b11111111111111110001100101110011;
assign LUT_4[5670] = 32'b11111111111111110111110100011111;
assign LUT_4[5671] = 32'b11111111111111110001000000010111;
assign LUT_4[5672] = 32'b11111111111111110100100101110100;
assign LUT_4[5673] = 32'b11111111111111101101110001101100;
assign LUT_4[5674] = 32'b11111111111111110100000000011000;
assign LUT_4[5675] = 32'b11111111111111101101001100010000;
assign LUT_4[5676] = 32'b11111111111111110001100110010000;
assign LUT_4[5677] = 32'b11111111111111101010110010001000;
assign LUT_4[5678] = 32'b11111111111111110001000000110100;
assign LUT_4[5679] = 32'b11111111111111101010001100101100;
assign LUT_4[5680] = 32'b11111111111111111001001011001101;
assign LUT_4[5681] = 32'b11111111111111110010010111000101;
assign LUT_4[5682] = 32'b11111111111111111000100101110001;
assign LUT_4[5683] = 32'b11111111111111110001110001101001;
assign LUT_4[5684] = 32'b11111111111111110110001011101001;
assign LUT_4[5685] = 32'b11111111111111101111010111100001;
assign LUT_4[5686] = 32'b11111111111111110101100110001101;
assign LUT_4[5687] = 32'b11111111111111101110110010000101;
assign LUT_4[5688] = 32'b11111111111111110010010111100010;
assign LUT_4[5689] = 32'b11111111111111101011100011011010;
assign LUT_4[5690] = 32'b11111111111111110001110010000110;
assign LUT_4[5691] = 32'b11111111111111101010111101111110;
assign LUT_4[5692] = 32'b11111111111111101111010111111110;
assign LUT_4[5693] = 32'b11111111111111101000100011110110;
assign LUT_4[5694] = 32'b11111111111111101110110010100010;
assign LUT_4[5695] = 32'b11111111111111100111111110011010;
assign LUT_4[5696] = 32'b11111111111111111110010101101100;
assign LUT_4[5697] = 32'b11111111111111110111100001100100;
assign LUT_4[5698] = 32'b11111111111111111101110000010000;
assign LUT_4[5699] = 32'b11111111111111110110111100001000;
assign LUT_4[5700] = 32'b11111111111111111011010110001000;
assign LUT_4[5701] = 32'b11111111111111110100100010000000;
assign LUT_4[5702] = 32'b11111111111111111010110000101100;
assign LUT_4[5703] = 32'b11111111111111110011111100100100;
assign LUT_4[5704] = 32'b11111111111111110111100010000001;
assign LUT_4[5705] = 32'b11111111111111110000101101111001;
assign LUT_4[5706] = 32'b11111111111111110110111100100101;
assign LUT_4[5707] = 32'b11111111111111110000001000011101;
assign LUT_4[5708] = 32'b11111111111111110100100010011101;
assign LUT_4[5709] = 32'b11111111111111101101101110010101;
assign LUT_4[5710] = 32'b11111111111111110011111101000001;
assign LUT_4[5711] = 32'b11111111111111101101001000111001;
assign LUT_4[5712] = 32'b11111111111111111100000111011010;
assign LUT_4[5713] = 32'b11111111111111110101010011010010;
assign LUT_4[5714] = 32'b11111111111111111011100001111110;
assign LUT_4[5715] = 32'b11111111111111110100101101110110;
assign LUT_4[5716] = 32'b11111111111111111001000111110110;
assign LUT_4[5717] = 32'b11111111111111110010010011101110;
assign LUT_4[5718] = 32'b11111111111111111000100010011010;
assign LUT_4[5719] = 32'b11111111111111110001101110010010;
assign LUT_4[5720] = 32'b11111111111111110101010011101111;
assign LUT_4[5721] = 32'b11111111111111101110011111100111;
assign LUT_4[5722] = 32'b11111111111111110100101110010011;
assign LUT_4[5723] = 32'b11111111111111101101111010001011;
assign LUT_4[5724] = 32'b11111111111111110010010100001011;
assign LUT_4[5725] = 32'b11111111111111101011100000000011;
assign LUT_4[5726] = 32'b11111111111111110001101110101111;
assign LUT_4[5727] = 32'b11111111111111101010111010100111;
assign LUT_4[5728] = 32'b11111111111111111100110000110011;
assign LUT_4[5729] = 32'b11111111111111110101111100101011;
assign LUT_4[5730] = 32'b11111111111111111100001011010111;
assign LUT_4[5731] = 32'b11111111111111110101010111001111;
assign LUT_4[5732] = 32'b11111111111111111001110001001111;
assign LUT_4[5733] = 32'b11111111111111110010111101000111;
assign LUT_4[5734] = 32'b11111111111111111001001011110011;
assign LUT_4[5735] = 32'b11111111111111110010010111101011;
assign LUT_4[5736] = 32'b11111111111111110101111101001000;
assign LUT_4[5737] = 32'b11111111111111101111001001000000;
assign LUT_4[5738] = 32'b11111111111111110101010111101100;
assign LUT_4[5739] = 32'b11111111111111101110100011100100;
assign LUT_4[5740] = 32'b11111111111111110010111101100100;
assign LUT_4[5741] = 32'b11111111111111101100001001011100;
assign LUT_4[5742] = 32'b11111111111111110010011000001000;
assign LUT_4[5743] = 32'b11111111111111101011100100000000;
assign LUT_4[5744] = 32'b11111111111111111010100010100001;
assign LUT_4[5745] = 32'b11111111111111110011101110011001;
assign LUT_4[5746] = 32'b11111111111111111001111101000101;
assign LUT_4[5747] = 32'b11111111111111110011001000111101;
assign LUT_4[5748] = 32'b11111111111111110111100010111101;
assign LUT_4[5749] = 32'b11111111111111110000101110110101;
assign LUT_4[5750] = 32'b11111111111111110110111101100001;
assign LUT_4[5751] = 32'b11111111111111110000001001011001;
assign LUT_4[5752] = 32'b11111111111111110011101110110110;
assign LUT_4[5753] = 32'b11111111111111101100111010101110;
assign LUT_4[5754] = 32'b11111111111111110011001001011010;
assign LUT_4[5755] = 32'b11111111111111101100010101010010;
assign LUT_4[5756] = 32'b11111111111111110000101111010010;
assign LUT_4[5757] = 32'b11111111111111101001111011001010;
assign LUT_4[5758] = 32'b11111111111111110000001001110110;
assign LUT_4[5759] = 32'b11111111111111101001010101101110;
assign LUT_4[5760] = 32'b11111111111111111111100100100000;
assign LUT_4[5761] = 32'b11111111111111111000110000011000;
assign LUT_4[5762] = 32'b11111111111111111110111111000100;
assign LUT_4[5763] = 32'b11111111111111111000001010111100;
assign LUT_4[5764] = 32'b11111111111111111100100100111100;
assign LUT_4[5765] = 32'b11111111111111110101110000110100;
assign LUT_4[5766] = 32'b11111111111111111011111111100000;
assign LUT_4[5767] = 32'b11111111111111110101001011011000;
assign LUT_4[5768] = 32'b11111111111111111000110000110101;
assign LUT_4[5769] = 32'b11111111111111110001111100101101;
assign LUT_4[5770] = 32'b11111111111111111000001011011001;
assign LUT_4[5771] = 32'b11111111111111110001010111010001;
assign LUT_4[5772] = 32'b11111111111111110101110001010001;
assign LUT_4[5773] = 32'b11111111111111101110111101001001;
assign LUT_4[5774] = 32'b11111111111111110101001011110101;
assign LUT_4[5775] = 32'b11111111111111101110010111101101;
assign LUT_4[5776] = 32'b11111111111111111101010110001110;
assign LUT_4[5777] = 32'b11111111111111110110100010000110;
assign LUT_4[5778] = 32'b11111111111111111100110000110010;
assign LUT_4[5779] = 32'b11111111111111110101111100101010;
assign LUT_4[5780] = 32'b11111111111111111010010110101010;
assign LUT_4[5781] = 32'b11111111111111110011100010100010;
assign LUT_4[5782] = 32'b11111111111111111001110001001110;
assign LUT_4[5783] = 32'b11111111111111110010111101000110;
assign LUT_4[5784] = 32'b11111111111111110110100010100011;
assign LUT_4[5785] = 32'b11111111111111101111101110011011;
assign LUT_4[5786] = 32'b11111111111111110101111101000111;
assign LUT_4[5787] = 32'b11111111111111101111001000111111;
assign LUT_4[5788] = 32'b11111111111111110011100010111111;
assign LUT_4[5789] = 32'b11111111111111101100101110110111;
assign LUT_4[5790] = 32'b11111111111111110010111101100011;
assign LUT_4[5791] = 32'b11111111111111101100001001011011;
assign LUT_4[5792] = 32'b11111111111111111101111111100111;
assign LUT_4[5793] = 32'b11111111111111110111001011011111;
assign LUT_4[5794] = 32'b11111111111111111101011010001011;
assign LUT_4[5795] = 32'b11111111111111110110100110000011;
assign LUT_4[5796] = 32'b11111111111111111011000000000011;
assign LUT_4[5797] = 32'b11111111111111110100001011111011;
assign LUT_4[5798] = 32'b11111111111111111010011010100111;
assign LUT_4[5799] = 32'b11111111111111110011100110011111;
assign LUT_4[5800] = 32'b11111111111111110111001011111100;
assign LUT_4[5801] = 32'b11111111111111110000010111110100;
assign LUT_4[5802] = 32'b11111111111111110110100110100000;
assign LUT_4[5803] = 32'b11111111111111101111110010011000;
assign LUT_4[5804] = 32'b11111111111111110100001100011000;
assign LUT_4[5805] = 32'b11111111111111101101011000010000;
assign LUT_4[5806] = 32'b11111111111111110011100110111100;
assign LUT_4[5807] = 32'b11111111111111101100110010110100;
assign LUT_4[5808] = 32'b11111111111111111011110001010101;
assign LUT_4[5809] = 32'b11111111111111110100111101001101;
assign LUT_4[5810] = 32'b11111111111111111011001011111001;
assign LUT_4[5811] = 32'b11111111111111110100010111110001;
assign LUT_4[5812] = 32'b11111111111111111000110001110001;
assign LUT_4[5813] = 32'b11111111111111110001111101101001;
assign LUT_4[5814] = 32'b11111111111111111000001100010101;
assign LUT_4[5815] = 32'b11111111111111110001011000001101;
assign LUT_4[5816] = 32'b11111111111111110100111101101010;
assign LUT_4[5817] = 32'b11111111111111101110001001100010;
assign LUT_4[5818] = 32'b11111111111111110100011000001110;
assign LUT_4[5819] = 32'b11111111111111101101100100000110;
assign LUT_4[5820] = 32'b11111111111111110001111110000110;
assign LUT_4[5821] = 32'b11111111111111101011001001111110;
assign LUT_4[5822] = 32'b11111111111111110001011000101010;
assign LUT_4[5823] = 32'b11111111111111101010100100100010;
assign LUT_4[5824] = 32'b00000000000000000000111011110100;
assign LUT_4[5825] = 32'b11111111111111111010000111101100;
assign LUT_4[5826] = 32'b00000000000000000000010110011000;
assign LUT_4[5827] = 32'b11111111111111111001100010010000;
assign LUT_4[5828] = 32'b11111111111111111101111100010000;
assign LUT_4[5829] = 32'b11111111111111110111001000001000;
assign LUT_4[5830] = 32'b11111111111111111101010110110100;
assign LUT_4[5831] = 32'b11111111111111110110100010101100;
assign LUT_4[5832] = 32'b11111111111111111010001000001001;
assign LUT_4[5833] = 32'b11111111111111110011010100000001;
assign LUT_4[5834] = 32'b11111111111111111001100010101101;
assign LUT_4[5835] = 32'b11111111111111110010101110100101;
assign LUT_4[5836] = 32'b11111111111111110111001000100101;
assign LUT_4[5837] = 32'b11111111111111110000010100011101;
assign LUT_4[5838] = 32'b11111111111111110110100011001001;
assign LUT_4[5839] = 32'b11111111111111101111101111000001;
assign LUT_4[5840] = 32'b11111111111111111110101101100010;
assign LUT_4[5841] = 32'b11111111111111110111111001011010;
assign LUT_4[5842] = 32'b11111111111111111110001000000110;
assign LUT_4[5843] = 32'b11111111111111110111010011111110;
assign LUT_4[5844] = 32'b11111111111111111011101101111110;
assign LUT_4[5845] = 32'b11111111111111110100111001110110;
assign LUT_4[5846] = 32'b11111111111111111011001000100010;
assign LUT_4[5847] = 32'b11111111111111110100010100011010;
assign LUT_4[5848] = 32'b11111111111111110111111001110111;
assign LUT_4[5849] = 32'b11111111111111110001000101101111;
assign LUT_4[5850] = 32'b11111111111111110111010100011011;
assign LUT_4[5851] = 32'b11111111111111110000100000010011;
assign LUT_4[5852] = 32'b11111111111111110100111010010011;
assign LUT_4[5853] = 32'b11111111111111101110000110001011;
assign LUT_4[5854] = 32'b11111111111111110100010100110111;
assign LUT_4[5855] = 32'b11111111111111101101100000101111;
assign LUT_4[5856] = 32'b11111111111111111111010110111011;
assign LUT_4[5857] = 32'b11111111111111111000100010110011;
assign LUT_4[5858] = 32'b11111111111111111110110001011111;
assign LUT_4[5859] = 32'b11111111111111110111111101010111;
assign LUT_4[5860] = 32'b11111111111111111100010111010111;
assign LUT_4[5861] = 32'b11111111111111110101100011001111;
assign LUT_4[5862] = 32'b11111111111111111011110001111011;
assign LUT_4[5863] = 32'b11111111111111110100111101110011;
assign LUT_4[5864] = 32'b11111111111111111000100011010000;
assign LUT_4[5865] = 32'b11111111111111110001101111001000;
assign LUT_4[5866] = 32'b11111111111111110111111101110100;
assign LUT_4[5867] = 32'b11111111111111110001001001101100;
assign LUT_4[5868] = 32'b11111111111111110101100011101100;
assign LUT_4[5869] = 32'b11111111111111101110101111100100;
assign LUT_4[5870] = 32'b11111111111111110100111110010000;
assign LUT_4[5871] = 32'b11111111111111101110001010001000;
assign LUT_4[5872] = 32'b11111111111111111101001000101001;
assign LUT_4[5873] = 32'b11111111111111110110010100100001;
assign LUT_4[5874] = 32'b11111111111111111100100011001101;
assign LUT_4[5875] = 32'b11111111111111110101101111000101;
assign LUT_4[5876] = 32'b11111111111111111010001001000101;
assign LUT_4[5877] = 32'b11111111111111110011010100111101;
assign LUT_4[5878] = 32'b11111111111111111001100011101001;
assign LUT_4[5879] = 32'b11111111111111110010101111100001;
assign LUT_4[5880] = 32'b11111111111111110110010100111110;
assign LUT_4[5881] = 32'b11111111111111101111100000110110;
assign LUT_4[5882] = 32'b11111111111111110101101111100010;
assign LUT_4[5883] = 32'b11111111111111101110111011011010;
assign LUT_4[5884] = 32'b11111111111111110011010101011010;
assign LUT_4[5885] = 32'b11111111111111101100100001010010;
assign LUT_4[5886] = 32'b11111111111111110010101111111110;
assign LUT_4[5887] = 32'b11111111111111101011111011110110;
assign LUT_4[5888] = 32'b00000000000000000001111001111011;
assign LUT_4[5889] = 32'b11111111111111111011000101110011;
assign LUT_4[5890] = 32'b00000000000000000001010100011111;
assign LUT_4[5891] = 32'b11111111111111111010100000010111;
assign LUT_4[5892] = 32'b11111111111111111110111010010111;
assign LUT_4[5893] = 32'b11111111111111111000000110001111;
assign LUT_4[5894] = 32'b11111111111111111110010100111011;
assign LUT_4[5895] = 32'b11111111111111110111100000110011;
assign LUT_4[5896] = 32'b11111111111111111011000110010000;
assign LUT_4[5897] = 32'b11111111111111110100010010001000;
assign LUT_4[5898] = 32'b11111111111111111010100000110100;
assign LUT_4[5899] = 32'b11111111111111110011101100101100;
assign LUT_4[5900] = 32'b11111111111111111000000110101100;
assign LUT_4[5901] = 32'b11111111111111110001010010100100;
assign LUT_4[5902] = 32'b11111111111111110111100001010000;
assign LUT_4[5903] = 32'b11111111111111110000101101001000;
assign LUT_4[5904] = 32'b11111111111111111111101011101001;
assign LUT_4[5905] = 32'b11111111111111111000110111100001;
assign LUT_4[5906] = 32'b11111111111111111111000110001101;
assign LUT_4[5907] = 32'b11111111111111111000010010000101;
assign LUT_4[5908] = 32'b11111111111111111100101100000101;
assign LUT_4[5909] = 32'b11111111111111110101110111111101;
assign LUT_4[5910] = 32'b11111111111111111100000110101001;
assign LUT_4[5911] = 32'b11111111111111110101010010100001;
assign LUT_4[5912] = 32'b11111111111111111000110111111110;
assign LUT_4[5913] = 32'b11111111111111110010000011110110;
assign LUT_4[5914] = 32'b11111111111111111000010010100010;
assign LUT_4[5915] = 32'b11111111111111110001011110011010;
assign LUT_4[5916] = 32'b11111111111111110101111000011010;
assign LUT_4[5917] = 32'b11111111111111101111000100010010;
assign LUT_4[5918] = 32'b11111111111111110101010010111110;
assign LUT_4[5919] = 32'b11111111111111101110011110110110;
assign LUT_4[5920] = 32'b00000000000000000000010101000010;
assign LUT_4[5921] = 32'b11111111111111111001100000111010;
assign LUT_4[5922] = 32'b11111111111111111111101111100110;
assign LUT_4[5923] = 32'b11111111111111111000111011011110;
assign LUT_4[5924] = 32'b11111111111111111101010101011110;
assign LUT_4[5925] = 32'b11111111111111110110100001010110;
assign LUT_4[5926] = 32'b11111111111111111100110000000010;
assign LUT_4[5927] = 32'b11111111111111110101111011111010;
assign LUT_4[5928] = 32'b11111111111111111001100001010111;
assign LUT_4[5929] = 32'b11111111111111110010101101001111;
assign LUT_4[5930] = 32'b11111111111111111000111011111011;
assign LUT_4[5931] = 32'b11111111111111110010000111110011;
assign LUT_4[5932] = 32'b11111111111111110110100001110011;
assign LUT_4[5933] = 32'b11111111111111101111101101101011;
assign LUT_4[5934] = 32'b11111111111111110101111100010111;
assign LUT_4[5935] = 32'b11111111111111101111001000001111;
assign LUT_4[5936] = 32'b11111111111111111110000110110000;
assign LUT_4[5937] = 32'b11111111111111110111010010101000;
assign LUT_4[5938] = 32'b11111111111111111101100001010100;
assign LUT_4[5939] = 32'b11111111111111110110101101001100;
assign LUT_4[5940] = 32'b11111111111111111011000111001100;
assign LUT_4[5941] = 32'b11111111111111110100010011000100;
assign LUT_4[5942] = 32'b11111111111111111010100001110000;
assign LUT_4[5943] = 32'b11111111111111110011101101101000;
assign LUT_4[5944] = 32'b11111111111111110111010011000101;
assign LUT_4[5945] = 32'b11111111111111110000011110111101;
assign LUT_4[5946] = 32'b11111111111111110110101101101001;
assign LUT_4[5947] = 32'b11111111111111101111111001100001;
assign LUT_4[5948] = 32'b11111111111111110100010011100001;
assign LUT_4[5949] = 32'b11111111111111101101011111011001;
assign LUT_4[5950] = 32'b11111111111111110011101110000101;
assign LUT_4[5951] = 32'b11111111111111101100111001111101;
assign LUT_4[5952] = 32'b00000000000000000011010001001111;
assign LUT_4[5953] = 32'b11111111111111111100011101000111;
assign LUT_4[5954] = 32'b00000000000000000010101011110011;
assign LUT_4[5955] = 32'b11111111111111111011110111101011;
assign LUT_4[5956] = 32'b00000000000000000000010001101011;
assign LUT_4[5957] = 32'b11111111111111111001011101100011;
assign LUT_4[5958] = 32'b11111111111111111111101100001111;
assign LUT_4[5959] = 32'b11111111111111111000111000000111;
assign LUT_4[5960] = 32'b11111111111111111100011101100100;
assign LUT_4[5961] = 32'b11111111111111110101101001011100;
assign LUT_4[5962] = 32'b11111111111111111011111000001000;
assign LUT_4[5963] = 32'b11111111111111110101000100000000;
assign LUT_4[5964] = 32'b11111111111111111001011110000000;
assign LUT_4[5965] = 32'b11111111111111110010101001111000;
assign LUT_4[5966] = 32'b11111111111111111000111000100100;
assign LUT_4[5967] = 32'b11111111111111110010000100011100;
assign LUT_4[5968] = 32'b00000000000000000001000010111101;
assign LUT_4[5969] = 32'b11111111111111111010001110110101;
assign LUT_4[5970] = 32'b00000000000000000000011101100001;
assign LUT_4[5971] = 32'b11111111111111111001101001011001;
assign LUT_4[5972] = 32'b11111111111111111110000011011001;
assign LUT_4[5973] = 32'b11111111111111110111001111010001;
assign LUT_4[5974] = 32'b11111111111111111101011101111101;
assign LUT_4[5975] = 32'b11111111111111110110101001110101;
assign LUT_4[5976] = 32'b11111111111111111010001111010010;
assign LUT_4[5977] = 32'b11111111111111110011011011001010;
assign LUT_4[5978] = 32'b11111111111111111001101001110110;
assign LUT_4[5979] = 32'b11111111111111110010110101101110;
assign LUT_4[5980] = 32'b11111111111111110111001111101110;
assign LUT_4[5981] = 32'b11111111111111110000011011100110;
assign LUT_4[5982] = 32'b11111111111111110110101010010010;
assign LUT_4[5983] = 32'b11111111111111101111110110001010;
assign LUT_4[5984] = 32'b00000000000000000001101100010110;
assign LUT_4[5985] = 32'b11111111111111111010111000001110;
assign LUT_4[5986] = 32'b00000000000000000001000110111010;
assign LUT_4[5987] = 32'b11111111111111111010010010110010;
assign LUT_4[5988] = 32'b11111111111111111110101100110010;
assign LUT_4[5989] = 32'b11111111111111110111111000101010;
assign LUT_4[5990] = 32'b11111111111111111110000111010110;
assign LUT_4[5991] = 32'b11111111111111110111010011001110;
assign LUT_4[5992] = 32'b11111111111111111010111000101011;
assign LUT_4[5993] = 32'b11111111111111110100000100100011;
assign LUT_4[5994] = 32'b11111111111111111010010011001111;
assign LUT_4[5995] = 32'b11111111111111110011011111000111;
assign LUT_4[5996] = 32'b11111111111111110111111001000111;
assign LUT_4[5997] = 32'b11111111111111110001000100111111;
assign LUT_4[5998] = 32'b11111111111111110111010011101011;
assign LUT_4[5999] = 32'b11111111111111110000011111100011;
assign LUT_4[6000] = 32'b11111111111111111111011110000100;
assign LUT_4[6001] = 32'b11111111111111111000101001111100;
assign LUT_4[6002] = 32'b11111111111111111110111000101000;
assign LUT_4[6003] = 32'b11111111111111111000000100100000;
assign LUT_4[6004] = 32'b11111111111111111100011110100000;
assign LUT_4[6005] = 32'b11111111111111110101101010011000;
assign LUT_4[6006] = 32'b11111111111111111011111001000100;
assign LUT_4[6007] = 32'b11111111111111110101000100111100;
assign LUT_4[6008] = 32'b11111111111111111000101010011001;
assign LUT_4[6009] = 32'b11111111111111110001110110010001;
assign LUT_4[6010] = 32'b11111111111111111000000100111101;
assign LUT_4[6011] = 32'b11111111111111110001010000110101;
assign LUT_4[6012] = 32'b11111111111111110101101010110101;
assign LUT_4[6013] = 32'b11111111111111101110110110101101;
assign LUT_4[6014] = 32'b11111111111111110101000101011001;
assign LUT_4[6015] = 32'b11111111111111101110010001010001;
assign LUT_4[6016] = 32'b00000000000000000100100000000011;
assign LUT_4[6017] = 32'b11111111111111111101101011111011;
assign LUT_4[6018] = 32'b00000000000000000011111010100111;
assign LUT_4[6019] = 32'b11111111111111111101000110011111;
assign LUT_4[6020] = 32'b00000000000000000001100000011111;
assign LUT_4[6021] = 32'b11111111111111111010101100010111;
assign LUT_4[6022] = 32'b00000000000000000000111011000011;
assign LUT_4[6023] = 32'b11111111111111111010000110111011;
assign LUT_4[6024] = 32'b11111111111111111101101100011000;
assign LUT_4[6025] = 32'b11111111111111110110111000010000;
assign LUT_4[6026] = 32'b11111111111111111101000110111100;
assign LUT_4[6027] = 32'b11111111111111110110010010110100;
assign LUT_4[6028] = 32'b11111111111111111010101100110100;
assign LUT_4[6029] = 32'b11111111111111110011111000101100;
assign LUT_4[6030] = 32'b11111111111111111010000111011000;
assign LUT_4[6031] = 32'b11111111111111110011010011010000;
assign LUT_4[6032] = 32'b00000000000000000010010001110001;
assign LUT_4[6033] = 32'b11111111111111111011011101101001;
assign LUT_4[6034] = 32'b00000000000000000001101100010101;
assign LUT_4[6035] = 32'b11111111111111111010111000001101;
assign LUT_4[6036] = 32'b11111111111111111111010010001101;
assign LUT_4[6037] = 32'b11111111111111111000011110000101;
assign LUT_4[6038] = 32'b11111111111111111110101100110001;
assign LUT_4[6039] = 32'b11111111111111110111111000101001;
assign LUT_4[6040] = 32'b11111111111111111011011110000110;
assign LUT_4[6041] = 32'b11111111111111110100101001111110;
assign LUT_4[6042] = 32'b11111111111111111010111000101010;
assign LUT_4[6043] = 32'b11111111111111110100000100100010;
assign LUT_4[6044] = 32'b11111111111111111000011110100010;
assign LUT_4[6045] = 32'b11111111111111110001101010011010;
assign LUT_4[6046] = 32'b11111111111111110111111001000110;
assign LUT_4[6047] = 32'b11111111111111110001000100111110;
assign LUT_4[6048] = 32'b00000000000000000010111011001010;
assign LUT_4[6049] = 32'b11111111111111111100000111000010;
assign LUT_4[6050] = 32'b00000000000000000010010101101110;
assign LUT_4[6051] = 32'b11111111111111111011100001100110;
assign LUT_4[6052] = 32'b11111111111111111111111011100110;
assign LUT_4[6053] = 32'b11111111111111111001000111011110;
assign LUT_4[6054] = 32'b11111111111111111111010110001010;
assign LUT_4[6055] = 32'b11111111111111111000100010000010;
assign LUT_4[6056] = 32'b11111111111111111100000111011111;
assign LUT_4[6057] = 32'b11111111111111110101010011010111;
assign LUT_4[6058] = 32'b11111111111111111011100010000011;
assign LUT_4[6059] = 32'b11111111111111110100101101111011;
assign LUT_4[6060] = 32'b11111111111111111001000111111011;
assign LUT_4[6061] = 32'b11111111111111110010010011110011;
assign LUT_4[6062] = 32'b11111111111111111000100010011111;
assign LUT_4[6063] = 32'b11111111111111110001101110010111;
assign LUT_4[6064] = 32'b00000000000000000000101100111000;
assign LUT_4[6065] = 32'b11111111111111111001111000110000;
assign LUT_4[6066] = 32'b00000000000000000000000111011100;
assign LUT_4[6067] = 32'b11111111111111111001010011010100;
assign LUT_4[6068] = 32'b11111111111111111101101101010100;
assign LUT_4[6069] = 32'b11111111111111110110111001001100;
assign LUT_4[6070] = 32'b11111111111111111101000111111000;
assign LUT_4[6071] = 32'b11111111111111110110010011110000;
assign LUT_4[6072] = 32'b11111111111111111001111001001101;
assign LUT_4[6073] = 32'b11111111111111110011000101000101;
assign LUT_4[6074] = 32'b11111111111111111001010011110001;
assign LUT_4[6075] = 32'b11111111111111110010011111101001;
assign LUT_4[6076] = 32'b11111111111111110110111001101001;
assign LUT_4[6077] = 32'b11111111111111110000000101100001;
assign LUT_4[6078] = 32'b11111111111111110110010100001101;
assign LUT_4[6079] = 32'b11111111111111101111100000000101;
assign LUT_4[6080] = 32'b00000000000000000101110111010111;
assign LUT_4[6081] = 32'b11111111111111111111000011001111;
assign LUT_4[6082] = 32'b00000000000000000101010001111011;
assign LUT_4[6083] = 32'b11111111111111111110011101110011;
assign LUT_4[6084] = 32'b00000000000000000010110111110011;
assign LUT_4[6085] = 32'b11111111111111111100000011101011;
assign LUT_4[6086] = 32'b00000000000000000010010010010111;
assign LUT_4[6087] = 32'b11111111111111111011011110001111;
assign LUT_4[6088] = 32'b11111111111111111111000011101100;
assign LUT_4[6089] = 32'b11111111111111111000001111100100;
assign LUT_4[6090] = 32'b11111111111111111110011110010000;
assign LUT_4[6091] = 32'b11111111111111110111101010001000;
assign LUT_4[6092] = 32'b11111111111111111100000100001000;
assign LUT_4[6093] = 32'b11111111111111110101010000000000;
assign LUT_4[6094] = 32'b11111111111111111011011110101100;
assign LUT_4[6095] = 32'b11111111111111110100101010100100;
assign LUT_4[6096] = 32'b00000000000000000011101001000101;
assign LUT_4[6097] = 32'b11111111111111111100110100111101;
assign LUT_4[6098] = 32'b00000000000000000011000011101001;
assign LUT_4[6099] = 32'b11111111111111111100001111100001;
assign LUT_4[6100] = 32'b00000000000000000000101001100001;
assign LUT_4[6101] = 32'b11111111111111111001110101011001;
assign LUT_4[6102] = 32'b00000000000000000000000100000101;
assign LUT_4[6103] = 32'b11111111111111111001001111111101;
assign LUT_4[6104] = 32'b11111111111111111100110101011010;
assign LUT_4[6105] = 32'b11111111111111110110000001010010;
assign LUT_4[6106] = 32'b11111111111111111100001111111110;
assign LUT_4[6107] = 32'b11111111111111110101011011110110;
assign LUT_4[6108] = 32'b11111111111111111001110101110110;
assign LUT_4[6109] = 32'b11111111111111110011000001101110;
assign LUT_4[6110] = 32'b11111111111111111001010000011010;
assign LUT_4[6111] = 32'b11111111111111110010011100010010;
assign LUT_4[6112] = 32'b00000000000000000100010010011110;
assign LUT_4[6113] = 32'b11111111111111111101011110010110;
assign LUT_4[6114] = 32'b00000000000000000011101101000010;
assign LUT_4[6115] = 32'b11111111111111111100111000111010;
assign LUT_4[6116] = 32'b00000000000000000001010010111010;
assign LUT_4[6117] = 32'b11111111111111111010011110110010;
assign LUT_4[6118] = 32'b00000000000000000000101101011110;
assign LUT_4[6119] = 32'b11111111111111111001111001010110;
assign LUT_4[6120] = 32'b11111111111111111101011110110011;
assign LUT_4[6121] = 32'b11111111111111110110101010101011;
assign LUT_4[6122] = 32'b11111111111111111100111001010111;
assign LUT_4[6123] = 32'b11111111111111110110000101001111;
assign LUT_4[6124] = 32'b11111111111111111010011111001111;
assign LUT_4[6125] = 32'b11111111111111110011101011000111;
assign LUT_4[6126] = 32'b11111111111111111001111001110011;
assign LUT_4[6127] = 32'b11111111111111110011000101101011;
assign LUT_4[6128] = 32'b00000000000000000010000100001100;
assign LUT_4[6129] = 32'b11111111111111111011010000000100;
assign LUT_4[6130] = 32'b00000000000000000001011110110000;
assign LUT_4[6131] = 32'b11111111111111111010101010101000;
assign LUT_4[6132] = 32'b11111111111111111111000100101000;
assign LUT_4[6133] = 32'b11111111111111111000010000100000;
assign LUT_4[6134] = 32'b11111111111111111110011111001100;
assign LUT_4[6135] = 32'b11111111111111110111101011000100;
assign LUT_4[6136] = 32'b11111111111111111011010000100001;
assign LUT_4[6137] = 32'b11111111111111110100011100011001;
assign LUT_4[6138] = 32'b11111111111111111010101011000101;
assign LUT_4[6139] = 32'b11111111111111110011110110111101;
assign LUT_4[6140] = 32'b11111111111111111000010000111101;
assign LUT_4[6141] = 32'b11111111111111110001011100110101;
assign LUT_4[6142] = 32'b11111111111111110111101011100001;
assign LUT_4[6143] = 32'b11111111111111110000110111011001;
assign LUT_4[6144] = 32'b11111111111111110111101110111011;
assign LUT_4[6145] = 32'b11111111111111110000111010110011;
assign LUT_4[6146] = 32'b11111111111111110111001001011111;
assign LUT_4[6147] = 32'b11111111111111110000010101010111;
assign LUT_4[6148] = 32'b11111111111111110100101111010111;
assign LUT_4[6149] = 32'b11111111111111101101111011001111;
assign LUT_4[6150] = 32'b11111111111111110100001001111011;
assign LUT_4[6151] = 32'b11111111111111101101010101110011;
assign LUT_4[6152] = 32'b11111111111111110000111011010000;
assign LUT_4[6153] = 32'b11111111111111101010000111001000;
assign LUT_4[6154] = 32'b11111111111111110000010101110100;
assign LUT_4[6155] = 32'b11111111111111101001100001101100;
assign LUT_4[6156] = 32'b11111111111111101101111011101100;
assign LUT_4[6157] = 32'b11111111111111100111000111100100;
assign LUT_4[6158] = 32'b11111111111111101101010110010000;
assign LUT_4[6159] = 32'b11111111111111100110100010001000;
assign LUT_4[6160] = 32'b11111111111111110101100000101001;
assign LUT_4[6161] = 32'b11111111111111101110101100100001;
assign LUT_4[6162] = 32'b11111111111111110100111011001101;
assign LUT_4[6163] = 32'b11111111111111101110000111000101;
assign LUT_4[6164] = 32'b11111111111111110010100001000101;
assign LUT_4[6165] = 32'b11111111111111101011101100111101;
assign LUT_4[6166] = 32'b11111111111111110001111011101001;
assign LUT_4[6167] = 32'b11111111111111101011000111100001;
assign LUT_4[6168] = 32'b11111111111111101110101100111110;
assign LUT_4[6169] = 32'b11111111111111100111111000110110;
assign LUT_4[6170] = 32'b11111111111111101110000111100010;
assign LUT_4[6171] = 32'b11111111111111100111010011011010;
assign LUT_4[6172] = 32'b11111111111111101011101101011010;
assign LUT_4[6173] = 32'b11111111111111100100111001010010;
assign LUT_4[6174] = 32'b11111111111111101011000111111110;
assign LUT_4[6175] = 32'b11111111111111100100010011110110;
assign LUT_4[6176] = 32'b11111111111111110110001010000010;
assign LUT_4[6177] = 32'b11111111111111101111010101111010;
assign LUT_4[6178] = 32'b11111111111111110101100100100110;
assign LUT_4[6179] = 32'b11111111111111101110110000011110;
assign LUT_4[6180] = 32'b11111111111111110011001010011110;
assign LUT_4[6181] = 32'b11111111111111101100010110010110;
assign LUT_4[6182] = 32'b11111111111111110010100101000010;
assign LUT_4[6183] = 32'b11111111111111101011110000111010;
assign LUT_4[6184] = 32'b11111111111111101111010110010111;
assign LUT_4[6185] = 32'b11111111111111101000100010001111;
assign LUT_4[6186] = 32'b11111111111111101110110000111011;
assign LUT_4[6187] = 32'b11111111111111100111111100110011;
assign LUT_4[6188] = 32'b11111111111111101100010110110011;
assign LUT_4[6189] = 32'b11111111111111100101100010101011;
assign LUT_4[6190] = 32'b11111111111111101011110001010111;
assign LUT_4[6191] = 32'b11111111111111100100111101001111;
assign LUT_4[6192] = 32'b11111111111111110011111011110000;
assign LUT_4[6193] = 32'b11111111111111101101000111101000;
assign LUT_4[6194] = 32'b11111111111111110011010110010100;
assign LUT_4[6195] = 32'b11111111111111101100100010001100;
assign LUT_4[6196] = 32'b11111111111111110000111100001100;
assign LUT_4[6197] = 32'b11111111111111101010001000000100;
assign LUT_4[6198] = 32'b11111111111111110000010110110000;
assign LUT_4[6199] = 32'b11111111111111101001100010101000;
assign LUT_4[6200] = 32'b11111111111111101101001000000101;
assign LUT_4[6201] = 32'b11111111111111100110010011111101;
assign LUT_4[6202] = 32'b11111111111111101100100010101001;
assign LUT_4[6203] = 32'b11111111111111100101101110100001;
assign LUT_4[6204] = 32'b11111111111111101010001000100001;
assign LUT_4[6205] = 32'b11111111111111100011010100011001;
assign LUT_4[6206] = 32'b11111111111111101001100011000101;
assign LUT_4[6207] = 32'b11111111111111100010101110111101;
assign LUT_4[6208] = 32'b11111111111111111001000110001111;
assign LUT_4[6209] = 32'b11111111111111110010010010000111;
assign LUT_4[6210] = 32'b11111111111111111000100000110011;
assign LUT_4[6211] = 32'b11111111111111110001101100101011;
assign LUT_4[6212] = 32'b11111111111111110110000110101011;
assign LUT_4[6213] = 32'b11111111111111101111010010100011;
assign LUT_4[6214] = 32'b11111111111111110101100001001111;
assign LUT_4[6215] = 32'b11111111111111101110101101000111;
assign LUT_4[6216] = 32'b11111111111111110010010010100100;
assign LUT_4[6217] = 32'b11111111111111101011011110011100;
assign LUT_4[6218] = 32'b11111111111111110001101101001000;
assign LUT_4[6219] = 32'b11111111111111101010111001000000;
assign LUT_4[6220] = 32'b11111111111111101111010011000000;
assign LUT_4[6221] = 32'b11111111111111101000011110111000;
assign LUT_4[6222] = 32'b11111111111111101110101101100100;
assign LUT_4[6223] = 32'b11111111111111100111111001011100;
assign LUT_4[6224] = 32'b11111111111111110110110111111101;
assign LUT_4[6225] = 32'b11111111111111110000000011110101;
assign LUT_4[6226] = 32'b11111111111111110110010010100001;
assign LUT_4[6227] = 32'b11111111111111101111011110011001;
assign LUT_4[6228] = 32'b11111111111111110011111000011001;
assign LUT_4[6229] = 32'b11111111111111101101000100010001;
assign LUT_4[6230] = 32'b11111111111111110011010010111101;
assign LUT_4[6231] = 32'b11111111111111101100011110110101;
assign LUT_4[6232] = 32'b11111111111111110000000100010010;
assign LUT_4[6233] = 32'b11111111111111101001010000001010;
assign LUT_4[6234] = 32'b11111111111111101111011110110110;
assign LUT_4[6235] = 32'b11111111111111101000101010101110;
assign LUT_4[6236] = 32'b11111111111111101101000100101110;
assign LUT_4[6237] = 32'b11111111111111100110010000100110;
assign LUT_4[6238] = 32'b11111111111111101100011111010010;
assign LUT_4[6239] = 32'b11111111111111100101101011001010;
assign LUT_4[6240] = 32'b11111111111111110111100001010110;
assign LUT_4[6241] = 32'b11111111111111110000101101001110;
assign LUT_4[6242] = 32'b11111111111111110110111011111010;
assign LUT_4[6243] = 32'b11111111111111110000000111110010;
assign LUT_4[6244] = 32'b11111111111111110100100001110010;
assign LUT_4[6245] = 32'b11111111111111101101101101101010;
assign LUT_4[6246] = 32'b11111111111111110011111100010110;
assign LUT_4[6247] = 32'b11111111111111101101001000001110;
assign LUT_4[6248] = 32'b11111111111111110000101101101011;
assign LUT_4[6249] = 32'b11111111111111101001111001100011;
assign LUT_4[6250] = 32'b11111111111111110000001000001111;
assign LUT_4[6251] = 32'b11111111111111101001010100000111;
assign LUT_4[6252] = 32'b11111111111111101101101110000111;
assign LUT_4[6253] = 32'b11111111111111100110111001111111;
assign LUT_4[6254] = 32'b11111111111111101101001000101011;
assign LUT_4[6255] = 32'b11111111111111100110010100100011;
assign LUT_4[6256] = 32'b11111111111111110101010011000100;
assign LUT_4[6257] = 32'b11111111111111101110011110111100;
assign LUT_4[6258] = 32'b11111111111111110100101101101000;
assign LUT_4[6259] = 32'b11111111111111101101111001100000;
assign LUT_4[6260] = 32'b11111111111111110010010011100000;
assign LUT_4[6261] = 32'b11111111111111101011011111011000;
assign LUT_4[6262] = 32'b11111111111111110001101110000100;
assign LUT_4[6263] = 32'b11111111111111101010111001111100;
assign LUT_4[6264] = 32'b11111111111111101110011111011001;
assign LUT_4[6265] = 32'b11111111111111100111101011010001;
assign LUT_4[6266] = 32'b11111111111111101101111001111101;
assign LUT_4[6267] = 32'b11111111111111100111000101110101;
assign LUT_4[6268] = 32'b11111111111111101011011111110101;
assign LUT_4[6269] = 32'b11111111111111100100101011101101;
assign LUT_4[6270] = 32'b11111111111111101010111010011001;
assign LUT_4[6271] = 32'b11111111111111100100000110010001;
assign LUT_4[6272] = 32'b11111111111111111010010101000011;
assign LUT_4[6273] = 32'b11111111111111110011100000111011;
assign LUT_4[6274] = 32'b11111111111111111001101111100111;
assign LUT_4[6275] = 32'b11111111111111110010111011011111;
assign LUT_4[6276] = 32'b11111111111111110111010101011111;
assign LUT_4[6277] = 32'b11111111111111110000100001010111;
assign LUT_4[6278] = 32'b11111111111111110110110000000011;
assign LUT_4[6279] = 32'b11111111111111101111111011111011;
assign LUT_4[6280] = 32'b11111111111111110011100001011000;
assign LUT_4[6281] = 32'b11111111111111101100101101010000;
assign LUT_4[6282] = 32'b11111111111111110010111011111100;
assign LUT_4[6283] = 32'b11111111111111101100000111110100;
assign LUT_4[6284] = 32'b11111111111111110000100001110100;
assign LUT_4[6285] = 32'b11111111111111101001101101101100;
assign LUT_4[6286] = 32'b11111111111111101111111100011000;
assign LUT_4[6287] = 32'b11111111111111101001001000010000;
assign LUT_4[6288] = 32'b11111111111111111000000110110001;
assign LUT_4[6289] = 32'b11111111111111110001010010101001;
assign LUT_4[6290] = 32'b11111111111111110111100001010101;
assign LUT_4[6291] = 32'b11111111111111110000101101001101;
assign LUT_4[6292] = 32'b11111111111111110101000111001101;
assign LUT_4[6293] = 32'b11111111111111101110010011000101;
assign LUT_4[6294] = 32'b11111111111111110100100001110001;
assign LUT_4[6295] = 32'b11111111111111101101101101101001;
assign LUT_4[6296] = 32'b11111111111111110001010011000110;
assign LUT_4[6297] = 32'b11111111111111101010011110111110;
assign LUT_4[6298] = 32'b11111111111111110000101101101010;
assign LUT_4[6299] = 32'b11111111111111101001111001100010;
assign LUT_4[6300] = 32'b11111111111111101110010011100010;
assign LUT_4[6301] = 32'b11111111111111100111011111011010;
assign LUT_4[6302] = 32'b11111111111111101101101110000110;
assign LUT_4[6303] = 32'b11111111111111100110111001111110;
assign LUT_4[6304] = 32'b11111111111111111000110000001010;
assign LUT_4[6305] = 32'b11111111111111110001111100000010;
assign LUT_4[6306] = 32'b11111111111111111000001010101110;
assign LUT_4[6307] = 32'b11111111111111110001010110100110;
assign LUT_4[6308] = 32'b11111111111111110101110000100110;
assign LUT_4[6309] = 32'b11111111111111101110111100011110;
assign LUT_4[6310] = 32'b11111111111111110101001011001010;
assign LUT_4[6311] = 32'b11111111111111101110010111000010;
assign LUT_4[6312] = 32'b11111111111111110001111100011111;
assign LUT_4[6313] = 32'b11111111111111101011001000010111;
assign LUT_4[6314] = 32'b11111111111111110001010111000011;
assign LUT_4[6315] = 32'b11111111111111101010100010111011;
assign LUT_4[6316] = 32'b11111111111111101110111100111011;
assign LUT_4[6317] = 32'b11111111111111101000001000110011;
assign LUT_4[6318] = 32'b11111111111111101110010111011111;
assign LUT_4[6319] = 32'b11111111111111100111100011010111;
assign LUT_4[6320] = 32'b11111111111111110110100001111000;
assign LUT_4[6321] = 32'b11111111111111101111101101110000;
assign LUT_4[6322] = 32'b11111111111111110101111100011100;
assign LUT_4[6323] = 32'b11111111111111101111001000010100;
assign LUT_4[6324] = 32'b11111111111111110011100010010100;
assign LUT_4[6325] = 32'b11111111111111101100101110001100;
assign LUT_4[6326] = 32'b11111111111111110010111100111000;
assign LUT_4[6327] = 32'b11111111111111101100001000110000;
assign LUT_4[6328] = 32'b11111111111111101111101110001101;
assign LUT_4[6329] = 32'b11111111111111101000111010000101;
assign LUT_4[6330] = 32'b11111111111111101111001000110001;
assign LUT_4[6331] = 32'b11111111111111101000010100101001;
assign LUT_4[6332] = 32'b11111111111111101100101110101001;
assign LUT_4[6333] = 32'b11111111111111100101111010100001;
assign LUT_4[6334] = 32'b11111111111111101100001001001101;
assign LUT_4[6335] = 32'b11111111111111100101010101000101;
assign LUT_4[6336] = 32'b11111111111111111011101100010111;
assign LUT_4[6337] = 32'b11111111111111110100111000001111;
assign LUT_4[6338] = 32'b11111111111111111011000110111011;
assign LUT_4[6339] = 32'b11111111111111110100010010110011;
assign LUT_4[6340] = 32'b11111111111111111000101100110011;
assign LUT_4[6341] = 32'b11111111111111110001111000101011;
assign LUT_4[6342] = 32'b11111111111111111000000111010111;
assign LUT_4[6343] = 32'b11111111111111110001010011001111;
assign LUT_4[6344] = 32'b11111111111111110100111000101100;
assign LUT_4[6345] = 32'b11111111111111101110000100100100;
assign LUT_4[6346] = 32'b11111111111111110100010011010000;
assign LUT_4[6347] = 32'b11111111111111101101011111001000;
assign LUT_4[6348] = 32'b11111111111111110001111001001000;
assign LUT_4[6349] = 32'b11111111111111101011000101000000;
assign LUT_4[6350] = 32'b11111111111111110001010011101100;
assign LUT_4[6351] = 32'b11111111111111101010011111100100;
assign LUT_4[6352] = 32'b11111111111111111001011110000101;
assign LUT_4[6353] = 32'b11111111111111110010101001111101;
assign LUT_4[6354] = 32'b11111111111111111000111000101001;
assign LUT_4[6355] = 32'b11111111111111110010000100100001;
assign LUT_4[6356] = 32'b11111111111111110110011110100001;
assign LUT_4[6357] = 32'b11111111111111101111101010011001;
assign LUT_4[6358] = 32'b11111111111111110101111001000101;
assign LUT_4[6359] = 32'b11111111111111101111000100111101;
assign LUT_4[6360] = 32'b11111111111111110010101010011010;
assign LUT_4[6361] = 32'b11111111111111101011110110010010;
assign LUT_4[6362] = 32'b11111111111111110010000100111110;
assign LUT_4[6363] = 32'b11111111111111101011010000110110;
assign LUT_4[6364] = 32'b11111111111111101111101010110110;
assign LUT_4[6365] = 32'b11111111111111101000110110101110;
assign LUT_4[6366] = 32'b11111111111111101111000101011010;
assign LUT_4[6367] = 32'b11111111111111101000010001010010;
assign LUT_4[6368] = 32'b11111111111111111010000111011110;
assign LUT_4[6369] = 32'b11111111111111110011010011010110;
assign LUT_4[6370] = 32'b11111111111111111001100010000010;
assign LUT_4[6371] = 32'b11111111111111110010101101111010;
assign LUT_4[6372] = 32'b11111111111111110111000111111010;
assign LUT_4[6373] = 32'b11111111111111110000010011110010;
assign LUT_4[6374] = 32'b11111111111111110110100010011110;
assign LUT_4[6375] = 32'b11111111111111101111101110010110;
assign LUT_4[6376] = 32'b11111111111111110011010011110011;
assign LUT_4[6377] = 32'b11111111111111101100011111101011;
assign LUT_4[6378] = 32'b11111111111111110010101110010111;
assign LUT_4[6379] = 32'b11111111111111101011111010001111;
assign LUT_4[6380] = 32'b11111111111111110000010100001111;
assign LUT_4[6381] = 32'b11111111111111101001100000000111;
assign LUT_4[6382] = 32'b11111111111111101111101110110011;
assign LUT_4[6383] = 32'b11111111111111101000111010101011;
assign LUT_4[6384] = 32'b11111111111111110111111001001100;
assign LUT_4[6385] = 32'b11111111111111110001000101000100;
assign LUT_4[6386] = 32'b11111111111111110111010011110000;
assign LUT_4[6387] = 32'b11111111111111110000011111101000;
assign LUT_4[6388] = 32'b11111111111111110100111001101000;
assign LUT_4[6389] = 32'b11111111111111101110000101100000;
assign LUT_4[6390] = 32'b11111111111111110100010100001100;
assign LUT_4[6391] = 32'b11111111111111101101100000000100;
assign LUT_4[6392] = 32'b11111111111111110001000101100001;
assign LUT_4[6393] = 32'b11111111111111101010010001011001;
assign LUT_4[6394] = 32'b11111111111111110000100000000101;
assign LUT_4[6395] = 32'b11111111111111101001101011111101;
assign LUT_4[6396] = 32'b11111111111111101110000101111101;
assign LUT_4[6397] = 32'b11111111111111100111010001110101;
assign LUT_4[6398] = 32'b11111111111111101101100000100001;
assign LUT_4[6399] = 32'b11111111111111100110101100011001;
assign LUT_4[6400] = 32'b11111111111111111100101010011110;
assign LUT_4[6401] = 32'b11111111111111110101110110010110;
assign LUT_4[6402] = 32'b11111111111111111100000101000010;
assign LUT_4[6403] = 32'b11111111111111110101010000111010;
assign LUT_4[6404] = 32'b11111111111111111001101010111010;
assign LUT_4[6405] = 32'b11111111111111110010110110110010;
assign LUT_4[6406] = 32'b11111111111111111001000101011110;
assign LUT_4[6407] = 32'b11111111111111110010010001010110;
assign LUT_4[6408] = 32'b11111111111111110101110110110011;
assign LUT_4[6409] = 32'b11111111111111101111000010101011;
assign LUT_4[6410] = 32'b11111111111111110101010001010111;
assign LUT_4[6411] = 32'b11111111111111101110011101001111;
assign LUT_4[6412] = 32'b11111111111111110010110111001111;
assign LUT_4[6413] = 32'b11111111111111101100000011000111;
assign LUT_4[6414] = 32'b11111111111111110010010001110011;
assign LUT_4[6415] = 32'b11111111111111101011011101101011;
assign LUT_4[6416] = 32'b11111111111111111010011100001100;
assign LUT_4[6417] = 32'b11111111111111110011101000000100;
assign LUT_4[6418] = 32'b11111111111111111001110110110000;
assign LUT_4[6419] = 32'b11111111111111110011000010101000;
assign LUT_4[6420] = 32'b11111111111111110111011100101000;
assign LUT_4[6421] = 32'b11111111111111110000101000100000;
assign LUT_4[6422] = 32'b11111111111111110110110111001100;
assign LUT_4[6423] = 32'b11111111111111110000000011000100;
assign LUT_4[6424] = 32'b11111111111111110011101000100001;
assign LUT_4[6425] = 32'b11111111111111101100110100011001;
assign LUT_4[6426] = 32'b11111111111111110011000011000101;
assign LUT_4[6427] = 32'b11111111111111101100001110111101;
assign LUT_4[6428] = 32'b11111111111111110000101000111101;
assign LUT_4[6429] = 32'b11111111111111101001110100110101;
assign LUT_4[6430] = 32'b11111111111111110000000011100001;
assign LUT_4[6431] = 32'b11111111111111101001001111011001;
assign LUT_4[6432] = 32'b11111111111111111011000101100101;
assign LUT_4[6433] = 32'b11111111111111110100010001011101;
assign LUT_4[6434] = 32'b11111111111111111010100000001001;
assign LUT_4[6435] = 32'b11111111111111110011101100000001;
assign LUT_4[6436] = 32'b11111111111111111000000110000001;
assign LUT_4[6437] = 32'b11111111111111110001010001111001;
assign LUT_4[6438] = 32'b11111111111111110111100000100101;
assign LUT_4[6439] = 32'b11111111111111110000101100011101;
assign LUT_4[6440] = 32'b11111111111111110100010001111010;
assign LUT_4[6441] = 32'b11111111111111101101011101110010;
assign LUT_4[6442] = 32'b11111111111111110011101100011110;
assign LUT_4[6443] = 32'b11111111111111101100111000010110;
assign LUT_4[6444] = 32'b11111111111111110001010010010110;
assign LUT_4[6445] = 32'b11111111111111101010011110001110;
assign LUT_4[6446] = 32'b11111111111111110000101100111010;
assign LUT_4[6447] = 32'b11111111111111101001111000110010;
assign LUT_4[6448] = 32'b11111111111111111000110111010011;
assign LUT_4[6449] = 32'b11111111111111110010000011001011;
assign LUT_4[6450] = 32'b11111111111111111000010001110111;
assign LUT_4[6451] = 32'b11111111111111110001011101101111;
assign LUT_4[6452] = 32'b11111111111111110101110111101111;
assign LUT_4[6453] = 32'b11111111111111101111000011100111;
assign LUT_4[6454] = 32'b11111111111111110101010010010011;
assign LUT_4[6455] = 32'b11111111111111101110011110001011;
assign LUT_4[6456] = 32'b11111111111111110010000011101000;
assign LUT_4[6457] = 32'b11111111111111101011001111100000;
assign LUT_4[6458] = 32'b11111111111111110001011110001100;
assign LUT_4[6459] = 32'b11111111111111101010101010000100;
assign LUT_4[6460] = 32'b11111111111111101111000100000100;
assign LUT_4[6461] = 32'b11111111111111101000001111111100;
assign LUT_4[6462] = 32'b11111111111111101110011110101000;
assign LUT_4[6463] = 32'b11111111111111100111101010100000;
assign LUT_4[6464] = 32'b11111111111111111110000001110010;
assign LUT_4[6465] = 32'b11111111111111110111001101101010;
assign LUT_4[6466] = 32'b11111111111111111101011100010110;
assign LUT_4[6467] = 32'b11111111111111110110101000001110;
assign LUT_4[6468] = 32'b11111111111111111011000010001110;
assign LUT_4[6469] = 32'b11111111111111110100001110000110;
assign LUT_4[6470] = 32'b11111111111111111010011100110010;
assign LUT_4[6471] = 32'b11111111111111110011101000101010;
assign LUT_4[6472] = 32'b11111111111111110111001110000111;
assign LUT_4[6473] = 32'b11111111111111110000011001111111;
assign LUT_4[6474] = 32'b11111111111111110110101000101011;
assign LUT_4[6475] = 32'b11111111111111101111110100100011;
assign LUT_4[6476] = 32'b11111111111111110100001110100011;
assign LUT_4[6477] = 32'b11111111111111101101011010011011;
assign LUT_4[6478] = 32'b11111111111111110011101001000111;
assign LUT_4[6479] = 32'b11111111111111101100110100111111;
assign LUT_4[6480] = 32'b11111111111111111011110011100000;
assign LUT_4[6481] = 32'b11111111111111110100111111011000;
assign LUT_4[6482] = 32'b11111111111111111011001110000100;
assign LUT_4[6483] = 32'b11111111111111110100011001111100;
assign LUT_4[6484] = 32'b11111111111111111000110011111100;
assign LUT_4[6485] = 32'b11111111111111110001111111110100;
assign LUT_4[6486] = 32'b11111111111111111000001110100000;
assign LUT_4[6487] = 32'b11111111111111110001011010011000;
assign LUT_4[6488] = 32'b11111111111111110100111111110101;
assign LUT_4[6489] = 32'b11111111111111101110001011101101;
assign LUT_4[6490] = 32'b11111111111111110100011010011001;
assign LUT_4[6491] = 32'b11111111111111101101100110010001;
assign LUT_4[6492] = 32'b11111111111111110010000000010001;
assign LUT_4[6493] = 32'b11111111111111101011001100001001;
assign LUT_4[6494] = 32'b11111111111111110001011010110101;
assign LUT_4[6495] = 32'b11111111111111101010100110101101;
assign LUT_4[6496] = 32'b11111111111111111100011100111001;
assign LUT_4[6497] = 32'b11111111111111110101101000110001;
assign LUT_4[6498] = 32'b11111111111111111011110111011101;
assign LUT_4[6499] = 32'b11111111111111110101000011010101;
assign LUT_4[6500] = 32'b11111111111111111001011101010101;
assign LUT_4[6501] = 32'b11111111111111110010101001001101;
assign LUT_4[6502] = 32'b11111111111111111000110111111001;
assign LUT_4[6503] = 32'b11111111111111110010000011110001;
assign LUT_4[6504] = 32'b11111111111111110101101001001110;
assign LUT_4[6505] = 32'b11111111111111101110110101000110;
assign LUT_4[6506] = 32'b11111111111111110101000011110010;
assign LUT_4[6507] = 32'b11111111111111101110001111101010;
assign LUT_4[6508] = 32'b11111111111111110010101001101010;
assign LUT_4[6509] = 32'b11111111111111101011110101100010;
assign LUT_4[6510] = 32'b11111111111111110010000100001110;
assign LUT_4[6511] = 32'b11111111111111101011010000000110;
assign LUT_4[6512] = 32'b11111111111111111010001110100111;
assign LUT_4[6513] = 32'b11111111111111110011011010011111;
assign LUT_4[6514] = 32'b11111111111111111001101001001011;
assign LUT_4[6515] = 32'b11111111111111110010110101000011;
assign LUT_4[6516] = 32'b11111111111111110111001111000011;
assign LUT_4[6517] = 32'b11111111111111110000011010111011;
assign LUT_4[6518] = 32'b11111111111111110110101001100111;
assign LUT_4[6519] = 32'b11111111111111101111110101011111;
assign LUT_4[6520] = 32'b11111111111111110011011010111100;
assign LUT_4[6521] = 32'b11111111111111101100100110110100;
assign LUT_4[6522] = 32'b11111111111111110010110101100000;
assign LUT_4[6523] = 32'b11111111111111101100000001011000;
assign LUT_4[6524] = 32'b11111111111111110000011011011000;
assign LUT_4[6525] = 32'b11111111111111101001100111010000;
assign LUT_4[6526] = 32'b11111111111111101111110101111100;
assign LUT_4[6527] = 32'b11111111111111101001000001110100;
assign LUT_4[6528] = 32'b11111111111111111111010000100110;
assign LUT_4[6529] = 32'b11111111111111111000011100011110;
assign LUT_4[6530] = 32'b11111111111111111110101011001010;
assign LUT_4[6531] = 32'b11111111111111110111110111000010;
assign LUT_4[6532] = 32'b11111111111111111100010001000010;
assign LUT_4[6533] = 32'b11111111111111110101011100111010;
assign LUT_4[6534] = 32'b11111111111111111011101011100110;
assign LUT_4[6535] = 32'b11111111111111110100110111011110;
assign LUT_4[6536] = 32'b11111111111111111000011100111011;
assign LUT_4[6537] = 32'b11111111111111110001101000110011;
assign LUT_4[6538] = 32'b11111111111111110111110111011111;
assign LUT_4[6539] = 32'b11111111111111110001000011010111;
assign LUT_4[6540] = 32'b11111111111111110101011101010111;
assign LUT_4[6541] = 32'b11111111111111101110101001001111;
assign LUT_4[6542] = 32'b11111111111111110100110111111011;
assign LUT_4[6543] = 32'b11111111111111101110000011110011;
assign LUT_4[6544] = 32'b11111111111111111101000010010100;
assign LUT_4[6545] = 32'b11111111111111110110001110001100;
assign LUT_4[6546] = 32'b11111111111111111100011100111000;
assign LUT_4[6547] = 32'b11111111111111110101101000110000;
assign LUT_4[6548] = 32'b11111111111111111010000010110000;
assign LUT_4[6549] = 32'b11111111111111110011001110101000;
assign LUT_4[6550] = 32'b11111111111111111001011101010100;
assign LUT_4[6551] = 32'b11111111111111110010101001001100;
assign LUT_4[6552] = 32'b11111111111111110110001110101001;
assign LUT_4[6553] = 32'b11111111111111101111011010100001;
assign LUT_4[6554] = 32'b11111111111111110101101001001101;
assign LUT_4[6555] = 32'b11111111111111101110110101000101;
assign LUT_4[6556] = 32'b11111111111111110011001111000101;
assign LUT_4[6557] = 32'b11111111111111101100011010111101;
assign LUT_4[6558] = 32'b11111111111111110010101001101001;
assign LUT_4[6559] = 32'b11111111111111101011110101100001;
assign LUT_4[6560] = 32'b11111111111111111101101011101101;
assign LUT_4[6561] = 32'b11111111111111110110110111100101;
assign LUT_4[6562] = 32'b11111111111111111101000110010001;
assign LUT_4[6563] = 32'b11111111111111110110010010001001;
assign LUT_4[6564] = 32'b11111111111111111010101100001001;
assign LUT_4[6565] = 32'b11111111111111110011111000000001;
assign LUT_4[6566] = 32'b11111111111111111010000110101101;
assign LUT_4[6567] = 32'b11111111111111110011010010100101;
assign LUT_4[6568] = 32'b11111111111111110110111000000010;
assign LUT_4[6569] = 32'b11111111111111110000000011111010;
assign LUT_4[6570] = 32'b11111111111111110110010010100110;
assign LUT_4[6571] = 32'b11111111111111101111011110011110;
assign LUT_4[6572] = 32'b11111111111111110011111000011110;
assign LUT_4[6573] = 32'b11111111111111101101000100010110;
assign LUT_4[6574] = 32'b11111111111111110011010011000010;
assign LUT_4[6575] = 32'b11111111111111101100011110111010;
assign LUT_4[6576] = 32'b11111111111111111011011101011011;
assign LUT_4[6577] = 32'b11111111111111110100101001010011;
assign LUT_4[6578] = 32'b11111111111111111010110111111111;
assign LUT_4[6579] = 32'b11111111111111110100000011110111;
assign LUT_4[6580] = 32'b11111111111111111000011101110111;
assign LUT_4[6581] = 32'b11111111111111110001101001101111;
assign LUT_4[6582] = 32'b11111111111111110111111000011011;
assign LUT_4[6583] = 32'b11111111111111110001000100010011;
assign LUT_4[6584] = 32'b11111111111111110100101001110000;
assign LUT_4[6585] = 32'b11111111111111101101110101101000;
assign LUT_4[6586] = 32'b11111111111111110100000100010100;
assign LUT_4[6587] = 32'b11111111111111101101010000001100;
assign LUT_4[6588] = 32'b11111111111111110001101010001100;
assign LUT_4[6589] = 32'b11111111111111101010110110000100;
assign LUT_4[6590] = 32'b11111111111111110001000100110000;
assign LUT_4[6591] = 32'b11111111111111101010010000101000;
assign LUT_4[6592] = 32'b00000000000000000000100111111010;
assign LUT_4[6593] = 32'b11111111111111111001110011110010;
assign LUT_4[6594] = 32'b00000000000000000000000010011110;
assign LUT_4[6595] = 32'b11111111111111111001001110010110;
assign LUT_4[6596] = 32'b11111111111111111101101000010110;
assign LUT_4[6597] = 32'b11111111111111110110110100001110;
assign LUT_4[6598] = 32'b11111111111111111101000010111010;
assign LUT_4[6599] = 32'b11111111111111110110001110110010;
assign LUT_4[6600] = 32'b11111111111111111001110100001111;
assign LUT_4[6601] = 32'b11111111111111110011000000000111;
assign LUT_4[6602] = 32'b11111111111111111001001110110011;
assign LUT_4[6603] = 32'b11111111111111110010011010101011;
assign LUT_4[6604] = 32'b11111111111111110110110100101011;
assign LUT_4[6605] = 32'b11111111111111110000000000100011;
assign LUT_4[6606] = 32'b11111111111111110110001111001111;
assign LUT_4[6607] = 32'b11111111111111101111011011000111;
assign LUT_4[6608] = 32'b11111111111111111110011001101000;
assign LUT_4[6609] = 32'b11111111111111110111100101100000;
assign LUT_4[6610] = 32'b11111111111111111101110100001100;
assign LUT_4[6611] = 32'b11111111111111110111000000000100;
assign LUT_4[6612] = 32'b11111111111111111011011010000100;
assign LUT_4[6613] = 32'b11111111111111110100100101111100;
assign LUT_4[6614] = 32'b11111111111111111010110100101000;
assign LUT_4[6615] = 32'b11111111111111110100000000100000;
assign LUT_4[6616] = 32'b11111111111111110111100101111101;
assign LUT_4[6617] = 32'b11111111111111110000110001110101;
assign LUT_4[6618] = 32'b11111111111111110111000000100001;
assign LUT_4[6619] = 32'b11111111111111110000001100011001;
assign LUT_4[6620] = 32'b11111111111111110100100110011001;
assign LUT_4[6621] = 32'b11111111111111101101110010010001;
assign LUT_4[6622] = 32'b11111111111111110100000000111101;
assign LUT_4[6623] = 32'b11111111111111101101001100110101;
assign LUT_4[6624] = 32'b11111111111111111111000011000001;
assign LUT_4[6625] = 32'b11111111111111111000001110111001;
assign LUT_4[6626] = 32'b11111111111111111110011101100101;
assign LUT_4[6627] = 32'b11111111111111110111101001011101;
assign LUT_4[6628] = 32'b11111111111111111100000011011101;
assign LUT_4[6629] = 32'b11111111111111110101001111010101;
assign LUT_4[6630] = 32'b11111111111111111011011110000001;
assign LUT_4[6631] = 32'b11111111111111110100101001111001;
assign LUT_4[6632] = 32'b11111111111111111000001111010110;
assign LUT_4[6633] = 32'b11111111111111110001011011001110;
assign LUT_4[6634] = 32'b11111111111111110111101001111010;
assign LUT_4[6635] = 32'b11111111111111110000110101110010;
assign LUT_4[6636] = 32'b11111111111111110101001111110010;
assign LUT_4[6637] = 32'b11111111111111101110011011101010;
assign LUT_4[6638] = 32'b11111111111111110100101010010110;
assign LUT_4[6639] = 32'b11111111111111101101110110001110;
assign LUT_4[6640] = 32'b11111111111111111100110100101111;
assign LUT_4[6641] = 32'b11111111111111110110000000100111;
assign LUT_4[6642] = 32'b11111111111111111100001111010011;
assign LUT_4[6643] = 32'b11111111111111110101011011001011;
assign LUT_4[6644] = 32'b11111111111111111001110101001011;
assign LUT_4[6645] = 32'b11111111111111110011000001000011;
assign LUT_4[6646] = 32'b11111111111111111001001111101111;
assign LUT_4[6647] = 32'b11111111111111110010011011100111;
assign LUT_4[6648] = 32'b11111111111111110110000001000100;
assign LUT_4[6649] = 32'b11111111111111101111001100111100;
assign LUT_4[6650] = 32'b11111111111111110101011011101000;
assign LUT_4[6651] = 32'b11111111111111101110100111100000;
assign LUT_4[6652] = 32'b11111111111111110011000001100000;
assign LUT_4[6653] = 32'b11111111111111101100001101011000;
assign LUT_4[6654] = 32'b11111111111111110010011100000100;
assign LUT_4[6655] = 32'b11111111111111101011100111111100;
assign LUT_4[6656] = 32'b11111111111111110110110011000011;
assign LUT_4[6657] = 32'b11111111111111101111111110111011;
assign LUT_4[6658] = 32'b11111111111111110110001101100111;
assign LUT_4[6659] = 32'b11111111111111101111011001011111;
assign LUT_4[6660] = 32'b11111111111111110011110011011111;
assign LUT_4[6661] = 32'b11111111111111101100111111010111;
assign LUT_4[6662] = 32'b11111111111111110011001110000011;
assign LUT_4[6663] = 32'b11111111111111101100011001111011;
assign LUT_4[6664] = 32'b11111111111111101111111111011000;
assign LUT_4[6665] = 32'b11111111111111101001001011010000;
assign LUT_4[6666] = 32'b11111111111111101111011001111100;
assign LUT_4[6667] = 32'b11111111111111101000100101110100;
assign LUT_4[6668] = 32'b11111111111111101100111111110100;
assign LUT_4[6669] = 32'b11111111111111100110001011101100;
assign LUT_4[6670] = 32'b11111111111111101100011010011000;
assign LUT_4[6671] = 32'b11111111111111100101100110010000;
assign LUT_4[6672] = 32'b11111111111111110100100100110001;
assign LUT_4[6673] = 32'b11111111111111101101110000101001;
assign LUT_4[6674] = 32'b11111111111111110011111111010101;
assign LUT_4[6675] = 32'b11111111111111101101001011001101;
assign LUT_4[6676] = 32'b11111111111111110001100101001101;
assign LUT_4[6677] = 32'b11111111111111101010110001000101;
assign LUT_4[6678] = 32'b11111111111111110000111111110001;
assign LUT_4[6679] = 32'b11111111111111101010001011101001;
assign LUT_4[6680] = 32'b11111111111111101101110001000110;
assign LUT_4[6681] = 32'b11111111111111100110111100111110;
assign LUT_4[6682] = 32'b11111111111111101101001011101010;
assign LUT_4[6683] = 32'b11111111111111100110010111100010;
assign LUT_4[6684] = 32'b11111111111111101010110001100010;
assign LUT_4[6685] = 32'b11111111111111100011111101011010;
assign LUT_4[6686] = 32'b11111111111111101010001100000110;
assign LUT_4[6687] = 32'b11111111111111100011010111111110;
assign LUT_4[6688] = 32'b11111111111111110101001110001010;
assign LUT_4[6689] = 32'b11111111111111101110011010000010;
assign LUT_4[6690] = 32'b11111111111111110100101000101110;
assign LUT_4[6691] = 32'b11111111111111101101110100100110;
assign LUT_4[6692] = 32'b11111111111111110010001110100110;
assign LUT_4[6693] = 32'b11111111111111101011011010011110;
assign LUT_4[6694] = 32'b11111111111111110001101001001010;
assign LUT_4[6695] = 32'b11111111111111101010110101000010;
assign LUT_4[6696] = 32'b11111111111111101110011010011111;
assign LUT_4[6697] = 32'b11111111111111100111100110010111;
assign LUT_4[6698] = 32'b11111111111111101101110101000011;
assign LUT_4[6699] = 32'b11111111111111100111000000111011;
assign LUT_4[6700] = 32'b11111111111111101011011010111011;
assign LUT_4[6701] = 32'b11111111111111100100100110110011;
assign LUT_4[6702] = 32'b11111111111111101010110101011111;
assign LUT_4[6703] = 32'b11111111111111100100000001010111;
assign LUT_4[6704] = 32'b11111111111111110010111111111000;
assign LUT_4[6705] = 32'b11111111111111101100001011110000;
assign LUT_4[6706] = 32'b11111111111111110010011010011100;
assign LUT_4[6707] = 32'b11111111111111101011100110010100;
assign LUT_4[6708] = 32'b11111111111111110000000000010100;
assign LUT_4[6709] = 32'b11111111111111101001001100001100;
assign LUT_4[6710] = 32'b11111111111111101111011010111000;
assign LUT_4[6711] = 32'b11111111111111101000100110110000;
assign LUT_4[6712] = 32'b11111111111111101100001100001101;
assign LUT_4[6713] = 32'b11111111111111100101011000000101;
assign LUT_4[6714] = 32'b11111111111111101011100110110001;
assign LUT_4[6715] = 32'b11111111111111100100110010101001;
assign LUT_4[6716] = 32'b11111111111111101001001100101001;
assign LUT_4[6717] = 32'b11111111111111100010011000100001;
assign LUT_4[6718] = 32'b11111111111111101000100111001101;
assign LUT_4[6719] = 32'b11111111111111100001110011000101;
assign LUT_4[6720] = 32'b11111111111111111000001010010111;
assign LUT_4[6721] = 32'b11111111111111110001010110001111;
assign LUT_4[6722] = 32'b11111111111111110111100100111011;
assign LUT_4[6723] = 32'b11111111111111110000110000110011;
assign LUT_4[6724] = 32'b11111111111111110101001010110011;
assign LUT_4[6725] = 32'b11111111111111101110010110101011;
assign LUT_4[6726] = 32'b11111111111111110100100101010111;
assign LUT_4[6727] = 32'b11111111111111101101110001001111;
assign LUT_4[6728] = 32'b11111111111111110001010110101100;
assign LUT_4[6729] = 32'b11111111111111101010100010100100;
assign LUT_4[6730] = 32'b11111111111111110000110001010000;
assign LUT_4[6731] = 32'b11111111111111101001111101001000;
assign LUT_4[6732] = 32'b11111111111111101110010111001000;
assign LUT_4[6733] = 32'b11111111111111100111100011000000;
assign LUT_4[6734] = 32'b11111111111111101101110001101100;
assign LUT_4[6735] = 32'b11111111111111100110111101100100;
assign LUT_4[6736] = 32'b11111111111111110101111100000101;
assign LUT_4[6737] = 32'b11111111111111101111000111111101;
assign LUT_4[6738] = 32'b11111111111111110101010110101001;
assign LUT_4[6739] = 32'b11111111111111101110100010100001;
assign LUT_4[6740] = 32'b11111111111111110010111100100001;
assign LUT_4[6741] = 32'b11111111111111101100001000011001;
assign LUT_4[6742] = 32'b11111111111111110010010111000101;
assign LUT_4[6743] = 32'b11111111111111101011100010111101;
assign LUT_4[6744] = 32'b11111111111111101111001000011010;
assign LUT_4[6745] = 32'b11111111111111101000010100010010;
assign LUT_4[6746] = 32'b11111111111111101110100010111110;
assign LUT_4[6747] = 32'b11111111111111100111101110110110;
assign LUT_4[6748] = 32'b11111111111111101100001000110110;
assign LUT_4[6749] = 32'b11111111111111100101010100101110;
assign LUT_4[6750] = 32'b11111111111111101011100011011010;
assign LUT_4[6751] = 32'b11111111111111100100101111010010;
assign LUT_4[6752] = 32'b11111111111111110110100101011110;
assign LUT_4[6753] = 32'b11111111111111101111110001010110;
assign LUT_4[6754] = 32'b11111111111111110110000000000010;
assign LUT_4[6755] = 32'b11111111111111101111001011111010;
assign LUT_4[6756] = 32'b11111111111111110011100101111010;
assign LUT_4[6757] = 32'b11111111111111101100110001110010;
assign LUT_4[6758] = 32'b11111111111111110011000000011110;
assign LUT_4[6759] = 32'b11111111111111101100001100010110;
assign LUT_4[6760] = 32'b11111111111111101111110001110011;
assign LUT_4[6761] = 32'b11111111111111101000111101101011;
assign LUT_4[6762] = 32'b11111111111111101111001100010111;
assign LUT_4[6763] = 32'b11111111111111101000011000001111;
assign LUT_4[6764] = 32'b11111111111111101100110010001111;
assign LUT_4[6765] = 32'b11111111111111100101111110000111;
assign LUT_4[6766] = 32'b11111111111111101100001100110011;
assign LUT_4[6767] = 32'b11111111111111100101011000101011;
assign LUT_4[6768] = 32'b11111111111111110100010111001100;
assign LUT_4[6769] = 32'b11111111111111101101100011000100;
assign LUT_4[6770] = 32'b11111111111111110011110001110000;
assign LUT_4[6771] = 32'b11111111111111101100111101101000;
assign LUT_4[6772] = 32'b11111111111111110001010111101000;
assign LUT_4[6773] = 32'b11111111111111101010100011100000;
assign LUT_4[6774] = 32'b11111111111111110000110010001100;
assign LUT_4[6775] = 32'b11111111111111101001111110000100;
assign LUT_4[6776] = 32'b11111111111111101101100011100001;
assign LUT_4[6777] = 32'b11111111111111100110101111011001;
assign LUT_4[6778] = 32'b11111111111111101100111110000101;
assign LUT_4[6779] = 32'b11111111111111100110001001111101;
assign LUT_4[6780] = 32'b11111111111111101010100011111101;
assign LUT_4[6781] = 32'b11111111111111100011101111110101;
assign LUT_4[6782] = 32'b11111111111111101001111110100001;
assign LUT_4[6783] = 32'b11111111111111100011001010011001;
assign LUT_4[6784] = 32'b11111111111111111001011001001011;
assign LUT_4[6785] = 32'b11111111111111110010100101000011;
assign LUT_4[6786] = 32'b11111111111111111000110011101111;
assign LUT_4[6787] = 32'b11111111111111110001111111100111;
assign LUT_4[6788] = 32'b11111111111111110110011001100111;
assign LUT_4[6789] = 32'b11111111111111101111100101011111;
assign LUT_4[6790] = 32'b11111111111111110101110100001011;
assign LUT_4[6791] = 32'b11111111111111101111000000000011;
assign LUT_4[6792] = 32'b11111111111111110010100101100000;
assign LUT_4[6793] = 32'b11111111111111101011110001011000;
assign LUT_4[6794] = 32'b11111111111111110010000000000100;
assign LUT_4[6795] = 32'b11111111111111101011001011111100;
assign LUT_4[6796] = 32'b11111111111111101111100101111100;
assign LUT_4[6797] = 32'b11111111111111101000110001110100;
assign LUT_4[6798] = 32'b11111111111111101111000000100000;
assign LUT_4[6799] = 32'b11111111111111101000001100011000;
assign LUT_4[6800] = 32'b11111111111111110111001010111001;
assign LUT_4[6801] = 32'b11111111111111110000010110110001;
assign LUT_4[6802] = 32'b11111111111111110110100101011101;
assign LUT_4[6803] = 32'b11111111111111101111110001010101;
assign LUT_4[6804] = 32'b11111111111111110100001011010101;
assign LUT_4[6805] = 32'b11111111111111101101010111001101;
assign LUT_4[6806] = 32'b11111111111111110011100101111001;
assign LUT_4[6807] = 32'b11111111111111101100110001110001;
assign LUT_4[6808] = 32'b11111111111111110000010111001110;
assign LUT_4[6809] = 32'b11111111111111101001100011000110;
assign LUT_4[6810] = 32'b11111111111111101111110001110010;
assign LUT_4[6811] = 32'b11111111111111101000111101101010;
assign LUT_4[6812] = 32'b11111111111111101101010111101010;
assign LUT_4[6813] = 32'b11111111111111100110100011100010;
assign LUT_4[6814] = 32'b11111111111111101100110010001110;
assign LUT_4[6815] = 32'b11111111111111100101111110000110;
assign LUT_4[6816] = 32'b11111111111111110111110100010010;
assign LUT_4[6817] = 32'b11111111111111110001000000001010;
assign LUT_4[6818] = 32'b11111111111111110111001110110110;
assign LUT_4[6819] = 32'b11111111111111110000011010101110;
assign LUT_4[6820] = 32'b11111111111111110100110100101110;
assign LUT_4[6821] = 32'b11111111111111101110000000100110;
assign LUT_4[6822] = 32'b11111111111111110100001111010010;
assign LUT_4[6823] = 32'b11111111111111101101011011001010;
assign LUT_4[6824] = 32'b11111111111111110001000000100111;
assign LUT_4[6825] = 32'b11111111111111101010001100011111;
assign LUT_4[6826] = 32'b11111111111111110000011011001011;
assign LUT_4[6827] = 32'b11111111111111101001100111000011;
assign LUT_4[6828] = 32'b11111111111111101110000001000011;
assign LUT_4[6829] = 32'b11111111111111100111001100111011;
assign LUT_4[6830] = 32'b11111111111111101101011011100111;
assign LUT_4[6831] = 32'b11111111111111100110100111011111;
assign LUT_4[6832] = 32'b11111111111111110101100110000000;
assign LUT_4[6833] = 32'b11111111111111101110110001111000;
assign LUT_4[6834] = 32'b11111111111111110101000000100100;
assign LUT_4[6835] = 32'b11111111111111101110001100011100;
assign LUT_4[6836] = 32'b11111111111111110010100110011100;
assign LUT_4[6837] = 32'b11111111111111101011110010010100;
assign LUT_4[6838] = 32'b11111111111111110010000001000000;
assign LUT_4[6839] = 32'b11111111111111101011001100111000;
assign LUT_4[6840] = 32'b11111111111111101110110010010101;
assign LUT_4[6841] = 32'b11111111111111100111111110001101;
assign LUT_4[6842] = 32'b11111111111111101110001100111001;
assign LUT_4[6843] = 32'b11111111111111100111011000110001;
assign LUT_4[6844] = 32'b11111111111111101011110010110001;
assign LUT_4[6845] = 32'b11111111111111100100111110101001;
assign LUT_4[6846] = 32'b11111111111111101011001101010101;
assign LUT_4[6847] = 32'b11111111111111100100011001001101;
assign LUT_4[6848] = 32'b11111111111111111010110000011111;
assign LUT_4[6849] = 32'b11111111111111110011111100010111;
assign LUT_4[6850] = 32'b11111111111111111010001011000011;
assign LUT_4[6851] = 32'b11111111111111110011010110111011;
assign LUT_4[6852] = 32'b11111111111111110111110000111011;
assign LUT_4[6853] = 32'b11111111111111110000111100110011;
assign LUT_4[6854] = 32'b11111111111111110111001011011111;
assign LUT_4[6855] = 32'b11111111111111110000010111010111;
assign LUT_4[6856] = 32'b11111111111111110011111100110100;
assign LUT_4[6857] = 32'b11111111111111101101001000101100;
assign LUT_4[6858] = 32'b11111111111111110011010111011000;
assign LUT_4[6859] = 32'b11111111111111101100100011010000;
assign LUT_4[6860] = 32'b11111111111111110000111101010000;
assign LUT_4[6861] = 32'b11111111111111101010001001001000;
assign LUT_4[6862] = 32'b11111111111111110000010111110100;
assign LUT_4[6863] = 32'b11111111111111101001100011101100;
assign LUT_4[6864] = 32'b11111111111111111000100010001101;
assign LUT_4[6865] = 32'b11111111111111110001101110000101;
assign LUT_4[6866] = 32'b11111111111111110111111100110001;
assign LUT_4[6867] = 32'b11111111111111110001001000101001;
assign LUT_4[6868] = 32'b11111111111111110101100010101001;
assign LUT_4[6869] = 32'b11111111111111101110101110100001;
assign LUT_4[6870] = 32'b11111111111111110100111101001101;
assign LUT_4[6871] = 32'b11111111111111101110001001000101;
assign LUT_4[6872] = 32'b11111111111111110001101110100010;
assign LUT_4[6873] = 32'b11111111111111101010111010011010;
assign LUT_4[6874] = 32'b11111111111111110001001001000110;
assign LUT_4[6875] = 32'b11111111111111101010010100111110;
assign LUT_4[6876] = 32'b11111111111111101110101110111110;
assign LUT_4[6877] = 32'b11111111111111100111111010110110;
assign LUT_4[6878] = 32'b11111111111111101110001001100010;
assign LUT_4[6879] = 32'b11111111111111100111010101011010;
assign LUT_4[6880] = 32'b11111111111111111001001011100110;
assign LUT_4[6881] = 32'b11111111111111110010010111011110;
assign LUT_4[6882] = 32'b11111111111111111000100110001010;
assign LUT_4[6883] = 32'b11111111111111110001110010000010;
assign LUT_4[6884] = 32'b11111111111111110110001100000010;
assign LUT_4[6885] = 32'b11111111111111101111010111111010;
assign LUT_4[6886] = 32'b11111111111111110101100110100110;
assign LUT_4[6887] = 32'b11111111111111101110110010011110;
assign LUT_4[6888] = 32'b11111111111111110010010111111011;
assign LUT_4[6889] = 32'b11111111111111101011100011110011;
assign LUT_4[6890] = 32'b11111111111111110001110010011111;
assign LUT_4[6891] = 32'b11111111111111101010111110010111;
assign LUT_4[6892] = 32'b11111111111111101111011000010111;
assign LUT_4[6893] = 32'b11111111111111101000100100001111;
assign LUT_4[6894] = 32'b11111111111111101110110010111011;
assign LUT_4[6895] = 32'b11111111111111100111111110110011;
assign LUT_4[6896] = 32'b11111111111111110110111101010100;
assign LUT_4[6897] = 32'b11111111111111110000001001001100;
assign LUT_4[6898] = 32'b11111111111111110110010111111000;
assign LUT_4[6899] = 32'b11111111111111101111100011110000;
assign LUT_4[6900] = 32'b11111111111111110011111101110000;
assign LUT_4[6901] = 32'b11111111111111101101001001101000;
assign LUT_4[6902] = 32'b11111111111111110011011000010100;
assign LUT_4[6903] = 32'b11111111111111101100100100001100;
assign LUT_4[6904] = 32'b11111111111111110000001001101001;
assign LUT_4[6905] = 32'b11111111111111101001010101100001;
assign LUT_4[6906] = 32'b11111111111111101111100100001101;
assign LUT_4[6907] = 32'b11111111111111101000110000000101;
assign LUT_4[6908] = 32'b11111111111111101101001010000101;
assign LUT_4[6909] = 32'b11111111111111100110010101111101;
assign LUT_4[6910] = 32'b11111111111111101100100100101001;
assign LUT_4[6911] = 32'b11111111111111100101110000100001;
assign LUT_4[6912] = 32'b11111111111111111011101110100110;
assign LUT_4[6913] = 32'b11111111111111110100111010011110;
assign LUT_4[6914] = 32'b11111111111111111011001001001010;
assign LUT_4[6915] = 32'b11111111111111110100010101000010;
assign LUT_4[6916] = 32'b11111111111111111000101111000010;
assign LUT_4[6917] = 32'b11111111111111110001111010111010;
assign LUT_4[6918] = 32'b11111111111111111000001001100110;
assign LUT_4[6919] = 32'b11111111111111110001010101011110;
assign LUT_4[6920] = 32'b11111111111111110100111010111011;
assign LUT_4[6921] = 32'b11111111111111101110000110110011;
assign LUT_4[6922] = 32'b11111111111111110100010101011111;
assign LUT_4[6923] = 32'b11111111111111101101100001010111;
assign LUT_4[6924] = 32'b11111111111111110001111011010111;
assign LUT_4[6925] = 32'b11111111111111101011000111001111;
assign LUT_4[6926] = 32'b11111111111111110001010101111011;
assign LUT_4[6927] = 32'b11111111111111101010100001110011;
assign LUT_4[6928] = 32'b11111111111111111001100000010100;
assign LUT_4[6929] = 32'b11111111111111110010101100001100;
assign LUT_4[6930] = 32'b11111111111111111000111010111000;
assign LUT_4[6931] = 32'b11111111111111110010000110110000;
assign LUT_4[6932] = 32'b11111111111111110110100000110000;
assign LUT_4[6933] = 32'b11111111111111101111101100101000;
assign LUT_4[6934] = 32'b11111111111111110101111011010100;
assign LUT_4[6935] = 32'b11111111111111101111000111001100;
assign LUT_4[6936] = 32'b11111111111111110010101100101001;
assign LUT_4[6937] = 32'b11111111111111101011111000100001;
assign LUT_4[6938] = 32'b11111111111111110010000111001101;
assign LUT_4[6939] = 32'b11111111111111101011010011000101;
assign LUT_4[6940] = 32'b11111111111111101111101101000101;
assign LUT_4[6941] = 32'b11111111111111101000111000111101;
assign LUT_4[6942] = 32'b11111111111111101111000111101001;
assign LUT_4[6943] = 32'b11111111111111101000010011100001;
assign LUT_4[6944] = 32'b11111111111111111010001001101101;
assign LUT_4[6945] = 32'b11111111111111110011010101100101;
assign LUT_4[6946] = 32'b11111111111111111001100100010001;
assign LUT_4[6947] = 32'b11111111111111110010110000001001;
assign LUT_4[6948] = 32'b11111111111111110111001010001001;
assign LUT_4[6949] = 32'b11111111111111110000010110000001;
assign LUT_4[6950] = 32'b11111111111111110110100100101101;
assign LUT_4[6951] = 32'b11111111111111101111110000100101;
assign LUT_4[6952] = 32'b11111111111111110011010110000010;
assign LUT_4[6953] = 32'b11111111111111101100100001111010;
assign LUT_4[6954] = 32'b11111111111111110010110000100110;
assign LUT_4[6955] = 32'b11111111111111101011111100011110;
assign LUT_4[6956] = 32'b11111111111111110000010110011110;
assign LUT_4[6957] = 32'b11111111111111101001100010010110;
assign LUT_4[6958] = 32'b11111111111111101111110001000010;
assign LUT_4[6959] = 32'b11111111111111101000111100111010;
assign LUT_4[6960] = 32'b11111111111111110111111011011011;
assign LUT_4[6961] = 32'b11111111111111110001000111010011;
assign LUT_4[6962] = 32'b11111111111111110111010101111111;
assign LUT_4[6963] = 32'b11111111111111110000100001110111;
assign LUT_4[6964] = 32'b11111111111111110100111011110111;
assign LUT_4[6965] = 32'b11111111111111101110000111101111;
assign LUT_4[6966] = 32'b11111111111111110100010110011011;
assign LUT_4[6967] = 32'b11111111111111101101100010010011;
assign LUT_4[6968] = 32'b11111111111111110001000111110000;
assign LUT_4[6969] = 32'b11111111111111101010010011101000;
assign LUT_4[6970] = 32'b11111111111111110000100010010100;
assign LUT_4[6971] = 32'b11111111111111101001101110001100;
assign LUT_4[6972] = 32'b11111111111111101110001000001100;
assign LUT_4[6973] = 32'b11111111111111100111010100000100;
assign LUT_4[6974] = 32'b11111111111111101101100010110000;
assign LUT_4[6975] = 32'b11111111111111100110101110101000;
assign LUT_4[6976] = 32'b11111111111111111101000101111010;
assign LUT_4[6977] = 32'b11111111111111110110010001110010;
assign LUT_4[6978] = 32'b11111111111111111100100000011110;
assign LUT_4[6979] = 32'b11111111111111110101101100010110;
assign LUT_4[6980] = 32'b11111111111111111010000110010110;
assign LUT_4[6981] = 32'b11111111111111110011010010001110;
assign LUT_4[6982] = 32'b11111111111111111001100000111010;
assign LUT_4[6983] = 32'b11111111111111110010101100110010;
assign LUT_4[6984] = 32'b11111111111111110110010010001111;
assign LUT_4[6985] = 32'b11111111111111101111011110000111;
assign LUT_4[6986] = 32'b11111111111111110101101100110011;
assign LUT_4[6987] = 32'b11111111111111101110111000101011;
assign LUT_4[6988] = 32'b11111111111111110011010010101011;
assign LUT_4[6989] = 32'b11111111111111101100011110100011;
assign LUT_4[6990] = 32'b11111111111111110010101101001111;
assign LUT_4[6991] = 32'b11111111111111101011111001000111;
assign LUT_4[6992] = 32'b11111111111111111010110111101000;
assign LUT_4[6993] = 32'b11111111111111110100000011100000;
assign LUT_4[6994] = 32'b11111111111111111010010010001100;
assign LUT_4[6995] = 32'b11111111111111110011011110000100;
assign LUT_4[6996] = 32'b11111111111111110111111000000100;
assign LUT_4[6997] = 32'b11111111111111110001000011111100;
assign LUT_4[6998] = 32'b11111111111111110111010010101000;
assign LUT_4[6999] = 32'b11111111111111110000011110100000;
assign LUT_4[7000] = 32'b11111111111111110100000011111101;
assign LUT_4[7001] = 32'b11111111111111101101001111110101;
assign LUT_4[7002] = 32'b11111111111111110011011110100001;
assign LUT_4[7003] = 32'b11111111111111101100101010011001;
assign LUT_4[7004] = 32'b11111111111111110001000100011001;
assign LUT_4[7005] = 32'b11111111111111101010010000010001;
assign LUT_4[7006] = 32'b11111111111111110000011110111101;
assign LUT_4[7007] = 32'b11111111111111101001101010110101;
assign LUT_4[7008] = 32'b11111111111111111011100001000001;
assign LUT_4[7009] = 32'b11111111111111110100101100111001;
assign LUT_4[7010] = 32'b11111111111111111010111011100101;
assign LUT_4[7011] = 32'b11111111111111110100000111011101;
assign LUT_4[7012] = 32'b11111111111111111000100001011101;
assign LUT_4[7013] = 32'b11111111111111110001101101010101;
assign LUT_4[7014] = 32'b11111111111111110111111100000001;
assign LUT_4[7015] = 32'b11111111111111110001000111111001;
assign LUT_4[7016] = 32'b11111111111111110100101101010110;
assign LUT_4[7017] = 32'b11111111111111101101111001001110;
assign LUT_4[7018] = 32'b11111111111111110100000111111010;
assign LUT_4[7019] = 32'b11111111111111101101010011110010;
assign LUT_4[7020] = 32'b11111111111111110001101101110010;
assign LUT_4[7021] = 32'b11111111111111101010111001101010;
assign LUT_4[7022] = 32'b11111111111111110001001000010110;
assign LUT_4[7023] = 32'b11111111111111101010010100001110;
assign LUT_4[7024] = 32'b11111111111111111001010010101111;
assign LUT_4[7025] = 32'b11111111111111110010011110100111;
assign LUT_4[7026] = 32'b11111111111111111000101101010011;
assign LUT_4[7027] = 32'b11111111111111110001111001001011;
assign LUT_4[7028] = 32'b11111111111111110110010011001011;
assign LUT_4[7029] = 32'b11111111111111101111011111000011;
assign LUT_4[7030] = 32'b11111111111111110101101101101111;
assign LUT_4[7031] = 32'b11111111111111101110111001100111;
assign LUT_4[7032] = 32'b11111111111111110010011111000100;
assign LUT_4[7033] = 32'b11111111111111101011101010111100;
assign LUT_4[7034] = 32'b11111111111111110001111001101000;
assign LUT_4[7035] = 32'b11111111111111101011000101100000;
assign LUT_4[7036] = 32'b11111111111111101111011111100000;
assign LUT_4[7037] = 32'b11111111111111101000101011011000;
assign LUT_4[7038] = 32'b11111111111111101110111010000100;
assign LUT_4[7039] = 32'b11111111111111101000000101111100;
assign LUT_4[7040] = 32'b11111111111111111110010100101110;
assign LUT_4[7041] = 32'b11111111111111110111100000100110;
assign LUT_4[7042] = 32'b11111111111111111101101111010010;
assign LUT_4[7043] = 32'b11111111111111110110111011001010;
assign LUT_4[7044] = 32'b11111111111111111011010101001010;
assign LUT_4[7045] = 32'b11111111111111110100100001000010;
assign LUT_4[7046] = 32'b11111111111111111010101111101110;
assign LUT_4[7047] = 32'b11111111111111110011111011100110;
assign LUT_4[7048] = 32'b11111111111111110111100001000011;
assign LUT_4[7049] = 32'b11111111111111110000101100111011;
assign LUT_4[7050] = 32'b11111111111111110110111011100111;
assign LUT_4[7051] = 32'b11111111111111110000000111011111;
assign LUT_4[7052] = 32'b11111111111111110100100001011111;
assign LUT_4[7053] = 32'b11111111111111101101101101010111;
assign LUT_4[7054] = 32'b11111111111111110011111100000011;
assign LUT_4[7055] = 32'b11111111111111101101000111111011;
assign LUT_4[7056] = 32'b11111111111111111100000110011100;
assign LUT_4[7057] = 32'b11111111111111110101010010010100;
assign LUT_4[7058] = 32'b11111111111111111011100001000000;
assign LUT_4[7059] = 32'b11111111111111110100101100111000;
assign LUT_4[7060] = 32'b11111111111111111001000110111000;
assign LUT_4[7061] = 32'b11111111111111110010010010110000;
assign LUT_4[7062] = 32'b11111111111111111000100001011100;
assign LUT_4[7063] = 32'b11111111111111110001101101010100;
assign LUT_4[7064] = 32'b11111111111111110101010010110001;
assign LUT_4[7065] = 32'b11111111111111101110011110101001;
assign LUT_4[7066] = 32'b11111111111111110100101101010101;
assign LUT_4[7067] = 32'b11111111111111101101111001001101;
assign LUT_4[7068] = 32'b11111111111111110010010011001101;
assign LUT_4[7069] = 32'b11111111111111101011011111000101;
assign LUT_4[7070] = 32'b11111111111111110001101101110001;
assign LUT_4[7071] = 32'b11111111111111101010111001101001;
assign LUT_4[7072] = 32'b11111111111111111100101111110101;
assign LUT_4[7073] = 32'b11111111111111110101111011101101;
assign LUT_4[7074] = 32'b11111111111111111100001010011001;
assign LUT_4[7075] = 32'b11111111111111110101010110010001;
assign LUT_4[7076] = 32'b11111111111111111001110000010001;
assign LUT_4[7077] = 32'b11111111111111110010111100001001;
assign LUT_4[7078] = 32'b11111111111111111001001010110101;
assign LUT_4[7079] = 32'b11111111111111110010010110101101;
assign LUT_4[7080] = 32'b11111111111111110101111100001010;
assign LUT_4[7081] = 32'b11111111111111101111001000000010;
assign LUT_4[7082] = 32'b11111111111111110101010110101110;
assign LUT_4[7083] = 32'b11111111111111101110100010100110;
assign LUT_4[7084] = 32'b11111111111111110010111100100110;
assign LUT_4[7085] = 32'b11111111111111101100001000011110;
assign LUT_4[7086] = 32'b11111111111111110010010111001010;
assign LUT_4[7087] = 32'b11111111111111101011100011000010;
assign LUT_4[7088] = 32'b11111111111111111010100001100011;
assign LUT_4[7089] = 32'b11111111111111110011101101011011;
assign LUT_4[7090] = 32'b11111111111111111001111100000111;
assign LUT_4[7091] = 32'b11111111111111110011000111111111;
assign LUT_4[7092] = 32'b11111111111111110111100001111111;
assign LUT_4[7093] = 32'b11111111111111110000101101110111;
assign LUT_4[7094] = 32'b11111111111111110110111100100011;
assign LUT_4[7095] = 32'b11111111111111110000001000011011;
assign LUT_4[7096] = 32'b11111111111111110011101101111000;
assign LUT_4[7097] = 32'b11111111111111101100111001110000;
assign LUT_4[7098] = 32'b11111111111111110011001000011100;
assign LUT_4[7099] = 32'b11111111111111101100010100010100;
assign LUT_4[7100] = 32'b11111111111111110000101110010100;
assign LUT_4[7101] = 32'b11111111111111101001111010001100;
assign LUT_4[7102] = 32'b11111111111111110000001000111000;
assign LUT_4[7103] = 32'b11111111111111101001010100110000;
assign LUT_4[7104] = 32'b11111111111111111111101100000010;
assign LUT_4[7105] = 32'b11111111111111111000110111111010;
assign LUT_4[7106] = 32'b11111111111111111111000110100110;
assign LUT_4[7107] = 32'b11111111111111111000010010011110;
assign LUT_4[7108] = 32'b11111111111111111100101100011110;
assign LUT_4[7109] = 32'b11111111111111110101111000010110;
assign LUT_4[7110] = 32'b11111111111111111100000111000010;
assign LUT_4[7111] = 32'b11111111111111110101010010111010;
assign LUT_4[7112] = 32'b11111111111111111000111000010111;
assign LUT_4[7113] = 32'b11111111111111110010000100001111;
assign LUT_4[7114] = 32'b11111111111111111000010010111011;
assign LUT_4[7115] = 32'b11111111111111110001011110110011;
assign LUT_4[7116] = 32'b11111111111111110101111000110011;
assign LUT_4[7117] = 32'b11111111111111101111000100101011;
assign LUT_4[7118] = 32'b11111111111111110101010011010111;
assign LUT_4[7119] = 32'b11111111111111101110011111001111;
assign LUT_4[7120] = 32'b11111111111111111101011101110000;
assign LUT_4[7121] = 32'b11111111111111110110101001101000;
assign LUT_4[7122] = 32'b11111111111111111100111000010100;
assign LUT_4[7123] = 32'b11111111111111110110000100001100;
assign LUT_4[7124] = 32'b11111111111111111010011110001100;
assign LUT_4[7125] = 32'b11111111111111110011101010000100;
assign LUT_4[7126] = 32'b11111111111111111001111000110000;
assign LUT_4[7127] = 32'b11111111111111110011000100101000;
assign LUT_4[7128] = 32'b11111111111111110110101010000101;
assign LUT_4[7129] = 32'b11111111111111101111110101111101;
assign LUT_4[7130] = 32'b11111111111111110110000100101001;
assign LUT_4[7131] = 32'b11111111111111101111010000100001;
assign LUT_4[7132] = 32'b11111111111111110011101010100001;
assign LUT_4[7133] = 32'b11111111111111101100110110011001;
assign LUT_4[7134] = 32'b11111111111111110011000101000101;
assign LUT_4[7135] = 32'b11111111111111101100010000111101;
assign LUT_4[7136] = 32'b11111111111111111110000111001001;
assign LUT_4[7137] = 32'b11111111111111110111010011000001;
assign LUT_4[7138] = 32'b11111111111111111101100001101101;
assign LUT_4[7139] = 32'b11111111111111110110101101100101;
assign LUT_4[7140] = 32'b11111111111111111011000111100101;
assign LUT_4[7141] = 32'b11111111111111110100010011011101;
assign LUT_4[7142] = 32'b11111111111111111010100010001001;
assign LUT_4[7143] = 32'b11111111111111110011101110000001;
assign LUT_4[7144] = 32'b11111111111111110111010011011110;
assign LUT_4[7145] = 32'b11111111111111110000011111010110;
assign LUT_4[7146] = 32'b11111111111111110110101110000010;
assign LUT_4[7147] = 32'b11111111111111101111111001111010;
assign LUT_4[7148] = 32'b11111111111111110100010011111010;
assign LUT_4[7149] = 32'b11111111111111101101011111110010;
assign LUT_4[7150] = 32'b11111111111111110011101110011110;
assign LUT_4[7151] = 32'b11111111111111101100111010010110;
assign LUT_4[7152] = 32'b11111111111111111011111000110111;
assign LUT_4[7153] = 32'b11111111111111110101000100101111;
assign LUT_4[7154] = 32'b11111111111111111011010011011011;
assign LUT_4[7155] = 32'b11111111111111110100011111010011;
assign LUT_4[7156] = 32'b11111111111111111000111001010011;
assign LUT_4[7157] = 32'b11111111111111110010000101001011;
assign LUT_4[7158] = 32'b11111111111111111000010011110111;
assign LUT_4[7159] = 32'b11111111111111110001011111101111;
assign LUT_4[7160] = 32'b11111111111111110101000101001100;
assign LUT_4[7161] = 32'b11111111111111101110010001000100;
assign LUT_4[7162] = 32'b11111111111111110100011111110000;
assign LUT_4[7163] = 32'b11111111111111101101101011101000;
assign LUT_4[7164] = 32'b11111111111111110010000101101000;
assign LUT_4[7165] = 32'b11111111111111101011010001100000;
assign LUT_4[7166] = 32'b11111111111111110001100000001100;
assign LUT_4[7167] = 32'b11111111111111101010101100000100;
assign LUT_4[7168] = 32'b11111111111111111001011001011010;
assign LUT_4[7169] = 32'b11111111111111110010100101010010;
assign LUT_4[7170] = 32'b11111111111111111000110011111110;
assign LUT_4[7171] = 32'b11111111111111110001111111110110;
assign LUT_4[7172] = 32'b11111111111111110110011001110110;
assign LUT_4[7173] = 32'b11111111111111101111100101101110;
assign LUT_4[7174] = 32'b11111111111111110101110100011010;
assign LUT_4[7175] = 32'b11111111111111101111000000010010;
assign LUT_4[7176] = 32'b11111111111111110010100101101111;
assign LUT_4[7177] = 32'b11111111111111101011110001100111;
assign LUT_4[7178] = 32'b11111111111111110010000000010011;
assign LUT_4[7179] = 32'b11111111111111101011001100001011;
assign LUT_4[7180] = 32'b11111111111111101111100110001011;
assign LUT_4[7181] = 32'b11111111111111101000110010000011;
assign LUT_4[7182] = 32'b11111111111111101111000000101111;
assign LUT_4[7183] = 32'b11111111111111101000001100100111;
assign LUT_4[7184] = 32'b11111111111111110111001011001000;
assign LUT_4[7185] = 32'b11111111111111110000010111000000;
assign LUT_4[7186] = 32'b11111111111111110110100101101100;
assign LUT_4[7187] = 32'b11111111111111101111110001100100;
assign LUT_4[7188] = 32'b11111111111111110100001011100100;
assign LUT_4[7189] = 32'b11111111111111101101010111011100;
assign LUT_4[7190] = 32'b11111111111111110011100110001000;
assign LUT_4[7191] = 32'b11111111111111101100110010000000;
assign LUT_4[7192] = 32'b11111111111111110000010111011101;
assign LUT_4[7193] = 32'b11111111111111101001100011010101;
assign LUT_4[7194] = 32'b11111111111111101111110010000001;
assign LUT_4[7195] = 32'b11111111111111101000111101111001;
assign LUT_4[7196] = 32'b11111111111111101101010111111001;
assign LUT_4[7197] = 32'b11111111111111100110100011110001;
assign LUT_4[7198] = 32'b11111111111111101100110010011101;
assign LUT_4[7199] = 32'b11111111111111100101111110010101;
assign LUT_4[7200] = 32'b11111111111111110111110100100001;
assign LUT_4[7201] = 32'b11111111111111110001000000011001;
assign LUT_4[7202] = 32'b11111111111111110111001111000101;
assign LUT_4[7203] = 32'b11111111111111110000011010111101;
assign LUT_4[7204] = 32'b11111111111111110100110100111101;
assign LUT_4[7205] = 32'b11111111111111101110000000110101;
assign LUT_4[7206] = 32'b11111111111111110100001111100001;
assign LUT_4[7207] = 32'b11111111111111101101011011011001;
assign LUT_4[7208] = 32'b11111111111111110001000000110110;
assign LUT_4[7209] = 32'b11111111111111101010001100101110;
assign LUT_4[7210] = 32'b11111111111111110000011011011010;
assign LUT_4[7211] = 32'b11111111111111101001100111010010;
assign LUT_4[7212] = 32'b11111111111111101110000001010010;
assign LUT_4[7213] = 32'b11111111111111100111001101001010;
assign LUT_4[7214] = 32'b11111111111111101101011011110110;
assign LUT_4[7215] = 32'b11111111111111100110100111101110;
assign LUT_4[7216] = 32'b11111111111111110101100110001111;
assign LUT_4[7217] = 32'b11111111111111101110110010000111;
assign LUT_4[7218] = 32'b11111111111111110101000000110011;
assign LUT_4[7219] = 32'b11111111111111101110001100101011;
assign LUT_4[7220] = 32'b11111111111111110010100110101011;
assign LUT_4[7221] = 32'b11111111111111101011110010100011;
assign LUT_4[7222] = 32'b11111111111111110010000001001111;
assign LUT_4[7223] = 32'b11111111111111101011001101000111;
assign LUT_4[7224] = 32'b11111111111111101110110010100100;
assign LUT_4[7225] = 32'b11111111111111100111111110011100;
assign LUT_4[7226] = 32'b11111111111111101110001101001000;
assign LUT_4[7227] = 32'b11111111111111100111011001000000;
assign LUT_4[7228] = 32'b11111111111111101011110011000000;
assign LUT_4[7229] = 32'b11111111111111100100111110111000;
assign LUT_4[7230] = 32'b11111111111111101011001101100100;
assign LUT_4[7231] = 32'b11111111111111100100011001011100;
assign LUT_4[7232] = 32'b11111111111111111010110000101110;
assign LUT_4[7233] = 32'b11111111111111110011111100100110;
assign LUT_4[7234] = 32'b11111111111111111010001011010010;
assign LUT_4[7235] = 32'b11111111111111110011010111001010;
assign LUT_4[7236] = 32'b11111111111111110111110001001010;
assign LUT_4[7237] = 32'b11111111111111110000111101000010;
assign LUT_4[7238] = 32'b11111111111111110111001011101110;
assign LUT_4[7239] = 32'b11111111111111110000010111100110;
assign LUT_4[7240] = 32'b11111111111111110011111101000011;
assign LUT_4[7241] = 32'b11111111111111101101001000111011;
assign LUT_4[7242] = 32'b11111111111111110011010111100111;
assign LUT_4[7243] = 32'b11111111111111101100100011011111;
assign LUT_4[7244] = 32'b11111111111111110000111101011111;
assign LUT_4[7245] = 32'b11111111111111101010001001010111;
assign LUT_4[7246] = 32'b11111111111111110000011000000011;
assign LUT_4[7247] = 32'b11111111111111101001100011111011;
assign LUT_4[7248] = 32'b11111111111111111000100010011100;
assign LUT_4[7249] = 32'b11111111111111110001101110010100;
assign LUT_4[7250] = 32'b11111111111111110111111101000000;
assign LUT_4[7251] = 32'b11111111111111110001001000111000;
assign LUT_4[7252] = 32'b11111111111111110101100010111000;
assign LUT_4[7253] = 32'b11111111111111101110101110110000;
assign LUT_4[7254] = 32'b11111111111111110100111101011100;
assign LUT_4[7255] = 32'b11111111111111101110001001010100;
assign LUT_4[7256] = 32'b11111111111111110001101110110001;
assign LUT_4[7257] = 32'b11111111111111101010111010101001;
assign LUT_4[7258] = 32'b11111111111111110001001001010101;
assign LUT_4[7259] = 32'b11111111111111101010010101001101;
assign LUT_4[7260] = 32'b11111111111111101110101111001101;
assign LUT_4[7261] = 32'b11111111111111100111111011000101;
assign LUT_4[7262] = 32'b11111111111111101110001001110001;
assign LUT_4[7263] = 32'b11111111111111100111010101101001;
assign LUT_4[7264] = 32'b11111111111111111001001011110101;
assign LUT_4[7265] = 32'b11111111111111110010010111101101;
assign LUT_4[7266] = 32'b11111111111111111000100110011001;
assign LUT_4[7267] = 32'b11111111111111110001110010010001;
assign LUT_4[7268] = 32'b11111111111111110110001100010001;
assign LUT_4[7269] = 32'b11111111111111101111011000001001;
assign LUT_4[7270] = 32'b11111111111111110101100110110101;
assign LUT_4[7271] = 32'b11111111111111101110110010101101;
assign LUT_4[7272] = 32'b11111111111111110010011000001010;
assign LUT_4[7273] = 32'b11111111111111101011100100000010;
assign LUT_4[7274] = 32'b11111111111111110001110010101110;
assign LUT_4[7275] = 32'b11111111111111101010111110100110;
assign LUT_4[7276] = 32'b11111111111111101111011000100110;
assign LUT_4[7277] = 32'b11111111111111101000100100011110;
assign LUT_4[7278] = 32'b11111111111111101110110011001010;
assign LUT_4[7279] = 32'b11111111111111100111111111000010;
assign LUT_4[7280] = 32'b11111111111111110110111101100011;
assign LUT_4[7281] = 32'b11111111111111110000001001011011;
assign LUT_4[7282] = 32'b11111111111111110110011000000111;
assign LUT_4[7283] = 32'b11111111111111101111100011111111;
assign LUT_4[7284] = 32'b11111111111111110011111101111111;
assign LUT_4[7285] = 32'b11111111111111101101001001110111;
assign LUT_4[7286] = 32'b11111111111111110011011000100011;
assign LUT_4[7287] = 32'b11111111111111101100100100011011;
assign LUT_4[7288] = 32'b11111111111111110000001001111000;
assign LUT_4[7289] = 32'b11111111111111101001010101110000;
assign LUT_4[7290] = 32'b11111111111111101111100100011100;
assign LUT_4[7291] = 32'b11111111111111101000110000010100;
assign LUT_4[7292] = 32'b11111111111111101101001010010100;
assign LUT_4[7293] = 32'b11111111111111100110010110001100;
assign LUT_4[7294] = 32'b11111111111111101100100100111000;
assign LUT_4[7295] = 32'b11111111111111100101110000110000;
assign LUT_4[7296] = 32'b11111111111111111011111111100010;
assign LUT_4[7297] = 32'b11111111111111110101001011011010;
assign LUT_4[7298] = 32'b11111111111111111011011010000110;
assign LUT_4[7299] = 32'b11111111111111110100100101111110;
assign LUT_4[7300] = 32'b11111111111111111000111111111110;
assign LUT_4[7301] = 32'b11111111111111110010001011110110;
assign LUT_4[7302] = 32'b11111111111111111000011010100010;
assign LUT_4[7303] = 32'b11111111111111110001100110011010;
assign LUT_4[7304] = 32'b11111111111111110101001011110111;
assign LUT_4[7305] = 32'b11111111111111101110010111101111;
assign LUT_4[7306] = 32'b11111111111111110100100110011011;
assign LUT_4[7307] = 32'b11111111111111101101110010010011;
assign LUT_4[7308] = 32'b11111111111111110010001100010011;
assign LUT_4[7309] = 32'b11111111111111101011011000001011;
assign LUT_4[7310] = 32'b11111111111111110001100110110111;
assign LUT_4[7311] = 32'b11111111111111101010110010101111;
assign LUT_4[7312] = 32'b11111111111111111001110001010000;
assign LUT_4[7313] = 32'b11111111111111110010111101001000;
assign LUT_4[7314] = 32'b11111111111111111001001011110100;
assign LUT_4[7315] = 32'b11111111111111110010010111101100;
assign LUT_4[7316] = 32'b11111111111111110110110001101100;
assign LUT_4[7317] = 32'b11111111111111101111111101100100;
assign LUT_4[7318] = 32'b11111111111111110110001100010000;
assign LUT_4[7319] = 32'b11111111111111101111011000001000;
assign LUT_4[7320] = 32'b11111111111111110010111101100101;
assign LUT_4[7321] = 32'b11111111111111101100001001011101;
assign LUT_4[7322] = 32'b11111111111111110010011000001001;
assign LUT_4[7323] = 32'b11111111111111101011100100000001;
assign LUT_4[7324] = 32'b11111111111111101111111110000001;
assign LUT_4[7325] = 32'b11111111111111101001001001111001;
assign LUT_4[7326] = 32'b11111111111111101111011000100101;
assign LUT_4[7327] = 32'b11111111111111101000100100011101;
assign LUT_4[7328] = 32'b11111111111111111010011010101001;
assign LUT_4[7329] = 32'b11111111111111110011100110100001;
assign LUT_4[7330] = 32'b11111111111111111001110101001101;
assign LUT_4[7331] = 32'b11111111111111110011000001000101;
assign LUT_4[7332] = 32'b11111111111111110111011011000101;
assign LUT_4[7333] = 32'b11111111111111110000100110111101;
assign LUT_4[7334] = 32'b11111111111111110110110101101001;
assign LUT_4[7335] = 32'b11111111111111110000000001100001;
assign LUT_4[7336] = 32'b11111111111111110011100110111110;
assign LUT_4[7337] = 32'b11111111111111101100110010110110;
assign LUT_4[7338] = 32'b11111111111111110011000001100010;
assign LUT_4[7339] = 32'b11111111111111101100001101011010;
assign LUT_4[7340] = 32'b11111111111111110000100111011010;
assign LUT_4[7341] = 32'b11111111111111101001110011010010;
assign LUT_4[7342] = 32'b11111111111111110000000001111110;
assign LUT_4[7343] = 32'b11111111111111101001001101110110;
assign LUT_4[7344] = 32'b11111111111111111000001100010111;
assign LUT_4[7345] = 32'b11111111111111110001011000001111;
assign LUT_4[7346] = 32'b11111111111111110111100110111011;
assign LUT_4[7347] = 32'b11111111111111110000110010110011;
assign LUT_4[7348] = 32'b11111111111111110101001100110011;
assign LUT_4[7349] = 32'b11111111111111101110011000101011;
assign LUT_4[7350] = 32'b11111111111111110100100111010111;
assign LUT_4[7351] = 32'b11111111111111101101110011001111;
assign LUT_4[7352] = 32'b11111111111111110001011000101100;
assign LUT_4[7353] = 32'b11111111111111101010100100100100;
assign LUT_4[7354] = 32'b11111111111111110000110011010000;
assign LUT_4[7355] = 32'b11111111111111101001111111001000;
assign LUT_4[7356] = 32'b11111111111111101110011001001000;
assign LUT_4[7357] = 32'b11111111111111100111100101000000;
assign LUT_4[7358] = 32'b11111111111111101101110011101100;
assign LUT_4[7359] = 32'b11111111111111100110111111100100;
assign LUT_4[7360] = 32'b11111111111111111101010110110110;
assign LUT_4[7361] = 32'b11111111111111110110100010101110;
assign LUT_4[7362] = 32'b11111111111111111100110001011010;
assign LUT_4[7363] = 32'b11111111111111110101111101010010;
assign LUT_4[7364] = 32'b11111111111111111010010111010010;
assign LUT_4[7365] = 32'b11111111111111110011100011001010;
assign LUT_4[7366] = 32'b11111111111111111001110001110110;
assign LUT_4[7367] = 32'b11111111111111110010111101101110;
assign LUT_4[7368] = 32'b11111111111111110110100011001011;
assign LUT_4[7369] = 32'b11111111111111101111101111000011;
assign LUT_4[7370] = 32'b11111111111111110101111101101111;
assign LUT_4[7371] = 32'b11111111111111101111001001100111;
assign LUT_4[7372] = 32'b11111111111111110011100011100111;
assign LUT_4[7373] = 32'b11111111111111101100101111011111;
assign LUT_4[7374] = 32'b11111111111111110010111110001011;
assign LUT_4[7375] = 32'b11111111111111101100001010000011;
assign LUT_4[7376] = 32'b11111111111111111011001000100100;
assign LUT_4[7377] = 32'b11111111111111110100010100011100;
assign LUT_4[7378] = 32'b11111111111111111010100011001000;
assign LUT_4[7379] = 32'b11111111111111110011101111000000;
assign LUT_4[7380] = 32'b11111111111111111000001001000000;
assign LUT_4[7381] = 32'b11111111111111110001010100111000;
assign LUT_4[7382] = 32'b11111111111111110111100011100100;
assign LUT_4[7383] = 32'b11111111111111110000101111011100;
assign LUT_4[7384] = 32'b11111111111111110100010100111001;
assign LUT_4[7385] = 32'b11111111111111101101100000110001;
assign LUT_4[7386] = 32'b11111111111111110011101111011101;
assign LUT_4[7387] = 32'b11111111111111101100111011010101;
assign LUT_4[7388] = 32'b11111111111111110001010101010101;
assign LUT_4[7389] = 32'b11111111111111101010100001001101;
assign LUT_4[7390] = 32'b11111111111111110000101111111001;
assign LUT_4[7391] = 32'b11111111111111101001111011110001;
assign LUT_4[7392] = 32'b11111111111111111011110001111101;
assign LUT_4[7393] = 32'b11111111111111110100111101110101;
assign LUT_4[7394] = 32'b11111111111111111011001100100001;
assign LUT_4[7395] = 32'b11111111111111110100011000011001;
assign LUT_4[7396] = 32'b11111111111111111000110010011001;
assign LUT_4[7397] = 32'b11111111111111110001111110010001;
assign LUT_4[7398] = 32'b11111111111111111000001100111101;
assign LUT_4[7399] = 32'b11111111111111110001011000110101;
assign LUT_4[7400] = 32'b11111111111111110100111110010010;
assign LUT_4[7401] = 32'b11111111111111101110001010001010;
assign LUT_4[7402] = 32'b11111111111111110100011000110110;
assign LUT_4[7403] = 32'b11111111111111101101100100101110;
assign LUT_4[7404] = 32'b11111111111111110001111110101110;
assign LUT_4[7405] = 32'b11111111111111101011001010100110;
assign LUT_4[7406] = 32'b11111111111111110001011001010010;
assign LUT_4[7407] = 32'b11111111111111101010100101001010;
assign LUT_4[7408] = 32'b11111111111111111001100011101011;
assign LUT_4[7409] = 32'b11111111111111110010101111100011;
assign LUT_4[7410] = 32'b11111111111111111000111110001111;
assign LUT_4[7411] = 32'b11111111111111110010001010000111;
assign LUT_4[7412] = 32'b11111111111111110110100100000111;
assign LUT_4[7413] = 32'b11111111111111101111101111111111;
assign LUT_4[7414] = 32'b11111111111111110101111110101011;
assign LUT_4[7415] = 32'b11111111111111101111001010100011;
assign LUT_4[7416] = 32'b11111111111111110010110000000000;
assign LUT_4[7417] = 32'b11111111111111101011111011111000;
assign LUT_4[7418] = 32'b11111111111111110010001010100100;
assign LUT_4[7419] = 32'b11111111111111101011010110011100;
assign LUT_4[7420] = 32'b11111111111111101111110000011100;
assign LUT_4[7421] = 32'b11111111111111101000111100010100;
assign LUT_4[7422] = 32'b11111111111111101111001011000000;
assign LUT_4[7423] = 32'b11111111111111101000010110111000;
assign LUT_4[7424] = 32'b11111111111111111110010100111101;
assign LUT_4[7425] = 32'b11111111111111110111100000110101;
assign LUT_4[7426] = 32'b11111111111111111101101111100001;
assign LUT_4[7427] = 32'b11111111111111110110111011011001;
assign LUT_4[7428] = 32'b11111111111111111011010101011001;
assign LUT_4[7429] = 32'b11111111111111110100100001010001;
assign LUT_4[7430] = 32'b11111111111111111010101111111101;
assign LUT_4[7431] = 32'b11111111111111110011111011110101;
assign LUT_4[7432] = 32'b11111111111111110111100001010010;
assign LUT_4[7433] = 32'b11111111111111110000101101001010;
assign LUT_4[7434] = 32'b11111111111111110110111011110110;
assign LUT_4[7435] = 32'b11111111111111110000000111101110;
assign LUT_4[7436] = 32'b11111111111111110100100001101110;
assign LUT_4[7437] = 32'b11111111111111101101101101100110;
assign LUT_4[7438] = 32'b11111111111111110011111100010010;
assign LUT_4[7439] = 32'b11111111111111101101001000001010;
assign LUT_4[7440] = 32'b11111111111111111100000110101011;
assign LUT_4[7441] = 32'b11111111111111110101010010100011;
assign LUT_4[7442] = 32'b11111111111111111011100001001111;
assign LUT_4[7443] = 32'b11111111111111110100101101000111;
assign LUT_4[7444] = 32'b11111111111111111001000111000111;
assign LUT_4[7445] = 32'b11111111111111110010010010111111;
assign LUT_4[7446] = 32'b11111111111111111000100001101011;
assign LUT_4[7447] = 32'b11111111111111110001101101100011;
assign LUT_4[7448] = 32'b11111111111111110101010011000000;
assign LUT_4[7449] = 32'b11111111111111101110011110111000;
assign LUT_4[7450] = 32'b11111111111111110100101101100100;
assign LUT_4[7451] = 32'b11111111111111101101111001011100;
assign LUT_4[7452] = 32'b11111111111111110010010011011100;
assign LUT_4[7453] = 32'b11111111111111101011011111010100;
assign LUT_4[7454] = 32'b11111111111111110001101110000000;
assign LUT_4[7455] = 32'b11111111111111101010111001111000;
assign LUT_4[7456] = 32'b11111111111111111100110000000100;
assign LUT_4[7457] = 32'b11111111111111110101111011111100;
assign LUT_4[7458] = 32'b11111111111111111100001010101000;
assign LUT_4[7459] = 32'b11111111111111110101010110100000;
assign LUT_4[7460] = 32'b11111111111111111001110000100000;
assign LUT_4[7461] = 32'b11111111111111110010111100011000;
assign LUT_4[7462] = 32'b11111111111111111001001011000100;
assign LUT_4[7463] = 32'b11111111111111110010010110111100;
assign LUT_4[7464] = 32'b11111111111111110101111100011001;
assign LUT_4[7465] = 32'b11111111111111101111001000010001;
assign LUT_4[7466] = 32'b11111111111111110101010110111101;
assign LUT_4[7467] = 32'b11111111111111101110100010110101;
assign LUT_4[7468] = 32'b11111111111111110010111100110101;
assign LUT_4[7469] = 32'b11111111111111101100001000101101;
assign LUT_4[7470] = 32'b11111111111111110010010111011001;
assign LUT_4[7471] = 32'b11111111111111101011100011010001;
assign LUT_4[7472] = 32'b11111111111111111010100001110010;
assign LUT_4[7473] = 32'b11111111111111110011101101101010;
assign LUT_4[7474] = 32'b11111111111111111001111100010110;
assign LUT_4[7475] = 32'b11111111111111110011001000001110;
assign LUT_4[7476] = 32'b11111111111111110111100010001110;
assign LUT_4[7477] = 32'b11111111111111110000101110000110;
assign LUT_4[7478] = 32'b11111111111111110110111100110010;
assign LUT_4[7479] = 32'b11111111111111110000001000101010;
assign LUT_4[7480] = 32'b11111111111111110011101110000111;
assign LUT_4[7481] = 32'b11111111111111101100111001111111;
assign LUT_4[7482] = 32'b11111111111111110011001000101011;
assign LUT_4[7483] = 32'b11111111111111101100010100100011;
assign LUT_4[7484] = 32'b11111111111111110000101110100011;
assign LUT_4[7485] = 32'b11111111111111101001111010011011;
assign LUT_4[7486] = 32'b11111111111111110000001001000111;
assign LUT_4[7487] = 32'b11111111111111101001010100111111;
assign LUT_4[7488] = 32'b11111111111111111111101100010001;
assign LUT_4[7489] = 32'b11111111111111111000111000001001;
assign LUT_4[7490] = 32'b11111111111111111111000110110101;
assign LUT_4[7491] = 32'b11111111111111111000010010101101;
assign LUT_4[7492] = 32'b11111111111111111100101100101101;
assign LUT_4[7493] = 32'b11111111111111110101111000100101;
assign LUT_4[7494] = 32'b11111111111111111100000111010001;
assign LUT_4[7495] = 32'b11111111111111110101010011001001;
assign LUT_4[7496] = 32'b11111111111111111000111000100110;
assign LUT_4[7497] = 32'b11111111111111110010000100011110;
assign LUT_4[7498] = 32'b11111111111111111000010011001010;
assign LUT_4[7499] = 32'b11111111111111110001011111000010;
assign LUT_4[7500] = 32'b11111111111111110101111001000010;
assign LUT_4[7501] = 32'b11111111111111101111000100111010;
assign LUT_4[7502] = 32'b11111111111111110101010011100110;
assign LUT_4[7503] = 32'b11111111111111101110011111011110;
assign LUT_4[7504] = 32'b11111111111111111101011101111111;
assign LUT_4[7505] = 32'b11111111111111110110101001110111;
assign LUT_4[7506] = 32'b11111111111111111100111000100011;
assign LUT_4[7507] = 32'b11111111111111110110000100011011;
assign LUT_4[7508] = 32'b11111111111111111010011110011011;
assign LUT_4[7509] = 32'b11111111111111110011101010010011;
assign LUT_4[7510] = 32'b11111111111111111001111000111111;
assign LUT_4[7511] = 32'b11111111111111110011000100110111;
assign LUT_4[7512] = 32'b11111111111111110110101010010100;
assign LUT_4[7513] = 32'b11111111111111101111110110001100;
assign LUT_4[7514] = 32'b11111111111111110110000100111000;
assign LUT_4[7515] = 32'b11111111111111101111010000110000;
assign LUT_4[7516] = 32'b11111111111111110011101010110000;
assign LUT_4[7517] = 32'b11111111111111101100110110101000;
assign LUT_4[7518] = 32'b11111111111111110011000101010100;
assign LUT_4[7519] = 32'b11111111111111101100010001001100;
assign LUT_4[7520] = 32'b11111111111111111110000111011000;
assign LUT_4[7521] = 32'b11111111111111110111010011010000;
assign LUT_4[7522] = 32'b11111111111111111101100001111100;
assign LUT_4[7523] = 32'b11111111111111110110101101110100;
assign LUT_4[7524] = 32'b11111111111111111011000111110100;
assign LUT_4[7525] = 32'b11111111111111110100010011101100;
assign LUT_4[7526] = 32'b11111111111111111010100010011000;
assign LUT_4[7527] = 32'b11111111111111110011101110010000;
assign LUT_4[7528] = 32'b11111111111111110111010011101101;
assign LUT_4[7529] = 32'b11111111111111110000011111100101;
assign LUT_4[7530] = 32'b11111111111111110110101110010001;
assign LUT_4[7531] = 32'b11111111111111101111111010001001;
assign LUT_4[7532] = 32'b11111111111111110100010100001001;
assign LUT_4[7533] = 32'b11111111111111101101100000000001;
assign LUT_4[7534] = 32'b11111111111111110011101110101101;
assign LUT_4[7535] = 32'b11111111111111101100111010100101;
assign LUT_4[7536] = 32'b11111111111111111011111001000110;
assign LUT_4[7537] = 32'b11111111111111110101000100111110;
assign LUT_4[7538] = 32'b11111111111111111011010011101010;
assign LUT_4[7539] = 32'b11111111111111110100011111100010;
assign LUT_4[7540] = 32'b11111111111111111000111001100010;
assign LUT_4[7541] = 32'b11111111111111110010000101011010;
assign LUT_4[7542] = 32'b11111111111111111000010100000110;
assign LUT_4[7543] = 32'b11111111111111110001011111111110;
assign LUT_4[7544] = 32'b11111111111111110101000101011011;
assign LUT_4[7545] = 32'b11111111111111101110010001010011;
assign LUT_4[7546] = 32'b11111111111111110100011111111111;
assign LUT_4[7547] = 32'b11111111111111101101101011110111;
assign LUT_4[7548] = 32'b11111111111111110010000101110111;
assign LUT_4[7549] = 32'b11111111111111101011010001101111;
assign LUT_4[7550] = 32'b11111111111111110001100000011011;
assign LUT_4[7551] = 32'b11111111111111101010101100010011;
assign LUT_4[7552] = 32'b00000000000000000000111011000101;
assign LUT_4[7553] = 32'b11111111111111111010000110111101;
assign LUT_4[7554] = 32'b00000000000000000000010101101001;
assign LUT_4[7555] = 32'b11111111111111111001100001100001;
assign LUT_4[7556] = 32'b11111111111111111101111011100001;
assign LUT_4[7557] = 32'b11111111111111110111000111011001;
assign LUT_4[7558] = 32'b11111111111111111101010110000101;
assign LUT_4[7559] = 32'b11111111111111110110100001111101;
assign LUT_4[7560] = 32'b11111111111111111010000111011010;
assign LUT_4[7561] = 32'b11111111111111110011010011010010;
assign LUT_4[7562] = 32'b11111111111111111001100001111110;
assign LUT_4[7563] = 32'b11111111111111110010101101110110;
assign LUT_4[7564] = 32'b11111111111111110111000111110110;
assign LUT_4[7565] = 32'b11111111111111110000010011101110;
assign LUT_4[7566] = 32'b11111111111111110110100010011010;
assign LUT_4[7567] = 32'b11111111111111101111101110010010;
assign LUT_4[7568] = 32'b11111111111111111110101100110011;
assign LUT_4[7569] = 32'b11111111111111110111111000101011;
assign LUT_4[7570] = 32'b11111111111111111110000111010111;
assign LUT_4[7571] = 32'b11111111111111110111010011001111;
assign LUT_4[7572] = 32'b11111111111111111011101101001111;
assign LUT_4[7573] = 32'b11111111111111110100111001000111;
assign LUT_4[7574] = 32'b11111111111111111011000111110011;
assign LUT_4[7575] = 32'b11111111111111110100010011101011;
assign LUT_4[7576] = 32'b11111111111111110111111001001000;
assign LUT_4[7577] = 32'b11111111111111110001000101000000;
assign LUT_4[7578] = 32'b11111111111111110111010011101100;
assign LUT_4[7579] = 32'b11111111111111110000011111100100;
assign LUT_4[7580] = 32'b11111111111111110100111001100100;
assign LUT_4[7581] = 32'b11111111111111101110000101011100;
assign LUT_4[7582] = 32'b11111111111111110100010100001000;
assign LUT_4[7583] = 32'b11111111111111101101100000000000;
assign LUT_4[7584] = 32'b11111111111111111111010110001100;
assign LUT_4[7585] = 32'b11111111111111111000100010000100;
assign LUT_4[7586] = 32'b11111111111111111110110000110000;
assign LUT_4[7587] = 32'b11111111111111110111111100101000;
assign LUT_4[7588] = 32'b11111111111111111100010110101000;
assign LUT_4[7589] = 32'b11111111111111110101100010100000;
assign LUT_4[7590] = 32'b11111111111111111011110001001100;
assign LUT_4[7591] = 32'b11111111111111110100111101000100;
assign LUT_4[7592] = 32'b11111111111111111000100010100001;
assign LUT_4[7593] = 32'b11111111111111110001101110011001;
assign LUT_4[7594] = 32'b11111111111111110111111101000101;
assign LUT_4[7595] = 32'b11111111111111110001001000111101;
assign LUT_4[7596] = 32'b11111111111111110101100010111101;
assign LUT_4[7597] = 32'b11111111111111101110101110110101;
assign LUT_4[7598] = 32'b11111111111111110100111101100001;
assign LUT_4[7599] = 32'b11111111111111101110001001011001;
assign LUT_4[7600] = 32'b11111111111111111101000111111010;
assign LUT_4[7601] = 32'b11111111111111110110010011110010;
assign LUT_4[7602] = 32'b11111111111111111100100010011110;
assign LUT_4[7603] = 32'b11111111111111110101101110010110;
assign LUT_4[7604] = 32'b11111111111111111010001000010110;
assign LUT_4[7605] = 32'b11111111111111110011010100001110;
assign LUT_4[7606] = 32'b11111111111111111001100010111010;
assign LUT_4[7607] = 32'b11111111111111110010101110110010;
assign LUT_4[7608] = 32'b11111111111111110110010100001111;
assign LUT_4[7609] = 32'b11111111111111101111100000000111;
assign LUT_4[7610] = 32'b11111111111111110101101110110011;
assign LUT_4[7611] = 32'b11111111111111101110111010101011;
assign LUT_4[7612] = 32'b11111111111111110011010100101011;
assign LUT_4[7613] = 32'b11111111111111101100100000100011;
assign LUT_4[7614] = 32'b11111111111111110010101111001111;
assign LUT_4[7615] = 32'b11111111111111101011111011000111;
assign LUT_4[7616] = 32'b00000000000000000010010010011001;
assign LUT_4[7617] = 32'b11111111111111111011011110010001;
assign LUT_4[7618] = 32'b00000000000000000001101100111101;
assign LUT_4[7619] = 32'b11111111111111111010111000110101;
assign LUT_4[7620] = 32'b11111111111111111111010010110101;
assign LUT_4[7621] = 32'b11111111111111111000011110101101;
assign LUT_4[7622] = 32'b11111111111111111110101101011001;
assign LUT_4[7623] = 32'b11111111111111110111111001010001;
assign LUT_4[7624] = 32'b11111111111111111011011110101110;
assign LUT_4[7625] = 32'b11111111111111110100101010100110;
assign LUT_4[7626] = 32'b11111111111111111010111001010010;
assign LUT_4[7627] = 32'b11111111111111110100000101001010;
assign LUT_4[7628] = 32'b11111111111111111000011111001010;
assign LUT_4[7629] = 32'b11111111111111110001101011000010;
assign LUT_4[7630] = 32'b11111111111111110111111001101110;
assign LUT_4[7631] = 32'b11111111111111110001000101100110;
assign LUT_4[7632] = 32'b00000000000000000000000100000111;
assign LUT_4[7633] = 32'b11111111111111111001001111111111;
assign LUT_4[7634] = 32'b11111111111111111111011110101011;
assign LUT_4[7635] = 32'b11111111111111111000101010100011;
assign LUT_4[7636] = 32'b11111111111111111101000100100011;
assign LUT_4[7637] = 32'b11111111111111110110010000011011;
assign LUT_4[7638] = 32'b11111111111111111100011111000111;
assign LUT_4[7639] = 32'b11111111111111110101101010111111;
assign LUT_4[7640] = 32'b11111111111111111001010000011100;
assign LUT_4[7641] = 32'b11111111111111110010011100010100;
assign LUT_4[7642] = 32'b11111111111111111000101011000000;
assign LUT_4[7643] = 32'b11111111111111110001110110111000;
assign LUT_4[7644] = 32'b11111111111111110110010000111000;
assign LUT_4[7645] = 32'b11111111111111101111011100110000;
assign LUT_4[7646] = 32'b11111111111111110101101011011100;
assign LUT_4[7647] = 32'b11111111111111101110110111010100;
assign LUT_4[7648] = 32'b00000000000000000000101101100000;
assign LUT_4[7649] = 32'b11111111111111111001111001011000;
assign LUT_4[7650] = 32'b00000000000000000000001000000100;
assign LUT_4[7651] = 32'b11111111111111111001010011111100;
assign LUT_4[7652] = 32'b11111111111111111101101101111100;
assign LUT_4[7653] = 32'b11111111111111110110111001110100;
assign LUT_4[7654] = 32'b11111111111111111101001000100000;
assign LUT_4[7655] = 32'b11111111111111110110010100011000;
assign LUT_4[7656] = 32'b11111111111111111001111001110101;
assign LUT_4[7657] = 32'b11111111111111110011000101101101;
assign LUT_4[7658] = 32'b11111111111111111001010100011001;
assign LUT_4[7659] = 32'b11111111111111110010100000010001;
assign LUT_4[7660] = 32'b11111111111111110110111010010001;
assign LUT_4[7661] = 32'b11111111111111110000000110001001;
assign LUT_4[7662] = 32'b11111111111111110110010100110101;
assign LUT_4[7663] = 32'b11111111111111101111100000101101;
assign LUT_4[7664] = 32'b11111111111111111110011111001110;
assign LUT_4[7665] = 32'b11111111111111110111101011000110;
assign LUT_4[7666] = 32'b11111111111111111101111001110010;
assign LUT_4[7667] = 32'b11111111111111110111000101101010;
assign LUT_4[7668] = 32'b11111111111111111011011111101010;
assign LUT_4[7669] = 32'b11111111111111110100101011100010;
assign LUT_4[7670] = 32'b11111111111111111010111010001110;
assign LUT_4[7671] = 32'b11111111111111110100000110000110;
assign LUT_4[7672] = 32'b11111111111111110111101011100011;
assign LUT_4[7673] = 32'b11111111111111110000110111011011;
assign LUT_4[7674] = 32'b11111111111111110111000110000111;
assign LUT_4[7675] = 32'b11111111111111110000010001111111;
assign LUT_4[7676] = 32'b11111111111111110100101011111111;
assign LUT_4[7677] = 32'b11111111111111101101110111110111;
assign LUT_4[7678] = 32'b11111111111111110100000110100011;
assign LUT_4[7679] = 32'b11111111111111101101010010011011;
assign LUT_4[7680] = 32'b11111111111111111000011101100010;
assign LUT_4[7681] = 32'b11111111111111110001101001011010;
assign LUT_4[7682] = 32'b11111111111111110111111000000110;
assign LUT_4[7683] = 32'b11111111111111110001000011111110;
assign LUT_4[7684] = 32'b11111111111111110101011101111110;
assign LUT_4[7685] = 32'b11111111111111101110101001110110;
assign LUT_4[7686] = 32'b11111111111111110100111000100010;
assign LUT_4[7687] = 32'b11111111111111101110000100011010;
assign LUT_4[7688] = 32'b11111111111111110001101001110111;
assign LUT_4[7689] = 32'b11111111111111101010110101101111;
assign LUT_4[7690] = 32'b11111111111111110001000100011011;
assign LUT_4[7691] = 32'b11111111111111101010010000010011;
assign LUT_4[7692] = 32'b11111111111111101110101010010011;
assign LUT_4[7693] = 32'b11111111111111100111110110001011;
assign LUT_4[7694] = 32'b11111111111111101110000100110111;
assign LUT_4[7695] = 32'b11111111111111100111010000101111;
assign LUT_4[7696] = 32'b11111111111111110110001111010000;
assign LUT_4[7697] = 32'b11111111111111101111011011001000;
assign LUT_4[7698] = 32'b11111111111111110101101001110100;
assign LUT_4[7699] = 32'b11111111111111101110110101101100;
assign LUT_4[7700] = 32'b11111111111111110011001111101100;
assign LUT_4[7701] = 32'b11111111111111101100011011100100;
assign LUT_4[7702] = 32'b11111111111111110010101010010000;
assign LUT_4[7703] = 32'b11111111111111101011110110001000;
assign LUT_4[7704] = 32'b11111111111111101111011011100101;
assign LUT_4[7705] = 32'b11111111111111101000100111011101;
assign LUT_4[7706] = 32'b11111111111111101110110110001001;
assign LUT_4[7707] = 32'b11111111111111101000000010000001;
assign LUT_4[7708] = 32'b11111111111111101100011100000001;
assign LUT_4[7709] = 32'b11111111111111100101100111111001;
assign LUT_4[7710] = 32'b11111111111111101011110110100101;
assign LUT_4[7711] = 32'b11111111111111100101000010011101;
assign LUT_4[7712] = 32'b11111111111111110110111000101001;
assign LUT_4[7713] = 32'b11111111111111110000000100100001;
assign LUT_4[7714] = 32'b11111111111111110110010011001101;
assign LUT_4[7715] = 32'b11111111111111101111011111000101;
assign LUT_4[7716] = 32'b11111111111111110011111001000101;
assign LUT_4[7717] = 32'b11111111111111101101000100111101;
assign LUT_4[7718] = 32'b11111111111111110011010011101001;
assign LUT_4[7719] = 32'b11111111111111101100011111100001;
assign LUT_4[7720] = 32'b11111111111111110000000100111110;
assign LUT_4[7721] = 32'b11111111111111101001010000110110;
assign LUT_4[7722] = 32'b11111111111111101111011111100010;
assign LUT_4[7723] = 32'b11111111111111101000101011011010;
assign LUT_4[7724] = 32'b11111111111111101101000101011010;
assign LUT_4[7725] = 32'b11111111111111100110010001010010;
assign LUT_4[7726] = 32'b11111111111111101100011111111110;
assign LUT_4[7727] = 32'b11111111111111100101101011110110;
assign LUT_4[7728] = 32'b11111111111111110100101010010111;
assign LUT_4[7729] = 32'b11111111111111101101110110001111;
assign LUT_4[7730] = 32'b11111111111111110100000100111011;
assign LUT_4[7731] = 32'b11111111111111101101010000110011;
assign LUT_4[7732] = 32'b11111111111111110001101010110011;
assign LUT_4[7733] = 32'b11111111111111101010110110101011;
assign LUT_4[7734] = 32'b11111111111111110001000101010111;
assign LUT_4[7735] = 32'b11111111111111101010010001001111;
assign LUT_4[7736] = 32'b11111111111111101101110110101100;
assign LUT_4[7737] = 32'b11111111111111100111000010100100;
assign LUT_4[7738] = 32'b11111111111111101101010001010000;
assign LUT_4[7739] = 32'b11111111111111100110011101001000;
assign LUT_4[7740] = 32'b11111111111111101010110111001000;
assign LUT_4[7741] = 32'b11111111111111100100000011000000;
assign LUT_4[7742] = 32'b11111111111111101010010001101100;
assign LUT_4[7743] = 32'b11111111111111100011011101100100;
assign LUT_4[7744] = 32'b11111111111111111001110100110110;
assign LUT_4[7745] = 32'b11111111111111110011000000101110;
assign LUT_4[7746] = 32'b11111111111111111001001111011010;
assign LUT_4[7747] = 32'b11111111111111110010011011010010;
assign LUT_4[7748] = 32'b11111111111111110110110101010010;
assign LUT_4[7749] = 32'b11111111111111110000000001001010;
assign LUT_4[7750] = 32'b11111111111111110110001111110110;
assign LUT_4[7751] = 32'b11111111111111101111011011101110;
assign LUT_4[7752] = 32'b11111111111111110011000001001011;
assign LUT_4[7753] = 32'b11111111111111101100001101000011;
assign LUT_4[7754] = 32'b11111111111111110010011011101111;
assign LUT_4[7755] = 32'b11111111111111101011100111100111;
assign LUT_4[7756] = 32'b11111111111111110000000001100111;
assign LUT_4[7757] = 32'b11111111111111101001001101011111;
assign LUT_4[7758] = 32'b11111111111111101111011100001011;
assign LUT_4[7759] = 32'b11111111111111101000101000000011;
assign LUT_4[7760] = 32'b11111111111111110111100110100100;
assign LUT_4[7761] = 32'b11111111111111110000110010011100;
assign LUT_4[7762] = 32'b11111111111111110111000001001000;
assign LUT_4[7763] = 32'b11111111111111110000001101000000;
assign LUT_4[7764] = 32'b11111111111111110100100111000000;
assign LUT_4[7765] = 32'b11111111111111101101110010111000;
assign LUT_4[7766] = 32'b11111111111111110100000001100100;
assign LUT_4[7767] = 32'b11111111111111101101001101011100;
assign LUT_4[7768] = 32'b11111111111111110000110010111001;
assign LUT_4[7769] = 32'b11111111111111101001111110110001;
assign LUT_4[7770] = 32'b11111111111111110000001101011101;
assign LUT_4[7771] = 32'b11111111111111101001011001010101;
assign LUT_4[7772] = 32'b11111111111111101101110011010101;
assign LUT_4[7773] = 32'b11111111111111100110111111001101;
assign LUT_4[7774] = 32'b11111111111111101101001101111001;
assign LUT_4[7775] = 32'b11111111111111100110011001110001;
assign LUT_4[7776] = 32'b11111111111111111000001111111101;
assign LUT_4[7777] = 32'b11111111111111110001011011110101;
assign LUT_4[7778] = 32'b11111111111111110111101010100001;
assign LUT_4[7779] = 32'b11111111111111110000110110011001;
assign LUT_4[7780] = 32'b11111111111111110101010000011001;
assign LUT_4[7781] = 32'b11111111111111101110011100010001;
assign LUT_4[7782] = 32'b11111111111111110100101010111101;
assign LUT_4[7783] = 32'b11111111111111101101110110110101;
assign LUT_4[7784] = 32'b11111111111111110001011100010010;
assign LUT_4[7785] = 32'b11111111111111101010101000001010;
assign LUT_4[7786] = 32'b11111111111111110000110110110110;
assign LUT_4[7787] = 32'b11111111111111101010000010101110;
assign LUT_4[7788] = 32'b11111111111111101110011100101110;
assign LUT_4[7789] = 32'b11111111111111100111101000100110;
assign LUT_4[7790] = 32'b11111111111111101101110111010010;
assign LUT_4[7791] = 32'b11111111111111100111000011001010;
assign LUT_4[7792] = 32'b11111111111111110110000001101011;
assign LUT_4[7793] = 32'b11111111111111101111001101100011;
assign LUT_4[7794] = 32'b11111111111111110101011100001111;
assign LUT_4[7795] = 32'b11111111111111101110101000000111;
assign LUT_4[7796] = 32'b11111111111111110011000010000111;
assign LUT_4[7797] = 32'b11111111111111101100001101111111;
assign LUT_4[7798] = 32'b11111111111111110010011100101011;
assign LUT_4[7799] = 32'b11111111111111101011101000100011;
assign LUT_4[7800] = 32'b11111111111111101111001110000000;
assign LUT_4[7801] = 32'b11111111111111101000011001111000;
assign LUT_4[7802] = 32'b11111111111111101110101000100100;
assign LUT_4[7803] = 32'b11111111111111100111110100011100;
assign LUT_4[7804] = 32'b11111111111111101100001110011100;
assign LUT_4[7805] = 32'b11111111111111100101011010010100;
assign LUT_4[7806] = 32'b11111111111111101011101001000000;
assign LUT_4[7807] = 32'b11111111111111100100110100111000;
assign LUT_4[7808] = 32'b11111111111111111011000011101010;
assign LUT_4[7809] = 32'b11111111111111110100001111100010;
assign LUT_4[7810] = 32'b11111111111111111010011110001110;
assign LUT_4[7811] = 32'b11111111111111110011101010000110;
assign LUT_4[7812] = 32'b11111111111111111000000100000110;
assign LUT_4[7813] = 32'b11111111111111110001001111111110;
assign LUT_4[7814] = 32'b11111111111111110111011110101010;
assign LUT_4[7815] = 32'b11111111111111110000101010100010;
assign LUT_4[7816] = 32'b11111111111111110100001111111111;
assign LUT_4[7817] = 32'b11111111111111101101011011110111;
assign LUT_4[7818] = 32'b11111111111111110011101010100011;
assign LUT_4[7819] = 32'b11111111111111101100110110011011;
assign LUT_4[7820] = 32'b11111111111111110001010000011011;
assign LUT_4[7821] = 32'b11111111111111101010011100010011;
assign LUT_4[7822] = 32'b11111111111111110000101010111111;
assign LUT_4[7823] = 32'b11111111111111101001110110110111;
assign LUT_4[7824] = 32'b11111111111111111000110101011000;
assign LUT_4[7825] = 32'b11111111111111110010000001010000;
assign LUT_4[7826] = 32'b11111111111111111000001111111100;
assign LUT_4[7827] = 32'b11111111111111110001011011110100;
assign LUT_4[7828] = 32'b11111111111111110101110101110100;
assign LUT_4[7829] = 32'b11111111111111101111000001101100;
assign LUT_4[7830] = 32'b11111111111111110101010000011000;
assign LUT_4[7831] = 32'b11111111111111101110011100010000;
assign LUT_4[7832] = 32'b11111111111111110010000001101101;
assign LUT_4[7833] = 32'b11111111111111101011001101100101;
assign LUT_4[7834] = 32'b11111111111111110001011100010001;
assign LUT_4[7835] = 32'b11111111111111101010101000001001;
assign LUT_4[7836] = 32'b11111111111111101111000010001001;
assign LUT_4[7837] = 32'b11111111111111101000001110000001;
assign LUT_4[7838] = 32'b11111111111111101110011100101101;
assign LUT_4[7839] = 32'b11111111111111100111101000100101;
assign LUT_4[7840] = 32'b11111111111111111001011110110001;
assign LUT_4[7841] = 32'b11111111111111110010101010101001;
assign LUT_4[7842] = 32'b11111111111111111000111001010101;
assign LUT_4[7843] = 32'b11111111111111110010000101001101;
assign LUT_4[7844] = 32'b11111111111111110110011111001101;
assign LUT_4[7845] = 32'b11111111111111101111101011000101;
assign LUT_4[7846] = 32'b11111111111111110101111001110001;
assign LUT_4[7847] = 32'b11111111111111101111000101101001;
assign LUT_4[7848] = 32'b11111111111111110010101011000110;
assign LUT_4[7849] = 32'b11111111111111101011110110111110;
assign LUT_4[7850] = 32'b11111111111111110010000101101010;
assign LUT_4[7851] = 32'b11111111111111101011010001100010;
assign LUT_4[7852] = 32'b11111111111111101111101011100010;
assign LUT_4[7853] = 32'b11111111111111101000110111011010;
assign LUT_4[7854] = 32'b11111111111111101111000110000110;
assign LUT_4[7855] = 32'b11111111111111101000010001111110;
assign LUT_4[7856] = 32'b11111111111111110111010000011111;
assign LUT_4[7857] = 32'b11111111111111110000011100010111;
assign LUT_4[7858] = 32'b11111111111111110110101011000011;
assign LUT_4[7859] = 32'b11111111111111101111110110111011;
assign LUT_4[7860] = 32'b11111111111111110100010000111011;
assign LUT_4[7861] = 32'b11111111111111101101011100110011;
assign LUT_4[7862] = 32'b11111111111111110011101011011111;
assign LUT_4[7863] = 32'b11111111111111101100110111010111;
assign LUT_4[7864] = 32'b11111111111111110000011100110100;
assign LUT_4[7865] = 32'b11111111111111101001101000101100;
assign LUT_4[7866] = 32'b11111111111111101111110111011000;
assign LUT_4[7867] = 32'b11111111111111101001000011010000;
assign LUT_4[7868] = 32'b11111111111111101101011101010000;
assign LUT_4[7869] = 32'b11111111111111100110101001001000;
assign LUT_4[7870] = 32'b11111111111111101100110111110100;
assign LUT_4[7871] = 32'b11111111111111100110000011101100;
assign LUT_4[7872] = 32'b11111111111111111100011010111110;
assign LUT_4[7873] = 32'b11111111111111110101100110110110;
assign LUT_4[7874] = 32'b11111111111111111011110101100010;
assign LUT_4[7875] = 32'b11111111111111110101000001011010;
assign LUT_4[7876] = 32'b11111111111111111001011011011010;
assign LUT_4[7877] = 32'b11111111111111110010100111010010;
assign LUT_4[7878] = 32'b11111111111111111000110101111110;
assign LUT_4[7879] = 32'b11111111111111110010000001110110;
assign LUT_4[7880] = 32'b11111111111111110101100111010011;
assign LUT_4[7881] = 32'b11111111111111101110110011001011;
assign LUT_4[7882] = 32'b11111111111111110101000001110111;
assign LUT_4[7883] = 32'b11111111111111101110001101101111;
assign LUT_4[7884] = 32'b11111111111111110010100111101111;
assign LUT_4[7885] = 32'b11111111111111101011110011100111;
assign LUT_4[7886] = 32'b11111111111111110010000010010011;
assign LUT_4[7887] = 32'b11111111111111101011001110001011;
assign LUT_4[7888] = 32'b11111111111111111010001100101100;
assign LUT_4[7889] = 32'b11111111111111110011011000100100;
assign LUT_4[7890] = 32'b11111111111111111001100111010000;
assign LUT_4[7891] = 32'b11111111111111110010110011001000;
assign LUT_4[7892] = 32'b11111111111111110111001101001000;
assign LUT_4[7893] = 32'b11111111111111110000011001000000;
assign LUT_4[7894] = 32'b11111111111111110110100111101100;
assign LUT_4[7895] = 32'b11111111111111101111110011100100;
assign LUT_4[7896] = 32'b11111111111111110011011001000001;
assign LUT_4[7897] = 32'b11111111111111101100100100111001;
assign LUT_4[7898] = 32'b11111111111111110010110011100101;
assign LUT_4[7899] = 32'b11111111111111101011111111011101;
assign LUT_4[7900] = 32'b11111111111111110000011001011101;
assign LUT_4[7901] = 32'b11111111111111101001100101010101;
assign LUT_4[7902] = 32'b11111111111111101111110100000001;
assign LUT_4[7903] = 32'b11111111111111101000111111111001;
assign LUT_4[7904] = 32'b11111111111111111010110110000101;
assign LUT_4[7905] = 32'b11111111111111110100000001111101;
assign LUT_4[7906] = 32'b11111111111111111010010000101001;
assign LUT_4[7907] = 32'b11111111111111110011011100100001;
assign LUT_4[7908] = 32'b11111111111111110111110110100001;
assign LUT_4[7909] = 32'b11111111111111110001000010011001;
assign LUT_4[7910] = 32'b11111111111111110111010001000101;
assign LUT_4[7911] = 32'b11111111111111110000011100111101;
assign LUT_4[7912] = 32'b11111111111111110100000010011010;
assign LUT_4[7913] = 32'b11111111111111101101001110010010;
assign LUT_4[7914] = 32'b11111111111111110011011100111110;
assign LUT_4[7915] = 32'b11111111111111101100101000110110;
assign LUT_4[7916] = 32'b11111111111111110001000010110110;
assign LUT_4[7917] = 32'b11111111111111101010001110101110;
assign LUT_4[7918] = 32'b11111111111111110000011101011010;
assign LUT_4[7919] = 32'b11111111111111101001101001010010;
assign LUT_4[7920] = 32'b11111111111111111000100111110011;
assign LUT_4[7921] = 32'b11111111111111110001110011101011;
assign LUT_4[7922] = 32'b11111111111111111000000010010111;
assign LUT_4[7923] = 32'b11111111111111110001001110001111;
assign LUT_4[7924] = 32'b11111111111111110101101000001111;
assign LUT_4[7925] = 32'b11111111111111101110110100000111;
assign LUT_4[7926] = 32'b11111111111111110101000010110011;
assign LUT_4[7927] = 32'b11111111111111101110001110101011;
assign LUT_4[7928] = 32'b11111111111111110001110100001000;
assign LUT_4[7929] = 32'b11111111111111101011000000000000;
assign LUT_4[7930] = 32'b11111111111111110001001110101100;
assign LUT_4[7931] = 32'b11111111111111101010011010100100;
assign LUT_4[7932] = 32'b11111111111111101110110100100100;
assign LUT_4[7933] = 32'b11111111111111101000000000011100;
assign LUT_4[7934] = 32'b11111111111111101110001111001000;
assign LUT_4[7935] = 32'b11111111111111100111011011000000;
assign LUT_4[7936] = 32'b11111111111111111101011001000101;
assign LUT_4[7937] = 32'b11111111111111110110100100111101;
assign LUT_4[7938] = 32'b11111111111111111100110011101001;
assign LUT_4[7939] = 32'b11111111111111110101111111100001;
assign LUT_4[7940] = 32'b11111111111111111010011001100001;
assign LUT_4[7941] = 32'b11111111111111110011100101011001;
assign LUT_4[7942] = 32'b11111111111111111001110100000101;
assign LUT_4[7943] = 32'b11111111111111110010111111111101;
assign LUT_4[7944] = 32'b11111111111111110110100101011010;
assign LUT_4[7945] = 32'b11111111111111101111110001010010;
assign LUT_4[7946] = 32'b11111111111111110101111111111110;
assign LUT_4[7947] = 32'b11111111111111101111001011110110;
assign LUT_4[7948] = 32'b11111111111111110011100101110110;
assign LUT_4[7949] = 32'b11111111111111101100110001101110;
assign LUT_4[7950] = 32'b11111111111111110011000000011010;
assign LUT_4[7951] = 32'b11111111111111101100001100010010;
assign LUT_4[7952] = 32'b11111111111111111011001010110011;
assign LUT_4[7953] = 32'b11111111111111110100010110101011;
assign LUT_4[7954] = 32'b11111111111111111010100101010111;
assign LUT_4[7955] = 32'b11111111111111110011110001001111;
assign LUT_4[7956] = 32'b11111111111111111000001011001111;
assign LUT_4[7957] = 32'b11111111111111110001010111000111;
assign LUT_4[7958] = 32'b11111111111111110111100101110011;
assign LUT_4[7959] = 32'b11111111111111110000110001101011;
assign LUT_4[7960] = 32'b11111111111111110100010111001000;
assign LUT_4[7961] = 32'b11111111111111101101100011000000;
assign LUT_4[7962] = 32'b11111111111111110011110001101100;
assign LUT_4[7963] = 32'b11111111111111101100111101100100;
assign LUT_4[7964] = 32'b11111111111111110001010111100100;
assign LUT_4[7965] = 32'b11111111111111101010100011011100;
assign LUT_4[7966] = 32'b11111111111111110000110010001000;
assign LUT_4[7967] = 32'b11111111111111101001111110000000;
assign LUT_4[7968] = 32'b11111111111111111011110100001100;
assign LUT_4[7969] = 32'b11111111111111110101000000000100;
assign LUT_4[7970] = 32'b11111111111111111011001110110000;
assign LUT_4[7971] = 32'b11111111111111110100011010101000;
assign LUT_4[7972] = 32'b11111111111111111000110100101000;
assign LUT_4[7973] = 32'b11111111111111110010000000100000;
assign LUT_4[7974] = 32'b11111111111111111000001111001100;
assign LUT_4[7975] = 32'b11111111111111110001011011000100;
assign LUT_4[7976] = 32'b11111111111111110101000000100001;
assign LUT_4[7977] = 32'b11111111111111101110001100011001;
assign LUT_4[7978] = 32'b11111111111111110100011011000101;
assign LUT_4[7979] = 32'b11111111111111101101100110111101;
assign LUT_4[7980] = 32'b11111111111111110010000000111101;
assign LUT_4[7981] = 32'b11111111111111101011001100110101;
assign LUT_4[7982] = 32'b11111111111111110001011011100001;
assign LUT_4[7983] = 32'b11111111111111101010100111011001;
assign LUT_4[7984] = 32'b11111111111111111001100101111010;
assign LUT_4[7985] = 32'b11111111111111110010110001110010;
assign LUT_4[7986] = 32'b11111111111111111001000000011110;
assign LUT_4[7987] = 32'b11111111111111110010001100010110;
assign LUT_4[7988] = 32'b11111111111111110110100110010110;
assign LUT_4[7989] = 32'b11111111111111101111110010001110;
assign LUT_4[7990] = 32'b11111111111111110110000000111010;
assign LUT_4[7991] = 32'b11111111111111101111001100110010;
assign LUT_4[7992] = 32'b11111111111111110010110010001111;
assign LUT_4[7993] = 32'b11111111111111101011111110000111;
assign LUT_4[7994] = 32'b11111111111111110010001100110011;
assign LUT_4[7995] = 32'b11111111111111101011011000101011;
assign LUT_4[7996] = 32'b11111111111111101111110010101011;
assign LUT_4[7997] = 32'b11111111111111101000111110100011;
assign LUT_4[7998] = 32'b11111111111111101111001101001111;
assign LUT_4[7999] = 32'b11111111111111101000011001000111;
assign LUT_4[8000] = 32'b11111111111111111110110000011001;
assign LUT_4[8001] = 32'b11111111111111110111111100010001;
assign LUT_4[8002] = 32'b11111111111111111110001010111101;
assign LUT_4[8003] = 32'b11111111111111110111010110110101;
assign LUT_4[8004] = 32'b11111111111111111011110000110101;
assign LUT_4[8005] = 32'b11111111111111110100111100101101;
assign LUT_4[8006] = 32'b11111111111111111011001011011001;
assign LUT_4[8007] = 32'b11111111111111110100010111010001;
assign LUT_4[8008] = 32'b11111111111111110111111100101110;
assign LUT_4[8009] = 32'b11111111111111110001001000100110;
assign LUT_4[8010] = 32'b11111111111111110111010111010010;
assign LUT_4[8011] = 32'b11111111111111110000100011001010;
assign LUT_4[8012] = 32'b11111111111111110100111101001010;
assign LUT_4[8013] = 32'b11111111111111101110001001000010;
assign LUT_4[8014] = 32'b11111111111111110100010111101110;
assign LUT_4[8015] = 32'b11111111111111101101100011100110;
assign LUT_4[8016] = 32'b11111111111111111100100010000111;
assign LUT_4[8017] = 32'b11111111111111110101101101111111;
assign LUT_4[8018] = 32'b11111111111111111011111100101011;
assign LUT_4[8019] = 32'b11111111111111110101001000100011;
assign LUT_4[8020] = 32'b11111111111111111001100010100011;
assign LUT_4[8021] = 32'b11111111111111110010101110011011;
assign LUT_4[8022] = 32'b11111111111111111000111101000111;
assign LUT_4[8023] = 32'b11111111111111110010001000111111;
assign LUT_4[8024] = 32'b11111111111111110101101110011100;
assign LUT_4[8025] = 32'b11111111111111101110111010010100;
assign LUT_4[8026] = 32'b11111111111111110101001001000000;
assign LUT_4[8027] = 32'b11111111111111101110010100111000;
assign LUT_4[8028] = 32'b11111111111111110010101110111000;
assign LUT_4[8029] = 32'b11111111111111101011111010110000;
assign LUT_4[8030] = 32'b11111111111111110010001001011100;
assign LUT_4[8031] = 32'b11111111111111101011010101010100;
assign LUT_4[8032] = 32'b11111111111111111101001011100000;
assign LUT_4[8033] = 32'b11111111111111110110010111011000;
assign LUT_4[8034] = 32'b11111111111111111100100110000100;
assign LUT_4[8035] = 32'b11111111111111110101110001111100;
assign LUT_4[8036] = 32'b11111111111111111010001011111100;
assign LUT_4[8037] = 32'b11111111111111110011010111110100;
assign LUT_4[8038] = 32'b11111111111111111001100110100000;
assign LUT_4[8039] = 32'b11111111111111110010110010011000;
assign LUT_4[8040] = 32'b11111111111111110110010111110101;
assign LUT_4[8041] = 32'b11111111111111101111100011101101;
assign LUT_4[8042] = 32'b11111111111111110101110010011001;
assign LUT_4[8043] = 32'b11111111111111101110111110010001;
assign LUT_4[8044] = 32'b11111111111111110011011000010001;
assign LUT_4[8045] = 32'b11111111111111101100100100001001;
assign LUT_4[8046] = 32'b11111111111111110010110010110101;
assign LUT_4[8047] = 32'b11111111111111101011111110101101;
assign LUT_4[8048] = 32'b11111111111111111010111101001110;
assign LUT_4[8049] = 32'b11111111111111110100001001000110;
assign LUT_4[8050] = 32'b11111111111111111010010111110010;
assign LUT_4[8051] = 32'b11111111111111110011100011101010;
assign LUT_4[8052] = 32'b11111111111111110111111101101010;
assign LUT_4[8053] = 32'b11111111111111110001001001100010;
assign LUT_4[8054] = 32'b11111111111111110111011000001110;
assign LUT_4[8055] = 32'b11111111111111110000100100000110;
assign LUT_4[8056] = 32'b11111111111111110100001001100011;
assign LUT_4[8057] = 32'b11111111111111101101010101011011;
assign LUT_4[8058] = 32'b11111111111111110011100100000111;
assign LUT_4[8059] = 32'b11111111111111101100101111111111;
assign LUT_4[8060] = 32'b11111111111111110001001001111111;
assign LUT_4[8061] = 32'b11111111111111101010010101110111;
assign LUT_4[8062] = 32'b11111111111111110000100100100011;
assign LUT_4[8063] = 32'b11111111111111101001110000011011;
assign LUT_4[8064] = 32'b11111111111111111111111111001101;
assign LUT_4[8065] = 32'b11111111111111111001001011000101;
assign LUT_4[8066] = 32'b11111111111111111111011001110001;
assign LUT_4[8067] = 32'b11111111111111111000100101101001;
assign LUT_4[8068] = 32'b11111111111111111100111111101001;
assign LUT_4[8069] = 32'b11111111111111110110001011100001;
assign LUT_4[8070] = 32'b11111111111111111100011010001101;
assign LUT_4[8071] = 32'b11111111111111110101100110000101;
assign LUT_4[8072] = 32'b11111111111111111001001011100010;
assign LUT_4[8073] = 32'b11111111111111110010010111011010;
assign LUT_4[8074] = 32'b11111111111111111000100110000110;
assign LUT_4[8075] = 32'b11111111111111110001110001111110;
assign LUT_4[8076] = 32'b11111111111111110110001011111110;
assign LUT_4[8077] = 32'b11111111111111101111010111110110;
assign LUT_4[8078] = 32'b11111111111111110101100110100010;
assign LUT_4[8079] = 32'b11111111111111101110110010011010;
assign LUT_4[8080] = 32'b11111111111111111101110000111011;
assign LUT_4[8081] = 32'b11111111111111110110111100110011;
assign LUT_4[8082] = 32'b11111111111111111101001011011111;
assign LUT_4[8083] = 32'b11111111111111110110010111010111;
assign LUT_4[8084] = 32'b11111111111111111010110001010111;
assign LUT_4[8085] = 32'b11111111111111110011111101001111;
assign LUT_4[8086] = 32'b11111111111111111010001011111011;
assign LUT_4[8087] = 32'b11111111111111110011010111110011;
assign LUT_4[8088] = 32'b11111111111111110110111101010000;
assign LUT_4[8089] = 32'b11111111111111110000001001001000;
assign LUT_4[8090] = 32'b11111111111111110110010111110100;
assign LUT_4[8091] = 32'b11111111111111101111100011101100;
assign LUT_4[8092] = 32'b11111111111111110011111101101100;
assign LUT_4[8093] = 32'b11111111111111101101001001100100;
assign LUT_4[8094] = 32'b11111111111111110011011000010000;
assign LUT_4[8095] = 32'b11111111111111101100100100001000;
assign LUT_4[8096] = 32'b11111111111111111110011010010100;
assign LUT_4[8097] = 32'b11111111111111110111100110001100;
assign LUT_4[8098] = 32'b11111111111111111101110100111000;
assign LUT_4[8099] = 32'b11111111111111110111000000110000;
assign LUT_4[8100] = 32'b11111111111111111011011010110000;
assign LUT_4[8101] = 32'b11111111111111110100100110101000;
assign LUT_4[8102] = 32'b11111111111111111010110101010100;
assign LUT_4[8103] = 32'b11111111111111110100000001001100;
assign LUT_4[8104] = 32'b11111111111111110111100110101001;
assign LUT_4[8105] = 32'b11111111111111110000110010100001;
assign LUT_4[8106] = 32'b11111111111111110111000001001101;
assign LUT_4[8107] = 32'b11111111111111110000001101000101;
assign LUT_4[8108] = 32'b11111111111111110100100111000101;
assign LUT_4[8109] = 32'b11111111111111101101110010111101;
assign LUT_4[8110] = 32'b11111111111111110100000001101001;
assign LUT_4[8111] = 32'b11111111111111101101001101100001;
assign LUT_4[8112] = 32'b11111111111111111100001100000010;
assign LUT_4[8113] = 32'b11111111111111110101010111111010;
assign LUT_4[8114] = 32'b11111111111111111011100110100110;
assign LUT_4[8115] = 32'b11111111111111110100110010011110;
assign LUT_4[8116] = 32'b11111111111111111001001100011110;
assign LUT_4[8117] = 32'b11111111111111110010011000010110;
assign LUT_4[8118] = 32'b11111111111111111000100111000010;
assign LUT_4[8119] = 32'b11111111111111110001110010111010;
assign LUT_4[8120] = 32'b11111111111111110101011000010111;
assign LUT_4[8121] = 32'b11111111111111101110100100001111;
assign LUT_4[8122] = 32'b11111111111111110100110010111011;
assign LUT_4[8123] = 32'b11111111111111101101111110110011;
assign LUT_4[8124] = 32'b11111111111111110010011000110011;
assign LUT_4[8125] = 32'b11111111111111101011100100101011;
assign LUT_4[8126] = 32'b11111111111111110001110011010111;
assign LUT_4[8127] = 32'b11111111111111101010111111001111;
assign LUT_4[8128] = 32'b00000000000000000001010110100001;
assign LUT_4[8129] = 32'b11111111111111111010100010011001;
assign LUT_4[8130] = 32'b00000000000000000000110001000101;
assign LUT_4[8131] = 32'b11111111111111111001111100111101;
assign LUT_4[8132] = 32'b11111111111111111110010110111101;
assign LUT_4[8133] = 32'b11111111111111110111100010110101;
assign LUT_4[8134] = 32'b11111111111111111101110001100001;
assign LUT_4[8135] = 32'b11111111111111110110111101011001;
assign LUT_4[8136] = 32'b11111111111111111010100010110110;
assign LUT_4[8137] = 32'b11111111111111110011101110101110;
assign LUT_4[8138] = 32'b11111111111111111001111101011010;
assign LUT_4[8139] = 32'b11111111111111110011001001010010;
assign LUT_4[8140] = 32'b11111111111111110111100011010010;
assign LUT_4[8141] = 32'b11111111111111110000101111001010;
assign LUT_4[8142] = 32'b11111111111111110110111101110110;
assign LUT_4[8143] = 32'b11111111111111110000001001101110;
assign LUT_4[8144] = 32'b11111111111111111111001000001111;
assign LUT_4[8145] = 32'b11111111111111111000010100000111;
assign LUT_4[8146] = 32'b11111111111111111110100010110011;
assign LUT_4[8147] = 32'b11111111111111110111101110101011;
assign LUT_4[8148] = 32'b11111111111111111100001000101011;
assign LUT_4[8149] = 32'b11111111111111110101010100100011;
assign LUT_4[8150] = 32'b11111111111111111011100011001111;
assign LUT_4[8151] = 32'b11111111111111110100101111000111;
assign LUT_4[8152] = 32'b11111111111111111000010100100100;
assign LUT_4[8153] = 32'b11111111111111110001100000011100;
assign LUT_4[8154] = 32'b11111111111111110111101111001000;
assign LUT_4[8155] = 32'b11111111111111110000111011000000;
assign LUT_4[8156] = 32'b11111111111111110101010101000000;
assign LUT_4[8157] = 32'b11111111111111101110100000111000;
assign LUT_4[8158] = 32'b11111111111111110100101111100100;
assign LUT_4[8159] = 32'b11111111111111101101111011011100;
assign LUT_4[8160] = 32'b11111111111111111111110001101000;
assign LUT_4[8161] = 32'b11111111111111111000111101100000;
assign LUT_4[8162] = 32'b11111111111111111111001100001100;
assign LUT_4[8163] = 32'b11111111111111111000011000000100;
assign LUT_4[8164] = 32'b11111111111111111100110010000100;
assign LUT_4[8165] = 32'b11111111111111110101111101111100;
assign LUT_4[8166] = 32'b11111111111111111100001100101000;
assign LUT_4[8167] = 32'b11111111111111110101011000100000;
assign LUT_4[8168] = 32'b11111111111111111000111101111101;
assign LUT_4[8169] = 32'b11111111111111110010001001110101;
assign LUT_4[8170] = 32'b11111111111111111000011000100001;
assign LUT_4[8171] = 32'b11111111111111110001100100011001;
assign LUT_4[8172] = 32'b11111111111111110101111110011001;
assign LUT_4[8173] = 32'b11111111111111101111001010010001;
assign LUT_4[8174] = 32'b11111111111111110101011000111101;
assign LUT_4[8175] = 32'b11111111111111101110100100110101;
assign LUT_4[8176] = 32'b11111111111111111101100011010110;
assign LUT_4[8177] = 32'b11111111111111110110101111001110;
assign LUT_4[8178] = 32'b11111111111111111100111101111010;
assign LUT_4[8179] = 32'b11111111111111110110001001110010;
assign LUT_4[8180] = 32'b11111111111111111010100011110010;
assign LUT_4[8181] = 32'b11111111111111110011101111101010;
assign LUT_4[8182] = 32'b11111111111111111001111110010110;
assign LUT_4[8183] = 32'b11111111111111110011001010001110;
assign LUT_4[8184] = 32'b11111111111111110110101111101011;
assign LUT_4[8185] = 32'b11111111111111101111111011100011;
assign LUT_4[8186] = 32'b11111111111111110110001010001111;
assign LUT_4[8187] = 32'b11111111111111101111010110000111;
assign LUT_4[8188] = 32'b11111111111111110011110000000111;
assign LUT_4[8189] = 32'b11111111111111101100111011111111;
assign LUT_4[8190] = 32'b11111111111111110011001010101011;
assign LUT_4[8191] = 32'b11111111111111101100010110100011;
assign LUT_4[8192] = 32'b00000000000000000110001111001100;
assign LUT_4[8193] = 32'b11111111111111111111011011000100;
assign LUT_4[8194] = 32'b00000000000000000101101001110000;
assign LUT_4[8195] = 32'b11111111111111111110110101101000;
assign LUT_4[8196] = 32'b00000000000000000011001111101000;
assign LUT_4[8197] = 32'b11111111111111111100011011100000;
assign LUT_4[8198] = 32'b00000000000000000010101010001100;
assign LUT_4[8199] = 32'b11111111111111111011110110000100;
assign LUT_4[8200] = 32'b11111111111111111111011011100001;
assign LUT_4[8201] = 32'b11111111111111111000100111011001;
assign LUT_4[8202] = 32'b11111111111111111110110110000101;
assign LUT_4[8203] = 32'b11111111111111111000000001111101;
assign LUT_4[8204] = 32'b11111111111111111100011011111101;
assign LUT_4[8205] = 32'b11111111111111110101100111110101;
assign LUT_4[8206] = 32'b11111111111111111011110110100001;
assign LUT_4[8207] = 32'b11111111111111110101000010011001;
assign LUT_4[8208] = 32'b00000000000000000100000000111010;
assign LUT_4[8209] = 32'b11111111111111111101001100110010;
assign LUT_4[8210] = 32'b00000000000000000011011011011110;
assign LUT_4[8211] = 32'b11111111111111111100100111010110;
assign LUT_4[8212] = 32'b00000000000000000001000001010110;
assign LUT_4[8213] = 32'b11111111111111111010001101001110;
assign LUT_4[8214] = 32'b00000000000000000000011011111010;
assign LUT_4[8215] = 32'b11111111111111111001100111110010;
assign LUT_4[8216] = 32'b11111111111111111101001101001111;
assign LUT_4[8217] = 32'b11111111111111110110011001000111;
assign LUT_4[8218] = 32'b11111111111111111100100111110011;
assign LUT_4[8219] = 32'b11111111111111110101110011101011;
assign LUT_4[8220] = 32'b11111111111111111010001101101011;
assign LUT_4[8221] = 32'b11111111111111110011011001100011;
assign LUT_4[8222] = 32'b11111111111111111001101000001111;
assign LUT_4[8223] = 32'b11111111111111110010110100000111;
assign LUT_4[8224] = 32'b00000000000000000100101010010011;
assign LUT_4[8225] = 32'b11111111111111111101110110001011;
assign LUT_4[8226] = 32'b00000000000000000100000100110111;
assign LUT_4[8227] = 32'b11111111111111111101010000101111;
assign LUT_4[8228] = 32'b00000000000000000001101010101111;
assign LUT_4[8229] = 32'b11111111111111111010110110100111;
assign LUT_4[8230] = 32'b00000000000000000001000101010011;
assign LUT_4[8231] = 32'b11111111111111111010010001001011;
assign LUT_4[8232] = 32'b11111111111111111101110110101000;
assign LUT_4[8233] = 32'b11111111111111110111000010100000;
assign LUT_4[8234] = 32'b11111111111111111101010001001100;
assign LUT_4[8235] = 32'b11111111111111110110011101000100;
assign LUT_4[8236] = 32'b11111111111111111010110111000100;
assign LUT_4[8237] = 32'b11111111111111110100000010111100;
assign LUT_4[8238] = 32'b11111111111111111010010001101000;
assign LUT_4[8239] = 32'b11111111111111110011011101100000;
assign LUT_4[8240] = 32'b00000000000000000010011100000001;
assign LUT_4[8241] = 32'b11111111111111111011100111111001;
assign LUT_4[8242] = 32'b00000000000000000001110110100101;
assign LUT_4[8243] = 32'b11111111111111111011000010011101;
assign LUT_4[8244] = 32'b11111111111111111111011100011101;
assign LUT_4[8245] = 32'b11111111111111111000101000010101;
assign LUT_4[8246] = 32'b11111111111111111110110111000001;
assign LUT_4[8247] = 32'b11111111111111111000000010111001;
assign LUT_4[8248] = 32'b11111111111111111011101000010110;
assign LUT_4[8249] = 32'b11111111111111110100110100001110;
assign LUT_4[8250] = 32'b11111111111111111011000010111010;
assign LUT_4[8251] = 32'b11111111111111110100001110110010;
assign LUT_4[8252] = 32'b11111111111111111000101000110010;
assign LUT_4[8253] = 32'b11111111111111110001110100101010;
assign LUT_4[8254] = 32'b11111111111111111000000011010110;
assign LUT_4[8255] = 32'b11111111111111110001001111001110;
assign LUT_4[8256] = 32'b00000000000000000111100110100000;
assign LUT_4[8257] = 32'b00000000000000000000110010011000;
assign LUT_4[8258] = 32'b00000000000000000111000001000100;
assign LUT_4[8259] = 32'b00000000000000000000001100111100;
assign LUT_4[8260] = 32'b00000000000000000100100110111100;
assign LUT_4[8261] = 32'b11111111111111111101110010110100;
assign LUT_4[8262] = 32'b00000000000000000100000001100000;
assign LUT_4[8263] = 32'b11111111111111111101001101011000;
assign LUT_4[8264] = 32'b00000000000000000000110010110101;
assign LUT_4[8265] = 32'b11111111111111111001111110101101;
assign LUT_4[8266] = 32'b00000000000000000000001101011001;
assign LUT_4[8267] = 32'b11111111111111111001011001010001;
assign LUT_4[8268] = 32'b11111111111111111101110011010001;
assign LUT_4[8269] = 32'b11111111111111110110111111001001;
assign LUT_4[8270] = 32'b11111111111111111101001101110101;
assign LUT_4[8271] = 32'b11111111111111110110011001101101;
assign LUT_4[8272] = 32'b00000000000000000101011000001110;
assign LUT_4[8273] = 32'b11111111111111111110100100000110;
assign LUT_4[8274] = 32'b00000000000000000100110010110010;
assign LUT_4[8275] = 32'b11111111111111111101111110101010;
assign LUT_4[8276] = 32'b00000000000000000010011000101010;
assign LUT_4[8277] = 32'b11111111111111111011100100100010;
assign LUT_4[8278] = 32'b00000000000000000001110011001110;
assign LUT_4[8279] = 32'b11111111111111111010111111000110;
assign LUT_4[8280] = 32'b11111111111111111110100100100011;
assign LUT_4[8281] = 32'b11111111111111110111110000011011;
assign LUT_4[8282] = 32'b11111111111111111101111111000111;
assign LUT_4[8283] = 32'b11111111111111110111001010111111;
assign LUT_4[8284] = 32'b11111111111111111011100100111111;
assign LUT_4[8285] = 32'b11111111111111110100110000110111;
assign LUT_4[8286] = 32'b11111111111111111010111111100011;
assign LUT_4[8287] = 32'b11111111111111110100001011011011;
assign LUT_4[8288] = 32'b00000000000000000110000001100111;
assign LUT_4[8289] = 32'b11111111111111111111001101011111;
assign LUT_4[8290] = 32'b00000000000000000101011100001011;
assign LUT_4[8291] = 32'b11111111111111111110101000000011;
assign LUT_4[8292] = 32'b00000000000000000011000010000011;
assign LUT_4[8293] = 32'b11111111111111111100001101111011;
assign LUT_4[8294] = 32'b00000000000000000010011100100111;
assign LUT_4[8295] = 32'b11111111111111111011101000011111;
assign LUT_4[8296] = 32'b11111111111111111111001101111100;
assign LUT_4[8297] = 32'b11111111111111111000011001110100;
assign LUT_4[8298] = 32'b11111111111111111110101000100000;
assign LUT_4[8299] = 32'b11111111111111110111110100011000;
assign LUT_4[8300] = 32'b11111111111111111100001110011000;
assign LUT_4[8301] = 32'b11111111111111110101011010010000;
assign LUT_4[8302] = 32'b11111111111111111011101000111100;
assign LUT_4[8303] = 32'b11111111111111110100110100110100;
assign LUT_4[8304] = 32'b00000000000000000011110011010101;
assign LUT_4[8305] = 32'b11111111111111111100111111001101;
assign LUT_4[8306] = 32'b00000000000000000011001101111001;
assign LUT_4[8307] = 32'b11111111111111111100011001110001;
assign LUT_4[8308] = 32'b00000000000000000000110011110001;
assign LUT_4[8309] = 32'b11111111111111111001111111101001;
assign LUT_4[8310] = 32'b00000000000000000000001110010101;
assign LUT_4[8311] = 32'b11111111111111111001011010001101;
assign LUT_4[8312] = 32'b11111111111111111100111111101010;
assign LUT_4[8313] = 32'b11111111111111110110001011100010;
assign LUT_4[8314] = 32'b11111111111111111100011010001110;
assign LUT_4[8315] = 32'b11111111111111110101100110000110;
assign LUT_4[8316] = 32'b11111111111111111010000000000110;
assign LUT_4[8317] = 32'b11111111111111110011001011111110;
assign LUT_4[8318] = 32'b11111111111111111001011010101010;
assign LUT_4[8319] = 32'b11111111111111110010100110100010;
assign LUT_4[8320] = 32'b00000000000000001000110101010100;
assign LUT_4[8321] = 32'b00000000000000000010000001001100;
assign LUT_4[8322] = 32'b00000000000000001000001111111000;
assign LUT_4[8323] = 32'b00000000000000000001011011110000;
assign LUT_4[8324] = 32'b00000000000000000101110101110000;
assign LUT_4[8325] = 32'b11111111111111111111000001101000;
assign LUT_4[8326] = 32'b00000000000000000101010000010100;
assign LUT_4[8327] = 32'b11111111111111111110011100001100;
assign LUT_4[8328] = 32'b00000000000000000010000001101001;
assign LUT_4[8329] = 32'b11111111111111111011001101100001;
assign LUT_4[8330] = 32'b00000000000000000001011100001101;
assign LUT_4[8331] = 32'b11111111111111111010101000000101;
assign LUT_4[8332] = 32'b11111111111111111111000010000101;
assign LUT_4[8333] = 32'b11111111111111111000001101111101;
assign LUT_4[8334] = 32'b11111111111111111110011100101001;
assign LUT_4[8335] = 32'b11111111111111110111101000100001;
assign LUT_4[8336] = 32'b00000000000000000110100111000010;
assign LUT_4[8337] = 32'b11111111111111111111110010111010;
assign LUT_4[8338] = 32'b00000000000000000110000001100110;
assign LUT_4[8339] = 32'b11111111111111111111001101011110;
assign LUT_4[8340] = 32'b00000000000000000011100111011110;
assign LUT_4[8341] = 32'b11111111111111111100110011010110;
assign LUT_4[8342] = 32'b00000000000000000011000010000010;
assign LUT_4[8343] = 32'b11111111111111111100001101111010;
assign LUT_4[8344] = 32'b11111111111111111111110011010111;
assign LUT_4[8345] = 32'b11111111111111111000111111001111;
assign LUT_4[8346] = 32'b11111111111111111111001101111011;
assign LUT_4[8347] = 32'b11111111111111111000011001110011;
assign LUT_4[8348] = 32'b11111111111111111100110011110011;
assign LUT_4[8349] = 32'b11111111111111110101111111101011;
assign LUT_4[8350] = 32'b11111111111111111100001110010111;
assign LUT_4[8351] = 32'b11111111111111110101011010001111;
assign LUT_4[8352] = 32'b00000000000000000111010000011011;
assign LUT_4[8353] = 32'b00000000000000000000011100010011;
assign LUT_4[8354] = 32'b00000000000000000110101010111111;
assign LUT_4[8355] = 32'b11111111111111111111110110110111;
assign LUT_4[8356] = 32'b00000000000000000100010000110111;
assign LUT_4[8357] = 32'b11111111111111111101011100101111;
assign LUT_4[8358] = 32'b00000000000000000011101011011011;
assign LUT_4[8359] = 32'b11111111111111111100110111010011;
assign LUT_4[8360] = 32'b00000000000000000000011100110000;
assign LUT_4[8361] = 32'b11111111111111111001101000101000;
assign LUT_4[8362] = 32'b11111111111111111111110111010100;
assign LUT_4[8363] = 32'b11111111111111111001000011001100;
assign LUT_4[8364] = 32'b11111111111111111101011101001100;
assign LUT_4[8365] = 32'b11111111111111110110101001000100;
assign LUT_4[8366] = 32'b11111111111111111100110111110000;
assign LUT_4[8367] = 32'b11111111111111110110000011101000;
assign LUT_4[8368] = 32'b00000000000000000101000010001001;
assign LUT_4[8369] = 32'b11111111111111111110001110000001;
assign LUT_4[8370] = 32'b00000000000000000100011100101101;
assign LUT_4[8371] = 32'b11111111111111111101101000100101;
assign LUT_4[8372] = 32'b00000000000000000010000010100101;
assign LUT_4[8373] = 32'b11111111111111111011001110011101;
assign LUT_4[8374] = 32'b00000000000000000001011101001001;
assign LUT_4[8375] = 32'b11111111111111111010101001000001;
assign LUT_4[8376] = 32'b11111111111111111110001110011110;
assign LUT_4[8377] = 32'b11111111111111110111011010010110;
assign LUT_4[8378] = 32'b11111111111111111101101001000010;
assign LUT_4[8379] = 32'b11111111111111110110110100111010;
assign LUT_4[8380] = 32'b11111111111111111011001110111010;
assign LUT_4[8381] = 32'b11111111111111110100011010110010;
assign LUT_4[8382] = 32'b11111111111111111010101001011110;
assign LUT_4[8383] = 32'b11111111111111110011110101010110;
assign LUT_4[8384] = 32'b00000000000000001010001100101000;
assign LUT_4[8385] = 32'b00000000000000000011011000100000;
assign LUT_4[8386] = 32'b00000000000000001001100111001100;
assign LUT_4[8387] = 32'b00000000000000000010110011000100;
assign LUT_4[8388] = 32'b00000000000000000111001101000100;
assign LUT_4[8389] = 32'b00000000000000000000011000111100;
assign LUT_4[8390] = 32'b00000000000000000110100111101000;
assign LUT_4[8391] = 32'b11111111111111111111110011100000;
assign LUT_4[8392] = 32'b00000000000000000011011000111101;
assign LUT_4[8393] = 32'b11111111111111111100100100110101;
assign LUT_4[8394] = 32'b00000000000000000010110011100001;
assign LUT_4[8395] = 32'b11111111111111111011111111011001;
assign LUT_4[8396] = 32'b00000000000000000000011001011001;
assign LUT_4[8397] = 32'b11111111111111111001100101010001;
assign LUT_4[8398] = 32'b11111111111111111111110011111101;
assign LUT_4[8399] = 32'b11111111111111111000111111110101;
assign LUT_4[8400] = 32'b00000000000000000111111110010110;
assign LUT_4[8401] = 32'b00000000000000000001001010001110;
assign LUT_4[8402] = 32'b00000000000000000111011000111010;
assign LUT_4[8403] = 32'b00000000000000000000100100110010;
assign LUT_4[8404] = 32'b00000000000000000100111110110010;
assign LUT_4[8405] = 32'b11111111111111111110001010101010;
assign LUT_4[8406] = 32'b00000000000000000100011001010110;
assign LUT_4[8407] = 32'b11111111111111111101100101001110;
assign LUT_4[8408] = 32'b00000000000000000001001010101011;
assign LUT_4[8409] = 32'b11111111111111111010010110100011;
assign LUT_4[8410] = 32'b00000000000000000000100101001111;
assign LUT_4[8411] = 32'b11111111111111111001110001000111;
assign LUT_4[8412] = 32'b11111111111111111110001011000111;
assign LUT_4[8413] = 32'b11111111111111110111010110111111;
assign LUT_4[8414] = 32'b11111111111111111101100101101011;
assign LUT_4[8415] = 32'b11111111111111110110110001100011;
assign LUT_4[8416] = 32'b00000000000000001000100111101111;
assign LUT_4[8417] = 32'b00000000000000000001110011100111;
assign LUT_4[8418] = 32'b00000000000000001000000010010011;
assign LUT_4[8419] = 32'b00000000000000000001001110001011;
assign LUT_4[8420] = 32'b00000000000000000101101000001011;
assign LUT_4[8421] = 32'b11111111111111111110110100000011;
assign LUT_4[8422] = 32'b00000000000000000101000010101111;
assign LUT_4[8423] = 32'b11111111111111111110001110100111;
assign LUT_4[8424] = 32'b00000000000000000001110100000100;
assign LUT_4[8425] = 32'b11111111111111111010111111111100;
assign LUT_4[8426] = 32'b00000000000000000001001110101000;
assign LUT_4[8427] = 32'b11111111111111111010011010100000;
assign LUT_4[8428] = 32'b11111111111111111110110100100000;
assign LUT_4[8429] = 32'b11111111111111111000000000011000;
assign LUT_4[8430] = 32'b11111111111111111110001111000100;
assign LUT_4[8431] = 32'b11111111111111110111011010111100;
assign LUT_4[8432] = 32'b00000000000000000110011001011101;
assign LUT_4[8433] = 32'b11111111111111111111100101010101;
assign LUT_4[8434] = 32'b00000000000000000101110100000001;
assign LUT_4[8435] = 32'b11111111111111111110111111111001;
assign LUT_4[8436] = 32'b00000000000000000011011001111001;
assign LUT_4[8437] = 32'b11111111111111111100100101110001;
assign LUT_4[8438] = 32'b00000000000000000010110100011101;
assign LUT_4[8439] = 32'b11111111111111111100000000010101;
assign LUT_4[8440] = 32'b11111111111111111111100101110010;
assign LUT_4[8441] = 32'b11111111111111111000110001101010;
assign LUT_4[8442] = 32'b11111111111111111111000000010110;
assign LUT_4[8443] = 32'b11111111111111111000001100001110;
assign LUT_4[8444] = 32'b11111111111111111100100110001110;
assign LUT_4[8445] = 32'b11111111111111110101110010000110;
assign LUT_4[8446] = 32'b11111111111111111100000000110010;
assign LUT_4[8447] = 32'b11111111111111110101001100101010;
assign LUT_4[8448] = 32'b00000000000000001011001010101111;
assign LUT_4[8449] = 32'b00000000000000000100010110100111;
assign LUT_4[8450] = 32'b00000000000000001010100101010011;
assign LUT_4[8451] = 32'b00000000000000000011110001001011;
assign LUT_4[8452] = 32'b00000000000000001000001011001011;
assign LUT_4[8453] = 32'b00000000000000000001010111000011;
assign LUT_4[8454] = 32'b00000000000000000111100101101111;
assign LUT_4[8455] = 32'b00000000000000000000110001100111;
assign LUT_4[8456] = 32'b00000000000000000100010111000100;
assign LUT_4[8457] = 32'b11111111111111111101100010111100;
assign LUT_4[8458] = 32'b00000000000000000011110001101000;
assign LUT_4[8459] = 32'b11111111111111111100111101100000;
assign LUT_4[8460] = 32'b00000000000000000001010111100000;
assign LUT_4[8461] = 32'b11111111111111111010100011011000;
assign LUT_4[8462] = 32'b00000000000000000000110010000100;
assign LUT_4[8463] = 32'b11111111111111111001111101111100;
assign LUT_4[8464] = 32'b00000000000000001000111100011101;
assign LUT_4[8465] = 32'b00000000000000000010001000010101;
assign LUT_4[8466] = 32'b00000000000000001000010111000001;
assign LUT_4[8467] = 32'b00000000000000000001100010111001;
assign LUT_4[8468] = 32'b00000000000000000101111100111001;
assign LUT_4[8469] = 32'b11111111111111111111001000110001;
assign LUT_4[8470] = 32'b00000000000000000101010111011101;
assign LUT_4[8471] = 32'b11111111111111111110100011010101;
assign LUT_4[8472] = 32'b00000000000000000010001000110010;
assign LUT_4[8473] = 32'b11111111111111111011010100101010;
assign LUT_4[8474] = 32'b00000000000000000001100011010110;
assign LUT_4[8475] = 32'b11111111111111111010101111001110;
assign LUT_4[8476] = 32'b11111111111111111111001001001110;
assign LUT_4[8477] = 32'b11111111111111111000010101000110;
assign LUT_4[8478] = 32'b11111111111111111110100011110010;
assign LUT_4[8479] = 32'b11111111111111110111101111101010;
assign LUT_4[8480] = 32'b00000000000000001001100101110110;
assign LUT_4[8481] = 32'b00000000000000000010110001101110;
assign LUT_4[8482] = 32'b00000000000000001001000000011010;
assign LUT_4[8483] = 32'b00000000000000000010001100010010;
assign LUT_4[8484] = 32'b00000000000000000110100110010010;
assign LUT_4[8485] = 32'b11111111111111111111110010001010;
assign LUT_4[8486] = 32'b00000000000000000110000000110110;
assign LUT_4[8487] = 32'b11111111111111111111001100101110;
assign LUT_4[8488] = 32'b00000000000000000010110010001011;
assign LUT_4[8489] = 32'b11111111111111111011111110000011;
assign LUT_4[8490] = 32'b00000000000000000010001100101111;
assign LUT_4[8491] = 32'b11111111111111111011011000100111;
assign LUT_4[8492] = 32'b11111111111111111111110010100111;
assign LUT_4[8493] = 32'b11111111111111111000111110011111;
assign LUT_4[8494] = 32'b11111111111111111111001101001011;
assign LUT_4[8495] = 32'b11111111111111111000011001000011;
assign LUT_4[8496] = 32'b00000000000000000111010111100100;
assign LUT_4[8497] = 32'b00000000000000000000100011011100;
assign LUT_4[8498] = 32'b00000000000000000110110010001000;
assign LUT_4[8499] = 32'b11111111111111111111111110000000;
assign LUT_4[8500] = 32'b00000000000000000100011000000000;
assign LUT_4[8501] = 32'b11111111111111111101100011111000;
assign LUT_4[8502] = 32'b00000000000000000011110010100100;
assign LUT_4[8503] = 32'b11111111111111111100111110011100;
assign LUT_4[8504] = 32'b00000000000000000000100011111001;
assign LUT_4[8505] = 32'b11111111111111111001101111110001;
assign LUT_4[8506] = 32'b11111111111111111111111110011101;
assign LUT_4[8507] = 32'b11111111111111111001001010010101;
assign LUT_4[8508] = 32'b11111111111111111101100100010101;
assign LUT_4[8509] = 32'b11111111111111110110110000001101;
assign LUT_4[8510] = 32'b11111111111111111100111110111001;
assign LUT_4[8511] = 32'b11111111111111110110001010110001;
assign LUT_4[8512] = 32'b00000000000000001100100010000011;
assign LUT_4[8513] = 32'b00000000000000000101101101111011;
assign LUT_4[8514] = 32'b00000000000000001011111100100111;
assign LUT_4[8515] = 32'b00000000000000000101001000011111;
assign LUT_4[8516] = 32'b00000000000000001001100010011111;
assign LUT_4[8517] = 32'b00000000000000000010101110010111;
assign LUT_4[8518] = 32'b00000000000000001000111101000011;
assign LUT_4[8519] = 32'b00000000000000000010001000111011;
assign LUT_4[8520] = 32'b00000000000000000101101110011000;
assign LUT_4[8521] = 32'b11111111111111111110111010010000;
assign LUT_4[8522] = 32'b00000000000000000101001000111100;
assign LUT_4[8523] = 32'b11111111111111111110010100110100;
assign LUT_4[8524] = 32'b00000000000000000010101110110100;
assign LUT_4[8525] = 32'b11111111111111111011111010101100;
assign LUT_4[8526] = 32'b00000000000000000010001001011000;
assign LUT_4[8527] = 32'b11111111111111111011010101010000;
assign LUT_4[8528] = 32'b00000000000000001010010011110001;
assign LUT_4[8529] = 32'b00000000000000000011011111101001;
assign LUT_4[8530] = 32'b00000000000000001001101110010101;
assign LUT_4[8531] = 32'b00000000000000000010111010001101;
assign LUT_4[8532] = 32'b00000000000000000111010100001101;
assign LUT_4[8533] = 32'b00000000000000000000100000000101;
assign LUT_4[8534] = 32'b00000000000000000110101110110001;
assign LUT_4[8535] = 32'b11111111111111111111111010101001;
assign LUT_4[8536] = 32'b00000000000000000011100000000110;
assign LUT_4[8537] = 32'b11111111111111111100101011111110;
assign LUT_4[8538] = 32'b00000000000000000010111010101010;
assign LUT_4[8539] = 32'b11111111111111111100000110100010;
assign LUT_4[8540] = 32'b00000000000000000000100000100010;
assign LUT_4[8541] = 32'b11111111111111111001101100011010;
assign LUT_4[8542] = 32'b11111111111111111111111011000110;
assign LUT_4[8543] = 32'b11111111111111111001000110111110;
assign LUT_4[8544] = 32'b00000000000000001010111101001010;
assign LUT_4[8545] = 32'b00000000000000000100001001000010;
assign LUT_4[8546] = 32'b00000000000000001010010111101110;
assign LUT_4[8547] = 32'b00000000000000000011100011100110;
assign LUT_4[8548] = 32'b00000000000000000111111101100110;
assign LUT_4[8549] = 32'b00000000000000000001001001011110;
assign LUT_4[8550] = 32'b00000000000000000111011000001010;
assign LUT_4[8551] = 32'b00000000000000000000100100000010;
assign LUT_4[8552] = 32'b00000000000000000100001001011111;
assign LUT_4[8553] = 32'b11111111111111111101010101010111;
assign LUT_4[8554] = 32'b00000000000000000011100100000011;
assign LUT_4[8555] = 32'b11111111111111111100101111111011;
assign LUT_4[8556] = 32'b00000000000000000001001001111011;
assign LUT_4[8557] = 32'b11111111111111111010010101110011;
assign LUT_4[8558] = 32'b00000000000000000000100100011111;
assign LUT_4[8559] = 32'b11111111111111111001110000010111;
assign LUT_4[8560] = 32'b00000000000000001000101110111000;
assign LUT_4[8561] = 32'b00000000000000000001111010110000;
assign LUT_4[8562] = 32'b00000000000000001000001001011100;
assign LUT_4[8563] = 32'b00000000000000000001010101010100;
assign LUT_4[8564] = 32'b00000000000000000101101111010100;
assign LUT_4[8565] = 32'b11111111111111111110111011001100;
assign LUT_4[8566] = 32'b00000000000000000101001001111000;
assign LUT_4[8567] = 32'b11111111111111111110010101110000;
assign LUT_4[8568] = 32'b00000000000000000001111011001101;
assign LUT_4[8569] = 32'b11111111111111111011000111000101;
assign LUT_4[8570] = 32'b00000000000000000001010101110001;
assign LUT_4[8571] = 32'b11111111111111111010100001101001;
assign LUT_4[8572] = 32'b11111111111111111110111011101001;
assign LUT_4[8573] = 32'b11111111111111111000000111100001;
assign LUT_4[8574] = 32'b11111111111111111110010110001101;
assign LUT_4[8575] = 32'b11111111111111110111100010000101;
assign LUT_4[8576] = 32'b00000000000000001101110000110111;
assign LUT_4[8577] = 32'b00000000000000000110111100101111;
assign LUT_4[8578] = 32'b00000000000000001101001011011011;
assign LUT_4[8579] = 32'b00000000000000000110010111010011;
assign LUT_4[8580] = 32'b00000000000000001010110001010011;
assign LUT_4[8581] = 32'b00000000000000000011111101001011;
assign LUT_4[8582] = 32'b00000000000000001010001011110111;
assign LUT_4[8583] = 32'b00000000000000000011010111101111;
assign LUT_4[8584] = 32'b00000000000000000110111101001100;
assign LUT_4[8585] = 32'b00000000000000000000001001000100;
assign LUT_4[8586] = 32'b00000000000000000110010111110000;
assign LUT_4[8587] = 32'b11111111111111111111100011101000;
assign LUT_4[8588] = 32'b00000000000000000011111101101000;
assign LUT_4[8589] = 32'b11111111111111111101001001100000;
assign LUT_4[8590] = 32'b00000000000000000011011000001100;
assign LUT_4[8591] = 32'b11111111111111111100100100000100;
assign LUT_4[8592] = 32'b00000000000000001011100010100101;
assign LUT_4[8593] = 32'b00000000000000000100101110011101;
assign LUT_4[8594] = 32'b00000000000000001010111101001001;
assign LUT_4[8595] = 32'b00000000000000000100001001000001;
assign LUT_4[8596] = 32'b00000000000000001000100011000001;
assign LUT_4[8597] = 32'b00000000000000000001101110111001;
assign LUT_4[8598] = 32'b00000000000000000111111101100101;
assign LUT_4[8599] = 32'b00000000000000000001001001011101;
assign LUT_4[8600] = 32'b00000000000000000100101110111010;
assign LUT_4[8601] = 32'b11111111111111111101111010110010;
assign LUT_4[8602] = 32'b00000000000000000100001001011110;
assign LUT_4[8603] = 32'b11111111111111111101010101010110;
assign LUT_4[8604] = 32'b00000000000000000001101111010110;
assign LUT_4[8605] = 32'b11111111111111111010111011001110;
assign LUT_4[8606] = 32'b00000000000000000001001001111010;
assign LUT_4[8607] = 32'b11111111111111111010010101110010;
assign LUT_4[8608] = 32'b00000000000000001100001011111110;
assign LUT_4[8609] = 32'b00000000000000000101010111110110;
assign LUT_4[8610] = 32'b00000000000000001011100110100010;
assign LUT_4[8611] = 32'b00000000000000000100110010011010;
assign LUT_4[8612] = 32'b00000000000000001001001100011010;
assign LUT_4[8613] = 32'b00000000000000000010011000010010;
assign LUT_4[8614] = 32'b00000000000000001000100110111110;
assign LUT_4[8615] = 32'b00000000000000000001110010110110;
assign LUT_4[8616] = 32'b00000000000000000101011000010011;
assign LUT_4[8617] = 32'b11111111111111111110100100001011;
assign LUT_4[8618] = 32'b00000000000000000100110010110111;
assign LUT_4[8619] = 32'b11111111111111111101111110101111;
assign LUT_4[8620] = 32'b00000000000000000010011000101111;
assign LUT_4[8621] = 32'b11111111111111111011100100100111;
assign LUT_4[8622] = 32'b00000000000000000001110011010011;
assign LUT_4[8623] = 32'b11111111111111111010111111001011;
assign LUT_4[8624] = 32'b00000000000000001001111101101100;
assign LUT_4[8625] = 32'b00000000000000000011001001100100;
assign LUT_4[8626] = 32'b00000000000000001001011000010000;
assign LUT_4[8627] = 32'b00000000000000000010100100001000;
assign LUT_4[8628] = 32'b00000000000000000110111110001000;
assign LUT_4[8629] = 32'b00000000000000000000001010000000;
assign LUT_4[8630] = 32'b00000000000000000110011000101100;
assign LUT_4[8631] = 32'b11111111111111111111100100100100;
assign LUT_4[8632] = 32'b00000000000000000011001010000001;
assign LUT_4[8633] = 32'b11111111111111111100010101111001;
assign LUT_4[8634] = 32'b00000000000000000010100100100101;
assign LUT_4[8635] = 32'b11111111111111111011110000011101;
assign LUT_4[8636] = 32'b00000000000000000000001010011101;
assign LUT_4[8637] = 32'b11111111111111111001010110010101;
assign LUT_4[8638] = 32'b11111111111111111111100101000001;
assign LUT_4[8639] = 32'b11111111111111111000110000111001;
assign LUT_4[8640] = 32'b00000000000000001111001000001011;
assign LUT_4[8641] = 32'b00000000000000001000010100000011;
assign LUT_4[8642] = 32'b00000000000000001110100010101111;
assign LUT_4[8643] = 32'b00000000000000000111101110100111;
assign LUT_4[8644] = 32'b00000000000000001100001000100111;
assign LUT_4[8645] = 32'b00000000000000000101010100011111;
assign LUT_4[8646] = 32'b00000000000000001011100011001011;
assign LUT_4[8647] = 32'b00000000000000000100101111000011;
assign LUT_4[8648] = 32'b00000000000000001000010100100000;
assign LUT_4[8649] = 32'b00000000000000000001100000011000;
assign LUT_4[8650] = 32'b00000000000000000111101111000100;
assign LUT_4[8651] = 32'b00000000000000000000111010111100;
assign LUT_4[8652] = 32'b00000000000000000101010100111100;
assign LUT_4[8653] = 32'b11111111111111111110100000110100;
assign LUT_4[8654] = 32'b00000000000000000100101111100000;
assign LUT_4[8655] = 32'b11111111111111111101111011011000;
assign LUT_4[8656] = 32'b00000000000000001100111001111001;
assign LUT_4[8657] = 32'b00000000000000000110000101110001;
assign LUT_4[8658] = 32'b00000000000000001100010100011101;
assign LUT_4[8659] = 32'b00000000000000000101100000010101;
assign LUT_4[8660] = 32'b00000000000000001001111010010101;
assign LUT_4[8661] = 32'b00000000000000000011000110001101;
assign LUT_4[8662] = 32'b00000000000000001001010100111001;
assign LUT_4[8663] = 32'b00000000000000000010100000110001;
assign LUT_4[8664] = 32'b00000000000000000110000110001110;
assign LUT_4[8665] = 32'b11111111111111111111010010000110;
assign LUT_4[8666] = 32'b00000000000000000101100000110010;
assign LUT_4[8667] = 32'b11111111111111111110101100101010;
assign LUT_4[8668] = 32'b00000000000000000011000110101010;
assign LUT_4[8669] = 32'b11111111111111111100010010100010;
assign LUT_4[8670] = 32'b00000000000000000010100001001110;
assign LUT_4[8671] = 32'b11111111111111111011101101000110;
assign LUT_4[8672] = 32'b00000000000000001101100011010010;
assign LUT_4[8673] = 32'b00000000000000000110101111001010;
assign LUT_4[8674] = 32'b00000000000000001100111101110110;
assign LUT_4[8675] = 32'b00000000000000000110001001101110;
assign LUT_4[8676] = 32'b00000000000000001010100011101110;
assign LUT_4[8677] = 32'b00000000000000000011101111100110;
assign LUT_4[8678] = 32'b00000000000000001001111110010010;
assign LUT_4[8679] = 32'b00000000000000000011001010001010;
assign LUT_4[8680] = 32'b00000000000000000110101111100111;
assign LUT_4[8681] = 32'b11111111111111111111111011011111;
assign LUT_4[8682] = 32'b00000000000000000110001010001011;
assign LUT_4[8683] = 32'b11111111111111111111010110000011;
assign LUT_4[8684] = 32'b00000000000000000011110000000011;
assign LUT_4[8685] = 32'b11111111111111111100111011111011;
assign LUT_4[8686] = 32'b00000000000000000011001010100111;
assign LUT_4[8687] = 32'b11111111111111111100010110011111;
assign LUT_4[8688] = 32'b00000000000000001011010101000000;
assign LUT_4[8689] = 32'b00000000000000000100100000111000;
assign LUT_4[8690] = 32'b00000000000000001010101111100100;
assign LUT_4[8691] = 32'b00000000000000000011111011011100;
assign LUT_4[8692] = 32'b00000000000000001000010101011100;
assign LUT_4[8693] = 32'b00000000000000000001100001010100;
assign LUT_4[8694] = 32'b00000000000000000111110000000000;
assign LUT_4[8695] = 32'b00000000000000000000111011111000;
assign LUT_4[8696] = 32'b00000000000000000100100001010101;
assign LUT_4[8697] = 32'b11111111111111111101101101001101;
assign LUT_4[8698] = 32'b00000000000000000011111011111001;
assign LUT_4[8699] = 32'b11111111111111111101000111110001;
assign LUT_4[8700] = 32'b00000000000000000001100001110001;
assign LUT_4[8701] = 32'b11111111111111111010101101101001;
assign LUT_4[8702] = 32'b00000000000000000000111100010101;
assign LUT_4[8703] = 32'b11111111111111111010001000001101;
assign LUT_4[8704] = 32'b00000000000000000101010011010100;
assign LUT_4[8705] = 32'b11111111111111111110011111001100;
assign LUT_4[8706] = 32'b00000000000000000100101101111000;
assign LUT_4[8707] = 32'b11111111111111111101111001110000;
assign LUT_4[8708] = 32'b00000000000000000010010011110000;
assign LUT_4[8709] = 32'b11111111111111111011011111101000;
assign LUT_4[8710] = 32'b00000000000000000001101110010100;
assign LUT_4[8711] = 32'b11111111111111111010111010001100;
assign LUT_4[8712] = 32'b11111111111111111110011111101001;
assign LUT_4[8713] = 32'b11111111111111110111101011100001;
assign LUT_4[8714] = 32'b11111111111111111101111010001101;
assign LUT_4[8715] = 32'b11111111111111110111000110000101;
assign LUT_4[8716] = 32'b11111111111111111011100000000101;
assign LUT_4[8717] = 32'b11111111111111110100101011111101;
assign LUT_4[8718] = 32'b11111111111111111010111010101001;
assign LUT_4[8719] = 32'b11111111111111110100000110100001;
assign LUT_4[8720] = 32'b00000000000000000011000101000010;
assign LUT_4[8721] = 32'b11111111111111111100010000111010;
assign LUT_4[8722] = 32'b00000000000000000010011111100110;
assign LUT_4[8723] = 32'b11111111111111111011101011011110;
assign LUT_4[8724] = 32'b00000000000000000000000101011110;
assign LUT_4[8725] = 32'b11111111111111111001010001010110;
assign LUT_4[8726] = 32'b11111111111111111111100000000010;
assign LUT_4[8727] = 32'b11111111111111111000101011111010;
assign LUT_4[8728] = 32'b11111111111111111100010001010111;
assign LUT_4[8729] = 32'b11111111111111110101011101001111;
assign LUT_4[8730] = 32'b11111111111111111011101011111011;
assign LUT_4[8731] = 32'b11111111111111110100110111110011;
assign LUT_4[8732] = 32'b11111111111111111001010001110011;
assign LUT_4[8733] = 32'b11111111111111110010011101101011;
assign LUT_4[8734] = 32'b11111111111111111000101100010111;
assign LUT_4[8735] = 32'b11111111111111110001111000001111;
assign LUT_4[8736] = 32'b00000000000000000011101110011011;
assign LUT_4[8737] = 32'b11111111111111111100111010010011;
assign LUT_4[8738] = 32'b00000000000000000011001000111111;
assign LUT_4[8739] = 32'b11111111111111111100010100110111;
assign LUT_4[8740] = 32'b00000000000000000000101110110111;
assign LUT_4[8741] = 32'b11111111111111111001111010101111;
assign LUT_4[8742] = 32'b00000000000000000000001001011011;
assign LUT_4[8743] = 32'b11111111111111111001010101010011;
assign LUT_4[8744] = 32'b11111111111111111100111010110000;
assign LUT_4[8745] = 32'b11111111111111110110000110101000;
assign LUT_4[8746] = 32'b11111111111111111100010101010100;
assign LUT_4[8747] = 32'b11111111111111110101100001001100;
assign LUT_4[8748] = 32'b11111111111111111001111011001100;
assign LUT_4[8749] = 32'b11111111111111110011000111000100;
assign LUT_4[8750] = 32'b11111111111111111001010101110000;
assign LUT_4[8751] = 32'b11111111111111110010100001101000;
assign LUT_4[8752] = 32'b00000000000000000001100000001001;
assign LUT_4[8753] = 32'b11111111111111111010101100000001;
assign LUT_4[8754] = 32'b00000000000000000000111010101101;
assign LUT_4[8755] = 32'b11111111111111111010000110100101;
assign LUT_4[8756] = 32'b11111111111111111110100000100101;
assign LUT_4[8757] = 32'b11111111111111110111101100011101;
assign LUT_4[8758] = 32'b11111111111111111101111011001001;
assign LUT_4[8759] = 32'b11111111111111110111000111000001;
assign LUT_4[8760] = 32'b11111111111111111010101100011110;
assign LUT_4[8761] = 32'b11111111111111110011111000010110;
assign LUT_4[8762] = 32'b11111111111111111010000111000010;
assign LUT_4[8763] = 32'b11111111111111110011010010111010;
assign LUT_4[8764] = 32'b11111111111111110111101100111010;
assign LUT_4[8765] = 32'b11111111111111110000111000110010;
assign LUT_4[8766] = 32'b11111111111111110111000111011110;
assign LUT_4[8767] = 32'b11111111111111110000010011010110;
assign LUT_4[8768] = 32'b00000000000000000110101010101000;
assign LUT_4[8769] = 32'b11111111111111111111110110100000;
assign LUT_4[8770] = 32'b00000000000000000110000101001100;
assign LUT_4[8771] = 32'b11111111111111111111010001000100;
assign LUT_4[8772] = 32'b00000000000000000011101011000100;
assign LUT_4[8773] = 32'b11111111111111111100110110111100;
assign LUT_4[8774] = 32'b00000000000000000011000101101000;
assign LUT_4[8775] = 32'b11111111111111111100010001100000;
assign LUT_4[8776] = 32'b11111111111111111111110110111101;
assign LUT_4[8777] = 32'b11111111111111111001000010110101;
assign LUT_4[8778] = 32'b11111111111111111111010001100001;
assign LUT_4[8779] = 32'b11111111111111111000011101011001;
assign LUT_4[8780] = 32'b11111111111111111100110111011001;
assign LUT_4[8781] = 32'b11111111111111110110000011010001;
assign LUT_4[8782] = 32'b11111111111111111100010001111101;
assign LUT_4[8783] = 32'b11111111111111110101011101110101;
assign LUT_4[8784] = 32'b00000000000000000100011100010110;
assign LUT_4[8785] = 32'b11111111111111111101101000001110;
assign LUT_4[8786] = 32'b00000000000000000011110110111010;
assign LUT_4[8787] = 32'b11111111111111111101000010110010;
assign LUT_4[8788] = 32'b00000000000000000001011100110010;
assign LUT_4[8789] = 32'b11111111111111111010101000101010;
assign LUT_4[8790] = 32'b00000000000000000000110111010110;
assign LUT_4[8791] = 32'b11111111111111111010000011001110;
assign LUT_4[8792] = 32'b11111111111111111101101000101011;
assign LUT_4[8793] = 32'b11111111111111110110110100100011;
assign LUT_4[8794] = 32'b11111111111111111101000011001111;
assign LUT_4[8795] = 32'b11111111111111110110001111000111;
assign LUT_4[8796] = 32'b11111111111111111010101001000111;
assign LUT_4[8797] = 32'b11111111111111110011110100111111;
assign LUT_4[8798] = 32'b11111111111111111010000011101011;
assign LUT_4[8799] = 32'b11111111111111110011001111100011;
assign LUT_4[8800] = 32'b00000000000000000101000101101111;
assign LUT_4[8801] = 32'b11111111111111111110010001100111;
assign LUT_4[8802] = 32'b00000000000000000100100000010011;
assign LUT_4[8803] = 32'b11111111111111111101101100001011;
assign LUT_4[8804] = 32'b00000000000000000010000110001011;
assign LUT_4[8805] = 32'b11111111111111111011010010000011;
assign LUT_4[8806] = 32'b00000000000000000001100000101111;
assign LUT_4[8807] = 32'b11111111111111111010101100100111;
assign LUT_4[8808] = 32'b11111111111111111110010010000100;
assign LUT_4[8809] = 32'b11111111111111110111011101111100;
assign LUT_4[8810] = 32'b11111111111111111101101100101000;
assign LUT_4[8811] = 32'b11111111111111110110111000100000;
assign LUT_4[8812] = 32'b11111111111111111011010010100000;
assign LUT_4[8813] = 32'b11111111111111110100011110011000;
assign LUT_4[8814] = 32'b11111111111111111010101101000100;
assign LUT_4[8815] = 32'b11111111111111110011111000111100;
assign LUT_4[8816] = 32'b00000000000000000010110111011101;
assign LUT_4[8817] = 32'b11111111111111111100000011010101;
assign LUT_4[8818] = 32'b00000000000000000010010010000001;
assign LUT_4[8819] = 32'b11111111111111111011011101111001;
assign LUT_4[8820] = 32'b11111111111111111111110111111001;
assign LUT_4[8821] = 32'b11111111111111111001000011110001;
assign LUT_4[8822] = 32'b11111111111111111111010010011101;
assign LUT_4[8823] = 32'b11111111111111111000011110010101;
assign LUT_4[8824] = 32'b11111111111111111100000011110010;
assign LUT_4[8825] = 32'b11111111111111110101001111101010;
assign LUT_4[8826] = 32'b11111111111111111011011110010110;
assign LUT_4[8827] = 32'b11111111111111110100101010001110;
assign LUT_4[8828] = 32'b11111111111111111001000100001110;
assign LUT_4[8829] = 32'b11111111111111110010010000000110;
assign LUT_4[8830] = 32'b11111111111111111000011110110010;
assign LUT_4[8831] = 32'b11111111111111110001101010101010;
assign LUT_4[8832] = 32'b00000000000000000111111001011100;
assign LUT_4[8833] = 32'b00000000000000000001000101010100;
assign LUT_4[8834] = 32'b00000000000000000111010100000000;
assign LUT_4[8835] = 32'b00000000000000000000011111111000;
assign LUT_4[8836] = 32'b00000000000000000100111001111000;
assign LUT_4[8837] = 32'b11111111111111111110000101110000;
assign LUT_4[8838] = 32'b00000000000000000100010100011100;
assign LUT_4[8839] = 32'b11111111111111111101100000010100;
assign LUT_4[8840] = 32'b00000000000000000001000101110001;
assign LUT_4[8841] = 32'b11111111111111111010010001101001;
assign LUT_4[8842] = 32'b00000000000000000000100000010101;
assign LUT_4[8843] = 32'b11111111111111111001101100001101;
assign LUT_4[8844] = 32'b11111111111111111110000110001101;
assign LUT_4[8845] = 32'b11111111111111110111010010000101;
assign LUT_4[8846] = 32'b11111111111111111101100000110001;
assign LUT_4[8847] = 32'b11111111111111110110101100101001;
assign LUT_4[8848] = 32'b00000000000000000101101011001010;
assign LUT_4[8849] = 32'b11111111111111111110110111000010;
assign LUT_4[8850] = 32'b00000000000000000101000101101110;
assign LUT_4[8851] = 32'b11111111111111111110010001100110;
assign LUT_4[8852] = 32'b00000000000000000010101011100110;
assign LUT_4[8853] = 32'b11111111111111111011110111011110;
assign LUT_4[8854] = 32'b00000000000000000010000110001010;
assign LUT_4[8855] = 32'b11111111111111111011010010000010;
assign LUT_4[8856] = 32'b11111111111111111110110111011111;
assign LUT_4[8857] = 32'b11111111111111111000000011010111;
assign LUT_4[8858] = 32'b11111111111111111110010010000011;
assign LUT_4[8859] = 32'b11111111111111110111011101111011;
assign LUT_4[8860] = 32'b11111111111111111011110111111011;
assign LUT_4[8861] = 32'b11111111111111110101000011110011;
assign LUT_4[8862] = 32'b11111111111111111011010010011111;
assign LUT_4[8863] = 32'b11111111111111110100011110010111;
assign LUT_4[8864] = 32'b00000000000000000110010100100011;
assign LUT_4[8865] = 32'b11111111111111111111100000011011;
assign LUT_4[8866] = 32'b00000000000000000101101111000111;
assign LUT_4[8867] = 32'b11111111111111111110111010111111;
assign LUT_4[8868] = 32'b00000000000000000011010100111111;
assign LUT_4[8869] = 32'b11111111111111111100100000110111;
assign LUT_4[8870] = 32'b00000000000000000010101111100011;
assign LUT_4[8871] = 32'b11111111111111111011111011011011;
assign LUT_4[8872] = 32'b11111111111111111111100000111000;
assign LUT_4[8873] = 32'b11111111111111111000101100110000;
assign LUT_4[8874] = 32'b11111111111111111110111011011100;
assign LUT_4[8875] = 32'b11111111111111111000000111010100;
assign LUT_4[8876] = 32'b11111111111111111100100001010100;
assign LUT_4[8877] = 32'b11111111111111110101101101001100;
assign LUT_4[8878] = 32'b11111111111111111011111011111000;
assign LUT_4[8879] = 32'b11111111111111110101000111110000;
assign LUT_4[8880] = 32'b00000000000000000100000110010001;
assign LUT_4[8881] = 32'b11111111111111111101010010001001;
assign LUT_4[8882] = 32'b00000000000000000011100000110101;
assign LUT_4[8883] = 32'b11111111111111111100101100101101;
assign LUT_4[8884] = 32'b00000000000000000001000110101101;
assign LUT_4[8885] = 32'b11111111111111111010010010100101;
assign LUT_4[8886] = 32'b00000000000000000000100001010001;
assign LUT_4[8887] = 32'b11111111111111111001101101001001;
assign LUT_4[8888] = 32'b11111111111111111101010010100110;
assign LUT_4[8889] = 32'b11111111111111110110011110011110;
assign LUT_4[8890] = 32'b11111111111111111100101101001010;
assign LUT_4[8891] = 32'b11111111111111110101111001000010;
assign LUT_4[8892] = 32'b11111111111111111010010011000010;
assign LUT_4[8893] = 32'b11111111111111110011011110111010;
assign LUT_4[8894] = 32'b11111111111111111001101101100110;
assign LUT_4[8895] = 32'b11111111111111110010111001011110;
assign LUT_4[8896] = 32'b00000000000000001001010000110000;
assign LUT_4[8897] = 32'b00000000000000000010011100101000;
assign LUT_4[8898] = 32'b00000000000000001000101011010100;
assign LUT_4[8899] = 32'b00000000000000000001110111001100;
assign LUT_4[8900] = 32'b00000000000000000110010001001100;
assign LUT_4[8901] = 32'b11111111111111111111011101000100;
assign LUT_4[8902] = 32'b00000000000000000101101011110000;
assign LUT_4[8903] = 32'b11111111111111111110110111101000;
assign LUT_4[8904] = 32'b00000000000000000010011101000101;
assign LUT_4[8905] = 32'b11111111111111111011101000111101;
assign LUT_4[8906] = 32'b00000000000000000001110111101001;
assign LUT_4[8907] = 32'b11111111111111111011000011100001;
assign LUT_4[8908] = 32'b11111111111111111111011101100001;
assign LUT_4[8909] = 32'b11111111111111111000101001011001;
assign LUT_4[8910] = 32'b11111111111111111110111000000101;
assign LUT_4[8911] = 32'b11111111111111111000000011111101;
assign LUT_4[8912] = 32'b00000000000000000111000010011110;
assign LUT_4[8913] = 32'b00000000000000000000001110010110;
assign LUT_4[8914] = 32'b00000000000000000110011101000010;
assign LUT_4[8915] = 32'b11111111111111111111101000111010;
assign LUT_4[8916] = 32'b00000000000000000100000010111010;
assign LUT_4[8917] = 32'b11111111111111111101001110110010;
assign LUT_4[8918] = 32'b00000000000000000011011101011110;
assign LUT_4[8919] = 32'b11111111111111111100101001010110;
assign LUT_4[8920] = 32'b00000000000000000000001110110011;
assign LUT_4[8921] = 32'b11111111111111111001011010101011;
assign LUT_4[8922] = 32'b11111111111111111111101001010111;
assign LUT_4[8923] = 32'b11111111111111111000110101001111;
assign LUT_4[8924] = 32'b11111111111111111101001111001111;
assign LUT_4[8925] = 32'b11111111111111110110011011000111;
assign LUT_4[8926] = 32'b11111111111111111100101001110011;
assign LUT_4[8927] = 32'b11111111111111110101110101101011;
assign LUT_4[8928] = 32'b00000000000000000111101011110111;
assign LUT_4[8929] = 32'b00000000000000000000110111101111;
assign LUT_4[8930] = 32'b00000000000000000111000110011011;
assign LUT_4[8931] = 32'b00000000000000000000010010010011;
assign LUT_4[8932] = 32'b00000000000000000100101100010011;
assign LUT_4[8933] = 32'b11111111111111111101111000001011;
assign LUT_4[8934] = 32'b00000000000000000100000110110111;
assign LUT_4[8935] = 32'b11111111111111111101010010101111;
assign LUT_4[8936] = 32'b00000000000000000000111000001100;
assign LUT_4[8937] = 32'b11111111111111111010000100000100;
assign LUT_4[8938] = 32'b00000000000000000000010010110000;
assign LUT_4[8939] = 32'b11111111111111111001011110101000;
assign LUT_4[8940] = 32'b11111111111111111101111000101000;
assign LUT_4[8941] = 32'b11111111111111110111000100100000;
assign LUT_4[8942] = 32'b11111111111111111101010011001100;
assign LUT_4[8943] = 32'b11111111111111110110011111000100;
assign LUT_4[8944] = 32'b00000000000000000101011101100101;
assign LUT_4[8945] = 32'b11111111111111111110101001011101;
assign LUT_4[8946] = 32'b00000000000000000100111000001001;
assign LUT_4[8947] = 32'b11111111111111111110000100000001;
assign LUT_4[8948] = 32'b00000000000000000010011110000001;
assign LUT_4[8949] = 32'b11111111111111111011101001111001;
assign LUT_4[8950] = 32'b00000000000000000001111000100101;
assign LUT_4[8951] = 32'b11111111111111111011000100011101;
assign LUT_4[8952] = 32'b11111111111111111110101001111010;
assign LUT_4[8953] = 32'b11111111111111110111110101110010;
assign LUT_4[8954] = 32'b11111111111111111110000100011110;
assign LUT_4[8955] = 32'b11111111111111110111010000010110;
assign LUT_4[8956] = 32'b11111111111111111011101010010110;
assign LUT_4[8957] = 32'b11111111111111110100110110001110;
assign LUT_4[8958] = 32'b11111111111111111011000100111010;
assign LUT_4[8959] = 32'b11111111111111110100010000110010;
assign LUT_4[8960] = 32'b00000000000000001010001110110111;
assign LUT_4[8961] = 32'b00000000000000000011011010101111;
assign LUT_4[8962] = 32'b00000000000000001001101001011011;
assign LUT_4[8963] = 32'b00000000000000000010110101010011;
assign LUT_4[8964] = 32'b00000000000000000111001111010011;
assign LUT_4[8965] = 32'b00000000000000000000011011001011;
assign LUT_4[8966] = 32'b00000000000000000110101001110111;
assign LUT_4[8967] = 32'b11111111111111111111110101101111;
assign LUT_4[8968] = 32'b00000000000000000011011011001100;
assign LUT_4[8969] = 32'b11111111111111111100100111000100;
assign LUT_4[8970] = 32'b00000000000000000010110101110000;
assign LUT_4[8971] = 32'b11111111111111111100000001101000;
assign LUT_4[8972] = 32'b00000000000000000000011011101000;
assign LUT_4[8973] = 32'b11111111111111111001100111100000;
assign LUT_4[8974] = 32'b11111111111111111111110110001100;
assign LUT_4[8975] = 32'b11111111111111111001000010000100;
assign LUT_4[8976] = 32'b00000000000000001000000000100101;
assign LUT_4[8977] = 32'b00000000000000000001001100011101;
assign LUT_4[8978] = 32'b00000000000000000111011011001001;
assign LUT_4[8979] = 32'b00000000000000000000100111000001;
assign LUT_4[8980] = 32'b00000000000000000101000001000001;
assign LUT_4[8981] = 32'b11111111111111111110001100111001;
assign LUT_4[8982] = 32'b00000000000000000100011011100101;
assign LUT_4[8983] = 32'b11111111111111111101100111011101;
assign LUT_4[8984] = 32'b00000000000000000001001100111010;
assign LUT_4[8985] = 32'b11111111111111111010011000110010;
assign LUT_4[8986] = 32'b00000000000000000000100111011110;
assign LUT_4[8987] = 32'b11111111111111111001110011010110;
assign LUT_4[8988] = 32'b11111111111111111110001101010110;
assign LUT_4[8989] = 32'b11111111111111110111011001001110;
assign LUT_4[8990] = 32'b11111111111111111101100111111010;
assign LUT_4[8991] = 32'b11111111111111110110110011110010;
assign LUT_4[8992] = 32'b00000000000000001000101001111110;
assign LUT_4[8993] = 32'b00000000000000000001110101110110;
assign LUT_4[8994] = 32'b00000000000000001000000100100010;
assign LUT_4[8995] = 32'b00000000000000000001010000011010;
assign LUT_4[8996] = 32'b00000000000000000101101010011010;
assign LUT_4[8997] = 32'b11111111111111111110110110010010;
assign LUT_4[8998] = 32'b00000000000000000101000100111110;
assign LUT_4[8999] = 32'b11111111111111111110010000110110;
assign LUT_4[9000] = 32'b00000000000000000001110110010011;
assign LUT_4[9001] = 32'b11111111111111111011000010001011;
assign LUT_4[9002] = 32'b00000000000000000001010000110111;
assign LUT_4[9003] = 32'b11111111111111111010011100101111;
assign LUT_4[9004] = 32'b11111111111111111110110110101111;
assign LUT_4[9005] = 32'b11111111111111111000000010100111;
assign LUT_4[9006] = 32'b11111111111111111110010001010011;
assign LUT_4[9007] = 32'b11111111111111110111011101001011;
assign LUT_4[9008] = 32'b00000000000000000110011011101100;
assign LUT_4[9009] = 32'b11111111111111111111100111100100;
assign LUT_4[9010] = 32'b00000000000000000101110110010000;
assign LUT_4[9011] = 32'b11111111111111111111000010001000;
assign LUT_4[9012] = 32'b00000000000000000011011100001000;
assign LUT_4[9013] = 32'b11111111111111111100101000000000;
assign LUT_4[9014] = 32'b00000000000000000010110110101100;
assign LUT_4[9015] = 32'b11111111111111111100000010100100;
assign LUT_4[9016] = 32'b11111111111111111111101000000001;
assign LUT_4[9017] = 32'b11111111111111111000110011111001;
assign LUT_4[9018] = 32'b11111111111111111111000010100101;
assign LUT_4[9019] = 32'b11111111111111111000001110011101;
assign LUT_4[9020] = 32'b11111111111111111100101000011101;
assign LUT_4[9021] = 32'b11111111111111110101110100010101;
assign LUT_4[9022] = 32'b11111111111111111100000011000001;
assign LUT_4[9023] = 32'b11111111111111110101001110111001;
assign LUT_4[9024] = 32'b00000000000000001011100110001011;
assign LUT_4[9025] = 32'b00000000000000000100110010000011;
assign LUT_4[9026] = 32'b00000000000000001011000000101111;
assign LUT_4[9027] = 32'b00000000000000000100001100100111;
assign LUT_4[9028] = 32'b00000000000000001000100110100111;
assign LUT_4[9029] = 32'b00000000000000000001110010011111;
assign LUT_4[9030] = 32'b00000000000000001000000001001011;
assign LUT_4[9031] = 32'b00000000000000000001001101000011;
assign LUT_4[9032] = 32'b00000000000000000100110010100000;
assign LUT_4[9033] = 32'b11111111111111111101111110011000;
assign LUT_4[9034] = 32'b00000000000000000100001101000100;
assign LUT_4[9035] = 32'b11111111111111111101011000111100;
assign LUT_4[9036] = 32'b00000000000000000001110010111100;
assign LUT_4[9037] = 32'b11111111111111111010111110110100;
assign LUT_4[9038] = 32'b00000000000000000001001101100000;
assign LUT_4[9039] = 32'b11111111111111111010011001011000;
assign LUT_4[9040] = 32'b00000000000000001001010111111001;
assign LUT_4[9041] = 32'b00000000000000000010100011110001;
assign LUT_4[9042] = 32'b00000000000000001000110010011101;
assign LUT_4[9043] = 32'b00000000000000000001111110010101;
assign LUT_4[9044] = 32'b00000000000000000110011000010101;
assign LUT_4[9045] = 32'b11111111111111111111100100001101;
assign LUT_4[9046] = 32'b00000000000000000101110010111001;
assign LUT_4[9047] = 32'b11111111111111111110111110110001;
assign LUT_4[9048] = 32'b00000000000000000010100100001110;
assign LUT_4[9049] = 32'b11111111111111111011110000000110;
assign LUT_4[9050] = 32'b00000000000000000001111110110010;
assign LUT_4[9051] = 32'b11111111111111111011001010101010;
assign LUT_4[9052] = 32'b11111111111111111111100100101010;
assign LUT_4[9053] = 32'b11111111111111111000110000100010;
assign LUT_4[9054] = 32'b11111111111111111110111111001110;
assign LUT_4[9055] = 32'b11111111111111111000001011000110;
assign LUT_4[9056] = 32'b00000000000000001010000001010010;
assign LUT_4[9057] = 32'b00000000000000000011001101001010;
assign LUT_4[9058] = 32'b00000000000000001001011011110110;
assign LUT_4[9059] = 32'b00000000000000000010100111101110;
assign LUT_4[9060] = 32'b00000000000000000111000001101110;
assign LUT_4[9061] = 32'b00000000000000000000001101100110;
assign LUT_4[9062] = 32'b00000000000000000110011100010010;
assign LUT_4[9063] = 32'b11111111111111111111101000001010;
assign LUT_4[9064] = 32'b00000000000000000011001101100111;
assign LUT_4[9065] = 32'b11111111111111111100011001011111;
assign LUT_4[9066] = 32'b00000000000000000010101000001011;
assign LUT_4[9067] = 32'b11111111111111111011110100000011;
assign LUT_4[9068] = 32'b00000000000000000000001110000011;
assign LUT_4[9069] = 32'b11111111111111111001011001111011;
assign LUT_4[9070] = 32'b11111111111111111111101000100111;
assign LUT_4[9071] = 32'b11111111111111111000110100011111;
assign LUT_4[9072] = 32'b00000000000000000111110011000000;
assign LUT_4[9073] = 32'b00000000000000000000111110111000;
assign LUT_4[9074] = 32'b00000000000000000111001101100100;
assign LUT_4[9075] = 32'b00000000000000000000011001011100;
assign LUT_4[9076] = 32'b00000000000000000100110011011100;
assign LUT_4[9077] = 32'b11111111111111111101111111010100;
assign LUT_4[9078] = 32'b00000000000000000100001110000000;
assign LUT_4[9079] = 32'b11111111111111111101011001111000;
assign LUT_4[9080] = 32'b00000000000000000000111111010101;
assign LUT_4[9081] = 32'b11111111111111111010001011001101;
assign LUT_4[9082] = 32'b00000000000000000000011001111001;
assign LUT_4[9083] = 32'b11111111111111111001100101110001;
assign LUT_4[9084] = 32'b11111111111111111101111111110001;
assign LUT_4[9085] = 32'b11111111111111110111001011101001;
assign LUT_4[9086] = 32'b11111111111111111101011010010101;
assign LUT_4[9087] = 32'b11111111111111110110100110001101;
assign LUT_4[9088] = 32'b00000000000000001100110100111111;
assign LUT_4[9089] = 32'b00000000000000000110000000110111;
assign LUT_4[9090] = 32'b00000000000000001100001111100011;
assign LUT_4[9091] = 32'b00000000000000000101011011011011;
assign LUT_4[9092] = 32'b00000000000000001001110101011011;
assign LUT_4[9093] = 32'b00000000000000000011000001010011;
assign LUT_4[9094] = 32'b00000000000000001001001111111111;
assign LUT_4[9095] = 32'b00000000000000000010011011110111;
assign LUT_4[9096] = 32'b00000000000000000110000001010100;
assign LUT_4[9097] = 32'b11111111111111111111001101001100;
assign LUT_4[9098] = 32'b00000000000000000101011011111000;
assign LUT_4[9099] = 32'b11111111111111111110100111110000;
assign LUT_4[9100] = 32'b00000000000000000011000001110000;
assign LUT_4[9101] = 32'b11111111111111111100001101101000;
assign LUT_4[9102] = 32'b00000000000000000010011100010100;
assign LUT_4[9103] = 32'b11111111111111111011101000001100;
assign LUT_4[9104] = 32'b00000000000000001010100110101101;
assign LUT_4[9105] = 32'b00000000000000000011110010100101;
assign LUT_4[9106] = 32'b00000000000000001010000001010001;
assign LUT_4[9107] = 32'b00000000000000000011001101001001;
assign LUT_4[9108] = 32'b00000000000000000111100111001001;
assign LUT_4[9109] = 32'b00000000000000000000110011000001;
assign LUT_4[9110] = 32'b00000000000000000111000001101101;
assign LUT_4[9111] = 32'b00000000000000000000001101100101;
assign LUT_4[9112] = 32'b00000000000000000011110011000010;
assign LUT_4[9113] = 32'b11111111111111111100111110111010;
assign LUT_4[9114] = 32'b00000000000000000011001101100110;
assign LUT_4[9115] = 32'b11111111111111111100011001011110;
assign LUT_4[9116] = 32'b00000000000000000000110011011110;
assign LUT_4[9117] = 32'b11111111111111111001111111010110;
assign LUT_4[9118] = 32'b00000000000000000000001110000010;
assign LUT_4[9119] = 32'b11111111111111111001011001111010;
assign LUT_4[9120] = 32'b00000000000000001011010000000110;
assign LUT_4[9121] = 32'b00000000000000000100011011111110;
assign LUT_4[9122] = 32'b00000000000000001010101010101010;
assign LUT_4[9123] = 32'b00000000000000000011110110100010;
assign LUT_4[9124] = 32'b00000000000000001000010000100010;
assign LUT_4[9125] = 32'b00000000000000000001011100011010;
assign LUT_4[9126] = 32'b00000000000000000111101011000110;
assign LUT_4[9127] = 32'b00000000000000000000110110111110;
assign LUT_4[9128] = 32'b00000000000000000100011100011011;
assign LUT_4[9129] = 32'b11111111111111111101101000010011;
assign LUT_4[9130] = 32'b00000000000000000011110110111111;
assign LUT_4[9131] = 32'b11111111111111111101000010110111;
assign LUT_4[9132] = 32'b00000000000000000001011100110111;
assign LUT_4[9133] = 32'b11111111111111111010101000101111;
assign LUT_4[9134] = 32'b00000000000000000000110111011011;
assign LUT_4[9135] = 32'b11111111111111111010000011010011;
assign LUT_4[9136] = 32'b00000000000000001001000001110100;
assign LUT_4[9137] = 32'b00000000000000000010001101101100;
assign LUT_4[9138] = 32'b00000000000000001000011100011000;
assign LUT_4[9139] = 32'b00000000000000000001101000010000;
assign LUT_4[9140] = 32'b00000000000000000110000010010000;
assign LUT_4[9141] = 32'b11111111111111111111001110001000;
assign LUT_4[9142] = 32'b00000000000000000101011100110100;
assign LUT_4[9143] = 32'b11111111111111111110101000101100;
assign LUT_4[9144] = 32'b00000000000000000010001110001001;
assign LUT_4[9145] = 32'b11111111111111111011011010000001;
assign LUT_4[9146] = 32'b00000000000000000001101000101101;
assign LUT_4[9147] = 32'b11111111111111111010110100100101;
assign LUT_4[9148] = 32'b11111111111111111111001110100101;
assign LUT_4[9149] = 32'b11111111111111111000011010011101;
assign LUT_4[9150] = 32'b11111111111111111110101001001001;
assign LUT_4[9151] = 32'b11111111111111110111110101000001;
assign LUT_4[9152] = 32'b00000000000000001110001100010011;
assign LUT_4[9153] = 32'b00000000000000000111011000001011;
assign LUT_4[9154] = 32'b00000000000000001101100110110111;
assign LUT_4[9155] = 32'b00000000000000000110110010101111;
assign LUT_4[9156] = 32'b00000000000000001011001100101111;
assign LUT_4[9157] = 32'b00000000000000000100011000100111;
assign LUT_4[9158] = 32'b00000000000000001010100111010011;
assign LUT_4[9159] = 32'b00000000000000000011110011001011;
assign LUT_4[9160] = 32'b00000000000000000111011000101000;
assign LUT_4[9161] = 32'b00000000000000000000100100100000;
assign LUT_4[9162] = 32'b00000000000000000110110011001100;
assign LUT_4[9163] = 32'b11111111111111111111111111000100;
assign LUT_4[9164] = 32'b00000000000000000100011001000100;
assign LUT_4[9165] = 32'b11111111111111111101100100111100;
assign LUT_4[9166] = 32'b00000000000000000011110011101000;
assign LUT_4[9167] = 32'b11111111111111111100111111100000;
assign LUT_4[9168] = 32'b00000000000000001011111110000001;
assign LUT_4[9169] = 32'b00000000000000000101001001111001;
assign LUT_4[9170] = 32'b00000000000000001011011000100101;
assign LUT_4[9171] = 32'b00000000000000000100100100011101;
assign LUT_4[9172] = 32'b00000000000000001000111110011101;
assign LUT_4[9173] = 32'b00000000000000000010001010010101;
assign LUT_4[9174] = 32'b00000000000000001000011001000001;
assign LUT_4[9175] = 32'b00000000000000000001100100111001;
assign LUT_4[9176] = 32'b00000000000000000101001010010110;
assign LUT_4[9177] = 32'b11111111111111111110010110001110;
assign LUT_4[9178] = 32'b00000000000000000100100100111010;
assign LUT_4[9179] = 32'b11111111111111111101110000110010;
assign LUT_4[9180] = 32'b00000000000000000010001010110010;
assign LUT_4[9181] = 32'b11111111111111111011010110101010;
assign LUT_4[9182] = 32'b00000000000000000001100101010110;
assign LUT_4[9183] = 32'b11111111111111111010110001001110;
assign LUT_4[9184] = 32'b00000000000000001100100111011010;
assign LUT_4[9185] = 32'b00000000000000000101110011010010;
assign LUT_4[9186] = 32'b00000000000000001100000001111110;
assign LUT_4[9187] = 32'b00000000000000000101001101110110;
assign LUT_4[9188] = 32'b00000000000000001001100111110110;
assign LUT_4[9189] = 32'b00000000000000000010110011101110;
assign LUT_4[9190] = 32'b00000000000000001001000010011010;
assign LUT_4[9191] = 32'b00000000000000000010001110010010;
assign LUT_4[9192] = 32'b00000000000000000101110011101111;
assign LUT_4[9193] = 32'b11111111111111111110111111100111;
assign LUT_4[9194] = 32'b00000000000000000101001110010011;
assign LUT_4[9195] = 32'b11111111111111111110011010001011;
assign LUT_4[9196] = 32'b00000000000000000010110100001011;
assign LUT_4[9197] = 32'b11111111111111111100000000000011;
assign LUT_4[9198] = 32'b00000000000000000010001110101111;
assign LUT_4[9199] = 32'b11111111111111111011011010100111;
assign LUT_4[9200] = 32'b00000000000000001010011001001000;
assign LUT_4[9201] = 32'b00000000000000000011100101000000;
assign LUT_4[9202] = 32'b00000000000000001001110011101100;
assign LUT_4[9203] = 32'b00000000000000000010111111100100;
assign LUT_4[9204] = 32'b00000000000000000111011001100100;
assign LUT_4[9205] = 32'b00000000000000000000100101011100;
assign LUT_4[9206] = 32'b00000000000000000110110100001000;
assign LUT_4[9207] = 32'b00000000000000000000000000000000;
assign LUT_4[9208] = 32'b00000000000000000011100101011101;
assign LUT_4[9209] = 32'b11111111111111111100110001010101;
assign LUT_4[9210] = 32'b00000000000000000011000000000001;
assign LUT_4[9211] = 32'b11111111111111111100001011111001;
assign LUT_4[9212] = 32'b00000000000000000000100101111001;
assign LUT_4[9213] = 32'b11111111111111111001110001110001;
assign LUT_4[9214] = 32'b00000000000000000000000000011101;
assign LUT_4[9215] = 32'b11111111111111111001001100010101;
assign LUT_4[9216] = 32'b00000000000000000111111001101011;
assign LUT_4[9217] = 32'b00000000000000000001000101100011;
assign LUT_4[9218] = 32'b00000000000000000111010100001111;
assign LUT_4[9219] = 32'b00000000000000000000100000000111;
assign LUT_4[9220] = 32'b00000000000000000100111010000111;
assign LUT_4[9221] = 32'b11111111111111111110000101111111;
assign LUT_4[9222] = 32'b00000000000000000100010100101011;
assign LUT_4[9223] = 32'b11111111111111111101100000100011;
assign LUT_4[9224] = 32'b00000000000000000001000110000000;
assign LUT_4[9225] = 32'b11111111111111111010010001111000;
assign LUT_4[9226] = 32'b00000000000000000000100000100100;
assign LUT_4[9227] = 32'b11111111111111111001101100011100;
assign LUT_4[9228] = 32'b11111111111111111110000110011100;
assign LUT_4[9229] = 32'b11111111111111110111010010010100;
assign LUT_4[9230] = 32'b11111111111111111101100001000000;
assign LUT_4[9231] = 32'b11111111111111110110101100111000;
assign LUT_4[9232] = 32'b00000000000000000101101011011001;
assign LUT_4[9233] = 32'b11111111111111111110110111010001;
assign LUT_4[9234] = 32'b00000000000000000101000101111101;
assign LUT_4[9235] = 32'b11111111111111111110010001110101;
assign LUT_4[9236] = 32'b00000000000000000010101011110101;
assign LUT_4[9237] = 32'b11111111111111111011110111101101;
assign LUT_4[9238] = 32'b00000000000000000010000110011001;
assign LUT_4[9239] = 32'b11111111111111111011010010010001;
assign LUT_4[9240] = 32'b11111111111111111110110111101110;
assign LUT_4[9241] = 32'b11111111111111111000000011100110;
assign LUT_4[9242] = 32'b11111111111111111110010010010010;
assign LUT_4[9243] = 32'b11111111111111110111011110001010;
assign LUT_4[9244] = 32'b11111111111111111011111000001010;
assign LUT_4[9245] = 32'b11111111111111110101000100000010;
assign LUT_4[9246] = 32'b11111111111111111011010010101110;
assign LUT_4[9247] = 32'b11111111111111110100011110100110;
assign LUT_4[9248] = 32'b00000000000000000110010100110010;
assign LUT_4[9249] = 32'b11111111111111111111100000101010;
assign LUT_4[9250] = 32'b00000000000000000101101111010110;
assign LUT_4[9251] = 32'b11111111111111111110111011001110;
assign LUT_4[9252] = 32'b00000000000000000011010101001110;
assign LUT_4[9253] = 32'b11111111111111111100100001000110;
assign LUT_4[9254] = 32'b00000000000000000010101111110010;
assign LUT_4[9255] = 32'b11111111111111111011111011101010;
assign LUT_4[9256] = 32'b11111111111111111111100001000111;
assign LUT_4[9257] = 32'b11111111111111111000101100111111;
assign LUT_4[9258] = 32'b11111111111111111110111011101011;
assign LUT_4[9259] = 32'b11111111111111111000000111100011;
assign LUT_4[9260] = 32'b11111111111111111100100001100011;
assign LUT_4[9261] = 32'b11111111111111110101101101011011;
assign LUT_4[9262] = 32'b11111111111111111011111100000111;
assign LUT_4[9263] = 32'b11111111111111110101000111111111;
assign LUT_4[9264] = 32'b00000000000000000100000110100000;
assign LUT_4[9265] = 32'b11111111111111111101010010011000;
assign LUT_4[9266] = 32'b00000000000000000011100001000100;
assign LUT_4[9267] = 32'b11111111111111111100101100111100;
assign LUT_4[9268] = 32'b00000000000000000001000110111100;
assign LUT_4[9269] = 32'b11111111111111111010010010110100;
assign LUT_4[9270] = 32'b00000000000000000000100001100000;
assign LUT_4[9271] = 32'b11111111111111111001101101011000;
assign LUT_4[9272] = 32'b11111111111111111101010010110101;
assign LUT_4[9273] = 32'b11111111111111110110011110101101;
assign LUT_4[9274] = 32'b11111111111111111100101101011001;
assign LUT_4[9275] = 32'b11111111111111110101111001010001;
assign LUT_4[9276] = 32'b11111111111111111010010011010001;
assign LUT_4[9277] = 32'b11111111111111110011011111001001;
assign LUT_4[9278] = 32'b11111111111111111001101101110101;
assign LUT_4[9279] = 32'b11111111111111110010111001101101;
assign LUT_4[9280] = 32'b00000000000000001001010000111111;
assign LUT_4[9281] = 32'b00000000000000000010011100110111;
assign LUT_4[9282] = 32'b00000000000000001000101011100011;
assign LUT_4[9283] = 32'b00000000000000000001110111011011;
assign LUT_4[9284] = 32'b00000000000000000110010001011011;
assign LUT_4[9285] = 32'b11111111111111111111011101010011;
assign LUT_4[9286] = 32'b00000000000000000101101011111111;
assign LUT_4[9287] = 32'b11111111111111111110110111110111;
assign LUT_4[9288] = 32'b00000000000000000010011101010100;
assign LUT_4[9289] = 32'b11111111111111111011101001001100;
assign LUT_4[9290] = 32'b00000000000000000001110111111000;
assign LUT_4[9291] = 32'b11111111111111111011000011110000;
assign LUT_4[9292] = 32'b11111111111111111111011101110000;
assign LUT_4[9293] = 32'b11111111111111111000101001101000;
assign LUT_4[9294] = 32'b11111111111111111110111000010100;
assign LUT_4[9295] = 32'b11111111111111111000000100001100;
assign LUT_4[9296] = 32'b00000000000000000111000010101101;
assign LUT_4[9297] = 32'b00000000000000000000001110100101;
assign LUT_4[9298] = 32'b00000000000000000110011101010001;
assign LUT_4[9299] = 32'b11111111111111111111101001001001;
assign LUT_4[9300] = 32'b00000000000000000100000011001001;
assign LUT_4[9301] = 32'b11111111111111111101001111000001;
assign LUT_4[9302] = 32'b00000000000000000011011101101101;
assign LUT_4[9303] = 32'b11111111111111111100101001100101;
assign LUT_4[9304] = 32'b00000000000000000000001111000010;
assign LUT_4[9305] = 32'b11111111111111111001011010111010;
assign LUT_4[9306] = 32'b11111111111111111111101001100110;
assign LUT_4[9307] = 32'b11111111111111111000110101011110;
assign LUT_4[9308] = 32'b11111111111111111101001111011110;
assign LUT_4[9309] = 32'b11111111111111110110011011010110;
assign LUT_4[9310] = 32'b11111111111111111100101010000010;
assign LUT_4[9311] = 32'b11111111111111110101110101111010;
assign LUT_4[9312] = 32'b00000000000000000111101100000110;
assign LUT_4[9313] = 32'b00000000000000000000110111111110;
assign LUT_4[9314] = 32'b00000000000000000111000110101010;
assign LUT_4[9315] = 32'b00000000000000000000010010100010;
assign LUT_4[9316] = 32'b00000000000000000100101100100010;
assign LUT_4[9317] = 32'b11111111111111111101111000011010;
assign LUT_4[9318] = 32'b00000000000000000100000111000110;
assign LUT_4[9319] = 32'b11111111111111111101010010111110;
assign LUT_4[9320] = 32'b00000000000000000000111000011011;
assign LUT_4[9321] = 32'b11111111111111111010000100010011;
assign LUT_4[9322] = 32'b00000000000000000000010010111111;
assign LUT_4[9323] = 32'b11111111111111111001011110110111;
assign LUT_4[9324] = 32'b11111111111111111101111000110111;
assign LUT_4[9325] = 32'b11111111111111110111000100101111;
assign LUT_4[9326] = 32'b11111111111111111101010011011011;
assign LUT_4[9327] = 32'b11111111111111110110011111010011;
assign LUT_4[9328] = 32'b00000000000000000101011101110100;
assign LUT_4[9329] = 32'b11111111111111111110101001101100;
assign LUT_4[9330] = 32'b00000000000000000100111000011000;
assign LUT_4[9331] = 32'b11111111111111111110000100010000;
assign LUT_4[9332] = 32'b00000000000000000010011110010000;
assign LUT_4[9333] = 32'b11111111111111111011101010001000;
assign LUT_4[9334] = 32'b00000000000000000001111000110100;
assign LUT_4[9335] = 32'b11111111111111111011000100101100;
assign LUT_4[9336] = 32'b11111111111111111110101010001001;
assign LUT_4[9337] = 32'b11111111111111110111110110000001;
assign LUT_4[9338] = 32'b11111111111111111110000100101101;
assign LUT_4[9339] = 32'b11111111111111110111010000100101;
assign LUT_4[9340] = 32'b11111111111111111011101010100101;
assign LUT_4[9341] = 32'b11111111111111110100110110011101;
assign LUT_4[9342] = 32'b11111111111111111011000101001001;
assign LUT_4[9343] = 32'b11111111111111110100010001000001;
assign LUT_4[9344] = 32'b00000000000000001010011111110011;
assign LUT_4[9345] = 32'b00000000000000000011101011101011;
assign LUT_4[9346] = 32'b00000000000000001001111010010111;
assign LUT_4[9347] = 32'b00000000000000000011000110001111;
assign LUT_4[9348] = 32'b00000000000000000111100000001111;
assign LUT_4[9349] = 32'b00000000000000000000101100000111;
assign LUT_4[9350] = 32'b00000000000000000110111010110011;
assign LUT_4[9351] = 32'b00000000000000000000000110101011;
assign LUT_4[9352] = 32'b00000000000000000011101100001000;
assign LUT_4[9353] = 32'b11111111111111111100111000000000;
assign LUT_4[9354] = 32'b00000000000000000011000110101100;
assign LUT_4[9355] = 32'b11111111111111111100010010100100;
assign LUT_4[9356] = 32'b00000000000000000000101100100100;
assign LUT_4[9357] = 32'b11111111111111111001111000011100;
assign LUT_4[9358] = 32'b00000000000000000000000111001000;
assign LUT_4[9359] = 32'b11111111111111111001010011000000;
assign LUT_4[9360] = 32'b00000000000000001000010001100001;
assign LUT_4[9361] = 32'b00000000000000000001011101011001;
assign LUT_4[9362] = 32'b00000000000000000111101100000101;
assign LUT_4[9363] = 32'b00000000000000000000110111111101;
assign LUT_4[9364] = 32'b00000000000000000101010001111101;
assign LUT_4[9365] = 32'b11111111111111111110011101110101;
assign LUT_4[9366] = 32'b00000000000000000100101100100001;
assign LUT_4[9367] = 32'b11111111111111111101111000011001;
assign LUT_4[9368] = 32'b00000000000000000001011101110110;
assign LUT_4[9369] = 32'b11111111111111111010101001101110;
assign LUT_4[9370] = 32'b00000000000000000000111000011010;
assign LUT_4[9371] = 32'b11111111111111111010000100010010;
assign LUT_4[9372] = 32'b11111111111111111110011110010010;
assign LUT_4[9373] = 32'b11111111111111110111101010001010;
assign LUT_4[9374] = 32'b11111111111111111101111000110110;
assign LUT_4[9375] = 32'b11111111111111110111000100101110;
assign LUT_4[9376] = 32'b00000000000000001000111010111010;
assign LUT_4[9377] = 32'b00000000000000000010000110110010;
assign LUT_4[9378] = 32'b00000000000000001000010101011110;
assign LUT_4[9379] = 32'b00000000000000000001100001010110;
assign LUT_4[9380] = 32'b00000000000000000101111011010110;
assign LUT_4[9381] = 32'b11111111111111111111000111001110;
assign LUT_4[9382] = 32'b00000000000000000101010101111010;
assign LUT_4[9383] = 32'b11111111111111111110100001110010;
assign LUT_4[9384] = 32'b00000000000000000010000111001111;
assign LUT_4[9385] = 32'b11111111111111111011010011000111;
assign LUT_4[9386] = 32'b00000000000000000001100001110011;
assign LUT_4[9387] = 32'b11111111111111111010101101101011;
assign LUT_4[9388] = 32'b11111111111111111111000111101011;
assign LUT_4[9389] = 32'b11111111111111111000010011100011;
assign LUT_4[9390] = 32'b11111111111111111110100010001111;
assign LUT_4[9391] = 32'b11111111111111110111101110000111;
assign LUT_4[9392] = 32'b00000000000000000110101100101000;
assign LUT_4[9393] = 32'b11111111111111111111111000100000;
assign LUT_4[9394] = 32'b00000000000000000110000111001100;
assign LUT_4[9395] = 32'b11111111111111111111010011000100;
assign LUT_4[9396] = 32'b00000000000000000011101101000100;
assign LUT_4[9397] = 32'b11111111111111111100111000111100;
assign LUT_4[9398] = 32'b00000000000000000011000111101000;
assign LUT_4[9399] = 32'b11111111111111111100010011100000;
assign LUT_4[9400] = 32'b11111111111111111111111000111101;
assign LUT_4[9401] = 32'b11111111111111111001000100110101;
assign LUT_4[9402] = 32'b11111111111111111111010011100001;
assign LUT_4[9403] = 32'b11111111111111111000011111011001;
assign LUT_4[9404] = 32'b11111111111111111100111001011001;
assign LUT_4[9405] = 32'b11111111111111110110000101010001;
assign LUT_4[9406] = 32'b11111111111111111100010011111101;
assign LUT_4[9407] = 32'b11111111111111110101011111110101;
assign LUT_4[9408] = 32'b00000000000000001011110111000111;
assign LUT_4[9409] = 32'b00000000000000000101000010111111;
assign LUT_4[9410] = 32'b00000000000000001011010001101011;
assign LUT_4[9411] = 32'b00000000000000000100011101100011;
assign LUT_4[9412] = 32'b00000000000000001000110111100011;
assign LUT_4[9413] = 32'b00000000000000000010000011011011;
assign LUT_4[9414] = 32'b00000000000000001000010010000111;
assign LUT_4[9415] = 32'b00000000000000000001011101111111;
assign LUT_4[9416] = 32'b00000000000000000101000011011100;
assign LUT_4[9417] = 32'b11111111111111111110001111010100;
assign LUT_4[9418] = 32'b00000000000000000100011110000000;
assign LUT_4[9419] = 32'b11111111111111111101101001111000;
assign LUT_4[9420] = 32'b00000000000000000010000011111000;
assign LUT_4[9421] = 32'b11111111111111111011001111110000;
assign LUT_4[9422] = 32'b00000000000000000001011110011100;
assign LUT_4[9423] = 32'b11111111111111111010101010010100;
assign LUT_4[9424] = 32'b00000000000000001001101000110101;
assign LUT_4[9425] = 32'b00000000000000000010110100101101;
assign LUT_4[9426] = 32'b00000000000000001001000011011001;
assign LUT_4[9427] = 32'b00000000000000000010001111010001;
assign LUT_4[9428] = 32'b00000000000000000110101001010001;
assign LUT_4[9429] = 32'b11111111111111111111110101001001;
assign LUT_4[9430] = 32'b00000000000000000110000011110101;
assign LUT_4[9431] = 32'b11111111111111111111001111101101;
assign LUT_4[9432] = 32'b00000000000000000010110101001010;
assign LUT_4[9433] = 32'b11111111111111111100000001000010;
assign LUT_4[9434] = 32'b00000000000000000010001111101110;
assign LUT_4[9435] = 32'b11111111111111111011011011100110;
assign LUT_4[9436] = 32'b11111111111111111111110101100110;
assign LUT_4[9437] = 32'b11111111111111111001000001011110;
assign LUT_4[9438] = 32'b11111111111111111111010000001010;
assign LUT_4[9439] = 32'b11111111111111111000011100000010;
assign LUT_4[9440] = 32'b00000000000000001010010010001110;
assign LUT_4[9441] = 32'b00000000000000000011011110000110;
assign LUT_4[9442] = 32'b00000000000000001001101100110010;
assign LUT_4[9443] = 32'b00000000000000000010111000101010;
assign LUT_4[9444] = 32'b00000000000000000111010010101010;
assign LUT_4[9445] = 32'b00000000000000000000011110100010;
assign LUT_4[9446] = 32'b00000000000000000110101101001110;
assign LUT_4[9447] = 32'b11111111111111111111111001000110;
assign LUT_4[9448] = 32'b00000000000000000011011110100011;
assign LUT_4[9449] = 32'b11111111111111111100101010011011;
assign LUT_4[9450] = 32'b00000000000000000010111001000111;
assign LUT_4[9451] = 32'b11111111111111111100000100111111;
assign LUT_4[9452] = 32'b00000000000000000000011110111111;
assign LUT_4[9453] = 32'b11111111111111111001101010110111;
assign LUT_4[9454] = 32'b11111111111111111111111001100011;
assign LUT_4[9455] = 32'b11111111111111111001000101011011;
assign LUT_4[9456] = 32'b00000000000000001000000011111100;
assign LUT_4[9457] = 32'b00000000000000000001001111110100;
assign LUT_4[9458] = 32'b00000000000000000111011110100000;
assign LUT_4[9459] = 32'b00000000000000000000101010011000;
assign LUT_4[9460] = 32'b00000000000000000101000100011000;
assign LUT_4[9461] = 32'b11111111111111111110010000010000;
assign LUT_4[9462] = 32'b00000000000000000100011110111100;
assign LUT_4[9463] = 32'b11111111111111111101101010110100;
assign LUT_4[9464] = 32'b00000000000000000001010000010001;
assign LUT_4[9465] = 32'b11111111111111111010011100001001;
assign LUT_4[9466] = 32'b00000000000000000000101010110101;
assign LUT_4[9467] = 32'b11111111111111111001110110101101;
assign LUT_4[9468] = 32'b11111111111111111110010000101101;
assign LUT_4[9469] = 32'b11111111111111110111011100100101;
assign LUT_4[9470] = 32'b11111111111111111101101011010001;
assign LUT_4[9471] = 32'b11111111111111110110110111001001;
assign LUT_4[9472] = 32'b00000000000000001100110101001110;
assign LUT_4[9473] = 32'b00000000000000000110000001000110;
assign LUT_4[9474] = 32'b00000000000000001100001111110010;
assign LUT_4[9475] = 32'b00000000000000000101011011101010;
assign LUT_4[9476] = 32'b00000000000000001001110101101010;
assign LUT_4[9477] = 32'b00000000000000000011000001100010;
assign LUT_4[9478] = 32'b00000000000000001001010000001110;
assign LUT_4[9479] = 32'b00000000000000000010011100000110;
assign LUT_4[9480] = 32'b00000000000000000110000001100011;
assign LUT_4[9481] = 32'b11111111111111111111001101011011;
assign LUT_4[9482] = 32'b00000000000000000101011100000111;
assign LUT_4[9483] = 32'b11111111111111111110100111111111;
assign LUT_4[9484] = 32'b00000000000000000011000001111111;
assign LUT_4[9485] = 32'b11111111111111111100001101110111;
assign LUT_4[9486] = 32'b00000000000000000010011100100011;
assign LUT_4[9487] = 32'b11111111111111111011101000011011;
assign LUT_4[9488] = 32'b00000000000000001010100110111100;
assign LUT_4[9489] = 32'b00000000000000000011110010110100;
assign LUT_4[9490] = 32'b00000000000000001010000001100000;
assign LUT_4[9491] = 32'b00000000000000000011001101011000;
assign LUT_4[9492] = 32'b00000000000000000111100111011000;
assign LUT_4[9493] = 32'b00000000000000000000110011010000;
assign LUT_4[9494] = 32'b00000000000000000111000001111100;
assign LUT_4[9495] = 32'b00000000000000000000001101110100;
assign LUT_4[9496] = 32'b00000000000000000011110011010001;
assign LUT_4[9497] = 32'b11111111111111111100111111001001;
assign LUT_4[9498] = 32'b00000000000000000011001101110101;
assign LUT_4[9499] = 32'b11111111111111111100011001101101;
assign LUT_4[9500] = 32'b00000000000000000000110011101101;
assign LUT_4[9501] = 32'b11111111111111111001111111100101;
assign LUT_4[9502] = 32'b00000000000000000000001110010001;
assign LUT_4[9503] = 32'b11111111111111111001011010001001;
assign LUT_4[9504] = 32'b00000000000000001011010000010101;
assign LUT_4[9505] = 32'b00000000000000000100011100001101;
assign LUT_4[9506] = 32'b00000000000000001010101010111001;
assign LUT_4[9507] = 32'b00000000000000000011110110110001;
assign LUT_4[9508] = 32'b00000000000000001000010000110001;
assign LUT_4[9509] = 32'b00000000000000000001011100101001;
assign LUT_4[9510] = 32'b00000000000000000111101011010101;
assign LUT_4[9511] = 32'b00000000000000000000110111001101;
assign LUT_4[9512] = 32'b00000000000000000100011100101010;
assign LUT_4[9513] = 32'b11111111111111111101101000100010;
assign LUT_4[9514] = 32'b00000000000000000011110111001110;
assign LUT_4[9515] = 32'b11111111111111111101000011000110;
assign LUT_4[9516] = 32'b00000000000000000001011101000110;
assign LUT_4[9517] = 32'b11111111111111111010101000111110;
assign LUT_4[9518] = 32'b00000000000000000000110111101010;
assign LUT_4[9519] = 32'b11111111111111111010000011100010;
assign LUT_4[9520] = 32'b00000000000000001001000010000011;
assign LUT_4[9521] = 32'b00000000000000000010001101111011;
assign LUT_4[9522] = 32'b00000000000000001000011100100111;
assign LUT_4[9523] = 32'b00000000000000000001101000011111;
assign LUT_4[9524] = 32'b00000000000000000110000010011111;
assign LUT_4[9525] = 32'b11111111111111111111001110010111;
assign LUT_4[9526] = 32'b00000000000000000101011101000011;
assign LUT_4[9527] = 32'b11111111111111111110101000111011;
assign LUT_4[9528] = 32'b00000000000000000010001110011000;
assign LUT_4[9529] = 32'b11111111111111111011011010010000;
assign LUT_4[9530] = 32'b00000000000000000001101000111100;
assign LUT_4[9531] = 32'b11111111111111111010110100110100;
assign LUT_4[9532] = 32'b11111111111111111111001110110100;
assign LUT_4[9533] = 32'b11111111111111111000011010101100;
assign LUT_4[9534] = 32'b11111111111111111110101001011000;
assign LUT_4[9535] = 32'b11111111111111110111110101010000;
assign LUT_4[9536] = 32'b00000000000000001110001100100010;
assign LUT_4[9537] = 32'b00000000000000000111011000011010;
assign LUT_4[9538] = 32'b00000000000000001101100111000110;
assign LUT_4[9539] = 32'b00000000000000000110110010111110;
assign LUT_4[9540] = 32'b00000000000000001011001100111110;
assign LUT_4[9541] = 32'b00000000000000000100011000110110;
assign LUT_4[9542] = 32'b00000000000000001010100111100010;
assign LUT_4[9543] = 32'b00000000000000000011110011011010;
assign LUT_4[9544] = 32'b00000000000000000111011000110111;
assign LUT_4[9545] = 32'b00000000000000000000100100101111;
assign LUT_4[9546] = 32'b00000000000000000110110011011011;
assign LUT_4[9547] = 32'b11111111111111111111111111010011;
assign LUT_4[9548] = 32'b00000000000000000100011001010011;
assign LUT_4[9549] = 32'b11111111111111111101100101001011;
assign LUT_4[9550] = 32'b00000000000000000011110011110111;
assign LUT_4[9551] = 32'b11111111111111111100111111101111;
assign LUT_4[9552] = 32'b00000000000000001011111110010000;
assign LUT_4[9553] = 32'b00000000000000000101001010001000;
assign LUT_4[9554] = 32'b00000000000000001011011000110100;
assign LUT_4[9555] = 32'b00000000000000000100100100101100;
assign LUT_4[9556] = 32'b00000000000000001000111110101100;
assign LUT_4[9557] = 32'b00000000000000000010001010100100;
assign LUT_4[9558] = 32'b00000000000000001000011001010000;
assign LUT_4[9559] = 32'b00000000000000000001100101001000;
assign LUT_4[9560] = 32'b00000000000000000101001010100101;
assign LUT_4[9561] = 32'b11111111111111111110010110011101;
assign LUT_4[9562] = 32'b00000000000000000100100101001001;
assign LUT_4[9563] = 32'b11111111111111111101110001000001;
assign LUT_4[9564] = 32'b00000000000000000010001011000001;
assign LUT_4[9565] = 32'b11111111111111111011010110111001;
assign LUT_4[9566] = 32'b00000000000000000001100101100101;
assign LUT_4[9567] = 32'b11111111111111111010110001011101;
assign LUT_4[9568] = 32'b00000000000000001100100111101001;
assign LUT_4[9569] = 32'b00000000000000000101110011100001;
assign LUT_4[9570] = 32'b00000000000000001100000010001101;
assign LUT_4[9571] = 32'b00000000000000000101001110000101;
assign LUT_4[9572] = 32'b00000000000000001001101000000101;
assign LUT_4[9573] = 32'b00000000000000000010110011111101;
assign LUT_4[9574] = 32'b00000000000000001001000010101001;
assign LUT_4[9575] = 32'b00000000000000000010001110100001;
assign LUT_4[9576] = 32'b00000000000000000101110011111110;
assign LUT_4[9577] = 32'b11111111111111111110111111110110;
assign LUT_4[9578] = 32'b00000000000000000101001110100010;
assign LUT_4[9579] = 32'b11111111111111111110011010011010;
assign LUT_4[9580] = 32'b00000000000000000010110100011010;
assign LUT_4[9581] = 32'b11111111111111111100000000010010;
assign LUT_4[9582] = 32'b00000000000000000010001110111110;
assign LUT_4[9583] = 32'b11111111111111111011011010110110;
assign LUT_4[9584] = 32'b00000000000000001010011001010111;
assign LUT_4[9585] = 32'b00000000000000000011100101001111;
assign LUT_4[9586] = 32'b00000000000000001001110011111011;
assign LUT_4[9587] = 32'b00000000000000000010111111110011;
assign LUT_4[9588] = 32'b00000000000000000111011001110011;
assign LUT_4[9589] = 32'b00000000000000000000100101101011;
assign LUT_4[9590] = 32'b00000000000000000110110100010111;
assign LUT_4[9591] = 32'b00000000000000000000000000001111;
assign LUT_4[9592] = 32'b00000000000000000011100101101100;
assign LUT_4[9593] = 32'b11111111111111111100110001100100;
assign LUT_4[9594] = 32'b00000000000000000011000000010000;
assign LUT_4[9595] = 32'b11111111111111111100001100001000;
assign LUT_4[9596] = 32'b00000000000000000000100110001000;
assign LUT_4[9597] = 32'b11111111111111111001110010000000;
assign LUT_4[9598] = 32'b00000000000000000000000000101100;
assign LUT_4[9599] = 32'b11111111111111111001001100100100;
assign LUT_4[9600] = 32'b00000000000000001111011011010110;
assign LUT_4[9601] = 32'b00000000000000001000100111001110;
assign LUT_4[9602] = 32'b00000000000000001110110101111010;
assign LUT_4[9603] = 32'b00000000000000001000000001110010;
assign LUT_4[9604] = 32'b00000000000000001100011011110010;
assign LUT_4[9605] = 32'b00000000000000000101100111101010;
assign LUT_4[9606] = 32'b00000000000000001011110110010110;
assign LUT_4[9607] = 32'b00000000000000000101000010001110;
assign LUT_4[9608] = 32'b00000000000000001000100111101011;
assign LUT_4[9609] = 32'b00000000000000000001110011100011;
assign LUT_4[9610] = 32'b00000000000000001000000010001111;
assign LUT_4[9611] = 32'b00000000000000000001001110000111;
assign LUT_4[9612] = 32'b00000000000000000101101000000111;
assign LUT_4[9613] = 32'b11111111111111111110110011111111;
assign LUT_4[9614] = 32'b00000000000000000101000010101011;
assign LUT_4[9615] = 32'b11111111111111111110001110100011;
assign LUT_4[9616] = 32'b00000000000000001101001101000100;
assign LUT_4[9617] = 32'b00000000000000000110011000111100;
assign LUT_4[9618] = 32'b00000000000000001100100111101000;
assign LUT_4[9619] = 32'b00000000000000000101110011100000;
assign LUT_4[9620] = 32'b00000000000000001010001101100000;
assign LUT_4[9621] = 32'b00000000000000000011011001011000;
assign LUT_4[9622] = 32'b00000000000000001001101000000100;
assign LUT_4[9623] = 32'b00000000000000000010110011111100;
assign LUT_4[9624] = 32'b00000000000000000110011001011001;
assign LUT_4[9625] = 32'b11111111111111111111100101010001;
assign LUT_4[9626] = 32'b00000000000000000101110011111101;
assign LUT_4[9627] = 32'b11111111111111111110111111110101;
assign LUT_4[9628] = 32'b00000000000000000011011001110101;
assign LUT_4[9629] = 32'b11111111111111111100100101101101;
assign LUT_4[9630] = 32'b00000000000000000010110100011001;
assign LUT_4[9631] = 32'b11111111111111111100000000010001;
assign LUT_4[9632] = 32'b00000000000000001101110110011101;
assign LUT_4[9633] = 32'b00000000000000000111000010010101;
assign LUT_4[9634] = 32'b00000000000000001101010001000001;
assign LUT_4[9635] = 32'b00000000000000000110011100111001;
assign LUT_4[9636] = 32'b00000000000000001010110110111001;
assign LUT_4[9637] = 32'b00000000000000000100000010110001;
assign LUT_4[9638] = 32'b00000000000000001010010001011101;
assign LUT_4[9639] = 32'b00000000000000000011011101010101;
assign LUT_4[9640] = 32'b00000000000000000111000010110010;
assign LUT_4[9641] = 32'b00000000000000000000001110101010;
assign LUT_4[9642] = 32'b00000000000000000110011101010110;
assign LUT_4[9643] = 32'b11111111111111111111101001001110;
assign LUT_4[9644] = 32'b00000000000000000100000011001110;
assign LUT_4[9645] = 32'b11111111111111111101001111000110;
assign LUT_4[9646] = 32'b00000000000000000011011101110010;
assign LUT_4[9647] = 32'b11111111111111111100101001101010;
assign LUT_4[9648] = 32'b00000000000000001011101000001011;
assign LUT_4[9649] = 32'b00000000000000000100110100000011;
assign LUT_4[9650] = 32'b00000000000000001011000010101111;
assign LUT_4[9651] = 32'b00000000000000000100001110100111;
assign LUT_4[9652] = 32'b00000000000000001000101000100111;
assign LUT_4[9653] = 32'b00000000000000000001110100011111;
assign LUT_4[9654] = 32'b00000000000000001000000011001011;
assign LUT_4[9655] = 32'b00000000000000000001001111000011;
assign LUT_4[9656] = 32'b00000000000000000100110100100000;
assign LUT_4[9657] = 32'b11111111111111111110000000011000;
assign LUT_4[9658] = 32'b00000000000000000100001111000100;
assign LUT_4[9659] = 32'b11111111111111111101011010111100;
assign LUT_4[9660] = 32'b00000000000000000001110100111100;
assign LUT_4[9661] = 32'b11111111111111111011000000110100;
assign LUT_4[9662] = 32'b00000000000000000001001111100000;
assign LUT_4[9663] = 32'b11111111111111111010011011011000;
assign LUT_4[9664] = 32'b00000000000000010000110010101010;
assign LUT_4[9665] = 32'b00000000000000001001111110100010;
assign LUT_4[9666] = 32'b00000000000000010000001101001110;
assign LUT_4[9667] = 32'b00000000000000001001011001000110;
assign LUT_4[9668] = 32'b00000000000000001101110011000110;
assign LUT_4[9669] = 32'b00000000000000000110111110111110;
assign LUT_4[9670] = 32'b00000000000000001101001101101010;
assign LUT_4[9671] = 32'b00000000000000000110011001100010;
assign LUT_4[9672] = 32'b00000000000000001001111110111111;
assign LUT_4[9673] = 32'b00000000000000000011001010110111;
assign LUT_4[9674] = 32'b00000000000000001001011001100011;
assign LUT_4[9675] = 32'b00000000000000000010100101011011;
assign LUT_4[9676] = 32'b00000000000000000110111111011011;
assign LUT_4[9677] = 32'b00000000000000000000001011010011;
assign LUT_4[9678] = 32'b00000000000000000110011001111111;
assign LUT_4[9679] = 32'b11111111111111111111100101110111;
assign LUT_4[9680] = 32'b00000000000000001110100100011000;
assign LUT_4[9681] = 32'b00000000000000000111110000010000;
assign LUT_4[9682] = 32'b00000000000000001101111110111100;
assign LUT_4[9683] = 32'b00000000000000000111001010110100;
assign LUT_4[9684] = 32'b00000000000000001011100100110100;
assign LUT_4[9685] = 32'b00000000000000000100110000101100;
assign LUT_4[9686] = 32'b00000000000000001010111111011000;
assign LUT_4[9687] = 32'b00000000000000000100001011010000;
assign LUT_4[9688] = 32'b00000000000000000111110000101101;
assign LUT_4[9689] = 32'b00000000000000000000111100100101;
assign LUT_4[9690] = 32'b00000000000000000111001011010001;
assign LUT_4[9691] = 32'b00000000000000000000010111001001;
assign LUT_4[9692] = 32'b00000000000000000100110001001001;
assign LUT_4[9693] = 32'b11111111111111111101111101000001;
assign LUT_4[9694] = 32'b00000000000000000100001011101101;
assign LUT_4[9695] = 32'b11111111111111111101010111100101;
assign LUT_4[9696] = 32'b00000000000000001111001101110001;
assign LUT_4[9697] = 32'b00000000000000001000011001101001;
assign LUT_4[9698] = 32'b00000000000000001110101000010101;
assign LUT_4[9699] = 32'b00000000000000000111110100001101;
assign LUT_4[9700] = 32'b00000000000000001100001110001101;
assign LUT_4[9701] = 32'b00000000000000000101011010000101;
assign LUT_4[9702] = 32'b00000000000000001011101000110001;
assign LUT_4[9703] = 32'b00000000000000000100110100101001;
assign LUT_4[9704] = 32'b00000000000000001000011010000110;
assign LUT_4[9705] = 32'b00000000000000000001100101111110;
assign LUT_4[9706] = 32'b00000000000000000111110100101010;
assign LUT_4[9707] = 32'b00000000000000000001000000100010;
assign LUT_4[9708] = 32'b00000000000000000101011010100010;
assign LUT_4[9709] = 32'b11111111111111111110100110011010;
assign LUT_4[9710] = 32'b00000000000000000100110101000110;
assign LUT_4[9711] = 32'b11111111111111111110000000111110;
assign LUT_4[9712] = 32'b00000000000000001100111111011111;
assign LUT_4[9713] = 32'b00000000000000000110001011010111;
assign LUT_4[9714] = 32'b00000000000000001100011010000011;
assign LUT_4[9715] = 32'b00000000000000000101100101111011;
assign LUT_4[9716] = 32'b00000000000000001001111111111011;
assign LUT_4[9717] = 32'b00000000000000000011001011110011;
assign LUT_4[9718] = 32'b00000000000000001001011010011111;
assign LUT_4[9719] = 32'b00000000000000000010100110010111;
assign LUT_4[9720] = 32'b00000000000000000110001011110100;
assign LUT_4[9721] = 32'b11111111111111111111010111101100;
assign LUT_4[9722] = 32'b00000000000000000101100110011000;
assign LUT_4[9723] = 32'b11111111111111111110110010010000;
assign LUT_4[9724] = 32'b00000000000000000011001100010000;
assign LUT_4[9725] = 32'b11111111111111111100011000001000;
assign LUT_4[9726] = 32'b00000000000000000010100110110100;
assign LUT_4[9727] = 32'b11111111111111111011110010101100;
assign LUT_4[9728] = 32'b00000000000000000110111101110011;
assign LUT_4[9729] = 32'b00000000000000000000001001101011;
assign LUT_4[9730] = 32'b00000000000000000110011000010111;
assign LUT_4[9731] = 32'b11111111111111111111100100001111;
assign LUT_4[9732] = 32'b00000000000000000011111110001111;
assign LUT_4[9733] = 32'b11111111111111111101001010000111;
assign LUT_4[9734] = 32'b00000000000000000011011000110011;
assign LUT_4[9735] = 32'b11111111111111111100100100101011;
assign LUT_4[9736] = 32'b00000000000000000000001010001000;
assign LUT_4[9737] = 32'b11111111111111111001010110000000;
assign LUT_4[9738] = 32'b11111111111111111111100100101100;
assign LUT_4[9739] = 32'b11111111111111111000110000100100;
assign LUT_4[9740] = 32'b11111111111111111101001010100100;
assign LUT_4[9741] = 32'b11111111111111110110010110011100;
assign LUT_4[9742] = 32'b11111111111111111100100101001000;
assign LUT_4[9743] = 32'b11111111111111110101110001000000;
assign LUT_4[9744] = 32'b00000000000000000100101111100001;
assign LUT_4[9745] = 32'b11111111111111111101111011011001;
assign LUT_4[9746] = 32'b00000000000000000100001010000101;
assign LUT_4[9747] = 32'b11111111111111111101010101111101;
assign LUT_4[9748] = 32'b00000000000000000001101111111101;
assign LUT_4[9749] = 32'b11111111111111111010111011110101;
assign LUT_4[9750] = 32'b00000000000000000001001010100001;
assign LUT_4[9751] = 32'b11111111111111111010010110011001;
assign LUT_4[9752] = 32'b11111111111111111101111011110110;
assign LUT_4[9753] = 32'b11111111111111110111000111101110;
assign LUT_4[9754] = 32'b11111111111111111101010110011010;
assign LUT_4[9755] = 32'b11111111111111110110100010010010;
assign LUT_4[9756] = 32'b11111111111111111010111100010010;
assign LUT_4[9757] = 32'b11111111111111110100001000001010;
assign LUT_4[9758] = 32'b11111111111111111010010110110110;
assign LUT_4[9759] = 32'b11111111111111110011100010101110;
assign LUT_4[9760] = 32'b00000000000000000101011000111010;
assign LUT_4[9761] = 32'b11111111111111111110100100110010;
assign LUT_4[9762] = 32'b00000000000000000100110011011110;
assign LUT_4[9763] = 32'b11111111111111111101111111010110;
assign LUT_4[9764] = 32'b00000000000000000010011001010110;
assign LUT_4[9765] = 32'b11111111111111111011100101001110;
assign LUT_4[9766] = 32'b00000000000000000001110011111010;
assign LUT_4[9767] = 32'b11111111111111111010111111110010;
assign LUT_4[9768] = 32'b11111111111111111110100101001111;
assign LUT_4[9769] = 32'b11111111111111110111110001000111;
assign LUT_4[9770] = 32'b11111111111111111101111111110011;
assign LUT_4[9771] = 32'b11111111111111110111001011101011;
assign LUT_4[9772] = 32'b11111111111111111011100101101011;
assign LUT_4[9773] = 32'b11111111111111110100110001100011;
assign LUT_4[9774] = 32'b11111111111111111011000000001111;
assign LUT_4[9775] = 32'b11111111111111110100001100000111;
assign LUT_4[9776] = 32'b00000000000000000011001010101000;
assign LUT_4[9777] = 32'b11111111111111111100010110100000;
assign LUT_4[9778] = 32'b00000000000000000010100101001100;
assign LUT_4[9779] = 32'b11111111111111111011110001000100;
assign LUT_4[9780] = 32'b00000000000000000000001011000100;
assign LUT_4[9781] = 32'b11111111111111111001010110111100;
assign LUT_4[9782] = 32'b11111111111111111111100101101000;
assign LUT_4[9783] = 32'b11111111111111111000110001100000;
assign LUT_4[9784] = 32'b11111111111111111100010110111101;
assign LUT_4[9785] = 32'b11111111111111110101100010110101;
assign LUT_4[9786] = 32'b11111111111111111011110001100001;
assign LUT_4[9787] = 32'b11111111111111110100111101011001;
assign LUT_4[9788] = 32'b11111111111111111001010111011001;
assign LUT_4[9789] = 32'b11111111111111110010100011010001;
assign LUT_4[9790] = 32'b11111111111111111000110001111101;
assign LUT_4[9791] = 32'b11111111111111110001111101110101;
assign LUT_4[9792] = 32'b00000000000000001000010101000111;
assign LUT_4[9793] = 32'b00000000000000000001100000111111;
assign LUT_4[9794] = 32'b00000000000000000111101111101011;
assign LUT_4[9795] = 32'b00000000000000000000111011100011;
assign LUT_4[9796] = 32'b00000000000000000101010101100011;
assign LUT_4[9797] = 32'b11111111111111111110100001011011;
assign LUT_4[9798] = 32'b00000000000000000100110000000111;
assign LUT_4[9799] = 32'b11111111111111111101111011111111;
assign LUT_4[9800] = 32'b00000000000000000001100001011100;
assign LUT_4[9801] = 32'b11111111111111111010101101010100;
assign LUT_4[9802] = 32'b00000000000000000000111100000000;
assign LUT_4[9803] = 32'b11111111111111111010000111111000;
assign LUT_4[9804] = 32'b11111111111111111110100001111000;
assign LUT_4[9805] = 32'b11111111111111110111101101110000;
assign LUT_4[9806] = 32'b11111111111111111101111100011100;
assign LUT_4[9807] = 32'b11111111111111110111001000010100;
assign LUT_4[9808] = 32'b00000000000000000110000110110101;
assign LUT_4[9809] = 32'b11111111111111111111010010101101;
assign LUT_4[9810] = 32'b00000000000000000101100001011001;
assign LUT_4[9811] = 32'b11111111111111111110101101010001;
assign LUT_4[9812] = 32'b00000000000000000011000111010001;
assign LUT_4[9813] = 32'b11111111111111111100010011001001;
assign LUT_4[9814] = 32'b00000000000000000010100001110101;
assign LUT_4[9815] = 32'b11111111111111111011101101101101;
assign LUT_4[9816] = 32'b11111111111111111111010011001010;
assign LUT_4[9817] = 32'b11111111111111111000011111000010;
assign LUT_4[9818] = 32'b11111111111111111110101101101110;
assign LUT_4[9819] = 32'b11111111111111110111111001100110;
assign LUT_4[9820] = 32'b11111111111111111100010011100110;
assign LUT_4[9821] = 32'b11111111111111110101011111011110;
assign LUT_4[9822] = 32'b11111111111111111011101110001010;
assign LUT_4[9823] = 32'b11111111111111110100111010000010;
assign LUT_4[9824] = 32'b00000000000000000110110000001110;
assign LUT_4[9825] = 32'b11111111111111111111111100000110;
assign LUT_4[9826] = 32'b00000000000000000110001010110010;
assign LUT_4[9827] = 32'b11111111111111111111010110101010;
assign LUT_4[9828] = 32'b00000000000000000011110000101010;
assign LUT_4[9829] = 32'b11111111111111111100111100100010;
assign LUT_4[9830] = 32'b00000000000000000011001011001110;
assign LUT_4[9831] = 32'b11111111111111111100010111000110;
assign LUT_4[9832] = 32'b11111111111111111111111100100011;
assign LUT_4[9833] = 32'b11111111111111111001001000011011;
assign LUT_4[9834] = 32'b11111111111111111111010111000111;
assign LUT_4[9835] = 32'b11111111111111111000100010111111;
assign LUT_4[9836] = 32'b11111111111111111100111100111111;
assign LUT_4[9837] = 32'b11111111111111110110001000110111;
assign LUT_4[9838] = 32'b11111111111111111100010111100011;
assign LUT_4[9839] = 32'b11111111111111110101100011011011;
assign LUT_4[9840] = 32'b00000000000000000100100001111100;
assign LUT_4[9841] = 32'b11111111111111111101101101110100;
assign LUT_4[9842] = 32'b00000000000000000011111100100000;
assign LUT_4[9843] = 32'b11111111111111111101001000011000;
assign LUT_4[9844] = 32'b00000000000000000001100010011000;
assign LUT_4[9845] = 32'b11111111111111111010101110010000;
assign LUT_4[9846] = 32'b00000000000000000000111100111100;
assign LUT_4[9847] = 32'b11111111111111111010001000110100;
assign LUT_4[9848] = 32'b11111111111111111101101110010001;
assign LUT_4[9849] = 32'b11111111111111110110111010001001;
assign LUT_4[9850] = 32'b11111111111111111101001000110101;
assign LUT_4[9851] = 32'b11111111111111110110010100101101;
assign LUT_4[9852] = 32'b11111111111111111010101110101101;
assign LUT_4[9853] = 32'b11111111111111110011111010100101;
assign LUT_4[9854] = 32'b11111111111111111010001001010001;
assign LUT_4[9855] = 32'b11111111111111110011010101001001;
assign LUT_4[9856] = 32'b00000000000000001001100011111011;
assign LUT_4[9857] = 32'b00000000000000000010101111110011;
assign LUT_4[9858] = 32'b00000000000000001000111110011111;
assign LUT_4[9859] = 32'b00000000000000000010001010010111;
assign LUT_4[9860] = 32'b00000000000000000110100100010111;
assign LUT_4[9861] = 32'b11111111111111111111110000001111;
assign LUT_4[9862] = 32'b00000000000000000101111110111011;
assign LUT_4[9863] = 32'b11111111111111111111001010110011;
assign LUT_4[9864] = 32'b00000000000000000010110000010000;
assign LUT_4[9865] = 32'b11111111111111111011111100001000;
assign LUT_4[9866] = 32'b00000000000000000010001010110100;
assign LUT_4[9867] = 32'b11111111111111111011010110101100;
assign LUT_4[9868] = 32'b11111111111111111111110000101100;
assign LUT_4[9869] = 32'b11111111111111111000111100100100;
assign LUT_4[9870] = 32'b11111111111111111111001011010000;
assign LUT_4[9871] = 32'b11111111111111111000010111001000;
assign LUT_4[9872] = 32'b00000000000000000111010101101001;
assign LUT_4[9873] = 32'b00000000000000000000100001100001;
assign LUT_4[9874] = 32'b00000000000000000110110000001101;
assign LUT_4[9875] = 32'b11111111111111111111111100000101;
assign LUT_4[9876] = 32'b00000000000000000100010110000101;
assign LUT_4[9877] = 32'b11111111111111111101100001111101;
assign LUT_4[9878] = 32'b00000000000000000011110000101001;
assign LUT_4[9879] = 32'b11111111111111111100111100100001;
assign LUT_4[9880] = 32'b00000000000000000000100001111110;
assign LUT_4[9881] = 32'b11111111111111111001101101110110;
assign LUT_4[9882] = 32'b11111111111111111111111100100010;
assign LUT_4[9883] = 32'b11111111111111111001001000011010;
assign LUT_4[9884] = 32'b11111111111111111101100010011010;
assign LUT_4[9885] = 32'b11111111111111110110101110010010;
assign LUT_4[9886] = 32'b11111111111111111100111100111110;
assign LUT_4[9887] = 32'b11111111111111110110001000110110;
assign LUT_4[9888] = 32'b00000000000000000111111111000010;
assign LUT_4[9889] = 32'b00000000000000000001001010111010;
assign LUT_4[9890] = 32'b00000000000000000111011001100110;
assign LUT_4[9891] = 32'b00000000000000000000100101011110;
assign LUT_4[9892] = 32'b00000000000000000100111111011110;
assign LUT_4[9893] = 32'b11111111111111111110001011010110;
assign LUT_4[9894] = 32'b00000000000000000100011010000010;
assign LUT_4[9895] = 32'b11111111111111111101100101111010;
assign LUT_4[9896] = 32'b00000000000000000001001011010111;
assign LUT_4[9897] = 32'b11111111111111111010010111001111;
assign LUT_4[9898] = 32'b00000000000000000000100101111011;
assign LUT_4[9899] = 32'b11111111111111111001110001110011;
assign LUT_4[9900] = 32'b11111111111111111110001011110011;
assign LUT_4[9901] = 32'b11111111111111110111010111101011;
assign LUT_4[9902] = 32'b11111111111111111101100110010111;
assign LUT_4[9903] = 32'b11111111111111110110110010001111;
assign LUT_4[9904] = 32'b00000000000000000101110000110000;
assign LUT_4[9905] = 32'b11111111111111111110111100101000;
assign LUT_4[9906] = 32'b00000000000000000101001011010100;
assign LUT_4[9907] = 32'b11111111111111111110010111001100;
assign LUT_4[9908] = 32'b00000000000000000010110001001100;
assign LUT_4[9909] = 32'b11111111111111111011111101000100;
assign LUT_4[9910] = 32'b00000000000000000010001011110000;
assign LUT_4[9911] = 32'b11111111111111111011010111101000;
assign LUT_4[9912] = 32'b11111111111111111110111101000101;
assign LUT_4[9913] = 32'b11111111111111111000001000111101;
assign LUT_4[9914] = 32'b11111111111111111110010111101001;
assign LUT_4[9915] = 32'b11111111111111110111100011100001;
assign LUT_4[9916] = 32'b11111111111111111011111101100001;
assign LUT_4[9917] = 32'b11111111111111110101001001011001;
assign LUT_4[9918] = 32'b11111111111111111011011000000101;
assign LUT_4[9919] = 32'b11111111111111110100100011111101;
assign LUT_4[9920] = 32'b00000000000000001010111011001111;
assign LUT_4[9921] = 32'b00000000000000000100000111000111;
assign LUT_4[9922] = 32'b00000000000000001010010101110011;
assign LUT_4[9923] = 32'b00000000000000000011100001101011;
assign LUT_4[9924] = 32'b00000000000000000111111011101011;
assign LUT_4[9925] = 32'b00000000000000000001000111100011;
assign LUT_4[9926] = 32'b00000000000000000111010110001111;
assign LUT_4[9927] = 32'b00000000000000000000100010000111;
assign LUT_4[9928] = 32'b00000000000000000100000111100100;
assign LUT_4[9929] = 32'b11111111111111111101010011011100;
assign LUT_4[9930] = 32'b00000000000000000011100010001000;
assign LUT_4[9931] = 32'b11111111111111111100101110000000;
assign LUT_4[9932] = 32'b00000000000000000001001000000000;
assign LUT_4[9933] = 32'b11111111111111111010010011111000;
assign LUT_4[9934] = 32'b00000000000000000000100010100100;
assign LUT_4[9935] = 32'b11111111111111111001101110011100;
assign LUT_4[9936] = 32'b00000000000000001000101100111101;
assign LUT_4[9937] = 32'b00000000000000000001111000110101;
assign LUT_4[9938] = 32'b00000000000000001000000111100001;
assign LUT_4[9939] = 32'b00000000000000000001010011011001;
assign LUT_4[9940] = 32'b00000000000000000101101101011001;
assign LUT_4[9941] = 32'b11111111111111111110111001010001;
assign LUT_4[9942] = 32'b00000000000000000101000111111101;
assign LUT_4[9943] = 32'b11111111111111111110010011110101;
assign LUT_4[9944] = 32'b00000000000000000001111001010010;
assign LUT_4[9945] = 32'b11111111111111111011000101001010;
assign LUT_4[9946] = 32'b00000000000000000001010011110110;
assign LUT_4[9947] = 32'b11111111111111111010011111101110;
assign LUT_4[9948] = 32'b11111111111111111110111001101110;
assign LUT_4[9949] = 32'b11111111111111111000000101100110;
assign LUT_4[9950] = 32'b11111111111111111110010100010010;
assign LUT_4[9951] = 32'b11111111111111110111100000001010;
assign LUT_4[9952] = 32'b00000000000000001001010110010110;
assign LUT_4[9953] = 32'b00000000000000000010100010001110;
assign LUT_4[9954] = 32'b00000000000000001000110000111010;
assign LUT_4[9955] = 32'b00000000000000000001111100110010;
assign LUT_4[9956] = 32'b00000000000000000110010110110010;
assign LUT_4[9957] = 32'b11111111111111111111100010101010;
assign LUT_4[9958] = 32'b00000000000000000101110001010110;
assign LUT_4[9959] = 32'b11111111111111111110111101001110;
assign LUT_4[9960] = 32'b00000000000000000010100010101011;
assign LUT_4[9961] = 32'b11111111111111111011101110100011;
assign LUT_4[9962] = 32'b00000000000000000001111101001111;
assign LUT_4[9963] = 32'b11111111111111111011001001000111;
assign LUT_4[9964] = 32'b11111111111111111111100011000111;
assign LUT_4[9965] = 32'b11111111111111111000101110111111;
assign LUT_4[9966] = 32'b11111111111111111110111101101011;
assign LUT_4[9967] = 32'b11111111111111111000001001100011;
assign LUT_4[9968] = 32'b00000000000000000111001000000100;
assign LUT_4[9969] = 32'b00000000000000000000010011111100;
assign LUT_4[9970] = 32'b00000000000000000110100010101000;
assign LUT_4[9971] = 32'b11111111111111111111101110100000;
assign LUT_4[9972] = 32'b00000000000000000100001000100000;
assign LUT_4[9973] = 32'b11111111111111111101010100011000;
assign LUT_4[9974] = 32'b00000000000000000011100011000100;
assign LUT_4[9975] = 32'b11111111111111111100101110111100;
assign LUT_4[9976] = 32'b00000000000000000000010100011001;
assign LUT_4[9977] = 32'b11111111111111111001100000010001;
assign LUT_4[9978] = 32'b11111111111111111111101110111101;
assign LUT_4[9979] = 32'b11111111111111111000111010110101;
assign LUT_4[9980] = 32'b11111111111111111101010100110101;
assign LUT_4[9981] = 32'b11111111111111110110100000101101;
assign LUT_4[9982] = 32'b11111111111111111100101111011001;
assign LUT_4[9983] = 32'b11111111111111110101111011010001;
assign LUT_4[9984] = 32'b00000000000000001011111001010110;
assign LUT_4[9985] = 32'b00000000000000000101000101001110;
assign LUT_4[9986] = 32'b00000000000000001011010011111010;
assign LUT_4[9987] = 32'b00000000000000000100011111110010;
assign LUT_4[9988] = 32'b00000000000000001000111001110010;
assign LUT_4[9989] = 32'b00000000000000000010000101101010;
assign LUT_4[9990] = 32'b00000000000000001000010100010110;
assign LUT_4[9991] = 32'b00000000000000000001100000001110;
assign LUT_4[9992] = 32'b00000000000000000101000101101011;
assign LUT_4[9993] = 32'b11111111111111111110010001100011;
assign LUT_4[9994] = 32'b00000000000000000100100000001111;
assign LUT_4[9995] = 32'b11111111111111111101101100000111;
assign LUT_4[9996] = 32'b00000000000000000010000110000111;
assign LUT_4[9997] = 32'b11111111111111111011010001111111;
assign LUT_4[9998] = 32'b00000000000000000001100000101011;
assign LUT_4[9999] = 32'b11111111111111111010101100100011;
assign LUT_4[10000] = 32'b00000000000000001001101011000100;
assign LUT_4[10001] = 32'b00000000000000000010110110111100;
assign LUT_4[10002] = 32'b00000000000000001001000101101000;
assign LUT_4[10003] = 32'b00000000000000000010010001100000;
assign LUT_4[10004] = 32'b00000000000000000110101011100000;
assign LUT_4[10005] = 32'b11111111111111111111110111011000;
assign LUT_4[10006] = 32'b00000000000000000110000110000100;
assign LUT_4[10007] = 32'b11111111111111111111010001111100;
assign LUT_4[10008] = 32'b00000000000000000010110111011001;
assign LUT_4[10009] = 32'b11111111111111111100000011010001;
assign LUT_4[10010] = 32'b00000000000000000010010001111101;
assign LUT_4[10011] = 32'b11111111111111111011011101110101;
assign LUT_4[10012] = 32'b11111111111111111111110111110101;
assign LUT_4[10013] = 32'b11111111111111111001000011101101;
assign LUT_4[10014] = 32'b11111111111111111111010010011001;
assign LUT_4[10015] = 32'b11111111111111111000011110010001;
assign LUT_4[10016] = 32'b00000000000000001010010100011101;
assign LUT_4[10017] = 32'b00000000000000000011100000010101;
assign LUT_4[10018] = 32'b00000000000000001001101111000001;
assign LUT_4[10019] = 32'b00000000000000000010111010111001;
assign LUT_4[10020] = 32'b00000000000000000111010100111001;
assign LUT_4[10021] = 32'b00000000000000000000100000110001;
assign LUT_4[10022] = 32'b00000000000000000110101111011101;
assign LUT_4[10023] = 32'b11111111111111111111111011010101;
assign LUT_4[10024] = 32'b00000000000000000011100000110010;
assign LUT_4[10025] = 32'b11111111111111111100101100101010;
assign LUT_4[10026] = 32'b00000000000000000010111011010110;
assign LUT_4[10027] = 32'b11111111111111111100000111001110;
assign LUT_4[10028] = 32'b00000000000000000000100001001110;
assign LUT_4[10029] = 32'b11111111111111111001101101000110;
assign LUT_4[10030] = 32'b11111111111111111111111011110010;
assign LUT_4[10031] = 32'b11111111111111111001000111101010;
assign LUT_4[10032] = 32'b00000000000000001000000110001011;
assign LUT_4[10033] = 32'b00000000000000000001010010000011;
assign LUT_4[10034] = 32'b00000000000000000111100000101111;
assign LUT_4[10035] = 32'b00000000000000000000101100100111;
assign LUT_4[10036] = 32'b00000000000000000101000110100111;
assign LUT_4[10037] = 32'b11111111111111111110010010011111;
assign LUT_4[10038] = 32'b00000000000000000100100001001011;
assign LUT_4[10039] = 32'b11111111111111111101101101000011;
assign LUT_4[10040] = 32'b00000000000000000001010010100000;
assign LUT_4[10041] = 32'b11111111111111111010011110011000;
assign LUT_4[10042] = 32'b00000000000000000000101101000100;
assign LUT_4[10043] = 32'b11111111111111111001111000111100;
assign LUT_4[10044] = 32'b11111111111111111110010010111100;
assign LUT_4[10045] = 32'b11111111111111110111011110110100;
assign LUT_4[10046] = 32'b11111111111111111101101101100000;
assign LUT_4[10047] = 32'b11111111111111110110111001011000;
assign LUT_4[10048] = 32'b00000000000000001101010000101010;
assign LUT_4[10049] = 32'b00000000000000000110011100100010;
assign LUT_4[10050] = 32'b00000000000000001100101011001110;
assign LUT_4[10051] = 32'b00000000000000000101110111000110;
assign LUT_4[10052] = 32'b00000000000000001010010001000110;
assign LUT_4[10053] = 32'b00000000000000000011011100111110;
assign LUT_4[10054] = 32'b00000000000000001001101011101010;
assign LUT_4[10055] = 32'b00000000000000000010110111100010;
assign LUT_4[10056] = 32'b00000000000000000110011100111111;
assign LUT_4[10057] = 32'b11111111111111111111101000110111;
assign LUT_4[10058] = 32'b00000000000000000101110111100011;
assign LUT_4[10059] = 32'b11111111111111111111000011011011;
assign LUT_4[10060] = 32'b00000000000000000011011101011011;
assign LUT_4[10061] = 32'b11111111111111111100101001010011;
assign LUT_4[10062] = 32'b00000000000000000010110111111111;
assign LUT_4[10063] = 32'b11111111111111111100000011110111;
assign LUT_4[10064] = 32'b00000000000000001011000010011000;
assign LUT_4[10065] = 32'b00000000000000000100001110010000;
assign LUT_4[10066] = 32'b00000000000000001010011100111100;
assign LUT_4[10067] = 32'b00000000000000000011101000110100;
assign LUT_4[10068] = 32'b00000000000000001000000010110100;
assign LUT_4[10069] = 32'b00000000000000000001001110101100;
assign LUT_4[10070] = 32'b00000000000000000111011101011000;
assign LUT_4[10071] = 32'b00000000000000000000101001010000;
assign LUT_4[10072] = 32'b00000000000000000100001110101101;
assign LUT_4[10073] = 32'b11111111111111111101011010100101;
assign LUT_4[10074] = 32'b00000000000000000011101001010001;
assign LUT_4[10075] = 32'b11111111111111111100110101001001;
assign LUT_4[10076] = 32'b00000000000000000001001111001001;
assign LUT_4[10077] = 32'b11111111111111111010011011000001;
assign LUT_4[10078] = 32'b00000000000000000000101001101101;
assign LUT_4[10079] = 32'b11111111111111111001110101100101;
assign LUT_4[10080] = 32'b00000000000000001011101011110001;
assign LUT_4[10081] = 32'b00000000000000000100110111101001;
assign LUT_4[10082] = 32'b00000000000000001011000110010101;
assign LUT_4[10083] = 32'b00000000000000000100010010001101;
assign LUT_4[10084] = 32'b00000000000000001000101100001101;
assign LUT_4[10085] = 32'b00000000000000000001111000000101;
assign LUT_4[10086] = 32'b00000000000000001000000110110001;
assign LUT_4[10087] = 32'b00000000000000000001010010101001;
assign LUT_4[10088] = 32'b00000000000000000100111000000110;
assign LUT_4[10089] = 32'b11111111111111111110000011111110;
assign LUT_4[10090] = 32'b00000000000000000100010010101010;
assign LUT_4[10091] = 32'b11111111111111111101011110100010;
assign LUT_4[10092] = 32'b00000000000000000001111000100010;
assign LUT_4[10093] = 32'b11111111111111111011000100011010;
assign LUT_4[10094] = 32'b00000000000000000001010011000110;
assign LUT_4[10095] = 32'b11111111111111111010011110111110;
assign LUT_4[10096] = 32'b00000000000000001001011101011111;
assign LUT_4[10097] = 32'b00000000000000000010101001010111;
assign LUT_4[10098] = 32'b00000000000000001000111000000011;
assign LUT_4[10099] = 32'b00000000000000000010000011111011;
assign LUT_4[10100] = 32'b00000000000000000110011101111011;
assign LUT_4[10101] = 32'b11111111111111111111101001110011;
assign LUT_4[10102] = 32'b00000000000000000101111000011111;
assign LUT_4[10103] = 32'b11111111111111111111000100010111;
assign LUT_4[10104] = 32'b00000000000000000010101001110100;
assign LUT_4[10105] = 32'b11111111111111111011110101101100;
assign LUT_4[10106] = 32'b00000000000000000010000100011000;
assign LUT_4[10107] = 32'b11111111111111111011010000010000;
assign LUT_4[10108] = 32'b11111111111111111111101010010000;
assign LUT_4[10109] = 32'b11111111111111111000110110001000;
assign LUT_4[10110] = 32'b11111111111111111111000100110100;
assign LUT_4[10111] = 32'b11111111111111111000010000101100;
assign LUT_4[10112] = 32'b00000000000000001110011111011110;
assign LUT_4[10113] = 32'b00000000000000000111101011010110;
assign LUT_4[10114] = 32'b00000000000000001101111010000010;
assign LUT_4[10115] = 32'b00000000000000000111000101111010;
assign LUT_4[10116] = 32'b00000000000000001011011111111010;
assign LUT_4[10117] = 32'b00000000000000000100101011110010;
assign LUT_4[10118] = 32'b00000000000000001010111010011110;
assign LUT_4[10119] = 32'b00000000000000000100000110010110;
assign LUT_4[10120] = 32'b00000000000000000111101011110011;
assign LUT_4[10121] = 32'b00000000000000000000110111101011;
assign LUT_4[10122] = 32'b00000000000000000111000110010111;
assign LUT_4[10123] = 32'b00000000000000000000010010001111;
assign LUT_4[10124] = 32'b00000000000000000100101100001111;
assign LUT_4[10125] = 32'b11111111111111111101111000000111;
assign LUT_4[10126] = 32'b00000000000000000100000110110011;
assign LUT_4[10127] = 32'b11111111111111111101010010101011;
assign LUT_4[10128] = 32'b00000000000000001100010001001100;
assign LUT_4[10129] = 32'b00000000000000000101011101000100;
assign LUT_4[10130] = 32'b00000000000000001011101011110000;
assign LUT_4[10131] = 32'b00000000000000000100110111101000;
assign LUT_4[10132] = 32'b00000000000000001001010001101000;
assign LUT_4[10133] = 32'b00000000000000000010011101100000;
assign LUT_4[10134] = 32'b00000000000000001000101100001100;
assign LUT_4[10135] = 32'b00000000000000000001111000000100;
assign LUT_4[10136] = 32'b00000000000000000101011101100001;
assign LUT_4[10137] = 32'b11111111111111111110101001011001;
assign LUT_4[10138] = 32'b00000000000000000100111000000101;
assign LUT_4[10139] = 32'b11111111111111111110000011111101;
assign LUT_4[10140] = 32'b00000000000000000010011101111101;
assign LUT_4[10141] = 32'b11111111111111111011101001110101;
assign LUT_4[10142] = 32'b00000000000000000001111000100001;
assign LUT_4[10143] = 32'b11111111111111111011000100011001;
assign LUT_4[10144] = 32'b00000000000000001100111010100101;
assign LUT_4[10145] = 32'b00000000000000000110000110011101;
assign LUT_4[10146] = 32'b00000000000000001100010101001001;
assign LUT_4[10147] = 32'b00000000000000000101100001000001;
assign LUT_4[10148] = 32'b00000000000000001001111011000001;
assign LUT_4[10149] = 32'b00000000000000000011000110111001;
assign LUT_4[10150] = 32'b00000000000000001001010101100101;
assign LUT_4[10151] = 32'b00000000000000000010100001011101;
assign LUT_4[10152] = 32'b00000000000000000110000110111010;
assign LUT_4[10153] = 32'b11111111111111111111010010110010;
assign LUT_4[10154] = 32'b00000000000000000101100001011110;
assign LUT_4[10155] = 32'b11111111111111111110101101010110;
assign LUT_4[10156] = 32'b00000000000000000011000111010110;
assign LUT_4[10157] = 32'b11111111111111111100010011001110;
assign LUT_4[10158] = 32'b00000000000000000010100001111010;
assign LUT_4[10159] = 32'b11111111111111111011101101110010;
assign LUT_4[10160] = 32'b00000000000000001010101100010011;
assign LUT_4[10161] = 32'b00000000000000000011111000001011;
assign LUT_4[10162] = 32'b00000000000000001010000110110111;
assign LUT_4[10163] = 32'b00000000000000000011010010101111;
assign LUT_4[10164] = 32'b00000000000000000111101100101111;
assign LUT_4[10165] = 32'b00000000000000000000111000100111;
assign LUT_4[10166] = 32'b00000000000000000111000111010011;
assign LUT_4[10167] = 32'b00000000000000000000010011001011;
assign LUT_4[10168] = 32'b00000000000000000011111000101000;
assign LUT_4[10169] = 32'b11111111111111111101000100100000;
assign LUT_4[10170] = 32'b00000000000000000011010011001100;
assign LUT_4[10171] = 32'b11111111111111111100011111000100;
assign LUT_4[10172] = 32'b00000000000000000000111001000100;
assign LUT_4[10173] = 32'b11111111111111111010000100111100;
assign LUT_4[10174] = 32'b00000000000000000000010011101000;
assign LUT_4[10175] = 32'b11111111111111111001011111100000;
assign LUT_4[10176] = 32'b00000000000000001111110110110010;
assign LUT_4[10177] = 32'b00000000000000001001000010101010;
assign LUT_4[10178] = 32'b00000000000000001111010001010110;
assign LUT_4[10179] = 32'b00000000000000001000011101001110;
assign LUT_4[10180] = 32'b00000000000000001100110111001110;
assign LUT_4[10181] = 32'b00000000000000000110000011000110;
assign LUT_4[10182] = 32'b00000000000000001100010001110010;
assign LUT_4[10183] = 32'b00000000000000000101011101101010;
assign LUT_4[10184] = 32'b00000000000000001001000011000111;
assign LUT_4[10185] = 32'b00000000000000000010001110111111;
assign LUT_4[10186] = 32'b00000000000000001000011101101011;
assign LUT_4[10187] = 32'b00000000000000000001101001100011;
assign LUT_4[10188] = 32'b00000000000000000110000011100011;
assign LUT_4[10189] = 32'b11111111111111111111001111011011;
assign LUT_4[10190] = 32'b00000000000000000101011110000111;
assign LUT_4[10191] = 32'b11111111111111111110101001111111;
assign LUT_4[10192] = 32'b00000000000000001101101000100000;
assign LUT_4[10193] = 32'b00000000000000000110110100011000;
assign LUT_4[10194] = 32'b00000000000000001101000011000100;
assign LUT_4[10195] = 32'b00000000000000000110001110111100;
assign LUT_4[10196] = 32'b00000000000000001010101000111100;
assign LUT_4[10197] = 32'b00000000000000000011110100110100;
assign LUT_4[10198] = 32'b00000000000000001010000011100000;
assign LUT_4[10199] = 32'b00000000000000000011001111011000;
assign LUT_4[10200] = 32'b00000000000000000110110100110101;
assign LUT_4[10201] = 32'b00000000000000000000000000101101;
assign LUT_4[10202] = 32'b00000000000000000110001111011001;
assign LUT_4[10203] = 32'b11111111111111111111011011010001;
assign LUT_4[10204] = 32'b00000000000000000011110101010001;
assign LUT_4[10205] = 32'b11111111111111111101000001001001;
assign LUT_4[10206] = 32'b00000000000000000011001111110101;
assign LUT_4[10207] = 32'b11111111111111111100011011101101;
assign LUT_4[10208] = 32'b00000000000000001110010001111001;
assign LUT_4[10209] = 32'b00000000000000000111011101110001;
assign LUT_4[10210] = 32'b00000000000000001101101100011101;
assign LUT_4[10211] = 32'b00000000000000000110111000010101;
assign LUT_4[10212] = 32'b00000000000000001011010010010101;
assign LUT_4[10213] = 32'b00000000000000000100011110001101;
assign LUT_4[10214] = 32'b00000000000000001010101100111001;
assign LUT_4[10215] = 32'b00000000000000000011111000110001;
assign LUT_4[10216] = 32'b00000000000000000111011110001110;
assign LUT_4[10217] = 32'b00000000000000000000101010000110;
assign LUT_4[10218] = 32'b00000000000000000110111000110010;
assign LUT_4[10219] = 32'b00000000000000000000000100101010;
assign LUT_4[10220] = 32'b00000000000000000100011110101010;
assign LUT_4[10221] = 32'b11111111111111111101101010100010;
assign LUT_4[10222] = 32'b00000000000000000011111001001110;
assign LUT_4[10223] = 32'b11111111111111111101000101000110;
assign LUT_4[10224] = 32'b00000000000000001100000011100111;
assign LUT_4[10225] = 32'b00000000000000000101001111011111;
assign LUT_4[10226] = 32'b00000000000000001011011110001011;
assign LUT_4[10227] = 32'b00000000000000000100101010000011;
assign LUT_4[10228] = 32'b00000000000000001001000100000011;
assign LUT_4[10229] = 32'b00000000000000000010001111111011;
assign LUT_4[10230] = 32'b00000000000000001000011110100111;
assign LUT_4[10231] = 32'b00000000000000000001101010011111;
assign LUT_4[10232] = 32'b00000000000000000101001111111100;
assign LUT_4[10233] = 32'b11111111111111111110011011110100;
assign LUT_4[10234] = 32'b00000000000000000100101010100000;
assign LUT_4[10235] = 32'b11111111111111111101110110011000;
assign LUT_4[10236] = 32'b00000000000000000010010000011000;
assign LUT_4[10237] = 32'b11111111111111111011011100010000;
assign LUT_4[10238] = 32'b00000000000000000001101010111100;
assign LUT_4[10239] = 32'b11111111111111111010110110110100;
assign LUT_4[10240] = 32'b00000000000000000001101110010110;
assign LUT_4[10241] = 32'b11111111111111111010111010001110;
assign LUT_4[10242] = 32'b00000000000000000001001000111010;
assign LUT_4[10243] = 32'b11111111111111111010010100110010;
assign LUT_4[10244] = 32'b11111111111111111110101110110010;
assign LUT_4[10245] = 32'b11111111111111110111111010101010;
assign LUT_4[10246] = 32'b11111111111111111110001001010110;
assign LUT_4[10247] = 32'b11111111111111110111010101001110;
assign LUT_4[10248] = 32'b11111111111111111010111010101011;
assign LUT_4[10249] = 32'b11111111111111110100000110100011;
assign LUT_4[10250] = 32'b11111111111111111010010101001111;
assign LUT_4[10251] = 32'b11111111111111110011100001000111;
assign LUT_4[10252] = 32'b11111111111111110111111011000111;
assign LUT_4[10253] = 32'b11111111111111110001000110111111;
assign LUT_4[10254] = 32'b11111111111111110111010101101011;
assign LUT_4[10255] = 32'b11111111111111110000100001100011;
assign LUT_4[10256] = 32'b11111111111111111111100000000100;
assign LUT_4[10257] = 32'b11111111111111111000101011111100;
assign LUT_4[10258] = 32'b11111111111111111110111010101000;
assign LUT_4[10259] = 32'b11111111111111111000000110100000;
assign LUT_4[10260] = 32'b11111111111111111100100000100000;
assign LUT_4[10261] = 32'b11111111111111110101101100011000;
assign LUT_4[10262] = 32'b11111111111111111011111011000100;
assign LUT_4[10263] = 32'b11111111111111110101000110111100;
assign LUT_4[10264] = 32'b11111111111111111000101100011001;
assign LUT_4[10265] = 32'b11111111111111110001111000010001;
assign LUT_4[10266] = 32'b11111111111111111000000110111101;
assign LUT_4[10267] = 32'b11111111111111110001010010110101;
assign LUT_4[10268] = 32'b11111111111111110101101100110101;
assign LUT_4[10269] = 32'b11111111111111101110111000101101;
assign LUT_4[10270] = 32'b11111111111111110101000111011001;
assign LUT_4[10271] = 32'b11111111111111101110010011010001;
assign LUT_4[10272] = 32'b00000000000000000000001001011101;
assign LUT_4[10273] = 32'b11111111111111111001010101010101;
assign LUT_4[10274] = 32'b11111111111111111111100100000001;
assign LUT_4[10275] = 32'b11111111111111111000101111111001;
assign LUT_4[10276] = 32'b11111111111111111101001001111001;
assign LUT_4[10277] = 32'b11111111111111110110010101110001;
assign LUT_4[10278] = 32'b11111111111111111100100100011101;
assign LUT_4[10279] = 32'b11111111111111110101110000010101;
assign LUT_4[10280] = 32'b11111111111111111001010101110010;
assign LUT_4[10281] = 32'b11111111111111110010100001101010;
assign LUT_4[10282] = 32'b11111111111111111000110000010110;
assign LUT_4[10283] = 32'b11111111111111110001111100001110;
assign LUT_4[10284] = 32'b11111111111111110110010110001110;
assign LUT_4[10285] = 32'b11111111111111101111100010000110;
assign LUT_4[10286] = 32'b11111111111111110101110000110010;
assign LUT_4[10287] = 32'b11111111111111101110111100101010;
assign LUT_4[10288] = 32'b11111111111111111101111011001011;
assign LUT_4[10289] = 32'b11111111111111110111000111000011;
assign LUT_4[10290] = 32'b11111111111111111101010101101111;
assign LUT_4[10291] = 32'b11111111111111110110100001100111;
assign LUT_4[10292] = 32'b11111111111111111010111011100111;
assign LUT_4[10293] = 32'b11111111111111110100000111011111;
assign LUT_4[10294] = 32'b11111111111111111010010110001011;
assign LUT_4[10295] = 32'b11111111111111110011100010000011;
assign LUT_4[10296] = 32'b11111111111111110111000111100000;
assign LUT_4[10297] = 32'b11111111111111110000010011011000;
assign LUT_4[10298] = 32'b11111111111111110110100010000100;
assign LUT_4[10299] = 32'b11111111111111101111101101111100;
assign LUT_4[10300] = 32'b11111111111111110100000111111100;
assign LUT_4[10301] = 32'b11111111111111101101010011110100;
assign LUT_4[10302] = 32'b11111111111111110011100010100000;
assign LUT_4[10303] = 32'b11111111111111101100101110011000;
assign LUT_4[10304] = 32'b00000000000000000011000101101010;
assign LUT_4[10305] = 32'b11111111111111111100010001100010;
assign LUT_4[10306] = 32'b00000000000000000010100000001110;
assign LUT_4[10307] = 32'b11111111111111111011101100000110;
assign LUT_4[10308] = 32'b00000000000000000000000110000110;
assign LUT_4[10309] = 32'b11111111111111111001010001111110;
assign LUT_4[10310] = 32'b11111111111111111111100000101010;
assign LUT_4[10311] = 32'b11111111111111111000101100100010;
assign LUT_4[10312] = 32'b11111111111111111100010001111111;
assign LUT_4[10313] = 32'b11111111111111110101011101110111;
assign LUT_4[10314] = 32'b11111111111111111011101100100011;
assign LUT_4[10315] = 32'b11111111111111110100111000011011;
assign LUT_4[10316] = 32'b11111111111111111001010010011011;
assign LUT_4[10317] = 32'b11111111111111110010011110010011;
assign LUT_4[10318] = 32'b11111111111111111000101100111111;
assign LUT_4[10319] = 32'b11111111111111110001111000110111;
assign LUT_4[10320] = 32'b00000000000000000000110111011000;
assign LUT_4[10321] = 32'b11111111111111111010000011010000;
assign LUT_4[10322] = 32'b00000000000000000000010001111100;
assign LUT_4[10323] = 32'b11111111111111111001011101110100;
assign LUT_4[10324] = 32'b11111111111111111101110111110100;
assign LUT_4[10325] = 32'b11111111111111110111000011101100;
assign LUT_4[10326] = 32'b11111111111111111101010010011000;
assign LUT_4[10327] = 32'b11111111111111110110011110010000;
assign LUT_4[10328] = 32'b11111111111111111010000011101101;
assign LUT_4[10329] = 32'b11111111111111110011001111100101;
assign LUT_4[10330] = 32'b11111111111111111001011110010001;
assign LUT_4[10331] = 32'b11111111111111110010101010001001;
assign LUT_4[10332] = 32'b11111111111111110111000100001001;
assign LUT_4[10333] = 32'b11111111111111110000010000000001;
assign LUT_4[10334] = 32'b11111111111111110110011110101101;
assign LUT_4[10335] = 32'b11111111111111101111101010100101;
assign LUT_4[10336] = 32'b00000000000000000001100000110001;
assign LUT_4[10337] = 32'b11111111111111111010101100101001;
assign LUT_4[10338] = 32'b00000000000000000000111011010101;
assign LUT_4[10339] = 32'b11111111111111111010000111001101;
assign LUT_4[10340] = 32'b11111111111111111110100001001101;
assign LUT_4[10341] = 32'b11111111111111110111101101000101;
assign LUT_4[10342] = 32'b11111111111111111101111011110001;
assign LUT_4[10343] = 32'b11111111111111110111000111101001;
assign LUT_4[10344] = 32'b11111111111111111010101101000110;
assign LUT_4[10345] = 32'b11111111111111110011111000111110;
assign LUT_4[10346] = 32'b11111111111111111010000111101010;
assign LUT_4[10347] = 32'b11111111111111110011010011100010;
assign LUT_4[10348] = 32'b11111111111111110111101101100010;
assign LUT_4[10349] = 32'b11111111111111110000111001011010;
assign LUT_4[10350] = 32'b11111111111111110111001000000110;
assign LUT_4[10351] = 32'b11111111111111110000010011111110;
assign LUT_4[10352] = 32'b11111111111111111111010010011111;
assign LUT_4[10353] = 32'b11111111111111111000011110010111;
assign LUT_4[10354] = 32'b11111111111111111110101101000011;
assign LUT_4[10355] = 32'b11111111111111110111111000111011;
assign LUT_4[10356] = 32'b11111111111111111100010010111011;
assign LUT_4[10357] = 32'b11111111111111110101011110110011;
assign LUT_4[10358] = 32'b11111111111111111011101101011111;
assign LUT_4[10359] = 32'b11111111111111110100111001010111;
assign LUT_4[10360] = 32'b11111111111111111000011110110100;
assign LUT_4[10361] = 32'b11111111111111110001101010101100;
assign LUT_4[10362] = 32'b11111111111111110111111001011000;
assign LUT_4[10363] = 32'b11111111111111110001000101010000;
assign LUT_4[10364] = 32'b11111111111111110101011111010000;
assign LUT_4[10365] = 32'b11111111111111101110101011001000;
assign LUT_4[10366] = 32'b11111111111111110100111001110100;
assign LUT_4[10367] = 32'b11111111111111101110000101101100;
assign LUT_4[10368] = 32'b00000000000000000100010100011110;
assign LUT_4[10369] = 32'b11111111111111111101100000010110;
assign LUT_4[10370] = 32'b00000000000000000011101111000010;
assign LUT_4[10371] = 32'b11111111111111111100111010111010;
assign LUT_4[10372] = 32'b00000000000000000001010100111010;
assign LUT_4[10373] = 32'b11111111111111111010100000110010;
assign LUT_4[10374] = 32'b00000000000000000000101111011110;
assign LUT_4[10375] = 32'b11111111111111111001111011010110;
assign LUT_4[10376] = 32'b11111111111111111101100000110011;
assign LUT_4[10377] = 32'b11111111111111110110101100101011;
assign LUT_4[10378] = 32'b11111111111111111100111011010111;
assign LUT_4[10379] = 32'b11111111111111110110000111001111;
assign LUT_4[10380] = 32'b11111111111111111010100001001111;
assign LUT_4[10381] = 32'b11111111111111110011101101000111;
assign LUT_4[10382] = 32'b11111111111111111001111011110011;
assign LUT_4[10383] = 32'b11111111111111110011000111101011;
assign LUT_4[10384] = 32'b00000000000000000010000110001100;
assign LUT_4[10385] = 32'b11111111111111111011010010000100;
assign LUT_4[10386] = 32'b00000000000000000001100000110000;
assign LUT_4[10387] = 32'b11111111111111111010101100101000;
assign LUT_4[10388] = 32'b11111111111111111111000110101000;
assign LUT_4[10389] = 32'b11111111111111111000010010100000;
assign LUT_4[10390] = 32'b11111111111111111110100001001100;
assign LUT_4[10391] = 32'b11111111111111110111101101000100;
assign LUT_4[10392] = 32'b11111111111111111011010010100001;
assign LUT_4[10393] = 32'b11111111111111110100011110011001;
assign LUT_4[10394] = 32'b11111111111111111010101101000101;
assign LUT_4[10395] = 32'b11111111111111110011111000111101;
assign LUT_4[10396] = 32'b11111111111111111000010010111101;
assign LUT_4[10397] = 32'b11111111111111110001011110110101;
assign LUT_4[10398] = 32'b11111111111111110111101101100001;
assign LUT_4[10399] = 32'b11111111111111110000111001011001;
assign LUT_4[10400] = 32'b00000000000000000010101111100101;
assign LUT_4[10401] = 32'b11111111111111111011111011011101;
assign LUT_4[10402] = 32'b00000000000000000010001010001001;
assign LUT_4[10403] = 32'b11111111111111111011010110000001;
assign LUT_4[10404] = 32'b11111111111111111111110000000001;
assign LUT_4[10405] = 32'b11111111111111111000111011111001;
assign LUT_4[10406] = 32'b11111111111111111111001010100101;
assign LUT_4[10407] = 32'b11111111111111111000010110011101;
assign LUT_4[10408] = 32'b11111111111111111011111011111010;
assign LUT_4[10409] = 32'b11111111111111110101000111110010;
assign LUT_4[10410] = 32'b11111111111111111011010110011110;
assign LUT_4[10411] = 32'b11111111111111110100100010010110;
assign LUT_4[10412] = 32'b11111111111111111000111100010110;
assign LUT_4[10413] = 32'b11111111111111110010001000001110;
assign LUT_4[10414] = 32'b11111111111111111000010110111010;
assign LUT_4[10415] = 32'b11111111111111110001100010110010;
assign LUT_4[10416] = 32'b00000000000000000000100001010011;
assign LUT_4[10417] = 32'b11111111111111111001101101001011;
assign LUT_4[10418] = 32'b11111111111111111111111011110111;
assign LUT_4[10419] = 32'b11111111111111111001000111101111;
assign LUT_4[10420] = 32'b11111111111111111101100001101111;
assign LUT_4[10421] = 32'b11111111111111110110101101100111;
assign LUT_4[10422] = 32'b11111111111111111100111100010011;
assign LUT_4[10423] = 32'b11111111111111110110001000001011;
assign LUT_4[10424] = 32'b11111111111111111001101101101000;
assign LUT_4[10425] = 32'b11111111111111110010111001100000;
assign LUT_4[10426] = 32'b11111111111111111001001000001100;
assign LUT_4[10427] = 32'b11111111111111110010010100000100;
assign LUT_4[10428] = 32'b11111111111111110110101110000100;
assign LUT_4[10429] = 32'b11111111111111101111111001111100;
assign LUT_4[10430] = 32'b11111111111111110110001000101000;
assign LUT_4[10431] = 32'b11111111111111101111010100100000;
assign LUT_4[10432] = 32'b00000000000000000101101011110010;
assign LUT_4[10433] = 32'b11111111111111111110110111101010;
assign LUT_4[10434] = 32'b00000000000000000101000110010110;
assign LUT_4[10435] = 32'b11111111111111111110010010001110;
assign LUT_4[10436] = 32'b00000000000000000010101100001110;
assign LUT_4[10437] = 32'b11111111111111111011111000000110;
assign LUT_4[10438] = 32'b00000000000000000010000110110010;
assign LUT_4[10439] = 32'b11111111111111111011010010101010;
assign LUT_4[10440] = 32'b11111111111111111110111000000111;
assign LUT_4[10441] = 32'b11111111111111111000000011111111;
assign LUT_4[10442] = 32'b11111111111111111110010010101011;
assign LUT_4[10443] = 32'b11111111111111110111011110100011;
assign LUT_4[10444] = 32'b11111111111111111011111000100011;
assign LUT_4[10445] = 32'b11111111111111110101000100011011;
assign LUT_4[10446] = 32'b11111111111111111011010011000111;
assign LUT_4[10447] = 32'b11111111111111110100011110111111;
assign LUT_4[10448] = 32'b00000000000000000011011101100000;
assign LUT_4[10449] = 32'b11111111111111111100101001011000;
assign LUT_4[10450] = 32'b00000000000000000010111000000100;
assign LUT_4[10451] = 32'b11111111111111111100000011111100;
assign LUT_4[10452] = 32'b00000000000000000000011101111100;
assign LUT_4[10453] = 32'b11111111111111111001101001110100;
assign LUT_4[10454] = 32'b11111111111111111111111000100000;
assign LUT_4[10455] = 32'b11111111111111111001000100011000;
assign LUT_4[10456] = 32'b11111111111111111100101001110101;
assign LUT_4[10457] = 32'b11111111111111110101110101101101;
assign LUT_4[10458] = 32'b11111111111111111100000100011001;
assign LUT_4[10459] = 32'b11111111111111110101010000010001;
assign LUT_4[10460] = 32'b11111111111111111001101010010001;
assign LUT_4[10461] = 32'b11111111111111110010110110001001;
assign LUT_4[10462] = 32'b11111111111111111001000100110101;
assign LUT_4[10463] = 32'b11111111111111110010010000101101;
assign LUT_4[10464] = 32'b00000000000000000100000110111001;
assign LUT_4[10465] = 32'b11111111111111111101010010110001;
assign LUT_4[10466] = 32'b00000000000000000011100001011101;
assign LUT_4[10467] = 32'b11111111111111111100101101010101;
assign LUT_4[10468] = 32'b00000000000000000001000111010101;
assign LUT_4[10469] = 32'b11111111111111111010010011001101;
assign LUT_4[10470] = 32'b00000000000000000000100001111001;
assign LUT_4[10471] = 32'b11111111111111111001101101110001;
assign LUT_4[10472] = 32'b11111111111111111101010011001110;
assign LUT_4[10473] = 32'b11111111111111110110011111000110;
assign LUT_4[10474] = 32'b11111111111111111100101101110010;
assign LUT_4[10475] = 32'b11111111111111110101111001101010;
assign LUT_4[10476] = 32'b11111111111111111010010011101010;
assign LUT_4[10477] = 32'b11111111111111110011011111100010;
assign LUT_4[10478] = 32'b11111111111111111001101110001110;
assign LUT_4[10479] = 32'b11111111111111110010111010000110;
assign LUT_4[10480] = 32'b00000000000000000001111000100111;
assign LUT_4[10481] = 32'b11111111111111111011000100011111;
assign LUT_4[10482] = 32'b00000000000000000001010011001011;
assign LUT_4[10483] = 32'b11111111111111111010011111000011;
assign LUT_4[10484] = 32'b11111111111111111110111001000011;
assign LUT_4[10485] = 32'b11111111111111111000000100111011;
assign LUT_4[10486] = 32'b11111111111111111110010011100111;
assign LUT_4[10487] = 32'b11111111111111110111011111011111;
assign LUT_4[10488] = 32'b11111111111111111011000100111100;
assign LUT_4[10489] = 32'b11111111111111110100010000110100;
assign LUT_4[10490] = 32'b11111111111111111010011111100000;
assign LUT_4[10491] = 32'b11111111111111110011101011011000;
assign LUT_4[10492] = 32'b11111111111111111000000101011000;
assign LUT_4[10493] = 32'b11111111111111110001010001010000;
assign LUT_4[10494] = 32'b11111111111111110111011111111100;
assign LUT_4[10495] = 32'b11111111111111110000101011110100;
assign LUT_4[10496] = 32'b00000000000000000110101001111001;
assign LUT_4[10497] = 32'b11111111111111111111110101110001;
assign LUT_4[10498] = 32'b00000000000000000110000100011101;
assign LUT_4[10499] = 32'b11111111111111111111010000010101;
assign LUT_4[10500] = 32'b00000000000000000011101010010101;
assign LUT_4[10501] = 32'b11111111111111111100110110001101;
assign LUT_4[10502] = 32'b00000000000000000011000100111001;
assign LUT_4[10503] = 32'b11111111111111111100010000110001;
assign LUT_4[10504] = 32'b11111111111111111111110110001110;
assign LUT_4[10505] = 32'b11111111111111111001000010000110;
assign LUT_4[10506] = 32'b11111111111111111111010000110010;
assign LUT_4[10507] = 32'b11111111111111111000011100101010;
assign LUT_4[10508] = 32'b11111111111111111100110110101010;
assign LUT_4[10509] = 32'b11111111111111110110000010100010;
assign LUT_4[10510] = 32'b11111111111111111100010001001110;
assign LUT_4[10511] = 32'b11111111111111110101011101000110;
assign LUT_4[10512] = 32'b00000000000000000100011011100111;
assign LUT_4[10513] = 32'b11111111111111111101100111011111;
assign LUT_4[10514] = 32'b00000000000000000011110110001011;
assign LUT_4[10515] = 32'b11111111111111111101000010000011;
assign LUT_4[10516] = 32'b00000000000000000001011100000011;
assign LUT_4[10517] = 32'b11111111111111111010100111111011;
assign LUT_4[10518] = 32'b00000000000000000000110110100111;
assign LUT_4[10519] = 32'b11111111111111111010000010011111;
assign LUT_4[10520] = 32'b11111111111111111101100111111100;
assign LUT_4[10521] = 32'b11111111111111110110110011110100;
assign LUT_4[10522] = 32'b11111111111111111101000010100000;
assign LUT_4[10523] = 32'b11111111111111110110001110011000;
assign LUT_4[10524] = 32'b11111111111111111010101000011000;
assign LUT_4[10525] = 32'b11111111111111110011110100010000;
assign LUT_4[10526] = 32'b11111111111111111010000010111100;
assign LUT_4[10527] = 32'b11111111111111110011001110110100;
assign LUT_4[10528] = 32'b00000000000000000101000101000000;
assign LUT_4[10529] = 32'b11111111111111111110010000111000;
assign LUT_4[10530] = 32'b00000000000000000100011111100100;
assign LUT_4[10531] = 32'b11111111111111111101101011011100;
assign LUT_4[10532] = 32'b00000000000000000010000101011100;
assign LUT_4[10533] = 32'b11111111111111111011010001010100;
assign LUT_4[10534] = 32'b00000000000000000001100000000000;
assign LUT_4[10535] = 32'b11111111111111111010101011111000;
assign LUT_4[10536] = 32'b11111111111111111110010001010101;
assign LUT_4[10537] = 32'b11111111111111110111011101001101;
assign LUT_4[10538] = 32'b11111111111111111101101011111001;
assign LUT_4[10539] = 32'b11111111111111110110110111110001;
assign LUT_4[10540] = 32'b11111111111111111011010001110001;
assign LUT_4[10541] = 32'b11111111111111110100011101101001;
assign LUT_4[10542] = 32'b11111111111111111010101100010101;
assign LUT_4[10543] = 32'b11111111111111110011111000001101;
assign LUT_4[10544] = 32'b00000000000000000010110110101110;
assign LUT_4[10545] = 32'b11111111111111111100000010100110;
assign LUT_4[10546] = 32'b00000000000000000010010001010010;
assign LUT_4[10547] = 32'b11111111111111111011011101001010;
assign LUT_4[10548] = 32'b11111111111111111111110111001010;
assign LUT_4[10549] = 32'b11111111111111111001000011000010;
assign LUT_4[10550] = 32'b11111111111111111111010001101110;
assign LUT_4[10551] = 32'b11111111111111111000011101100110;
assign LUT_4[10552] = 32'b11111111111111111100000011000011;
assign LUT_4[10553] = 32'b11111111111111110101001110111011;
assign LUT_4[10554] = 32'b11111111111111111011011101100111;
assign LUT_4[10555] = 32'b11111111111111110100101001011111;
assign LUT_4[10556] = 32'b11111111111111111001000011011111;
assign LUT_4[10557] = 32'b11111111111111110010001111010111;
assign LUT_4[10558] = 32'b11111111111111111000011110000011;
assign LUT_4[10559] = 32'b11111111111111110001101001111011;
assign LUT_4[10560] = 32'b00000000000000001000000001001101;
assign LUT_4[10561] = 32'b00000000000000000001001101000101;
assign LUT_4[10562] = 32'b00000000000000000111011011110001;
assign LUT_4[10563] = 32'b00000000000000000000100111101001;
assign LUT_4[10564] = 32'b00000000000000000101000001101001;
assign LUT_4[10565] = 32'b11111111111111111110001101100001;
assign LUT_4[10566] = 32'b00000000000000000100011100001101;
assign LUT_4[10567] = 32'b11111111111111111101101000000101;
assign LUT_4[10568] = 32'b00000000000000000001001101100010;
assign LUT_4[10569] = 32'b11111111111111111010011001011010;
assign LUT_4[10570] = 32'b00000000000000000000101000000110;
assign LUT_4[10571] = 32'b11111111111111111001110011111110;
assign LUT_4[10572] = 32'b11111111111111111110001101111110;
assign LUT_4[10573] = 32'b11111111111111110111011001110110;
assign LUT_4[10574] = 32'b11111111111111111101101000100010;
assign LUT_4[10575] = 32'b11111111111111110110110100011010;
assign LUT_4[10576] = 32'b00000000000000000101110010111011;
assign LUT_4[10577] = 32'b11111111111111111110111110110011;
assign LUT_4[10578] = 32'b00000000000000000101001101011111;
assign LUT_4[10579] = 32'b11111111111111111110011001010111;
assign LUT_4[10580] = 32'b00000000000000000010110011010111;
assign LUT_4[10581] = 32'b11111111111111111011111111001111;
assign LUT_4[10582] = 32'b00000000000000000010001101111011;
assign LUT_4[10583] = 32'b11111111111111111011011001110011;
assign LUT_4[10584] = 32'b11111111111111111110111111010000;
assign LUT_4[10585] = 32'b11111111111111111000001011001000;
assign LUT_4[10586] = 32'b11111111111111111110011001110100;
assign LUT_4[10587] = 32'b11111111111111110111100101101100;
assign LUT_4[10588] = 32'b11111111111111111011111111101100;
assign LUT_4[10589] = 32'b11111111111111110101001011100100;
assign LUT_4[10590] = 32'b11111111111111111011011010010000;
assign LUT_4[10591] = 32'b11111111111111110100100110001000;
assign LUT_4[10592] = 32'b00000000000000000110011100010100;
assign LUT_4[10593] = 32'b11111111111111111111101000001100;
assign LUT_4[10594] = 32'b00000000000000000101110110111000;
assign LUT_4[10595] = 32'b11111111111111111111000010110000;
assign LUT_4[10596] = 32'b00000000000000000011011100110000;
assign LUT_4[10597] = 32'b11111111111111111100101000101000;
assign LUT_4[10598] = 32'b00000000000000000010110111010100;
assign LUT_4[10599] = 32'b11111111111111111100000011001100;
assign LUT_4[10600] = 32'b11111111111111111111101000101001;
assign LUT_4[10601] = 32'b11111111111111111000110100100001;
assign LUT_4[10602] = 32'b11111111111111111111000011001101;
assign LUT_4[10603] = 32'b11111111111111111000001111000101;
assign LUT_4[10604] = 32'b11111111111111111100101001000101;
assign LUT_4[10605] = 32'b11111111111111110101110100111101;
assign LUT_4[10606] = 32'b11111111111111111100000011101001;
assign LUT_4[10607] = 32'b11111111111111110101001111100001;
assign LUT_4[10608] = 32'b00000000000000000100001110000010;
assign LUT_4[10609] = 32'b11111111111111111101011001111010;
assign LUT_4[10610] = 32'b00000000000000000011101000100110;
assign LUT_4[10611] = 32'b11111111111111111100110100011110;
assign LUT_4[10612] = 32'b00000000000000000001001110011110;
assign LUT_4[10613] = 32'b11111111111111111010011010010110;
assign LUT_4[10614] = 32'b00000000000000000000101001000010;
assign LUT_4[10615] = 32'b11111111111111111001110100111010;
assign LUT_4[10616] = 32'b11111111111111111101011010010111;
assign LUT_4[10617] = 32'b11111111111111110110100110001111;
assign LUT_4[10618] = 32'b11111111111111111100110100111011;
assign LUT_4[10619] = 32'b11111111111111110110000000110011;
assign LUT_4[10620] = 32'b11111111111111111010011010110011;
assign LUT_4[10621] = 32'b11111111111111110011100110101011;
assign LUT_4[10622] = 32'b11111111111111111001110101010111;
assign LUT_4[10623] = 32'b11111111111111110011000001001111;
assign LUT_4[10624] = 32'b00000000000000001001010000000001;
assign LUT_4[10625] = 32'b00000000000000000010011011111001;
assign LUT_4[10626] = 32'b00000000000000001000101010100101;
assign LUT_4[10627] = 32'b00000000000000000001110110011101;
assign LUT_4[10628] = 32'b00000000000000000110010000011101;
assign LUT_4[10629] = 32'b11111111111111111111011100010101;
assign LUT_4[10630] = 32'b00000000000000000101101011000001;
assign LUT_4[10631] = 32'b11111111111111111110110110111001;
assign LUT_4[10632] = 32'b00000000000000000010011100010110;
assign LUT_4[10633] = 32'b11111111111111111011101000001110;
assign LUT_4[10634] = 32'b00000000000000000001110110111010;
assign LUT_4[10635] = 32'b11111111111111111011000010110010;
assign LUT_4[10636] = 32'b11111111111111111111011100110010;
assign LUT_4[10637] = 32'b11111111111111111000101000101010;
assign LUT_4[10638] = 32'b11111111111111111110110111010110;
assign LUT_4[10639] = 32'b11111111111111111000000011001110;
assign LUT_4[10640] = 32'b00000000000000000111000001101111;
assign LUT_4[10641] = 32'b00000000000000000000001101100111;
assign LUT_4[10642] = 32'b00000000000000000110011100010011;
assign LUT_4[10643] = 32'b11111111111111111111101000001011;
assign LUT_4[10644] = 32'b00000000000000000100000010001011;
assign LUT_4[10645] = 32'b11111111111111111101001110000011;
assign LUT_4[10646] = 32'b00000000000000000011011100101111;
assign LUT_4[10647] = 32'b11111111111111111100101000100111;
assign LUT_4[10648] = 32'b00000000000000000000001110000100;
assign LUT_4[10649] = 32'b11111111111111111001011001111100;
assign LUT_4[10650] = 32'b11111111111111111111101000101000;
assign LUT_4[10651] = 32'b11111111111111111000110100100000;
assign LUT_4[10652] = 32'b11111111111111111101001110100000;
assign LUT_4[10653] = 32'b11111111111111110110011010011000;
assign LUT_4[10654] = 32'b11111111111111111100101001000100;
assign LUT_4[10655] = 32'b11111111111111110101110100111100;
assign LUT_4[10656] = 32'b00000000000000000111101011001000;
assign LUT_4[10657] = 32'b00000000000000000000110111000000;
assign LUT_4[10658] = 32'b00000000000000000111000101101100;
assign LUT_4[10659] = 32'b00000000000000000000010001100100;
assign LUT_4[10660] = 32'b00000000000000000100101011100100;
assign LUT_4[10661] = 32'b11111111111111111101110111011100;
assign LUT_4[10662] = 32'b00000000000000000100000110001000;
assign LUT_4[10663] = 32'b11111111111111111101010010000000;
assign LUT_4[10664] = 32'b00000000000000000000110111011101;
assign LUT_4[10665] = 32'b11111111111111111010000011010101;
assign LUT_4[10666] = 32'b00000000000000000000010010000001;
assign LUT_4[10667] = 32'b11111111111111111001011101111001;
assign LUT_4[10668] = 32'b11111111111111111101110111111001;
assign LUT_4[10669] = 32'b11111111111111110111000011110001;
assign LUT_4[10670] = 32'b11111111111111111101010010011101;
assign LUT_4[10671] = 32'b11111111111111110110011110010101;
assign LUT_4[10672] = 32'b00000000000000000101011100110110;
assign LUT_4[10673] = 32'b11111111111111111110101000101110;
assign LUT_4[10674] = 32'b00000000000000000100110111011010;
assign LUT_4[10675] = 32'b11111111111111111110000011010010;
assign LUT_4[10676] = 32'b00000000000000000010011101010010;
assign LUT_4[10677] = 32'b11111111111111111011101001001010;
assign LUT_4[10678] = 32'b00000000000000000001110111110110;
assign LUT_4[10679] = 32'b11111111111111111011000011101110;
assign LUT_4[10680] = 32'b11111111111111111110101001001011;
assign LUT_4[10681] = 32'b11111111111111110111110101000011;
assign LUT_4[10682] = 32'b11111111111111111110000011101111;
assign LUT_4[10683] = 32'b11111111111111110111001111100111;
assign LUT_4[10684] = 32'b11111111111111111011101001100111;
assign LUT_4[10685] = 32'b11111111111111110100110101011111;
assign LUT_4[10686] = 32'b11111111111111111011000100001011;
assign LUT_4[10687] = 32'b11111111111111110100010000000011;
assign LUT_4[10688] = 32'b00000000000000001010100111010101;
assign LUT_4[10689] = 32'b00000000000000000011110011001101;
assign LUT_4[10690] = 32'b00000000000000001010000001111001;
assign LUT_4[10691] = 32'b00000000000000000011001101110001;
assign LUT_4[10692] = 32'b00000000000000000111100111110001;
assign LUT_4[10693] = 32'b00000000000000000000110011101001;
assign LUT_4[10694] = 32'b00000000000000000111000010010101;
assign LUT_4[10695] = 32'b00000000000000000000001110001101;
assign LUT_4[10696] = 32'b00000000000000000011110011101010;
assign LUT_4[10697] = 32'b11111111111111111100111111100010;
assign LUT_4[10698] = 32'b00000000000000000011001110001110;
assign LUT_4[10699] = 32'b11111111111111111100011010000110;
assign LUT_4[10700] = 32'b00000000000000000000110100000110;
assign LUT_4[10701] = 32'b11111111111111111001111111111110;
assign LUT_4[10702] = 32'b00000000000000000000001110101010;
assign LUT_4[10703] = 32'b11111111111111111001011010100010;
assign LUT_4[10704] = 32'b00000000000000001000011001000011;
assign LUT_4[10705] = 32'b00000000000000000001100100111011;
assign LUT_4[10706] = 32'b00000000000000000111110011100111;
assign LUT_4[10707] = 32'b00000000000000000000111111011111;
assign LUT_4[10708] = 32'b00000000000000000101011001011111;
assign LUT_4[10709] = 32'b11111111111111111110100101010111;
assign LUT_4[10710] = 32'b00000000000000000100110100000011;
assign LUT_4[10711] = 32'b11111111111111111101111111111011;
assign LUT_4[10712] = 32'b00000000000000000001100101011000;
assign LUT_4[10713] = 32'b11111111111111111010110001010000;
assign LUT_4[10714] = 32'b00000000000000000000111111111100;
assign LUT_4[10715] = 32'b11111111111111111010001011110100;
assign LUT_4[10716] = 32'b11111111111111111110100101110100;
assign LUT_4[10717] = 32'b11111111111111110111110001101100;
assign LUT_4[10718] = 32'b11111111111111111110000000011000;
assign LUT_4[10719] = 32'b11111111111111110111001100010000;
assign LUT_4[10720] = 32'b00000000000000001001000010011100;
assign LUT_4[10721] = 32'b00000000000000000010001110010100;
assign LUT_4[10722] = 32'b00000000000000001000011101000000;
assign LUT_4[10723] = 32'b00000000000000000001101000111000;
assign LUT_4[10724] = 32'b00000000000000000110000010111000;
assign LUT_4[10725] = 32'b11111111111111111111001110110000;
assign LUT_4[10726] = 32'b00000000000000000101011101011100;
assign LUT_4[10727] = 32'b11111111111111111110101001010100;
assign LUT_4[10728] = 32'b00000000000000000010001110110001;
assign LUT_4[10729] = 32'b11111111111111111011011010101001;
assign LUT_4[10730] = 32'b00000000000000000001101001010101;
assign LUT_4[10731] = 32'b11111111111111111010110101001101;
assign LUT_4[10732] = 32'b11111111111111111111001111001101;
assign LUT_4[10733] = 32'b11111111111111111000011011000101;
assign LUT_4[10734] = 32'b11111111111111111110101001110001;
assign LUT_4[10735] = 32'b11111111111111110111110101101001;
assign LUT_4[10736] = 32'b00000000000000000110110100001010;
assign LUT_4[10737] = 32'b00000000000000000000000000000010;
assign LUT_4[10738] = 32'b00000000000000000110001110101110;
assign LUT_4[10739] = 32'b11111111111111111111011010100110;
assign LUT_4[10740] = 32'b00000000000000000011110100100110;
assign LUT_4[10741] = 32'b11111111111111111101000000011110;
assign LUT_4[10742] = 32'b00000000000000000011001111001010;
assign LUT_4[10743] = 32'b11111111111111111100011011000010;
assign LUT_4[10744] = 32'b00000000000000000000000000011111;
assign LUT_4[10745] = 32'b11111111111111111001001100010111;
assign LUT_4[10746] = 32'b11111111111111111111011011000011;
assign LUT_4[10747] = 32'b11111111111111111000100110111011;
assign LUT_4[10748] = 32'b11111111111111111101000000111011;
assign LUT_4[10749] = 32'b11111111111111110110001100110011;
assign LUT_4[10750] = 32'b11111111111111111100011011011111;
assign LUT_4[10751] = 32'b11111111111111110101100111010111;
assign LUT_4[10752] = 32'b00000000000000000000110010011110;
assign LUT_4[10753] = 32'b11111111111111111001111110010110;
assign LUT_4[10754] = 32'b00000000000000000000001101000010;
assign LUT_4[10755] = 32'b11111111111111111001011000111010;
assign LUT_4[10756] = 32'b11111111111111111101110010111010;
assign LUT_4[10757] = 32'b11111111111111110110111110110010;
assign LUT_4[10758] = 32'b11111111111111111101001101011110;
assign LUT_4[10759] = 32'b11111111111111110110011001010110;
assign LUT_4[10760] = 32'b11111111111111111001111110110011;
assign LUT_4[10761] = 32'b11111111111111110011001010101011;
assign LUT_4[10762] = 32'b11111111111111111001011001010111;
assign LUT_4[10763] = 32'b11111111111111110010100101001111;
assign LUT_4[10764] = 32'b11111111111111110110111111001111;
assign LUT_4[10765] = 32'b11111111111111110000001011000111;
assign LUT_4[10766] = 32'b11111111111111110110011001110011;
assign LUT_4[10767] = 32'b11111111111111101111100101101011;
assign LUT_4[10768] = 32'b11111111111111111110100100001100;
assign LUT_4[10769] = 32'b11111111111111110111110000000100;
assign LUT_4[10770] = 32'b11111111111111111101111110110000;
assign LUT_4[10771] = 32'b11111111111111110111001010101000;
assign LUT_4[10772] = 32'b11111111111111111011100100101000;
assign LUT_4[10773] = 32'b11111111111111110100110000100000;
assign LUT_4[10774] = 32'b11111111111111111010111111001100;
assign LUT_4[10775] = 32'b11111111111111110100001011000100;
assign LUT_4[10776] = 32'b11111111111111110111110000100001;
assign LUT_4[10777] = 32'b11111111111111110000111100011001;
assign LUT_4[10778] = 32'b11111111111111110111001011000101;
assign LUT_4[10779] = 32'b11111111111111110000010110111101;
assign LUT_4[10780] = 32'b11111111111111110100110000111101;
assign LUT_4[10781] = 32'b11111111111111101101111100110101;
assign LUT_4[10782] = 32'b11111111111111110100001011100001;
assign LUT_4[10783] = 32'b11111111111111101101010111011001;
assign LUT_4[10784] = 32'b11111111111111111111001101100101;
assign LUT_4[10785] = 32'b11111111111111111000011001011101;
assign LUT_4[10786] = 32'b11111111111111111110101000001001;
assign LUT_4[10787] = 32'b11111111111111110111110100000001;
assign LUT_4[10788] = 32'b11111111111111111100001110000001;
assign LUT_4[10789] = 32'b11111111111111110101011001111001;
assign LUT_4[10790] = 32'b11111111111111111011101000100101;
assign LUT_4[10791] = 32'b11111111111111110100110100011101;
assign LUT_4[10792] = 32'b11111111111111111000011001111010;
assign LUT_4[10793] = 32'b11111111111111110001100101110010;
assign LUT_4[10794] = 32'b11111111111111110111110100011110;
assign LUT_4[10795] = 32'b11111111111111110001000000010110;
assign LUT_4[10796] = 32'b11111111111111110101011010010110;
assign LUT_4[10797] = 32'b11111111111111101110100110001110;
assign LUT_4[10798] = 32'b11111111111111110100110100111010;
assign LUT_4[10799] = 32'b11111111111111101110000000110010;
assign LUT_4[10800] = 32'b11111111111111111100111111010011;
assign LUT_4[10801] = 32'b11111111111111110110001011001011;
assign LUT_4[10802] = 32'b11111111111111111100011001110111;
assign LUT_4[10803] = 32'b11111111111111110101100101101111;
assign LUT_4[10804] = 32'b11111111111111111001111111101111;
assign LUT_4[10805] = 32'b11111111111111110011001011100111;
assign LUT_4[10806] = 32'b11111111111111111001011010010011;
assign LUT_4[10807] = 32'b11111111111111110010100110001011;
assign LUT_4[10808] = 32'b11111111111111110110001011101000;
assign LUT_4[10809] = 32'b11111111111111101111010111100000;
assign LUT_4[10810] = 32'b11111111111111110101100110001100;
assign LUT_4[10811] = 32'b11111111111111101110110010000100;
assign LUT_4[10812] = 32'b11111111111111110011001100000100;
assign LUT_4[10813] = 32'b11111111111111101100010111111100;
assign LUT_4[10814] = 32'b11111111111111110010100110101000;
assign LUT_4[10815] = 32'b11111111111111101011110010100000;
assign LUT_4[10816] = 32'b00000000000000000010001001110010;
assign LUT_4[10817] = 32'b11111111111111111011010101101010;
assign LUT_4[10818] = 32'b00000000000000000001100100010110;
assign LUT_4[10819] = 32'b11111111111111111010110000001110;
assign LUT_4[10820] = 32'b11111111111111111111001010001110;
assign LUT_4[10821] = 32'b11111111111111111000010110000110;
assign LUT_4[10822] = 32'b11111111111111111110100100110010;
assign LUT_4[10823] = 32'b11111111111111110111110000101010;
assign LUT_4[10824] = 32'b11111111111111111011010110000111;
assign LUT_4[10825] = 32'b11111111111111110100100001111111;
assign LUT_4[10826] = 32'b11111111111111111010110000101011;
assign LUT_4[10827] = 32'b11111111111111110011111100100011;
assign LUT_4[10828] = 32'b11111111111111111000010110100011;
assign LUT_4[10829] = 32'b11111111111111110001100010011011;
assign LUT_4[10830] = 32'b11111111111111110111110001000111;
assign LUT_4[10831] = 32'b11111111111111110000111100111111;
assign LUT_4[10832] = 32'b11111111111111111111111011100000;
assign LUT_4[10833] = 32'b11111111111111111001000111011000;
assign LUT_4[10834] = 32'b11111111111111111111010110000100;
assign LUT_4[10835] = 32'b11111111111111111000100001111100;
assign LUT_4[10836] = 32'b11111111111111111100111011111100;
assign LUT_4[10837] = 32'b11111111111111110110000111110100;
assign LUT_4[10838] = 32'b11111111111111111100010110100000;
assign LUT_4[10839] = 32'b11111111111111110101100010011000;
assign LUT_4[10840] = 32'b11111111111111111001000111110101;
assign LUT_4[10841] = 32'b11111111111111110010010011101101;
assign LUT_4[10842] = 32'b11111111111111111000100010011001;
assign LUT_4[10843] = 32'b11111111111111110001101110010001;
assign LUT_4[10844] = 32'b11111111111111110110001000010001;
assign LUT_4[10845] = 32'b11111111111111101111010100001001;
assign LUT_4[10846] = 32'b11111111111111110101100010110101;
assign LUT_4[10847] = 32'b11111111111111101110101110101101;
assign LUT_4[10848] = 32'b00000000000000000000100100111001;
assign LUT_4[10849] = 32'b11111111111111111001110000110001;
assign LUT_4[10850] = 32'b11111111111111111111111111011101;
assign LUT_4[10851] = 32'b11111111111111111001001011010101;
assign LUT_4[10852] = 32'b11111111111111111101100101010101;
assign LUT_4[10853] = 32'b11111111111111110110110001001101;
assign LUT_4[10854] = 32'b11111111111111111100111111111001;
assign LUT_4[10855] = 32'b11111111111111110110001011110001;
assign LUT_4[10856] = 32'b11111111111111111001110001001110;
assign LUT_4[10857] = 32'b11111111111111110010111101000110;
assign LUT_4[10858] = 32'b11111111111111111001001011110010;
assign LUT_4[10859] = 32'b11111111111111110010010111101010;
assign LUT_4[10860] = 32'b11111111111111110110110001101010;
assign LUT_4[10861] = 32'b11111111111111101111111101100010;
assign LUT_4[10862] = 32'b11111111111111110110001100001110;
assign LUT_4[10863] = 32'b11111111111111101111011000000110;
assign LUT_4[10864] = 32'b11111111111111111110010110100111;
assign LUT_4[10865] = 32'b11111111111111110111100010011111;
assign LUT_4[10866] = 32'b11111111111111111101110001001011;
assign LUT_4[10867] = 32'b11111111111111110110111101000011;
assign LUT_4[10868] = 32'b11111111111111111011010111000011;
assign LUT_4[10869] = 32'b11111111111111110100100010111011;
assign LUT_4[10870] = 32'b11111111111111111010110001100111;
assign LUT_4[10871] = 32'b11111111111111110011111101011111;
assign LUT_4[10872] = 32'b11111111111111110111100010111100;
assign LUT_4[10873] = 32'b11111111111111110000101110110100;
assign LUT_4[10874] = 32'b11111111111111110110111101100000;
assign LUT_4[10875] = 32'b11111111111111110000001001011000;
assign LUT_4[10876] = 32'b11111111111111110100100011011000;
assign LUT_4[10877] = 32'b11111111111111101101101111010000;
assign LUT_4[10878] = 32'b11111111111111110011111101111100;
assign LUT_4[10879] = 32'b11111111111111101101001001110100;
assign LUT_4[10880] = 32'b00000000000000000011011000100110;
assign LUT_4[10881] = 32'b11111111111111111100100100011110;
assign LUT_4[10882] = 32'b00000000000000000010110011001010;
assign LUT_4[10883] = 32'b11111111111111111011111111000010;
assign LUT_4[10884] = 32'b00000000000000000000011001000010;
assign LUT_4[10885] = 32'b11111111111111111001100100111010;
assign LUT_4[10886] = 32'b11111111111111111111110011100110;
assign LUT_4[10887] = 32'b11111111111111111000111111011110;
assign LUT_4[10888] = 32'b11111111111111111100100100111011;
assign LUT_4[10889] = 32'b11111111111111110101110000110011;
assign LUT_4[10890] = 32'b11111111111111111011111111011111;
assign LUT_4[10891] = 32'b11111111111111110101001011010111;
assign LUT_4[10892] = 32'b11111111111111111001100101010111;
assign LUT_4[10893] = 32'b11111111111111110010110001001111;
assign LUT_4[10894] = 32'b11111111111111111000111111111011;
assign LUT_4[10895] = 32'b11111111111111110010001011110011;
assign LUT_4[10896] = 32'b00000000000000000001001010010100;
assign LUT_4[10897] = 32'b11111111111111111010010110001100;
assign LUT_4[10898] = 32'b00000000000000000000100100111000;
assign LUT_4[10899] = 32'b11111111111111111001110000110000;
assign LUT_4[10900] = 32'b11111111111111111110001010110000;
assign LUT_4[10901] = 32'b11111111111111110111010110101000;
assign LUT_4[10902] = 32'b11111111111111111101100101010100;
assign LUT_4[10903] = 32'b11111111111111110110110001001100;
assign LUT_4[10904] = 32'b11111111111111111010010110101001;
assign LUT_4[10905] = 32'b11111111111111110011100010100001;
assign LUT_4[10906] = 32'b11111111111111111001110001001101;
assign LUT_4[10907] = 32'b11111111111111110010111101000101;
assign LUT_4[10908] = 32'b11111111111111110111010111000101;
assign LUT_4[10909] = 32'b11111111111111110000100010111101;
assign LUT_4[10910] = 32'b11111111111111110110110001101001;
assign LUT_4[10911] = 32'b11111111111111101111111101100001;
assign LUT_4[10912] = 32'b00000000000000000001110011101101;
assign LUT_4[10913] = 32'b11111111111111111010111111100101;
assign LUT_4[10914] = 32'b00000000000000000001001110010001;
assign LUT_4[10915] = 32'b11111111111111111010011010001001;
assign LUT_4[10916] = 32'b11111111111111111110110100001001;
assign LUT_4[10917] = 32'b11111111111111111000000000000001;
assign LUT_4[10918] = 32'b11111111111111111110001110101101;
assign LUT_4[10919] = 32'b11111111111111110111011010100101;
assign LUT_4[10920] = 32'b11111111111111111011000000000010;
assign LUT_4[10921] = 32'b11111111111111110100001011111010;
assign LUT_4[10922] = 32'b11111111111111111010011010100110;
assign LUT_4[10923] = 32'b11111111111111110011100110011110;
assign LUT_4[10924] = 32'b11111111111111111000000000011110;
assign LUT_4[10925] = 32'b11111111111111110001001100010110;
assign LUT_4[10926] = 32'b11111111111111110111011011000010;
assign LUT_4[10927] = 32'b11111111111111110000100110111010;
assign LUT_4[10928] = 32'b11111111111111111111100101011011;
assign LUT_4[10929] = 32'b11111111111111111000110001010011;
assign LUT_4[10930] = 32'b11111111111111111110111111111111;
assign LUT_4[10931] = 32'b11111111111111111000001011110111;
assign LUT_4[10932] = 32'b11111111111111111100100101110111;
assign LUT_4[10933] = 32'b11111111111111110101110001101111;
assign LUT_4[10934] = 32'b11111111111111111100000000011011;
assign LUT_4[10935] = 32'b11111111111111110101001100010011;
assign LUT_4[10936] = 32'b11111111111111111000110001110000;
assign LUT_4[10937] = 32'b11111111111111110001111101101000;
assign LUT_4[10938] = 32'b11111111111111111000001100010100;
assign LUT_4[10939] = 32'b11111111111111110001011000001100;
assign LUT_4[10940] = 32'b11111111111111110101110010001100;
assign LUT_4[10941] = 32'b11111111111111101110111110000100;
assign LUT_4[10942] = 32'b11111111111111110101001100110000;
assign LUT_4[10943] = 32'b11111111111111101110011000101000;
assign LUT_4[10944] = 32'b00000000000000000100101111111010;
assign LUT_4[10945] = 32'b11111111111111111101111011110010;
assign LUT_4[10946] = 32'b00000000000000000100001010011110;
assign LUT_4[10947] = 32'b11111111111111111101010110010110;
assign LUT_4[10948] = 32'b00000000000000000001110000010110;
assign LUT_4[10949] = 32'b11111111111111111010111100001110;
assign LUT_4[10950] = 32'b00000000000000000001001010111010;
assign LUT_4[10951] = 32'b11111111111111111010010110110010;
assign LUT_4[10952] = 32'b11111111111111111101111100001111;
assign LUT_4[10953] = 32'b11111111111111110111001000000111;
assign LUT_4[10954] = 32'b11111111111111111101010110110011;
assign LUT_4[10955] = 32'b11111111111111110110100010101011;
assign LUT_4[10956] = 32'b11111111111111111010111100101011;
assign LUT_4[10957] = 32'b11111111111111110100001000100011;
assign LUT_4[10958] = 32'b11111111111111111010010111001111;
assign LUT_4[10959] = 32'b11111111111111110011100011000111;
assign LUT_4[10960] = 32'b00000000000000000010100001101000;
assign LUT_4[10961] = 32'b11111111111111111011101101100000;
assign LUT_4[10962] = 32'b00000000000000000001111100001100;
assign LUT_4[10963] = 32'b11111111111111111011001000000100;
assign LUT_4[10964] = 32'b11111111111111111111100010000100;
assign LUT_4[10965] = 32'b11111111111111111000101101111100;
assign LUT_4[10966] = 32'b11111111111111111110111100101000;
assign LUT_4[10967] = 32'b11111111111111111000001000100000;
assign LUT_4[10968] = 32'b11111111111111111011101101111101;
assign LUT_4[10969] = 32'b11111111111111110100111001110101;
assign LUT_4[10970] = 32'b11111111111111111011001000100001;
assign LUT_4[10971] = 32'b11111111111111110100010100011001;
assign LUT_4[10972] = 32'b11111111111111111000101110011001;
assign LUT_4[10973] = 32'b11111111111111110001111010010001;
assign LUT_4[10974] = 32'b11111111111111111000001000111101;
assign LUT_4[10975] = 32'b11111111111111110001010100110101;
assign LUT_4[10976] = 32'b00000000000000000011001011000001;
assign LUT_4[10977] = 32'b11111111111111111100010110111001;
assign LUT_4[10978] = 32'b00000000000000000010100101100101;
assign LUT_4[10979] = 32'b11111111111111111011110001011101;
assign LUT_4[10980] = 32'b00000000000000000000001011011101;
assign LUT_4[10981] = 32'b11111111111111111001010111010101;
assign LUT_4[10982] = 32'b11111111111111111111100110000001;
assign LUT_4[10983] = 32'b11111111111111111000110001111001;
assign LUT_4[10984] = 32'b11111111111111111100010111010110;
assign LUT_4[10985] = 32'b11111111111111110101100011001110;
assign LUT_4[10986] = 32'b11111111111111111011110001111010;
assign LUT_4[10987] = 32'b11111111111111110100111101110010;
assign LUT_4[10988] = 32'b11111111111111111001010111110010;
assign LUT_4[10989] = 32'b11111111111111110010100011101010;
assign LUT_4[10990] = 32'b11111111111111111000110010010110;
assign LUT_4[10991] = 32'b11111111111111110001111110001110;
assign LUT_4[10992] = 32'b00000000000000000000111100101111;
assign LUT_4[10993] = 32'b11111111111111111010001000100111;
assign LUT_4[10994] = 32'b00000000000000000000010111010011;
assign LUT_4[10995] = 32'b11111111111111111001100011001011;
assign LUT_4[10996] = 32'b11111111111111111101111101001011;
assign LUT_4[10997] = 32'b11111111111111110111001001000011;
assign LUT_4[10998] = 32'b11111111111111111101010111101111;
assign LUT_4[10999] = 32'b11111111111111110110100011100111;
assign LUT_4[11000] = 32'b11111111111111111010001001000100;
assign LUT_4[11001] = 32'b11111111111111110011010100111100;
assign LUT_4[11002] = 32'b11111111111111111001100011101000;
assign LUT_4[11003] = 32'b11111111111111110010101111100000;
assign LUT_4[11004] = 32'b11111111111111110111001001100000;
assign LUT_4[11005] = 32'b11111111111111110000010101011000;
assign LUT_4[11006] = 32'b11111111111111110110100100000100;
assign LUT_4[11007] = 32'b11111111111111101111101111111100;
assign LUT_4[11008] = 32'b00000000000000000101101110000001;
assign LUT_4[11009] = 32'b11111111111111111110111001111001;
assign LUT_4[11010] = 32'b00000000000000000101001000100101;
assign LUT_4[11011] = 32'b11111111111111111110010100011101;
assign LUT_4[11012] = 32'b00000000000000000010101110011101;
assign LUT_4[11013] = 32'b11111111111111111011111010010101;
assign LUT_4[11014] = 32'b00000000000000000010001001000001;
assign LUT_4[11015] = 32'b11111111111111111011010100111001;
assign LUT_4[11016] = 32'b11111111111111111110111010010110;
assign LUT_4[11017] = 32'b11111111111111111000000110001110;
assign LUT_4[11018] = 32'b11111111111111111110010100111010;
assign LUT_4[11019] = 32'b11111111111111110111100000110010;
assign LUT_4[11020] = 32'b11111111111111111011111010110010;
assign LUT_4[11021] = 32'b11111111111111110101000110101010;
assign LUT_4[11022] = 32'b11111111111111111011010101010110;
assign LUT_4[11023] = 32'b11111111111111110100100001001110;
assign LUT_4[11024] = 32'b00000000000000000011011111101111;
assign LUT_4[11025] = 32'b11111111111111111100101011100111;
assign LUT_4[11026] = 32'b00000000000000000010111010010011;
assign LUT_4[11027] = 32'b11111111111111111100000110001011;
assign LUT_4[11028] = 32'b00000000000000000000100000001011;
assign LUT_4[11029] = 32'b11111111111111111001101100000011;
assign LUT_4[11030] = 32'b11111111111111111111111010101111;
assign LUT_4[11031] = 32'b11111111111111111001000110100111;
assign LUT_4[11032] = 32'b11111111111111111100101100000100;
assign LUT_4[11033] = 32'b11111111111111110101110111111100;
assign LUT_4[11034] = 32'b11111111111111111100000110101000;
assign LUT_4[11035] = 32'b11111111111111110101010010100000;
assign LUT_4[11036] = 32'b11111111111111111001101100100000;
assign LUT_4[11037] = 32'b11111111111111110010111000011000;
assign LUT_4[11038] = 32'b11111111111111111001000111000100;
assign LUT_4[11039] = 32'b11111111111111110010010010111100;
assign LUT_4[11040] = 32'b00000000000000000100001001001000;
assign LUT_4[11041] = 32'b11111111111111111101010101000000;
assign LUT_4[11042] = 32'b00000000000000000011100011101100;
assign LUT_4[11043] = 32'b11111111111111111100101111100100;
assign LUT_4[11044] = 32'b00000000000000000001001001100100;
assign LUT_4[11045] = 32'b11111111111111111010010101011100;
assign LUT_4[11046] = 32'b00000000000000000000100100001000;
assign LUT_4[11047] = 32'b11111111111111111001110000000000;
assign LUT_4[11048] = 32'b11111111111111111101010101011101;
assign LUT_4[11049] = 32'b11111111111111110110100001010101;
assign LUT_4[11050] = 32'b11111111111111111100110000000001;
assign LUT_4[11051] = 32'b11111111111111110101111011111001;
assign LUT_4[11052] = 32'b11111111111111111010010101111001;
assign LUT_4[11053] = 32'b11111111111111110011100001110001;
assign LUT_4[11054] = 32'b11111111111111111001110000011101;
assign LUT_4[11055] = 32'b11111111111111110010111100010101;
assign LUT_4[11056] = 32'b00000000000000000001111010110110;
assign LUT_4[11057] = 32'b11111111111111111011000110101110;
assign LUT_4[11058] = 32'b00000000000000000001010101011010;
assign LUT_4[11059] = 32'b11111111111111111010100001010010;
assign LUT_4[11060] = 32'b11111111111111111110111011010010;
assign LUT_4[11061] = 32'b11111111111111111000000111001010;
assign LUT_4[11062] = 32'b11111111111111111110010101110110;
assign LUT_4[11063] = 32'b11111111111111110111100001101110;
assign LUT_4[11064] = 32'b11111111111111111011000111001011;
assign LUT_4[11065] = 32'b11111111111111110100010011000011;
assign LUT_4[11066] = 32'b11111111111111111010100001101111;
assign LUT_4[11067] = 32'b11111111111111110011101101100111;
assign LUT_4[11068] = 32'b11111111111111111000000111100111;
assign LUT_4[11069] = 32'b11111111111111110001010011011111;
assign LUT_4[11070] = 32'b11111111111111110111100010001011;
assign LUT_4[11071] = 32'b11111111111111110000101110000011;
assign LUT_4[11072] = 32'b00000000000000000111000101010101;
assign LUT_4[11073] = 32'b00000000000000000000010001001101;
assign LUT_4[11074] = 32'b00000000000000000110011111111001;
assign LUT_4[11075] = 32'b11111111111111111111101011110001;
assign LUT_4[11076] = 32'b00000000000000000100000101110001;
assign LUT_4[11077] = 32'b11111111111111111101010001101001;
assign LUT_4[11078] = 32'b00000000000000000011100000010101;
assign LUT_4[11079] = 32'b11111111111111111100101100001101;
assign LUT_4[11080] = 32'b00000000000000000000010001101010;
assign LUT_4[11081] = 32'b11111111111111111001011101100010;
assign LUT_4[11082] = 32'b11111111111111111111101100001110;
assign LUT_4[11083] = 32'b11111111111111111000111000000110;
assign LUT_4[11084] = 32'b11111111111111111101010010000110;
assign LUT_4[11085] = 32'b11111111111111110110011101111110;
assign LUT_4[11086] = 32'b11111111111111111100101100101010;
assign LUT_4[11087] = 32'b11111111111111110101111000100010;
assign LUT_4[11088] = 32'b00000000000000000100110111000011;
assign LUT_4[11089] = 32'b11111111111111111110000010111011;
assign LUT_4[11090] = 32'b00000000000000000100010001100111;
assign LUT_4[11091] = 32'b11111111111111111101011101011111;
assign LUT_4[11092] = 32'b00000000000000000001110111011111;
assign LUT_4[11093] = 32'b11111111111111111011000011010111;
assign LUT_4[11094] = 32'b00000000000000000001010010000011;
assign LUT_4[11095] = 32'b11111111111111111010011101111011;
assign LUT_4[11096] = 32'b11111111111111111110000011011000;
assign LUT_4[11097] = 32'b11111111111111110111001111010000;
assign LUT_4[11098] = 32'b11111111111111111101011101111100;
assign LUT_4[11099] = 32'b11111111111111110110101001110100;
assign LUT_4[11100] = 32'b11111111111111111011000011110100;
assign LUT_4[11101] = 32'b11111111111111110100001111101100;
assign LUT_4[11102] = 32'b11111111111111111010011110011000;
assign LUT_4[11103] = 32'b11111111111111110011101010010000;
assign LUT_4[11104] = 32'b00000000000000000101100000011100;
assign LUT_4[11105] = 32'b11111111111111111110101100010100;
assign LUT_4[11106] = 32'b00000000000000000100111011000000;
assign LUT_4[11107] = 32'b11111111111111111110000110111000;
assign LUT_4[11108] = 32'b00000000000000000010100000111000;
assign LUT_4[11109] = 32'b11111111111111111011101100110000;
assign LUT_4[11110] = 32'b00000000000000000001111011011100;
assign LUT_4[11111] = 32'b11111111111111111011000111010100;
assign LUT_4[11112] = 32'b11111111111111111110101100110001;
assign LUT_4[11113] = 32'b11111111111111110111111000101001;
assign LUT_4[11114] = 32'b11111111111111111110000111010101;
assign LUT_4[11115] = 32'b11111111111111110111010011001101;
assign LUT_4[11116] = 32'b11111111111111111011101101001101;
assign LUT_4[11117] = 32'b11111111111111110100111001000101;
assign LUT_4[11118] = 32'b11111111111111111011000111110001;
assign LUT_4[11119] = 32'b11111111111111110100010011101001;
assign LUT_4[11120] = 32'b00000000000000000011010010001010;
assign LUT_4[11121] = 32'b11111111111111111100011110000010;
assign LUT_4[11122] = 32'b00000000000000000010101100101110;
assign LUT_4[11123] = 32'b11111111111111111011111000100110;
assign LUT_4[11124] = 32'b00000000000000000000010010100110;
assign LUT_4[11125] = 32'b11111111111111111001011110011110;
assign LUT_4[11126] = 32'b11111111111111111111101101001010;
assign LUT_4[11127] = 32'b11111111111111111000111001000010;
assign LUT_4[11128] = 32'b11111111111111111100011110011111;
assign LUT_4[11129] = 32'b11111111111111110101101010010111;
assign LUT_4[11130] = 32'b11111111111111111011111001000011;
assign LUT_4[11131] = 32'b11111111111111110101000100111011;
assign LUT_4[11132] = 32'b11111111111111111001011110111011;
assign LUT_4[11133] = 32'b11111111111111110010101010110011;
assign LUT_4[11134] = 32'b11111111111111111000111001011111;
assign LUT_4[11135] = 32'b11111111111111110010000101010111;
assign LUT_4[11136] = 32'b00000000000000001000010100001001;
assign LUT_4[11137] = 32'b00000000000000000001100000000001;
assign LUT_4[11138] = 32'b00000000000000000111101110101101;
assign LUT_4[11139] = 32'b00000000000000000000111010100101;
assign LUT_4[11140] = 32'b00000000000000000101010100100101;
assign LUT_4[11141] = 32'b11111111111111111110100000011101;
assign LUT_4[11142] = 32'b00000000000000000100101111001001;
assign LUT_4[11143] = 32'b11111111111111111101111011000001;
assign LUT_4[11144] = 32'b00000000000000000001100000011110;
assign LUT_4[11145] = 32'b11111111111111111010101100010110;
assign LUT_4[11146] = 32'b00000000000000000000111011000010;
assign LUT_4[11147] = 32'b11111111111111111010000110111010;
assign LUT_4[11148] = 32'b11111111111111111110100000111010;
assign LUT_4[11149] = 32'b11111111111111110111101100110010;
assign LUT_4[11150] = 32'b11111111111111111101111011011110;
assign LUT_4[11151] = 32'b11111111111111110111000111010110;
assign LUT_4[11152] = 32'b00000000000000000110000101110111;
assign LUT_4[11153] = 32'b11111111111111111111010001101111;
assign LUT_4[11154] = 32'b00000000000000000101100000011011;
assign LUT_4[11155] = 32'b11111111111111111110101100010011;
assign LUT_4[11156] = 32'b00000000000000000011000110010011;
assign LUT_4[11157] = 32'b11111111111111111100010010001011;
assign LUT_4[11158] = 32'b00000000000000000010100000110111;
assign LUT_4[11159] = 32'b11111111111111111011101100101111;
assign LUT_4[11160] = 32'b11111111111111111111010010001100;
assign LUT_4[11161] = 32'b11111111111111111000011110000100;
assign LUT_4[11162] = 32'b11111111111111111110101100110000;
assign LUT_4[11163] = 32'b11111111111111110111111000101000;
assign LUT_4[11164] = 32'b11111111111111111100010010101000;
assign LUT_4[11165] = 32'b11111111111111110101011110100000;
assign LUT_4[11166] = 32'b11111111111111111011101101001100;
assign LUT_4[11167] = 32'b11111111111111110100111001000100;
assign LUT_4[11168] = 32'b00000000000000000110101111010000;
assign LUT_4[11169] = 32'b11111111111111111111111011001000;
assign LUT_4[11170] = 32'b00000000000000000110001001110100;
assign LUT_4[11171] = 32'b11111111111111111111010101101100;
assign LUT_4[11172] = 32'b00000000000000000011101111101100;
assign LUT_4[11173] = 32'b11111111111111111100111011100100;
assign LUT_4[11174] = 32'b00000000000000000011001010010000;
assign LUT_4[11175] = 32'b11111111111111111100010110001000;
assign LUT_4[11176] = 32'b11111111111111111111111011100101;
assign LUT_4[11177] = 32'b11111111111111111001000111011101;
assign LUT_4[11178] = 32'b11111111111111111111010110001001;
assign LUT_4[11179] = 32'b11111111111111111000100010000001;
assign LUT_4[11180] = 32'b11111111111111111100111100000001;
assign LUT_4[11181] = 32'b11111111111111110110000111111001;
assign LUT_4[11182] = 32'b11111111111111111100010110100101;
assign LUT_4[11183] = 32'b11111111111111110101100010011101;
assign LUT_4[11184] = 32'b00000000000000000100100000111110;
assign LUT_4[11185] = 32'b11111111111111111101101100110110;
assign LUT_4[11186] = 32'b00000000000000000011111011100010;
assign LUT_4[11187] = 32'b11111111111111111101000111011010;
assign LUT_4[11188] = 32'b00000000000000000001100001011010;
assign LUT_4[11189] = 32'b11111111111111111010101101010010;
assign LUT_4[11190] = 32'b00000000000000000000111011111110;
assign LUT_4[11191] = 32'b11111111111111111010000111110110;
assign LUT_4[11192] = 32'b11111111111111111101101101010011;
assign LUT_4[11193] = 32'b11111111111111110110111001001011;
assign LUT_4[11194] = 32'b11111111111111111101000111110111;
assign LUT_4[11195] = 32'b11111111111111110110010011101111;
assign LUT_4[11196] = 32'b11111111111111111010101101101111;
assign LUT_4[11197] = 32'b11111111111111110011111001100111;
assign LUT_4[11198] = 32'b11111111111111111010001000010011;
assign LUT_4[11199] = 32'b11111111111111110011010100001011;
assign LUT_4[11200] = 32'b00000000000000001001101011011101;
assign LUT_4[11201] = 32'b00000000000000000010110111010101;
assign LUT_4[11202] = 32'b00000000000000001001000110000001;
assign LUT_4[11203] = 32'b00000000000000000010010001111001;
assign LUT_4[11204] = 32'b00000000000000000110101011111001;
assign LUT_4[11205] = 32'b11111111111111111111110111110001;
assign LUT_4[11206] = 32'b00000000000000000110000110011101;
assign LUT_4[11207] = 32'b11111111111111111111010010010101;
assign LUT_4[11208] = 32'b00000000000000000010110111110010;
assign LUT_4[11209] = 32'b11111111111111111100000011101010;
assign LUT_4[11210] = 32'b00000000000000000010010010010110;
assign LUT_4[11211] = 32'b11111111111111111011011110001110;
assign LUT_4[11212] = 32'b11111111111111111111111000001110;
assign LUT_4[11213] = 32'b11111111111111111001000100000110;
assign LUT_4[11214] = 32'b11111111111111111111010010110010;
assign LUT_4[11215] = 32'b11111111111111111000011110101010;
assign LUT_4[11216] = 32'b00000000000000000111011101001011;
assign LUT_4[11217] = 32'b00000000000000000000101001000011;
assign LUT_4[11218] = 32'b00000000000000000110110111101111;
assign LUT_4[11219] = 32'b00000000000000000000000011100111;
assign LUT_4[11220] = 32'b00000000000000000100011101100111;
assign LUT_4[11221] = 32'b11111111111111111101101001011111;
assign LUT_4[11222] = 32'b00000000000000000011111000001011;
assign LUT_4[11223] = 32'b11111111111111111101000100000011;
assign LUT_4[11224] = 32'b00000000000000000000101001100000;
assign LUT_4[11225] = 32'b11111111111111111001110101011000;
assign LUT_4[11226] = 32'b00000000000000000000000100000100;
assign LUT_4[11227] = 32'b11111111111111111001001111111100;
assign LUT_4[11228] = 32'b11111111111111111101101001111100;
assign LUT_4[11229] = 32'b11111111111111110110110101110100;
assign LUT_4[11230] = 32'b11111111111111111101000100100000;
assign LUT_4[11231] = 32'b11111111111111110110010000011000;
assign LUT_4[11232] = 32'b00000000000000001000000110100100;
assign LUT_4[11233] = 32'b00000000000000000001010010011100;
assign LUT_4[11234] = 32'b00000000000000000111100001001000;
assign LUT_4[11235] = 32'b00000000000000000000101101000000;
assign LUT_4[11236] = 32'b00000000000000000101000111000000;
assign LUT_4[11237] = 32'b11111111111111111110010010111000;
assign LUT_4[11238] = 32'b00000000000000000100100001100100;
assign LUT_4[11239] = 32'b11111111111111111101101101011100;
assign LUT_4[11240] = 32'b00000000000000000001010010111001;
assign LUT_4[11241] = 32'b11111111111111111010011110110001;
assign LUT_4[11242] = 32'b00000000000000000000101101011101;
assign LUT_4[11243] = 32'b11111111111111111001111001010101;
assign LUT_4[11244] = 32'b11111111111111111110010011010101;
assign LUT_4[11245] = 32'b11111111111111110111011111001101;
assign LUT_4[11246] = 32'b11111111111111111101101101111001;
assign LUT_4[11247] = 32'b11111111111111110110111001110001;
assign LUT_4[11248] = 32'b00000000000000000101111000010010;
assign LUT_4[11249] = 32'b11111111111111111111000100001010;
assign LUT_4[11250] = 32'b00000000000000000101010010110110;
assign LUT_4[11251] = 32'b11111111111111111110011110101110;
assign LUT_4[11252] = 32'b00000000000000000010111000101110;
assign LUT_4[11253] = 32'b11111111111111111100000100100110;
assign LUT_4[11254] = 32'b00000000000000000010010011010010;
assign LUT_4[11255] = 32'b11111111111111111011011111001010;
assign LUT_4[11256] = 32'b11111111111111111111000100100111;
assign LUT_4[11257] = 32'b11111111111111111000010000011111;
assign LUT_4[11258] = 32'b11111111111111111110011111001011;
assign LUT_4[11259] = 32'b11111111111111110111101011000011;
assign LUT_4[11260] = 32'b11111111111111111100000101000011;
assign LUT_4[11261] = 32'b11111111111111110101010000111011;
assign LUT_4[11262] = 32'b11111111111111111011011111100111;
assign LUT_4[11263] = 32'b11111111111111110100101011011111;
assign LUT_4[11264] = 32'b00000000000000000011011000110101;
assign LUT_4[11265] = 32'b11111111111111111100100100101101;
assign LUT_4[11266] = 32'b00000000000000000010110011011001;
assign LUT_4[11267] = 32'b11111111111111111011111111010001;
assign LUT_4[11268] = 32'b00000000000000000000011001010001;
assign LUT_4[11269] = 32'b11111111111111111001100101001001;
assign LUT_4[11270] = 32'b11111111111111111111110011110101;
assign LUT_4[11271] = 32'b11111111111111111000111111101101;
assign LUT_4[11272] = 32'b11111111111111111100100101001010;
assign LUT_4[11273] = 32'b11111111111111110101110001000010;
assign LUT_4[11274] = 32'b11111111111111111011111111101110;
assign LUT_4[11275] = 32'b11111111111111110101001011100110;
assign LUT_4[11276] = 32'b11111111111111111001100101100110;
assign LUT_4[11277] = 32'b11111111111111110010110001011110;
assign LUT_4[11278] = 32'b11111111111111111001000000001010;
assign LUT_4[11279] = 32'b11111111111111110010001100000010;
assign LUT_4[11280] = 32'b00000000000000000001001010100011;
assign LUT_4[11281] = 32'b11111111111111111010010110011011;
assign LUT_4[11282] = 32'b00000000000000000000100101000111;
assign LUT_4[11283] = 32'b11111111111111111001110000111111;
assign LUT_4[11284] = 32'b11111111111111111110001010111111;
assign LUT_4[11285] = 32'b11111111111111110111010110110111;
assign LUT_4[11286] = 32'b11111111111111111101100101100011;
assign LUT_4[11287] = 32'b11111111111111110110110001011011;
assign LUT_4[11288] = 32'b11111111111111111010010110111000;
assign LUT_4[11289] = 32'b11111111111111110011100010110000;
assign LUT_4[11290] = 32'b11111111111111111001110001011100;
assign LUT_4[11291] = 32'b11111111111111110010111101010100;
assign LUT_4[11292] = 32'b11111111111111110111010111010100;
assign LUT_4[11293] = 32'b11111111111111110000100011001100;
assign LUT_4[11294] = 32'b11111111111111110110110001111000;
assign LUT_4[11295] = 32'b11111111111111101111111101110000;
assign LUT_4[11296] = 32'b00000000000000000001110011111100;
assign LUT_4[11297] = 32'b11111111111111111010111111110100;
assign LUT_4[11298] = 32'b00000000000000000001001110100000;
assign LUT_4[11299] = 32'b11111111111111111010011010011000;
assign LUT_4[11300] = 32'b11111111111111111110110100011000;
assign LUT_4[11301] = 32'b11111111111111111000000000010000;
assign LUT_4[11302] = 32'b11111111111111111110001110111100;
assign LUT_4[11303] = 32'b11111111111111110111011010110100;
assign LUT_4[11304] = 32'b11111111111111111011000000010001;
assign LUT_4[11305] = 32'b11111111111111110100001100001001;
assign LUT_4[11306] = 32'b11111111111111111010011010110101;
assign LUT_4[11307] = 32'b11111111111111110011100110101101;
assign LUT_4[11308] = 32'b11111111111111111000000000101101;
assign LUT_4[11309] = 32'b11111111111111110001001100100101;
assign LUT_4[11310] = 32'b11111111111111110111011011010001;
assign LUT_4[11311] = 32'b11111111111111110000100111001001;
assign LUT_4[11312] = 32'b11111111111111111111100101101010;
assign LUT_4[11313] = 32'b11111111111111111000110001100010;
assign LUT_4[11314] = 32'b11111111111111111111000000001110;
assign LUT_4[11315] = 32'b11111111111111111000001100000110;
assign LUT_4[11316] = 32'b11111111111111111100100110000110;
assign LUT_4[11317] = 32'b11111111111111110101110001111110;
assign LUT_4[11318] = 32'b11111111111111111100000000101010;
assign LUT_4[11319] = 32'b11111111111111110101001100100010;
assign LUT_4[11320] = 32'b11111111111111111000110001111111;
assign LUT_4[11321] = 32'b11111111111111110001111101110111;
assign LUT_4[11322] = 32'b11111111111111111000001100100011;
assign LUT_4[11323] = 32'b11111111111111110001011000011011;
assign LUT_4[11324] = 32'b11111111111111110101110010011011;
assign LUT_4[11325] = 32'b11111111111111101110111110010011;
assign LUT_4[11326] = 32'b11111111111111110101001100111111;
assign LUT_4[11327] = 32'b11111111111111101110011000110111;
assign LUT_4[11328] = 32'b00000000000000000100110000001001;
assign LUT_4[11329] = 32'b11111111111111111101111100000001;
assign LUT_4[11330] = 32'b00000000000000000100001010101101;
assign LUT_4[11331] = 32'b11111111111111111101010110100101;
assign LUT_4[11332] = 32'b00000000000000000001110000100101;
assign LUT_4[11333] = 32'b11111111111111111010111100011101;
assign LUT_4[11334] = 32'b00000000000000000001001011001001;
assign LUT_4[11335] = 32'b11111111111111111010010111000001;
assign LUT_4[11336] = 32'b11111111111111111101111100011110;
assign LUT_4[11337] = 32'b11111111111111110111001000010110;
assign LUT_4[11338] = 32'b11111111111111111101010111000010;
assign LUT_4[11339] = 32'b11111111111111110110100010111010;
assign LUT_4[11340] = 32'b11111111111111111010111100111010;
assign LUT_4[11341] = 32'b11111111111111110100001000110010;
assign LUT_4[11342] = 32'b11111111111111111010010111011110;
assign LUT_4[11343] = 32'b11111111111111110011100011010110;
assign LUT_4[11344] = 32'b00000000000000000010100001110111;
assign LUT_4[11345] = 32'b11111111111111111011101101101111;
assign LUT_4[11346] = 32'b00000000000000000001111100011011;
assign LUT_4[11347] = 32'b11111111111111111011001000010011;
assign LUT_4[11348] = 32'b11111111111111111111100010010011;
assign LUT_4[11349] = 32'b11111111111111111000101110001011;
assign LUT_4[11350] = 32'b11111111111111111110111100110111;
assign LUT_4[11351] = 32'b11111111111111111000001000101111;
assign LUT_4[11352] = 32'b11111111111111111011101110001100;
assign LUT_4[11353] = 32'b11111111111111110100111010000100;
assign LUT_4[11354] = 32'b11111111111111111011001000110000;
assign LUT_4[11355] = 32'b11111111111111110100010100101000;
assign LUT_4[11356] = 32'b11111111111111111000101110101000;
assign LUT_4[11357] = 32'b11111111111111110001111010100000;
assign LUT_4[11358] = 32'b11111111111111111000001001001100;
assign LUT_4[11359] = 32'b11111111111111110001010101000100;
assign LUT_4[11360] = 32'b00000000000000000011001011010000;
assign LUT_4[11361] = 32'b11111111111111111100010111001000;
assign LUT_4[11362] = 32'b00000000000000000010100101110100;
assign LUT_4[11363] = 32'b11111111111111111011110001101100;
assign LUT_4[11364] = 32'b00000000000000000000001011101100;
assign LUT_4[11365] = 32'b11111111111111111001010111100100;
assign LUT_4[11366] = 32'b11111111111111111111100110010000;
assign LUT_4[11367] = 32'b11111111111111111000110010001000;
assign LUT_4[11368] = 32'b11111111111111111100010111100101;
assign LUT_4[11369] = 32'b11111111111111110101100011011101;
assign LUT_4[11370] = 32'b11111111111111111011110010001001;
assign LUT_4[11371] = 32'b11111111111111110100111110000001;
assign LUT_4[11372] = 32'b11111111111111111001011000000001;
assign LUT_4[11373] = 32'b11111111111111110010100011111001;
assign LUT_4[11374] = 32'b11111111111111111000110010100101;
assign LUT_4[11375] = 32'b11111111111111110001111110011101;
assign LUT_4[11376] = 32'b00000000000000000000111100111110;
assign LUT_4[11377] = 32'b11111111111111111010001000110110;
assign LUT_4[11378] = 32'b00000000000000000000010111100010;
assign LUT_4[11379] = 32'b11111111111111111001100011011010;
assign LUT_4[11380] = 32'b11111111111111111101111101011010;
assign LUT_4[11381] = 32'b11111111111111110111001001010010;
assign LUT_4[11382] = 32'b11111111111111111101010111111110;
assign LUT_4[11383] = 32'b11111111111111110110100011110110;
assign LUT_4[11384] = 32'b11111111111111111010001001010011;
assign LUT_4[11385] = 32'b11111111111111110011010101001011;
assign LUT_4[11386] = 32'b11111111111111111001100011110111;
assign LUT_4[11387] = 32'b11111111111111110010101111101111;
assign LUT_4[11388] = 32'b11111111111111110111001001101111;
assign LUT_4[11389] = 32'b11111111111111110000010101100111;
assign LUT_4[11390] = 32'b11111111111111110110100100010011;
assign LUT_4[11391] = 32'b11111111111111101111110000001011;
assign LUT_4[11392] = 32'b00000000000000000101111110111101;
assign LUT_4[11393] = 32'b11111111111111111111001010110101;
assign LUT_4[11394] = 32'b00000000000000000101011001100001;
assign LUT_4[11395] = 32'b11111111111111111110100101011001;
assign LUT_4[11396] = 32'b00000000000000000010111111011001;
assign LUT_4[11397] = 32'b11111111111111111100001011010001;
assign LUT_4[11398] = 32'b00000000000000000010011001111101;
assign LUT_4[11399] = 32'b11111111111111111011100101110101;
assign LUT_4[11400] = 32'b11111111111111111111001011010010;
assign LUT_4[11401] = 32'b11111111111111111000010111001010;
assign LUT_4[11402] = 32'b11111111111111111110100101110110;
assign LUT_4[11403] = 32'b11111111111111110111110001101110;
assign LUT_4[11404] = 32'b11111111111111111100001011101110;
assign LUT_4[11405] = 32'b11111111111111110101010111100110;
assign LUT_4[11406] = 32'b11111111111111111011100110010010;
assign LUT_4[11407] = 32'b11111111111111110100110010001010;
assign LUT_4[11408] = 32'b00000000000000000011110000101011;
assign LUT_4[11409] = 32'b11111111111111111100111100100011;
assign LUT_4[11410] = 32'b00000000000000000011001011001111;
assign LUT_4[11411] = 32'b11111111111111111100010111000111;
assign LUT_4[11412] = 32'b00000000000000000000110001000111;
assign LUT_4[11413] = 32'b11111111111111111001111100111111;
assign LUT_4[11414] = 32'b00000000000000000000001011101011;
assign LUT_4[11415] = 32'b11111111111111111001010111100011;
assign LUT_4[11416] = 32'b11111111111111111100111101000000;
assign LUT_4[11417] = 32'b11111111111111110110001000111000;
assign LUT_4[11418] = 32'b11111111111111111100010111100100;
assign LUT_4[11419] = 32'b11111111111111110101100011011100;
assign LUT_4[11420] = 32'b11111111111111111001111101011100;
assign LUT_4[11421] = 32'b11111111111111110011001001010100;
assign LUT_4[11422] = 32'b11111111111111111001011000000000;
assign LUT_4[11423] = 32'b11111111111111110010100011111000;
assign LUT_4[11424] = 32'b00000000000000000100011010000100;
assign LUT_4[11425] = 32'b11111111111111111101100101111100;
assign LUT_4[11426] = 32'b00000000000000000011110100101000;
assign LUT_4[11427] = 32'b11111111111111111101000000100000;
assign LUT_4[11428] = 32'b00000000000000000001011010100000;
assign LUT_4[11429] = 32'b11111111111111111010100110011000;
assign LUT_4[11430] = 32'b00000000000000000000110101000100;
assign LUT_4[11431] = 32'b11111111111111111010000000111100;
assign LUT_4[11432] = 32'b11111111111111111101100110011001;
assign LUT_4[11433] = 32'b11111111111111110110110010010001;
assign LUT_4[11434] = 32'b11111111111111111101000000111101;
assign LUT_4[11435] = 32'b11111111111111110110001100110101;
assign LUT_4[11436] = 32'b11111111111111111010100110110101;
assign LUT_4[11437] = 32'b11111111111111110011110010101101;
assign LUT_4[11438] = 32'b11111111111111111010000001011001;
assign LUT_4[11439] = 32'b11111111111111110011001101010001;
assign LUT_4[11440] = 32'b00000000000000000010001011110010;
assign LUT_4[11441] = 32'b11111111111111111011010111101010;
assign LUT_4[11442] = 32'b00000000000000000001100110010110;
assign LUT_4[11443] = 32'b11111111111111111010110010001110;
assign LUT_4[11444] = 32'b11111111111111111111001100001110;
assign LUT_4[11445] = 32'b11111111111111111000011000000110;
assign LUT_4[11446] = 32'b11111111111111111110100110110010;
assign LUT_4[11447] = 32'b11111111111111110111110010101010;
assign LUT_4[11448] = 32'b11111111111111111011011000000111;
assign LUT_4[11449] = 32'b11111111111111110100100011111111;
assign LUT_4[11450] = 32'b11111111111111111010110010101011;
assign LUT_4[11451] = 32'b11111111111111110011111110100011;
assign LUT_4[11452] = 32'b11111111111111111000011000100011;
assign LUT_4[11453] = 32'b11111111111111110001100100011011;
assign LUT_4[11454] = 32'b11111111111111110111110011000111;
assign LUT_4[11455] = 32'b11111111111111110000111110111111;
assign LUT_4[11456] = 32'b00000000000000000111010110010001;
assign LUT_4[11457] = 32'b00000000000000000000100010001001;
assign LUT_4[11458] = 32'b00000000000000000110110000110101;
assign LUT_4[11459] = 32'b11111111111111111111111100101101;
assign LUT_4[11460] = 32'b00000000000000000100010110101101;
assign LUT_4[11461] = 32'b11111111111111111101100010100101;
assign LUT_4[11462] = 32'b00000000000000000011110001010001;
assign LUT_4[11463] = 32'b11111111111111111100111101001001;
assign LUT_4[11464] = 32'b00000000000000000000100010100110;
assign LUT_4[11465] = 32'b11111111111111111001101110011110;
assign LUT_4[11466] = 32'b11111111111111111111111101001010;
assign LUT_4[11467] = 32'b11111111111111111001001001000010;
assign LUT_4[11468] = 32'b11111111111111111101100011000010;
assign LUT_4[11469] = 32'b11111111111111110110101110111010;
assign LUT_4[11470] = 32'b11111111111111111100111101100110;
assign LUT_4[11471] = 32'b11111111111111110110001001011110;
assign LUT_4[11472] = 32'b00000000000000000101000111111111;
assign LUT_4[11473] = 32'b11111111111111111110010011110111;
assign LUT_4[11474] = 32'b00000000000000000100100010100011;
assign LUT_4[11475] = 32'b11111111111111111101101110011011;
assign LUT_4[11476] = 32'b00000000000000000010001000011011;
assign LUT_4[11477] = 32'b11111111111111111011010100010011;
assign LUT_4[11478] = 32'b00000000000000000001100010111111;
assign LUT_4[11479] = 32'b11111111111111111010101110110111;
assign LUT_4[11480] = 32'b11111111111111111110010100010100;
assign LUT_4[11481] = 32'b11111111111111110111100000001100;
assign LUT_4[11482] = 32'b11111111111111111101101110111000;
assign LUT_4[11483] = 32'b11111111111111110110111010110000;
assign LUT_4[11484] = 32'b11111111111111111011010100110000;
assign LUT_4[11485] = 32'b11111111111111110100100000101000;
assign LUT_4[11486] = 32'b11111111111111111010101111010100;
assign LUT_4[11487] = 32'b11111111111111110011111011001100;
assign LUT_4[11488] = 32'b00000000000000000101110001011000;
assign LUT_4[11489] = 32'b11111111111111111110111101010000;
assign LUT_4[11490] = 32'b00000000000000000101001011111100;
assign LUT_4[11491] = 32'b11111111111111111110010111110100;
assign LUT_4[11492] = 32'b00000000000000000010110001110100;
assign LUT_4[11493] = 32'b11111111111111111011111101101100;
assign LUT_4[11494] = 32'b00000000000000000010001100011000;
assign LUT_4[11495] = 32'b11111111111111111011011000010000;
assign LUT_4[11496] = 32'b11111111111111111110111101101101;
assign LUT_4[11497] = 32'b11111111111111111000001001100101;
assign LUT_4[11498] = 32'b11111111111111111110011000010001;
assign LUT_4[11499] = 32'b11111111111111110111100100001001;
assign LUT_4[11500] = 32'b11111111111111111011111110001001;
assign LUT_4[11501] = 32'b11111111111111110101001010000001;
assign LUT_4[11502] = 32'b11111111111111111011011000101101;
assign LUT_4[11503] = 32'b11111111111111110100100100100101;
assign LUT_4[11504] = 32'b00000000000000000011100011000110;
assign LUT_4[11505] = 32'b11111111111111111100101110111110;
assign LUT_4[11506] = 32'b00000000000000000010111101101010;
assign LUT_4[11507] = 32'b11111111111111111100001001100010;
assign LUT_4[11508] = 32'b00000000000000000000100011100010;
assign LUT_4[11509] = 32'b11111111111111111001101111011010;
assign LUT_4[11510] = 32'b11111111111111111111111110000110;
assign LUT_4[11511] = 32'b11111111111111111001001001111110;
assign LUT_4[11512] = 32'b11111111111111111100101111011011;
assign LUT_4[11513] = 32'b11111111111111110101111011010011;
assign LUT_4[11514] = 32'b11111111111111111100001001111111;
assign LUT_4[11515] = 32'b11111111111111110101010101110111;
assign LUT_4[11516] = 32'b11111111111111111001101111110111;
assign LUT_4[11517] = 32'b11111111111111110010111011101111;
assign LUT_4[11518] = 32'b11111111111111111001001010011011;
assign LUT_4[11519] = 32'b11111111111111110010010110010011;
assign LUT_4[11520] = 32'b00000000000000001000010100011000;
assign LUT_4[11521] = 32'b00000000000000000001100000010000;
assign LUT_4[11522] = 32'b00000000000000000111101110111100;
assign LUT_4[11523] = 32'b00000000000000000000111010110100;
assign LUT_4[11524] = 32'b00000000000000000101010100110100;
assign LUT_4[11525] = 32'b11111111111111111110100000101100;
assign LUT_4[11526] = 32'b00000000000000000100101111011000;
assign LUT_4[11527] = 32'b11111111111111111101111011010000;
assign LUT_4[11528] = 32'b00000000000000000001100000101101;
assign LUT_4[11529] = 32'b11111111111111111010101100100101;
assign LUT_4[11530] = 32'b00000000000000000000111011010001;
assign LUT_4[11531] = 32'b11111111111111111010000111001001;
assign LUT_4[11532] = 32'b11111111111111111110100001001001;
assign LUT_4[11533] = 32'b11111111111111110111101101000001;
assign LUT_4[11534] = 32'b11111111111111111101111011101101;
assign LUT_4[11535] = 32'b11111111111111110111000111100101;
assign LUT_4[11536] = 32'b00000000000000000110000110000110;
assign LUT_4[11537] = 32'b11111111111111111111010001111110;
assign LUT_4[11538] = 32'b00000000000000000101100000101010;
assign LUT_4[11539] = 32'b11111111111111111110101100100010;
assign LUT_4[11540] = 32'b00000000000000000011000110100010;
assign LUT_4[11541] = 32'b11111111111111111100010010011010;
assign LUT_4[11542] = 32'b00000000000000000010100001000110;
assign LUT_4[11543] = 32'b11111111111111111011101100111110;
assign LUT_4[11544] = 32'b11111111111111111111010010011011;
assign LUT_4[11545] = 32'b11111111111111111000011110010011;
assign LUT_4[11546] = 32'b11111111111111111110101100111111;
assign LUT_4[11547] = 32'b11111111111111110111111000110111;
assign LUT_4[11548] = 32'b11111111111111111100010010110111;
assign LUT_4[11549] = 32'b11111111111111110101011110101111;
assign LUT_4[11550] = 32'b11111111111111111011101101011011;
assign LUT_4[11551] = 32'b11111111111111110100111001010011;
assign LUT_4[11552] = 32'b00000000000000000110101111011111;
assign LUT_4[11553] = 32'b11111111111111111111111011010111;
assign LUT_4[11554] = 32'b00000000000000000110001010000011;
assign LUT_4[11555] = 32'b11111111111111111111010101111011;
assign LUT_4[11556] = 32'b00000000000000000011101111111011;
assign LUT_4[11557] = 32'b11111111111111111100111011110011;
assign LUT_4[11558] = 32'b00000000000000000011001010011111;
assign LUT_4[11559] = 32'b11111111111111111100010110010111;
assign LUT_4[11560] = 32'b11111111111111111111111011110100;
assign LUT_4[11561] = 32'b11111111111111111001000111101100;
assign LUT_4[11562] = 32'b11111111111111111111010110011000;
assign LUT_4[11563] = 32'b11111111111111111000100010010000;
assign LUT_4[11564] = 32'b11111111111111111100111100010000;
assign LUT_4[11565] = 32'b11111111111111110110001000001000;
assign LUT_4[11566] = 32'b11111111111111111100010110110100;
assign LUT_4[11567] = 32'b11111111111111110101100010101100;
assign LUT_4[11568] = 32'b00000000000000000100100001001101;
assign LUT_4[11569] = 32'b11111111111111111101101101000101;
assign LUT_4[11570] = 32'b00000000000000000011111011110001;
assign LUT_4[11571] = 32'b11111111111111111101000111101001;
assign LUT_4[11572] = 32'b00000000000000000001100001101001;
assign LUT_4[11573] = 32'b11111111111111111010101101100001;
assign LUT_4[11574] = 32'b00000000000000000000111100001101;
assign LUT_4[11575] = 32'b11111111111111111010001000000101;
assign LUT_4[11576] = 32'b11111111111111111101101101100010;
assign LUT_4[11577] = 32'b11111111111111110110111001011010;
assign LUT_4[11578] = 32'b11111111111111111101001000000110;
assign LUT_4[11579] = 32'b11111111111111110110010011111110;
assign LUT_4[11580] = 32'b11111111111111111010101101111110;
assign LUT_4[11581] = 32'b11111111111111110011111001110110;
assign LUT_4[11582] = 32'b11111111111111111010001000100010;
assign LUT_4[11583] = 32'b11111111111111110011010100011010;
assign LUT_4[11584] = 32'b00000000000000001001101011101100;
assign LUT_4[11585] = 32'b00000000000000000010110111100100;
assign LUT_4[11586] = 32'b00000000000000001001000110010000;
assign LUT_4[11587] = 32'b00000000000000000010010010001000;
assign LUT_4[11588] = 32'b00000000000000000110101100001000;
assign LUT_4[11589] = 32'b11111111111111111111111000000000;
assign LUT_4[11590] = 32'b00000000000000000110000110101100;
assign LUT_4[11591] = 32'b11111111111111111111010010100100;
assign LUT_4[11592] = 32'b00000000000000000010111000000001;
assign LUT_4[11593] = 32'b11111111111111111100000011111001;
assign LUT_4[11594] = 32'b00000000000000000010010010100101;
assign LUT_4[11595] = 32'b11111111111111111011011110011101;
assign LUT_4[11596] = 32'b11111111111111111111111000011101;
assign LUT_4[11597] = 32'b11111111111111111001000100010101;
assign LUT_4[11598] = 32'b11111111111111111111010011000001;
assign LUT_4[11599] = 32'b11111111111111111000011110111001;
assign LUT_4[11600] = 32'b00000000000000000111011101011010;
assign LUT_4[11601] = 32'b00000000000000000000101001010010;
assign LUT_4[11602] = 32'b00000000000000000110110111111110;
assign LUT_4[11603] = 32'b00000000000000000000000011110110;
assign LUT_4[11604] = 32'b00000000000000000100011101110110;
assign LUT_4[11605] = 32'b11111111111111111101101001101110;
assign LUT_4[11606] = 32'b00000000000000000011111000011010;
assign LUT_4[11607] = 32'b11111111111111111101000100010010;
assign LUT_4[11608] = 32'b00000000000000000000101001101111;
assign LUT_4[11609] = 32'b11111111111111111001110101100111;
assign LUT_4[11610] = 32'b00000000000000000000000100010011;
assign LUT_4[11611] = 32'b11111111111111111001010000001011;
assign LUT_4[11612] = 32'b11111111111111111101101010001011;
assign LUT_4[11613] = 32'b11111111111111110110110110000011;
assign LUT_4[11614] = 32'b11111111111111111101000100101111;
assign LUT_4[11615] = 32'b11111111111111110110010000100111;
assign LUT_4[11616] = 32'b00000000000000001000000110110011;
assign LUT_4[11617] = 32'b00000000000000000001010010101011;
assign LUT_4[11618] = 32'b00000000000000000111100001010111;
assign LUT_4[11619] = 32'b00000000000000000000101101001111;
assign LUT_4[11620] = 32'b00000000000000000101000111001111;
assign LUT_4[11621] = 32'b11111111111111111110010011000111;
assign LUT_4[11622] = 32'b00000000000000000100100001110011;
assign LUT_4[11623] = 32'b11111111111111111101101101101011;
assign LUT_4[11624] = 32'b00000000000000000001010011001000;
assign LUT_4[11625] = 32'b11111111111111111010011111000000;
assign LUT_4[11626] = 32'b00000000000000000000101101101100;
assign LUT_4[11627] = 32'b11111111111111111001111001100100;
assign LUT_4[11628] = 32'b11111111111111111110010011100100;
assign LUT_4[11629] = 32'b11111111111111110111011111011100;
assign LUT_4[11630] = 32'b11111111111111111101101110001000;
assign LUT_4[11631] = 32'b11111111111111110110111010000000;
assign LUT_4[11632] = 32'b00000000000000000101111000100001;
assign LUT_4[11633] = 32'b11111111111111111111000100011001;
assign LUT_4[11634] = 32'b00000000000000000101010011000101;
assign LUT_4[11635] = 32'b11111111111111111110011110111101;
assign LUT_4[11636] = 32'b00000000000000000010111000111101;
assign LUT_4[11637] = 32'b11111111111111111100000100110101;
assign LUT_4[11638] = 32'b00000000000000000010010011100001;
assign LUT_4[11639] = 32'b11111111111111111011011111011001;
assign LUT_4[11640] = 32'b11111111111111111111000100110110;
assign LUT_4[11641] = 32'b11111111111111111000010000101110;
assign LUT_4[11642] = 32'b11111111111111111110011111011010;
assign LUT_4[11643] = 32'b11111111111111110111101011010010;
assign LUT_4[11644] = 32'b11111111111111111100000101010010;
assign LUT_4[11645] = 32'b11111111111111110101010001001010;
assign LUT_4[11646] = 32'b11111111111111111011011111110110;
assign LUT_4[11647] = 32'b11111111111111110100101011101110;
assign LUT_4[11648] = 32'b00000000000000001010111010100000;
assign LUT_4[11649] = 32'b00000000000000000100000110011000;
assign LUT_4[11650] = 32'b00000000000000001010010101000100;
assign LUT_4[11651] = 32'b00000000000000000011100000111100;
assign LUT_4[11652] = 32'b00000000000000000111111010111100;
assign LUT_4[11653] = 32'b00000000000000000001000110110100;
assign LUT_4[11654] = 32'b00000000000000000111010101100000;
assign LUT_4[11655] = 32'b00000000000000000000100001011000;
assign LUT_4[11656] = 32'b00000000000000000100000110110101;
assign LUT_4[11657] = 32'b11111111111111111101010010101101;
assign LUT_4[11658] = 32'b00000000000000000011100001011001;
assign LUT_4[11659] = 32'b11111111111111111100101101010001;
assign LUT_4[11660] = 32'b00000000000000000001000111010001;
assign LUT_4[11661] = 32'b11111111111111111010010011001001;
assign LUT_4[11662] = 32'b00000000000000000000100001110101;
assign LUT_4[11663] = 32'b11111111111111111001101101101101;
assign LUT_4[11664] = 32'b00000000000000001000101100001110;
assign LUT_4[11665] = 32'b00000000000000000001111000000110;
assign LUT_4[11666] = 32'b00000000000000001000000110110010;
assign LUT_4[11667] = 32'b00000000000000000001010010101010;
assign LUT_4[11668] = 32'b00000000000000000101101100101010;
assign LUT_4[11669] = 32'b11111111111111111110111000100010;
assign LUT_4[11670] = 32'b00000000000000000101000111001110;
assign LUT_4[11671] = 32'b11111111111111111110010011000110;
assign LUT_4[11672] = 32'b00000000000000000001111000100011;
assign LUT_4[11673] = 32'b11111111111111111011000100011011;
assign LUT_4[11674] = 32'b00000000000000000001010011000111;
assign LUT_4[11675] = 32'b11111111111111111010011110111111;
assign LUT_4[11676] = 32'b11111111111111111110111000111111;
assign LUT_4[11677] = 32'b11111111111111111000000100110111;
assign LUT_4[11678] = 32'b11111111111111111110010011100011;
assign LUT_4[11679] = 32'b11111111111111110111011111011011;
assign LUT_4[11680] = 32'b00000000000000001001010101100111;
assign LUT_4[11681] = 32'b00000000000000000010100001011111;
assign LUT_4[11682] = 32'b00000000000000001000110000001011;
assign LUT_4[11683] = 32'b00000000000000000001111100000011;
assign LUT_4[11684] = 32'b00000000000000000110010110000011;
assign LUT_4[11685] = 32'b11111111111111111111100001111011;
assign LUT_4[11686] = 32'b00000000000000000101110000100111;
assign LUT_4[11687] = 32'b11111111111111111110111100011111;
assign LUT_4[11688] = 32'b00000000000000000010100001111100;
assign LUT_4[11689] = 32'b11111111111111111011101101110100;
assign LUT_4[11690] = 32'b00000000000000000001111100100000;
assign LUT_4[11691] = 32'b11111111111111111011001000011000;
assign LUT_4[11692] = 32'b11111111111111111111100010011000;
assign LUT_4[11693] = 32'b11111111111111111000101110010000;
assign LUT_4[11694] = 32'b11111111111111111110111100111100;
assign LUT_4[11695] = 32'b11111111111111111000001000110100;
assign LUT_4[11696] = 32'b00000000000000000111000111010101;
assign LUT_4[11697] = 32'b00000000000000000000010011001101;
assign LUT_4[11698] = 32'b00000000000000000110100001111001;
assign LUT_4[11699] = 32'b11111111111111111111101101110001;
assign LUT_4[11700] = 32'b00000000000000000100000111110001;
assign LUT_4[11701] = 32'b11111111111111111101010011101001;
assign LUT_4[11702] = 32'b00000000000000000011100010010101;
assign LUT_4[11703] = 32'b11111111111111111100101110001101;
assign LUT_4[11704] = 32'b00000000000000000000010011101010;
assign LUT_4[11705] = 32'b11111111111111111001011111100010;
assign LUT_4[11706] = 32'b11111111111111111111101110001110;
assign LUT_4[11707] = 32'b11111111111111111000111010000110;
assign LUT_4[11708] = 32'b11111111111111111101010100000110;
assign LUT_4[11709] = 32'b11111111111111110110011111111110;
assign LUT_4[11710] = 32'b11111111111111111100101110101010;
assign LUT_4[11711] = 32'b11111111111111110101111010100010;
assign LUT_4[11712] = 32'b00000000000000001100010001110100;
assign LUT_4[11713] = 32'b00000000000000000101011101101100;
assign LUT_4[11714] = 32'b00000000000000001011101100011000;
assign LUT_4[11715] = 32'b00000000000000000100111000010000;
assign LUT_4[11716] = 32'b00000000000000001001010010010000;
assign LUT_4[11717] = 32'b00000000000000000010011110001000;
assign LUT_4[11718] = 32'b00000000000000001000101100110100;
assign LUT_4[11719] = 32'b00000000000000000001111000101100;
assign LUT_4[11720] = 32'b00000000000000000101011110001001;
assign LUT_4[11721] = 32'b11111111111111111110101010000001;
assign LUT_4[11722] = 32'b00000000000000000100111000101101;
assign LUT_4[11723] = 32'b11111111111111111110000100100101;
assign LUT_4[11724] = 32'b00000000000000000010011110100101;
assign LUT_4[11725] = 32'b11111111111111111011101010011101;
assign LUT_4[11726] = 32'b00000000000000000001111001001001;
assign LUT_4[11727] = 32'b11111111111111111011000101000001;
assign LUT_4[11728] = 32'b00000000000000001010000011100010;
assign LUT_4[11729] = 32'b00000000000000000011001111011010;
assign LUT_4[11730] = 32'b00000000000000001001011110000110;
assign LUT_4[11731] = 32'b00000000000000000010101001111110;
assign LUT_4[11732] = 32'b00000000000000000111000011111110;
assign LUT_4[11733] = 32'b00000000000000000000001111110110;
assign LUT_4[11734] = 32'b00000000000000000110011110100010;
assign LUT_4[11735] = 32'b11111111111111111111101010011010;
assign LUT_4[11736] = 32'b00000000000000000011001111110111;
assign LUT_4[11737] = 32'b11111111111111111100011011101111;
assign LUT_4[11738] = 32'b00000000000000000010101010011011;
assign LUT_4[11739] = 32'b11111111111111111011110110010011;
assign LUT_4[11740] = 32'b00000000000000000000010000010011;
assign LUT_4[11741] = 32'b11111111111111111001011100001011;
assign LUT_4[11742] = 32'b11111111111111111111101010110111;
assign LUT_4[11743] = 32'b11111111111111111000110110101111;
assign LUT_4[11744] = 32'b00000000000000001010101100111011;
assign LUT_4[11745] = 32'b00000000000000000011111000110011;
assign LUT_4[11746] = 32'b00000000000000001010000111011111;
assign LUT_4[11747] = 32'b00000000000000000011010011010111;
assign LUT_4[11748] = 32'b00000000000000000111101101010111;
assign LUT_4[11749] = 32'b00000000000000000000111001001111;
assign LUT_4[11750] = 32'b00000000000000000111000111111011;
assign LUT_4[11751] = 32'b00000000000000000000010011110011;
assign LUT_4[11752] = 32'b00000000000000000011111001010000;
assign LUT_4[11753] = 32'b11111111111111111101000101001000;
assign LUT_4[11754] = 32'b00000000000000000011010011110100;
assign LUT_4[11755] = 32'b11111111111111111100011111101100;
assign LUT_4[11756] = 32'b00000000000000000000111001101100;
assign LUT_4[11757] = 32'b11111111111111111010000101100100;
assign LUT_4[11758] = 32'b00000000000000000000010100010000;
assign LUT_4[11759] = 32'b11111111111111111001100000001000;
assign LUT_4[11760] = 32'b00000000000000001000011110101001;
assign LUT_4[11761] = 32'b00000000000000000001101010100001;
assign LUT_4[11762] = 32'b00000000000000000111111001001101;
assign LUT_4[11763] = 32'b00000000000000000001000101000101;
assign LUT_4[11764] = 32'b00000000000000000101011111000101;
assign LUT_4[11765] = 32'b11111111111111111110101010111101;
assign LUT_4[11766] = 32'b00000000000000000100111001101001;
assign LUT_4[11767] = 32'b11111111111111111110000101100001;
assign LUT_4[11768] = 32'b00000000000000000001101010111110;
assign LUT_4[11769] = 32'b11111111111111111010110110110110;
assign LUT_4[11770] = 32'b00000000000000000001000101100010;
assign LUT_4[11771] = 32'b11111111111111111010010001011010;
assign LUT_4[11772] = 32'b11111111111111111110101011011010;
assign LUT_4[11773] = 32'b11111111111111110111110111010010;
assign LUT_4[11774] = 32'b11111111111111111110000101111110;
assign LUT_4[11775] = 32'b11111111111111110111010001110110;
assign LUT_4[11776] = 32'b00000000000000000010011100111101;
assign LUT_4[11777] = 32'b11111111111111111011101000110101;
assign LUT_4[11778] = 32'b00000000000000000001110111100001;
assign LUT_4[11779] = 32'b11111111111111111011000011011001;
assign LUT_4[11780] = 32'b11111111111111111111011101011001;
assign LUT_4[11781] = 32'b11111111111111111000101001010001;
assign LUT_4[11782] = 32'b11111111111111111110110111111101;
assign LUT_4[11783] = 32'b11111111111111111000000011110101;
assign LUT_4[11784] = 32'b11111111111111111011101001010010;
assign LUT_4[11785] = 32'b11111111111111110100110101001010;
assign LUT_4[11786] = 32'b11111111111111111011000011110110;
assign LUT_4[11787] = 32'b11111111111111110100001111101110;
assign LUT_4[11788] = 32'b11111111111111111000101001101110;
assign LUT_4[11789] = 32'b11111111111111110001110101100110;
assign LUT_4[11790] = 32'b11111111111111111000000100010010;
assign LUT_4[11791] = 32'b11111111111111110001010000001010;
assign LUT_4[11792] = 32'b00000000000000000000001110101011;
assign LUT_4[11793] = 32'b11111111111111111001011010100011;
assign LUT_4[11794] = 32'b11111111111111111111101001001111;
assign LUT_4[11795] = 32'b11111111111111111000110101000111;
assign LUT_4[11796] = 32'b11111111111111111101001111000111;
assign LUT_4[11797] = 32'b11111111111111110110011010111111;
assign LUT_4[11798] = 32'b11111111111111111100101001101011;
assign LUT_4[11799] = 32'b11111111111111110101110101100011;
assign LUT_4[11800] = 32'b11111111111111111001011011000000;
assign LUT_4[11801] = 32'b11111111111111110010100110111000;
assign LUT_4[11802] = 32'b11111111111111111000110101100100;
assign LUT_4[11803] = 32'b11111111111111110010000001011100;
assign LUT_4[11804] = 32'b11111111111111110110011011011100;
assign LUT_4[11805] = 32'b11111111111111101111100111010100;
assign LUT_4[11806] = 32'b11111111111111110101110110000000;
assign LUT_4[11807] = 32'b11111111111111101111000001111000;
assign LUT_4[11808] = 32'b00000000000000000000111000000100;
assign LUT_4[11809] = 32'b11111111111111111010000011111100;
assign LUT_4[11810] = 32'b00000000000000000000010010101000;
assign LUT_4[11811] = 32'b11111111111111111001011110100000;
assign LUT_4[11812] = 32'b11111111111111111101111000100000;
assign LUT_4[11813] = 32'b11111111111111110111000100011000;
assign LUT_4[11814] = 32'b11111111111111111101010011000100;
assign LUT_4[11815] = 32'b11111111111111110110011110111100;
assign LUT_4[11816] = 32'b11111111111111111010000100011001;
assign LUT_4[11817] = 32'b11111111111111110011010000010001;
assign LUT_4[11818] = 32'b11111111111111111001011110111101;
assign LUT_4[11819] = 32'b11111111111111110010101010110101;
assign LUT_4[11820] = 32'b11111111111111110111000100110101;
assign LUT_4[11821] = 32'b11111111111111110000010000101101;
assign LUT_4[11822] = 32'b11111111111111110110011111011001;
assign LUT_4[11823] = 32'b11111111111111101111101011010001;
assign LUT_4[11824] = 32'b11111111111111111110101001110010;
assign LUT_4[11825] = 32'b11111111111111110111110101101010;
assign LUT_4[11826] = 32'b11111111111111111110000100010110;
assign LUT_4[11827] = 32'b11111111111111110111010000001110;
assign LUT_4[11828] = 32'b11111111111111111011101010001110;
assign LUT_4[11829] = 32'b11111111111111110100110110000110;
assign LUT_4[11830] = 32'b11111111111111111011000100110010;
assign LUT_4[11831] = 32'b11111111111111110100010000101010;
assign LUT_4[11832] = 32'b11111111111111110111110110000111;
assign LUT_4[11833] = 32'b11111111111111110001000001111111;
assign LUT_4[11834] = 32'b11111111111111110111010000101011;
assign LUT_4[11835] = 32'b11111111111111110000011100100011;
assign LUT_4[11836] = 32'b11111111111111110100110110100011;
assign LUT_4[11837] = 32'b11111111111111101110000010011011;
assign LUT_4[11838] = 32'b11111111111111110100010001000111;
assign LUT_4[11839] = 32'b11111111111111101101011100111111;
assign LUT_4[11840] = 32'b00000000000000000011110100010001;
assign LUT_4[11841] = 32'b11111111111111111101000000001001;
assign LUT_4[11842] = 32'b00000000000000000011001110110101;
assign LUT_4[11843] = 32'b11111111111111111100011010101101;
assign LUT_4[11844] = 32'b00000000000000000000110100101101;
assign LUT_4[11845] = 32'b11111111111111111010000000100101;
assign LUT_4[11846] = 32'b00000000000000000000001111010001;
assign LUT_4[11847] = 32'b11111111111111111001011011001001;
assign LUT_4[11848] = 32'b11111111111111111101000000100110;
assign LUT_4[11849] = 32'b11111111111111110110001100011110;
assign LUT_4[11850] = 32'b11111111111111111100011011001010;
assign LUT_4[11851] = 32'b11111111111111110101100111000010;
assign LUT_4[11852] = 32'b11111111111111111010000001000010;
assign LUT_4[11853] = 32'b11111111111111110011001100111010;
assign LUT_4[11854] = 32'b11111111111111111001011011100110;
assign LUT_4[11855] = 32'b11111111111111110010100111011110;
assign LUT_4[11856] = 32'b00000000000000000001100101111111;
assign LUT_4[11857] = 32'b11111111111111111010110001110111;
assign LUT_4[11858] = 32'b00000000000000000001000000100011;
assign LUT_4[11859] = 32'b11111111111111111010001100011011;
assign LUT_4[11860] = 32'b11111111111111111110100110011011;
assign LUT_4[11861] = 32'b11111111111111110111110010010011;
assign LUT_4[11862] = 32'b11111111111111111110000000111111;
assign LUT_4[11863] = 32'b11111111111111110111001100110111;
assign LUT_4[11864] = 32'b11111111111111111010110010010100;
assign LUT_4[11865] = 32'b11111111111111110011111110001100;
assign LUT_4[11866] = 32'b11111111111111111010001100111000;
assign LUT_4[11867] = 32'b11111111111111110011011000110000;
assign LUT_4[11868] = 32'b11111111111111110111110010110000;
assign LUT_4[11869] = 32'b11111111111111110000111110101000;
assign LUT_4[11870] = 32'b11111111111111110111001101010100;
assign LUT_4[11871] = 32'b11111111111111110000011001001100;
assign LUT_4[11872] = 32'b00000000000000000010001111011000;
assign LUT_4[11873] = 32'b11111111111111111011011011010000;
assign LUT_4[11874] = 32'b00000000000000000001101001111100;
assign LUT_4[11875] = 32'b11111111111111111010110101110100;
assign LUT_4[11876] = 32'b11111111111111111111001111110100;
assign LUT_4[11877] = 32'b11111111111111111000011011101100;
assign LUT_4[11878] = 32'b11111111111111111110101010011000;
assign LUT_4[11879] = 32'b11111111111111110111110110010000;
assign LUT_4[11880] = 32'b11111111111111111011011011101101;
assign LUT_4[11881] = 32'b11111111111111110100100111100101;
assign LUT_4[11882] = 32'b11111111111111111010110110010001;
assign LUT_4[11883] = 32'b11111111111111110100000010001001;
assign LUT_4[11884] = 32'b11111111111111111000011100001001;
assign LUT_4[11885] = 32'b11111111111111110001101000000001;
assign LUT_4[11886] = 32'b11111111111111110111110110101101;
assign LUT_4[11887] = 32'b11111111111111110001000010100101;
assign LUT_4[11888] = 32'b00000000000000000000000001000110;
assign LUT_4[11889] = 32'b11111111111111111001001100111110;
assign LUT_4[11890] = 32'b11111111111111111111011011101010;
assign LUT_4[11891] = 32'b11111111111111111000100111100010;
assign LUT_4[11892] = 32'b11111111111111111101000001100010;
assign LUT_4[11893] = 32'b11111111111111110110001101011010;
assign LUT_4[11894] = 32'b11111111111111111100011100000110;
assign LUT_4[11895] = 32'b11111111111111110101100111111110;
assign LUT_4[11896] = 32'b11111111111111111001001101011011;
assign LUT_4[11897] = 32'b11111111111111110010011001010011;
assign LUT_4[11898] = 32'b11111111111111111000100111111111;
assign LUT_4[11899] = 32'b11111111111111110001110011110111;
assign LUT_4[11900] = 32'b11111111111111110110001101110111;
assign LUT_4[11901] = 32'b11111111111111101111011001101111;
assign LUT_4[11902] = 32'b11111111111111110101101000011011;
assign LUT_4[11903] = 32'b11111111111111101110110100010011;
assign LUT_4[11904] = 32'b00000000000000000101000011000101;
assign LUT_4[11905] = 32'b11111111111111111110001110111101;
assign LUT_4[11906] = 32'b00000000000000000100011101101001;
assign LUT_4[11907] = 32'b11111111111111111101101001100001;
assign LUT_4[11908] = 32'b00000000000000000010000011100001;
assign LUT_4[11909] = 32'b11111111111111111011001111011001;
assign LUT_4[11910] = 32'b00000000000000000001011110000101;
assign LUT_4[11911] = 32'b11111111111111111010101001111101;
assign LUT_4[11912] = 32'b11111111111111111110001111011010;
assign LUT_4[11913] = 32'b11111111111111110111011011010010;
assign LUT_4[11914] = 32'b11111111111111111101101001111110;
assign LUT_4[11915] = 32'b11111111111111110110110101110110;
assign LUT_4[11916] = 32'b11111111111111111011001111110110;
assign LUT_4[11917] = 32'b11111111111111110100011011101110;
assign LUT_4[11918] = 32'b11111111111111111010101010011010;
assign LUT_4[11919] = 32'b11111111111111110011110110010010;
assign LUT_4[11920] = 32'b00000000000000000010110100110011;
assign LUT_4[11921] = 32'b11111111111111111100000000101011;
assign LUT_4[11922] = 32'b00000000000000000010001111010111;
assign LUT_4[11923] = 32'b11111111111111111011011011001111;
assign LUT_4[11924] = 32'b11111111111111111111110101001111;
assign LUT_4[11925] = 32'b11111111111111111001000001000111;
assign LUT_4[11926] = 32'b11111111111111111111001111110011;
assign LUT_4[11927] = 32'b11111111111111111000011011101011;
assign LUT_4[11928] = 32'b11111111111111111100000001001000;
assign LUT_4[11929] = 32'b11111111111111110101001101000000;
assign LUT_4[11930] = 32'b11111111111111111011011011101100;
assign LUT_4[11931] = 32'b11111111111111110100100111100100;
assign LUT_4[11932] = 32'b11111111111111111001000001100100;
assign LUT_4[11933] = 32'b11111111111111110010001101011100;
assign LUT_4[11934] = 32'b11111111111111111000011100001000;
assign LUT_4[11935] = 32'b11111111111111110001101000000000;
assign LUT_4[11936] = 32'b00000000000000000011011110001100;
assign LUT_4[11937] = 32'b11111111111111111100101010000100;
assign LUT_4[11938] = 32'b00000000000000000010111000110000;
assign LUT_4[11939] = 32'b11111111111111111100000100101000;
assign LUT_4[11940] = 32'b00000000000000000000011110101000;
assign LUT_4[11941] = 32'b11111111111111111001101010100000;
assign LUT_4[11942] = 32'b11111111111111111111111001001100;
assign LUT_4[11943] = 32'b11111111111111111001000101000100;
assign LUT_4[11944] = 32'b11111111111111111100101010100001;
assign LUT_4[11945] = 32'b11111111111111110101110110011001;
assign LUT_4[11946] = 32'b11111111111111111100000101000101;
assign LUT_4[11947] = 32'b11111111111111110101010000111101;
assign LUT_4[11948] = 32'b11111111111111111001101010111101;
assign LUT_4[11949] = 32'b11111111111111110010110110110101;
assign LUT_4[11950] = 32'b11111111111111111001000101100001;
assign LUT_4[11951] = 32'b11111111111111110010010001011001;
assign LUT_4[11952] = 32'b00000000000000000001001111111010;
assign LUT_4[11953] = 32'b11111111111111111010011011110010;
assign LUT_4[11954] = 32'b00000000000000000000101010011110;
assign LUT_4[11955] = 32'b11111111111111111001110110010110;
assign LUT_4[11956] = 32'b11111111111111111110010000010110;
assign LUT_4[11957] = 32'b11111111111111110111011100001110;
assign LUT_4[11958] = 32'b11111111111111111101101010111010;
assign LUT_4[11959] = 32'b11111111111111110110110110110010;
assign LUT_4[11960] = 32'b11111111111111111010011100001111;
assign LUT_4[11961] = 32'b11111111111111110011101000000111;
assign LUT_4[11962] = 32'b11111111111111111001110110110011;
assign LUT_4[11963] = 32'b11111111111111110011000010101011;
assign LUT_4[11964] = 32'b11111111111111110111011100101011;
assign LUT_4[11965] = 32'b11111111111111110000101000100011;
assign LUT_4[11966] = 32'b11111111111111110110110111001111;
assign LUT_4[11967] = 32'b11111111111111110000000011000111;
assign LUT_4[11968] = 32'b00000000000000000110011010011001;
assign LUT_4[11969] = 32'b11111111111111111111100110010001;
assign LUT_4[11970] = 32'b00000000000000000101110100111101;
assign LUT_4[11971] = 32'b11111111111111111111000000110101;
assign LUT_4[11972] = 32'b00000000000000000011011010110101;
assign LUT_4[11973] = 32'b11111111111111111100100110101101;
assign LUT_4[11974] = 32'b00000000000000000010110101011001;
assign LUT_4[11975] = 32'b11111111111111111100000001010001;
assign LUT_4[11976] = 32'b11111111111111111111100110101110;
assign LUT_4[11977] = 32'b11111111111111111000110010100110;
assign LUT_4[11978] = 32'b11111111111111111111000001010010;
assign LUT_4[11979] = 32'b11111111111111111000001101001010;
assign LUT_4[11980] = 32'b11111111111111111100100111001010;
assign LUT_4[11981] = 32'b11111111111111110101110011000010;
assign LUT_4[11982] = 32'b11111111111111111100000001101110;
assign LUT_4[11983] = 32'b11111111111111110101001101100110;
assign LUT_4[11984] = 32'b00000000000000000100001100000111;
assign LUT_4[11985] = 32'b11111111111111111101010111111111;
assign LUT_4[11986] = 32'b00000000000000000011100110101011;
assign LUT_4[11987] = 32'b11111111111111111100110010100011;
assign LUT_4[11988] = 32'b00000000000000000001001100100011;
assign LUT_4[11989] = 32'b11111111111111111010011000011011;
assign LUT_4[11990] = 32'b00000000000000000000100111000111;
assign LUT_4[11991] = 32'b11111111111111111001110010111111;
assign LUT_4[11992] = 32'b11111111111111111101011000011100;
assign LUT_4[11993] = 32'b11111111111111110110100100010100;
assign LUT_4[11994] = 32'b11111111111111111100110011000000;
assign LUT_4[11995] = 32'b11111111111111110101111110111000;
assign LUT_4[11996] = 32'b11111111111111111010011000111000;
assign LUT_4[11997] = 32'b11111111111111110011100100110000;
assign LUT_4[11998] = 32'b11111111111111111001110011011100;
assign LUT_4[11999] = 32'b11111111111111110010111111010100;
assign LUT_4[12000] = 32'b00000000000000000100110101100000;
assign LUT_4[12001] = 32'b11111111111111111110000001011000;
assign LUT_4[12002] = 32'b00000000000000000100010000000100;
assign LUT_4[12003] = 32'b11111111111111111101011011111100;
assign LUT_4[12004] = 32'b00000000000000000001110101111100;
assign LUT_4[12005] = 32'b11111111111111111011000001110100;
assign LUT_4[12006] = 32'b00000000000000000001010000100000;
assign LUT_4[12007] = 32'b11111111111111111010011100011000;
assign LUT_4[12008] = 32'b11111111111111111110000001110101;
assign LUT_4[12009] = 32'b11111111111111110111001101101101;
assign LUT_4[12010] = 32'b11111111111111111101011100011001;
assign LUT_4[12011] = 32'b11111111111111110110101000010001;
assign LUT_4[12012] = 32'b11111111111111111011000010010001;
assign LUT_4[12013] = 32'b11111111111111110100001110001001;
assign LUT_4[12014] = 32'b11111111111111111010011100110101;
assign LUT_4[12015] = 32'b11111111111111110011101000101101;
assign LUT_4[12016] = 32'b00000000000000000010100111001110;
assign LUT_4[12017] = 32'b11111111111111111011110011000110;
assign LUT_4[12018] = 32'b00000000000000000010000001110010;
assign LUT_4[12019] = 32'b11111111111111111011001101101010;
assign LUT_4[12020] = 32'b11111111111111111111100111101010;
assign LUT_4[12021] = 32'b11111111111111111000110011100010;
assign LUT_4[12022] = 32'b11111111111111111111000010001110;
assign LUT_4[12023] = 32'b11111111111111111000001110000110;
assign LUT_4[12024] = 32'b11111111111111111011110011100011;
assign LUT_4[12025] = 32'b11111111111111110100111111011011;
assign LUT_4[12026] = 32'b11111111111111111011001110000111;
assign LUT_4[12027] = 32'b11111111111111110100011001111111;
assign LUT_4[12028] = 32'b11111111111111111000110011111111;
assign LUT_4[12029] = 32'b11111111111111110001111111110111;
assign LUT_4[12030] = 32'b11111111111111111000001110100011;
assign LUT_4[12031] = 32'b11111111111111110001011010011011;
assign LUT_4[12032] = 32'b00000000000000000111011000100000;
assign LUT_4[12033] = 32'b00000000000000000000100100011000;
assign LUT_4[12034] = 32'b00000000000000000110110011000100;
assign LUT_4[12035] = 32'b11111111111111111111111110111100;
assign LUT_4[12036] = 32'b00000000000000000100011000111100;
assign LUT_4[12037] = 32'b11111111111111111101100100110100;
assign LUT_4[12038] = 32'b00000000000000000011110011100000;
assign LUT_4[12039] = 32'b11111111111111111100111111011000;
assign LUT_4[12040] = 32'b00000000000000000000100100110101;
assign LUT_4[12041] = 32'b11111111111111111001110000101101;
assign LUT_4[12042] = 32'b11111111111111111111111111011001;
assign LUT_4[12043] = 32'b11111111111111111001001011010001;
assign LUT_4[12044] = 32'b11111111111111111101100101010001;
assign LUT_4[12045] = 32'b11111111111111110110110001001001;
assign LUT_4[12046] = 32'b11111111111111111100111111110101;
assign LUT_4[12047] = 32'b11111111111111110110001011101101;
assign LUT_4[12048] = 32'b00000000000000000101001010001110;
assign LUT_4[12049] = 32'b11111111111111111110010110000110;
assign LUT_4[12050] = 32'b00000000000000000100100100110010;
assign LUT_4[12051] = 32'b11111111111111111101110000101010;
assign LUT_4[12052] = 32'b00000000000000000010001010101010;
assign LUT_4[12053] = 32'b11111111111111111011010110100010;
assign LUT_4[12054] = 32'b00000000000000000001100101001110;
assign LUT_4[12055] = 32'b11111111111111111010110001000110;
assign LUT_4[12056] = 32'b11111111111111111110010110100011;
assign LUT_4[12057] = 32'b11111111111111110111100010011011;
assign LUT_4[12058] = 32'b11111111111111111101110001000111;
assign LUT_4[12059] = 32'b11111111111111110110111100111111;
assign LUT_4[12060] = 32'b11111111111111111011010110111111;
assign LUT_4[12061] = 32'b11111111111111110100100010110111;
assign LUT_4[12062] = 32'b11111111111111111010110001100011;
assign LUT_4[12063] = 32'b11111111111111110011111101011011;
assign LUT_4[12064] = 32'b00000000000000000101110011100111;
assign LUT_4[12065] = 32'b11111111111111111110111111011111;
assign LUT_4[12066] = 32'b00000000000000000101001110001011;
assign LUT_4[12067] = 32'b11111111111111111110011010000011;
assign LUT_4[12068] = 32'b00000000000000000010110100000011;
assign LUT_4[12069] = 32'b11111111111111111011111111111011;
assign LUT_4[12070] = 32'b00000000000000000010001110100111;
assign LUT_4[12071] = 32'b11111111111111111011011010011111;
assign LUT_4[12072] = 32'b11111111111111111110111111111100;
assign LUT_4[12073] = 32'b11111111111111111000001011110100;
assign LUT_4[12074] = 32'b11111111111111111110011010100000;
assign LUT_4[12075] = 32'b11111111111111110111100110011000;
assign LUT_4[12076] = 32'b11111111111111111100000000011000;
assign LUT_4[12077] = 32'b11111111111111110101001100010000;
assign LUT_4[12078] = 32'b11111111111111111011011010111100;
assign LUT_4[12079] = 32'b11111111111111110100100110110100;
assign LUT_4[12080] = 32'b00000000000000000011100101010101;
assign LUT_4[12081] = 32'b11111111111111111100110001001101;
assign LUT_4[12082] = 32'b00000000000000000010111111111001;
assign LUT_4[12083] = 32'b11111111111111111100001011110001;
assign LUT_4[12084] = 32'b00000000000000000000100101110001;
assign LUT_4[12085] = 32'b11111111111111111001110001101001;
assign LUT_4[12086] = 32'b00000000000000000000000000010101;
assign LUT_4[12087] = 32'b11111111111111111001001100001101;
assign LUT_4[12088] = 32'b11111111111111111100110001101010;
assign LUT_4[12089] = 32'b11111111111111110101111101100010;
assign LUT_4[12090] = 32'b11111111111111111100001100001110;
assign LUT_4[12091] = 32'b11111111111111110101011000000110;
assign LUT_4[12092] = 32'b11111111111111111001110010000110;
assign LUT_4[12093] = 32'b11111111111111110010111101111110;
assign LUT_4[12094] = 32'b11111111111111111001001100101010;
assign LUT_4[12095] = 32'b11111111111111110010011000100010;
assign LUT_4[12096] = 32'b00000000000000001000101111110100;
assign LUT_4[12097] = 32'b00000000000000000001111011101100;
assign LUT_4[12098] = 32'b00000000000000001000001010011000;
assign LUT_4[12099] = 32'b00000000000000000001010110010000;
assign LUT_4[12100] = 32'b00000000000000000101110000010000;
assign LUT_4[12101] = 32'b11111111111111111110111100001000;
assign LUT_4[12102] = 32'b00000000000000000101001010110100;
assign LUT_4[12103] = 32'b11111111111111111110010110101100;
assign LUT_4[12104] = 32'b00000000000000000001111100001001;
assign LUT_4[12105] = 32'b11111111111111111011001000000001;
assign LUT_4[12106] = 32'b00000000000000000001010110101101;
assign LUT_4[12107] = 32'b11111111111111111010100010100101;
assign LUT_4[12108] = 32'b11111111111111111110111100100101;
assign LUT_4[12109] = 32'b11111111111111111000001000011101;
assign LUT_4[12110] = 32'b11111111111111111110010111001001;
assign LUT_4[12111] = 32'b11111111111111110111100011000001;
assign LUT_4[12112] = 32'b00000000000000000110100001100010;
assign LUT_4[12113] = 32'b11111111111111111111101101011010;
assign LUT_4[12114] = 32'b00000000000000000101111100000110;
assign LUT_4[12115] = 32'b11111111111111111111000111111110;
assign LUT_4[12116] = 32'b00000000000000000011100001111110;
assign LUT_4[12117] = 32'b11111111111111111100101101110110;
assign LUT_4[12118] = 32'b00000000000000000010111100100010;
assign LUT_4[12119] = 32'b11111111111111111100001000011010;
assign LUT_4[12120] = 32'b11111111111111111111101101110111;
assign LUT_4[12121] = 32'b11111111111111111000111001101111;
assign LUT_4[12122] = 32'b11111111111111111111001000011011;
assign LUT_4[12123] = 32'b11111111111111111000010100010011;
assign LUT_4[12124] = 32'b11111111111111111100101110010011;
assign LUT_4[12125] = 32'b11111111111111110101111010001011;
assign LUT_4[12126] = 32'b11111111111111111100001000110111;
assign LUT_4[12127] = 32'b11111111111111110101010100101111;
assign LUT_4[12128] = 32'b00000000000000000111001010111011;
assign LUT_4[12129] = 32'b00000000000000000000010110110011;
assign LUT_4[12130] = 32'b00000000000000000110100101011111;
assign LUT_4[12131] = 32'b11111111111111111111110001010111;
assign LUT_4[12132] = 32'b00000000000000000100001011010111;
assign LUT_4[12133] = 32'b11111111111111111101010111001111;
assign LUT_4[12134] = 32'b00000000000000000011100101111011;
assign LUT_4[12135] = 32'b11111111111111111100110001110011;
assign LUT_4[12136] = 32'b00000000000000000000010111010000;
assign LUT_4[12137] = 32'b11111111111111111001100011001000;
assign LUT_4[12138] = 32'b11111111111111111111110001110100;
assign LUT_4[12139] = 32'b11111111111111111000111101101100;
assign LUT_4[12140] = 32'b11111111111111111101010111101100;
assign LUT_4[12141] = 32'b11111111111111110110100011100100;
assign LUT_4[12142] = 32'b11111111111111111100110010010000;
assign LUT_4[12143] = 32'b11111111111111110101111110001000;
assign LUT_4[12144] = 32'b00000000000000000100111100101001;
assign LUT_4[12145] = 32'b11111111111111111110001000100001;
assign LUT_4[12146] = 32'b00000000000000000100010111001101;
assign LUT_4[12147] = 32'b11111111111111111101100011000101;
assign LUT_4[12148] = 32'b00000000000000000001111101000101;
assign LUT_4[12149] = 32'b11111111111111111011001000111101;
assign LUT_4[12150] = 32'b00000000000000000001010111101001;
assign LUT_4[12151] = 32'b11111111111111111010100011100001;
assign LUT_4[12152] = 32'b11111111111111111110001000111110;
assign LUT_4[12153] = 32'b11111111111111110111010100110110;
assign LUT_4[12154] = 32'b11111111111111111101100011100010;
assign LUT_4[12155] = 32'b11111111111111110110101111011010;
assign LUT_4[12156] = 32'b11111111111111111011001001011010;
assign LUT_4[12157] = 32'b11111111111111110100010101010010;
assign LUT_4[12158] = 32'b11111111111111111010100011111110;
assign LUT_4[12159] = 32'b11111111111111110011101111110110;
assign LUT_4[12160] = 32'b00000000000000001001111110101000;
assign LUT_4[12161] = 32'b00000000000000000011001010100000;
assign LUT_4[12162] = 32'b00000000000000001001011001001100;
assign LUT_4[12163] = 32'b00000000000000000010100101000100;
assign LUT_4[12164] = 32'b00000000000000000110111111000100;
assign LUT_4[12165] = 32'b00000000000000000000001010111100;
assign LUT_4[12166] = 32'b00000000000000000110011001101000;
assign LUT_4[12167] = 32'b11111111111111111111100101100000;
assign LUT_4[12168] = 32'b00000000000000000011001010111101;
assign LUT_4[12169] = 32'b11111111111111111100010110110101;
assign LUT_4[12170] = 32'b00000000000000000010100101100001;
assign LUT_4[12171] = 32'b11111111111111111011110001011001;
assign LUT_4[12172] = 32'b00000000000000000000001011011001;
assign LUT_4[12173] = 32'b11111111111111111001010111010001;
assign LUT_4[12174] = 32'b11111111111111111111100101111101;
assign LUT_4[12175] = 32'b11111111111111111000110001110101;
assign LUT_4[12176] = 32'b00000000000000000111110000010110;
assign LUT_4[12177] = 32'b00000000000000000000111100001110;
assign LUT_4[12178] = 32'b00000000000000000111001010111010;
assign LUT_4[12179] = 32'b00000000000000000000010110110010;
assign LUT_4[12180] = 32'b00000000000000000100110000110010;
assign LUT_4[12181] = 32'b11111111111111111101111100101010;
assign LUT_4[12182] = 32'b00000000000000000100001011010110;
assign LUT_4[12183] = 32'b11111111111111111101010111001110;
assign LUT_4[12184] = 32'b00000000000000000000111100101011;
assign LUT_4[12185] = 32'b11111111111111111010001000100011;
assign LUT_4[12186] = 32'b00000000000000000000010111001111;
assign LUT_4[12187] = 32'b11111111111111111001100011000111;
assign LUT_4[12188] = 32'b11111111111111111101111101000111;
assign LUT_4[12189] = 32'b11111111111111110111001000111111;
assign LUT_4[12190] = 32'b11111111111111111101010111101011;
assign LUT_4[12191] = 32'b11111111111111110110100011100011;
assign LUT_4[12192] = 32'b00000000000000001000011001101111;
assign LUT_4[12193] = 32'b00000000000000000001100101100111;
assign LUT_4[12194] = 32'b00000000000000000111110100010011;
assign LUT_4[12195] = 32'b00000000000000000001000000001011;
assign LUT_4[12196] = 32'b00000000000000000101011010001011;
assign LUT_4[12197] = 32'b11111111111111111110100110000011;
assign LUT_4[12198] = 32'b00000000000000000100110100101111;
assign LUT_4[12199] = 32'b11111111111111111110000000100111;
assign LUT_4[12200] = 32'b00000000000000000001100110000100;
assign LUT_4[12201] = 32'b11111111111111111010110001111100;
assign LUT_4[12202] = 32'b00000000000000000001000000101000;
assign LUT_4[12203] = 32'b11111111111111111010001100100000;
assign LUT_4[12204] = 32'b11111111111111111110100110100000;
assign LUT_4[12205] = 32'b11111111111111110111110010011000;
assign LUT_4[12206] = 32'b11111111111111111110000001000100;
assign LUT_4[12207] = 32'b11111111111111110111001100111100;
assign LUT_4[12208] = 32'b00000000000000000110001011011101;
assign LUT_4[12209] = 32'b11111111111111111111010111010101;
assign LUT_4[12210] = 32'b00000000000000000101100110000001;
assign LUT_4[12211] = 32'b11111111111111111110110001111001;
assign LUT_4[12212] = 32'b00000000000000000011001011111001;
assign LUT_4[12213] = 32'b11111111111111111100010111110001;
assign LUT_4[12214] = 32'b00000000000000000010100110011101;
assign LUT_4[12215] = 32'b11111111111111111011110010010101;
assign LUT_4[12216] = 32'b11111111111111111111010111110010;
assign LUT_4[12217] = 32'b11111111111111111000100011101010;
assign LUT_4[12218] = 32'b11111111111111111110110010010110;
assign LUT_4[12219] = 32'b11111111111111110111111110001110;
assign LUT_4[12220] = 32'b11111111111111111100011000001110;
assign LUT_4[12221] = 32'b11111111111111110101100100000110;
assign LUT_4[12222] = 32'b11111111111111111011110010110010;
assign LUT_4[12223] = 32'b11111111111111110100111110101010;
assign LUT_4[12224] = 32'b00000000000000001011010101111100;
assign LUT_4[12225] = 32'b00000000000000000100100001110100;
assign LUT_4[12226] = 32'b00000000000000001010110000100000;
assign LUT_4[12227] = 32'b00000000000000000011111100011000;
assign LUT_4[12228] = 32'b00000000000000001000010110011000;
assign LUT_4[12229] = 32'b00000000000000000001100010010000;
assign LUT_4[12230] = 32'b00000000000000000111110000111100;
assign LUT_4[12231] = 32'b00000000000000000000111100110100;
assign LUT_4[12232] = 32'b00000000000000000100100010010001;
assign LUT_4[12233] = 32'b11111111111111111101101110001001;
assign LUT_4[12234] = 32'b00000000000000000011111100110101;
assign LUT_4[12235] = 32'b11111111111111111101001000101101;
assign LUT_4[12236] = 32'b00000000000000000001100010101101;
assign LUT_4[12237] = 32'b11111111111111111010101110100101;
assign LUT_4[12238] = 32'b00000000000000000000111101010001;
assign LUT_4[12239] = 32'b11111111111111111010001001001001;
assign LUT_4[12240] = 32'b00000000000000001001000111101010;
assign LUT_4[12241] = 32'b00000000000000000010010011100010;
assign LUT_4[12242] = 32'b00000000000000001000100010001110;
assign LUT_4[12243] = 32'b00000000000000000001101110000110;
assign LUT_4[12244] = 32'b00000000000000000110001000000110;
assign LUT_4[12245] = 32'b11111111111111111111010011111110;
assign LUT_4[12246] = 32'b00000000000000000101100010101010;
assign LUT_4[12247] = 32'b11111111111111111110101110100010;
assign LUT_4[12248] = 32'b00000000000000000010010011111111;
assign LUT_4[12249] = 32'b11111111111111111011011111110111;
assign LUT_4[12250] = 32'b00000000000000000001101110100011;
assign LUT_4[12251] = 32'b11111111111111111010111010011011;
assign LUT_4[12252] = 32'b11111111111111111111010100011011;
assign LUT_4[12253] = 32'b11111111111111111000100000010011;
assign LUT_4[12254] = 32'b11111111111111111110101110111111;
assign LUT_4[12255] = 32'b11111111111111110111111010110111;
assign LUT_4[12256] = 32'b00000000000000001001110001000011;
assign LUT_4[12257] = 32'b00000000000000000010111100111011;
assign LUT_4[12258] = 32'b00000000000000001001001011100111;
assign LUT_4[12259] = 32'b00000000000000000010010111011111;
assign LUT_4[12260] = 32'b00000000000000000110110001011111;
assign LUT_4[12261] = 32'b11111111111111111111111101010111;
assign LUT_4[12262] = 32'b00000000000000000110001100000011;
assign LUT_4[12263] = 32'b11111111111111111111010111111011;
assign LUT_4[12264] = 32'b00000000000000000010111101011000;
assign LUT_4[12265] = 32'b11111111111111111100001001010000;
assign LUT_4[12266] = 32'b00000000000000000010010111111100;
assign LUT_4[12267] = 32'b11111111111111111011100011110100;
assign LUT_4[12268] = 32'b11111111111111111111111101110100;
assign LUT_4[12269] = 32'b11111111111111111001001001101100;
assign LUT_4[12270] = 32'b11111111111111111111011000011000;
assign LUT_4[12271] = 32'b11111111111111111000100100010000;
assign LUT_4[12272] = 32'b00000000000000000111100010110001;
assign LUT_4[12273] = 32'b00000000000000000000101110101001;
assign LUT_4[12274] = 32'b00000000000000000110111101010101;
assign LUT_4[12275] = 32'b00000000000000000000001001001101;
assign LUT_4[12276] = 32'b00000000000000000100100011001101;
assign LUT_4[12277] = 32'b11111111111111111101101111000101;
assign LUT_4[12278] = 32'b00000000000000000011111101110001;
assign LUT_4[12279] = 32'b11111111111111111101001001101001;
assign LUT_4[12280] = 32'b00000000000000000000101111000110;
assign LUT_4[12281] = 32'b11111111111111111001111010111110;
assign LUT_4[12282] = 32'b00000000000000000000001001101010;
assign LUT_4[12283] = 32'b11111111111111111001010101100010;
assign LUT_4[12284] = 32'b11111111111111111101101111100010;
assign LUT_4[12285] = 32'b11111111111111110110111011011010;
assign LUT_4[12286] = 32'b11111111111111111101001010000110;
assign LUT_4[12287] = 32'b11111111111111110110010101111110;
assign LUT_4[12288] = 32'b00000000000000000010011110111101;
assign LUT_4[12289] = 32'b11111111111111111011101010110101;
assign LUT_4[12290] = 32'b00000000000000000001111001100001;
assign LUT_4[12291] = 32'b11111111111111111011000101011001;
assign LUT_4[12292] = 32'b11111111111111111111011111011001;
assign LUT_4[12293] = 32'b11111111111111111000101011010001;
assign LUT_4[12294] = 32'b11111111111111111110111001111101;
assign LUT_4[12295] = 32'b11111111111111111000000101110101;
assign LUT_4[12296] = 32'b11111111111111111011101011010010;
assign LUT_4[12297] = 32'b11111111111111110100110111001010;
assign LUT_4[12298] = 32'b11111111111111111011000101110110;
assign LUT_4[12299] = 32'b11111111111111110100010001101110;
assign LUT_4[12300] = 32'b11111111111111111000101011101110;
assign LUT_4[12301] = 32'b11111111111111110001110111100110;
assign LUT_4[12302] = 32'b11111111111111111000000110010010;
assign LUT_4[12303] = 32'b11111111111111110001010010001010;
assign LUT_4[12304] = 32'b00000000000000000000010000101011;
assign LUT_4[12305] = 32'b11111111111111111001011100100011;
assign LUT_4[12306] = 32'b11111111111111111111101011001111;
assign LUT_4[12307] = 32'b11111111111111111000110111000111;
assign LUT_4[12308] = 32'b11111111111111111101010001000111;
assign LUT_4[12309] = 32'b11111111111111110110011100111111;
assign LUT_4[12310] = 32'b11111111111111111100101011101011;
assign LUT_4[12311] = 32'b11111111111111110101110111100011;
assign LUT_4[12312] = 32'b11111111111111111001011101000000;
assign LUT_4[12313] = 32'b11111111111111110010101000111000;
assign LUT_4[12314] = 32'b11111111111111111000110111100100;
assign LUT_4[12315] = 32'b11111111111111110010000011011100;
assign LUT_4[12316] = 32'b11111111111111110110011101011100;
assign LUT_4[12317] = 32'b11111111111111101111101001010100;
assign LUT_4[12318] = 32'b11111111111111110101111000000000;
assign LUT_4[12319] = 32'b11111111111111101111000011111000;
assign LUT_4[12320] = 32'b00000000000000000000111010000100;
assign LUT_4[12321] = 32'b11111111111111111010000101111100;
assign LUT_4[12322] = 32'b00000000000000000000010100101000;
assign LUT_4[12323] = 32'b11111111111111111001100000100000;
assign LUT_4[12324] = 32'b11111111111111111101111010100000;
assign LUT_4[12325] = 32'b11111111111111110111000110011000;
assign LUT_4[12326] = 32'b11111111111111111101010101000100;
assign LUT_4[12327] = 32'b11111111111111110110100000111100;
assign LUT_4[12328] = 32'b11111111111111111010000110011001;
assign LUT_4[12329] = 32'b11111111111111110011010010010001;
assign LUT_4[12330] = 32'b11111111111111111001100000111101;
assign LUT_4[12331] = 32'b11111111111111110010101100110101;
assign LUT_4[12332] = 32'b11111111111111110111000110110101;
assign LUT_4[12333] = 32'b11111111111111110000010010101101;
assign LUT_4[12334] = 32'b11111111111111110110100001011001;
assign LUT_4[12335] = 32'b11111111111111101111101101010001;
assign LUT_4[12336] = 32'b11111111111111111110101011110010;
assign LUT_4[12337] = 32'b11111111111111110111110111101010;
assign LUT_4[12338] = 32'b11111111111111111110000110010110;
assign LUT_4[12339] = 32'b11111111111111110111010010001110;
assign LUT_4[12340] = 32'b11111111111111111011101100001110;
assign LUT_4[12341] = 32'b11111111111111110100111000000110;
assign LUT_4[12342] = 32'b11111111111111111011000110110010;
assign LUT_4[12343] = 32'b11111111111111110100010010101010;
assign LUT_4[12344] = 32'b11111111111111110111111000000111;
assign LUT_4[12345] = 32'b11111111111111110001000011111111;
assign LUT_4[12346] = 32'b11111111111111110111010010101011;
assign LUT_4[12347] = 32'b11111111111111110000011110100011;
assign LUT_4[12348] = 32'b11111111111111110100111000100011;
assign LUT_4[12349] = 32'b11111111111111101110000100011011;
assign LUT_4[12350] = 32'b11111111111111110100010011000111;
assign LUT_4[12351] = 32'b11111111111111101101011110111111;
assign LUT_4[12352] = 32'b00000000000000000011110110010001;
assign LUT_4[12353] = 32'b11111111111111111101000010001001;
assign LUT_4[12354] = 32'b00000000000000000011010000110101;
assign LUT_4[12355] = 32'b11111111111111111100011100101101;
assign LUT_4[12356] = 32'b00000000000000000000110110101101;
assign LUT_4[12357] = 32'b11111111111111111010000010100101;
assign LUT_4[12358] = 32'b00000000000000000000010001010001;
assign LUT_4[12359] = 32'b11111111111111111001011101001001;
assign LUT_4[12360] = 32'b11111111111111111101000010100110;
assign LUT_4[12361] = 32'b11111111111111110110001110011110;
assign LUT_4[12362] = 32'b11111111111111111100011101001010;
assign LUT_4[12363] = 32'b11111111111111110101101001000010;
assign LUT_4[12364] = 32'b11111111111111111010000011000010;
assign LUT_4[12365] = 32'b11111111111111110011001110111010;
assign LUT_4[12366] = 32'b11111111111111111001011101100110;
assign LUT_4[12367] = 32'b11111111111111110010101001011110;
assign LUT_4[12368] = 32'b00000000000000000001100111111111;
assign LUT_4[12369] = 32'b11111111111111111010110011110111;
assign LUT_4[12370] = 32'b00000000000000000001000010100011;
assign LUT_4[12371] = 32'b11111111111111111010001110011011;
assign LUT_4[12372] = 32'b11111111111111111110101000011011;
assign LUT_4[12373] = 32'b11111111111111110111110100010011;
assign LUT_4[12374] = 32'b11111111111111111110000010111111;
assign LUT_4[12375] = 32'b11111111111111110111001110110111;
assign LUT_4[12376] = 32'b11111111111111111010110100010100;
assign LUT_4[12377] = 32'b11111111111111110100000000001100;
assign LUT_4[12378] = 32'b11111111111111111010001110111000;
assign LUT_4[12379] = 32'b11111111111111110011011010110000;
assign LUT_4[12380] = 32'b11111111111111110111110100110000;
assign LUT_4[12381] = 32'b11111111111111110001000000101000;
assign LUT_4[12382] = 32'b11111111111111110111001111010100;
assign LUT_4[12383] = 32'b11111111111111110000011011001100;
assign LUT_4[12384] = 32'b00000000000000000010010001011000;
assign LUT_4[12385] = 32'b11111111111111111011011101010000;
assign LUT_4[12386] = 32'b00000000000000000001101011111100;
assign LUT_4[12387] = 32'b11111111111111111010110111110100;
assign LUT_4[12388] = 32'b11111111111111111111010001110100;
assign LUT_4[12389] = 32'b11111111111111111000011101101100;
assign LUT_4[12390] = 32'b11111111111111111110101100011000;
assign LUT_4[12391] = 32'b11111111111111110111111000010000;
assign LUT_4[12392] = 32'b11111111111111111011011101101101;
assign LUT_4[12393] = 32'b11111111111111110100101001100101;
assign LUT_4[12394] = 32'b11111111111111111010111000010001;
assign LUT_4[12395] = 32'b11111111111111110100000100001001;
assign LUT_4[12396] = 32'b11111111111111111000011110001001;
assign LUT_4[12397] = 32'b11111111111111110001101010000001;
assign LUT_4[12398] = 32'b11111111111111110111111000101101;
assign LUT_4[12399] = 32'b11111111111111110001000100100101;
assign LUT_4[12400] = 32'b00000000000000000000000011000110;
assign LUT_4[12401] = 32'b11111111111111111001001110111110;
assign LUT_4[12402] = 32'b11111111111111111111011101101010;
assign LUT_4[12403] = 32'b11111111111111111000101001100010;
assign LUT_4[12404] = 32'b11111111111111111101000011100010;
assign LUT_4[12405] = 32'b11111111111111110110001111011010;
assign LUT_4[12406] = 32'b11111111111111111100011110000110;
assign LUT_4[12407] = 32'b11111111111111110101101001111110;
assign LUT_4[12408] = 32'b11111111111111111001001111011011;
assign LUT_4[12409] = 32'b11111111111111110010011011010011;
assign LUT_4[12410] = 32'b11111111111111111000101001111111;
assign LUT_4[12411] = 32'b11111111111111110001110101110111;
assign LUT_4[12412] = 32'b11111111111111110110001111110111;
assign LUT_4[12413] = 32'b11111111111111101111011011101111;
assign LUT_4[12414] = 32'b11111111111111110101101010011011;
assign LUT_4[12415] = 32'b11111111111111101110110110010011;
assign LUT_4[12416] = 32'b00000000000000000101000101000101;
assign LUT_4[12417] = 32'b11111111111111111110010000111101;
assign LUT_4[12418] = 32'b00000000000000000100011111101001;
assign LUT_4[12419] = 32'b11111111111111111101101011100001;
assign LUT_4[12420] = 32'b00000000000000000010000101100001;
assign LUT_4[12421] = 32'b11111111111111111011010001011001;
assign LUT_4[12422] = 32'b00000000000000000001100000000101;
assign LUT_4[12423] = 32'b11111111111111111010101011111101;
assign LUT_4[12424] = 32'b11111111111111111110010001011010;
assign LUT_4[12425] = 32'b11111111111111110111011101010010;
assign LUT_4[12426] = 32'b11111111111111111101101011111110;
assign LUT_4[12427] = 32'b11111111111111110110110111110110;
assign LUT_4[12428] = 32'b11111111111111111011010001110110;
assign LUT_4[12429] = 32'b11111111111111110100011101101110;
assign LUT_4[12430] = 32'b11111111111111111010101100011010;
assign LUT_4[12431] = 32'b11111111111111110011111000010010;
assign LUT_4[12432] = 32'b00000000000000000010110110110011;
assign LUT_4[12433] = 32'b11111111111111111100000010101011;
assign LUT_4[12434] = 32'b00000000000000000010010001010111;
assign LUT_4[12435] = 32'b11111111111111111011011101001111;
assign LUT_4[12436] = 32'b11111111111111111111110111001111;
assign LUT_4[12437] = 32'b11111111111111111001000011000111;
assign LUT_4[12438] = 32'b11111111111111111111010001110011;
assign LUT_4[12439] = 32'b11111111111111111000011101101011;
assign LUT_4[12440] = 32'b11111111111111111100000011001000;
assign LUT_4[12441] = 32'b11111111111111110101001111000000;
assign LUT_4[12442] = 32'b11111111111111111011011101101100;
assign LUT_4[12443] = 32'b11111111111111110100101001100100;
assign LUT_4[12444] = 32'b11111111111111111001000011100100;
assign LUT_4[12445] = 32'b11111111111111110010001111011100;
assign LUT_4[12446] = 32'b11111111111111111000011110001000;
assign LUT_4[12447] = 32'b11111111111111110001101010000000;
assign LUT_4[12448] = 32'b00000000000000000011100000001100;
assign LUT_4[12449] = 32'b11111111111111111100101100000100;
assign LUT_4[12450] = 32'b00000000000000000010111010110000;
assign LUT_4[12451] = 32'b11111111111111111100000110101000;
assign LUT_4[12452] = 32'b00000000000000000000100000101000;
assign LUT_4[12453] = 32'b11111111111111111001101100100000;
assign LUT_4[12454] = 32'b11111111111111111111111011001100;
assign LUT_4[12455] = 32'b11111111111111111001000111000100;
assign LUT_4[12456] = 32'b11111111111111111100101100100001;
assign LUT_4[12457] = 32'b11111111111111110101111000011001;
assign LUT_4[12458] = 32'b11111111111111111100000111000101;
assign LUT_4[12459] = 32'b11111111111111110101010010111101;
assign LUT_4[12460] = 32'b11111111111111111001101100111101;
assign LUT_4[12461] = 32'b11111111111111110010111000110101;
assign LUT_4[12462] = 32'b11111111111111111001000111100001;
assign LUT_4[12463] = 32'b11111111111111110010010011011001;
assign LUT_4[12464] = 32'b00000000000000000001010001111010;
assign LUT_4[12465] = 32'b11111111111111111010011101110010;
assign LUT_4[12466] = 32'b00000000000000000000101100011110;
assign LUT_4[12467] = 32'b11111111111111111001111000010110;
assign LUT_4[12468] = 32'b11111111111111111110010010010110;
assign LUT_4[12469] = 32'b11111111111111110111011110001110;
assign LUT_4[12470] = 32'b11111111111111111101101100111010;
assign LUT_4[12471] = 32'b11111111111111110110111000110010;
assign LUT_4[12472] = 32'b11111111111111111010011110001111;
assign LUT_4[12473] = 32'b11111111111111110011101010000111;
assign LUT_4[12474] = 32'b11111111111111111001111000110011;
assign LUT_4[12475] = 32'b11111111111111110011000100101011;
assign LUT_4[12476] = 32'b11111111111111110111011110101011;
assign LUT_4[12477] = 32'b11111111111111110000101010100011;
assign LUT_4[12478] = 32'b11111111111111110110111001001111;
assign LUT_4[12479] = 32'b11111111111111110000000101000111;
assign LUT_4[12480] = 32'b00000000000000000110011100011001;
assign LUT_4[12481] = 32'b11111111111111111111101000010001;
assign LUT_4[12482] = 32'b00000000000000000101110110111101;
assign LUT_4[12483] = 32'b11111111111111111111000010110101;
assign LUT_4[12484] = 32'b00000000000000000011011100110101;
assign LUT_4[12485] = 32'b11111111111111111100101000101101;
assign LUT_4[12486] = 32'b00000000000000000010110111011001;
assign LUT_4[12487] = 32'b11111111111111111100000011010001;
assign LUT_4[12488] = 32'b11111111111111111111101000101110;
assign LUT_4[12489] = 32'b11111111111111111000110100100110;
assign LUT_4[12490] = 32'b11111111111111111111000011010010;
assign LUT_4[12491] = 32'b11111111111111111000001111001010;
assign LUT_4[12492] = 32'b11111111111111111100101001001010;
assign LUT_4[12493] = 32'b11111111111111110101110101000010;
assign LUT_4[12494] = 32'b11111111111111111100000011101110;
assign LUT_4[12495] = 32'b11111111111111110101001111100110;
assign LUT_4[12496] = 32'b00000000000000000100001110000111;
assign LUT_4[12497] = 32'b11111111111111111101011001111111;
assign LUT_4[12498] = 32'b00000000000000000011101000101011;
assign LUT_4[12499] = 32'b11111111111111111100110100100011;
assign LUT_4[12500] = 32'b00000000000000000001001110100011;
assign LUT_4[12501] = 32'b11111111111111111010011010011011;
assign LUT_4[12502] = 32'b00000000000000000000101001000111;
assign LUT_4[12503] = 32'b11111111111111111001110100111111;
assign LUT_4[12504] = 32'b11111111111111111101011010011100;
assign LUT_4[12505] = 32'b11111111111111110110100110010100;
assign LUT_4[12506] = 32'b11111111111111111100110101000000;
assign LUT_4[12507] = 32'b11111111111111110110000000111000;
assign LUT_4[12508] = 32'b11111111111111111010011010111000;
assign LUT_4[12509] = 32'b11111111111111110011100110110000;
assign LUT_4[12510] = 32'b11111111111111111001110101011100;
assign LUT_4[12511] = 32'b11111111111111110011000001010100;
assign LUT_4[12512] = 32'b00000000000000000100110111100000;
assign LUT_4[12513] = 32'b11111111111111111110000011011000;
assign LUT_4[12514] = 32'b00000000000000000100010010000100;
assign LUT_4[12515] = 32'b11111111111111111101011101111100;
assign LUT_4[12516] = 32'b00000000000000000001110111111100;
assign LUT_4[12517] = 32'b11111111111111111011000011110100;
assign LUT_4[12518] = 32'b00000000000000000001010010100000;
assign LUT_4[12519] = 32'b11111111111111111010011110011000;
assign LUT_4[12520] = 32'b11111111111111111110000011110101;
assign LUT_4[12521] = 32'b11111111111111110111001111101101;
assign LUT_4[12522] = 32'b11111111111111111101011110011001;
assign LUT_4[12523] = 32'b11111111111111110110101010010001;
assign LUT_4[12524] = 32'b11111111111111111011000100010001;
assign LUT_4[12525] = 32'b11111111111111110100010000001001;
assign LUT_4[12526] = 32'b11111111111111111010011110110101;
assign LUT_4[12527] = 32'b11111111111111110011101010101101;
assign LUT_4[12528] = 32'b00000000000000000010101001001110;
assign LUT_4[12529] = 32'b11111111111111111011110101000110;
assign LUT_4[12530] = 32'b00000000000000000010000011110010;
assign LUT_4[12531] = 32'b11111111111111111011001111101010;
assign LUT_4[12532] = 32'b11111111111111111111101001101010;
assign LUT_4[12533] = 32'b11111111111111111000110101100010;
assign LUT_4[12534] = 32'b11111111111111111111000100001110;
assign LUT_4[12535] = 32'b11111111111111111000010000000110;
assign LUT_4[12536] = 32'b11111111111111111011110101100011;
assign LUT_4[12537] = 32'b11111111111111110101000001011011;
assign LUT_4[12538] = 32'b11111111111111111011010000000111;
assign LUT_4[12539] = 32'b11111111111111110100011011111111;
assign LUT_4[12540] = 32'b11111111111111111000110101111111;
assign LUT_4[12541] = 32'b11111111111111110010000001110111;
assign LUT_4[12542] = 32'b11111111111111111000010000100011;
assign LUT_4[12543] = 32'b11111111111111110001011100011011;
assign LUT_4[12544] = 32'b00000000000000000111011010100000;
assign LUT_4[12545] = 32'b00000000000000000000100110011000;
assign LUT_4[12546] = 32'b00000000000000000110110101000100;
assign LUT_4[12547] = 32'b00000000000000000000000000111100;
assign LUT_4[12548] = 32'b00000000000000000100011010111100;
assign LUT_4[12549] = 32'b11111111111111111101100110110100;
assign LUT_4[12550] = 32'b00000000000000000011110101100000;
assign LUT_4[12551] = 32'b11111111111111111101000001011000;
assign LUT_4[12552] = 32'b00000000000000000000100110110101;
assign LUT_4[12553] = 32'b11111111111111111001110010101101;
assign LUT_4[12554] = 32'b00000000000000000000000001011001;
assign LUT_4[12555] = 32'b11111111111111111001001101010001;
assign LUT_4[12556] = 32'b11111111111111111101100111010001;
assign LUT_4[12557] = 32'b11111111111111110110110011001001;
assign LUT_4[12558] = 32'b11111111111111111101000001110101;
assign LUT_4[12559] = 32'b11111111111111110110001101101101;
assign LUT_4[12560] = 32'b00000000000000000101001100001110;
assign LUT_4[12561] = 32'b11111111111111111110011000000110;
assign LUT_4[12562] = 32'b00000000000000000100100110110010;
assign LUT_4[12563] = 32'b11111111111111111101110010101010;
assign LUT_4[12564] = 32'b00000000000000000010001100101010;
assign LUT_4[12565] = 32'b11111111111111111011011000100010;
assign LUT_4[12566] = 32'b00000000000000000001100111001110;
assign LUT_4[12567] = 32'b11111111111111111010110011000110;
assign LUT_4[12568] = 32'b11111111111111111110011000100011;
assign LUT_4[12569] = 32'b11111111111111110111100100011011;
assign LUT_4[12570] = 32'b11111111111111111101110011000111;
assign LUT_4[12571] = 32'b11111111111111110110111110111111;
assign LUT_4[12572] = 32'b11111111111111111011011000111111;
assign LUT_4[12573] = 32'b11111111111111110100100100110111;
assign LUT_4[12574] = 32'b11111111111111111010110011100011;
assign LUT_4[12575] = 32'b11111111111111110011111111011011;
assign LUT_4[12576] = 32'b00000000000000000101110101100111;
assign LUT_4[12577] = 32'b11111111111111111111000001011111;
assign LUT_4[12578] = 32'b00000000000000000101010000001011;
assign LUT_4[12579] = 32'b11111111111111111110011100000011;
assign LUT_4[12580] = 32'b00000000000000000010110110000011;
assign LUT_4[12581] = 32'b11111111111111111100000001111011;
assign LUT_4[12582] = 32'b00000000000000000010010000100111;
assign LUT_4[12583] = 32'b11111111111111111011011100011111;
assign LUT_4[12584] = 32'b11111111111111111111000001111100;
assign LUT_4[12585] = 32'b11111111111111111000001101110100;
assign LUT_4[12586] = 32'b11111111111111111110011100100000;
assign LUT_4[12587] = 32'b11111111111111110111101000011000;
assign LUT_4[12588] = 32'b11111111111111111100000010011000;
assign LUT_4[12589] = 32'b11111111111111110101001110010000;
assign LUT_4[12590] = 32'b11111111111111111011011100111100;
assign LUT_4[12591] = 32'b11111111111111110100101000110100;
assign LUT_4[12592] = 32'b00000000000000000011100111010101;
assign LUT_4[12593] = 32'b11111111111111111100110011001101;
assign LUT_4[12594] = 32'b00000000000000000011000001111001;
assign LUT_4[12595] = 32'b11111111111111111100001101110001;
assign LUT_4[12596] = 32'b00000000000000000000100111110001;
assign LUT_4[12597] = 32'b11111111111111111001110011101001;
assign LUT_4[12598] = 32'b00000000000000000000000010010101;
assign LUT_4[12599] = 32'b11111111111111111001001110001101;
assign LUT_4[12600] = 32'b11111111111111111100110011101010;
assign LUT_4[12601] = 32'b11111111111111110101111111100010;
assign LUT_4[12602] = 32'b11111111111111111100001110001110;
assign LUT_4[12603] = 32'b11111111111111110101011010000110;
assign LUT_4[12604] = 32'b11111111111111111001110100000110;
assign LUT_4[12605] = 32'b11111111111111110010111111111110;
assign LUT_4[12606] = 32'b11111111111111111001001110101010;
assign LUT_4[12607] = 32'b11111111111111110010011010100010;
assign LUT_4[12608] = 32'b00000000000000001000110001110100;
assign LUT_4[12609] = 32'b00000000000000000001111101101100;
assign LUT_4[12610] = 32'b00000000000000001000001100011000;
assign LUT_4[12611] = 32'b00000000000000000001011000010000;
assign LUT_4[12612] = 32'b00000000000000000101110010010000;
assign LUT_4[12613] = 32'b11111111111111111110111110001000;
assign LUT_4[12614] = 32'b00000000000000000101001100110100;
assign LUT_4[12615] = 32'b11111111111111111110011000101100;
assign LUT_4[12616] = 32'b00000000000000000001111110001001;
assign LUT_4[12617] = 32'b11111111111111111011001010000001;
assign LUT_4[12618] = 32'b00000000000000000001011000101101;
assign LUT_4[12619] = 32'b11111111111111111010100100100101;
assign LUT_4[12620] = 32'b11111111111111111110111110100101;
assign LUT_4[12621] = 32'b11111111111111111000001010011101;
assign LUT_4[12622] = 32'b11111111111111111110011001001001;
assign LUT_4[12623] = 32'b11111111111111110111100101000001;
assign LUT_4[12624] = 32'b00000000000000000110100011100010;
assign LUT_4[12625] = 32'b11111111111111111111101111011010;
assign LUT_4[12626] = 32'b00000000000000000101111110000110;
assign LUT_4[12627] = 32'b11111111111111111111001001111110;
assign LUT_4[12628] = 32'b00000000000000000011100011111110;
assign LUT_4[12629] = 32'b11111111111111111100101111110110;
assign LUT_4[12630] = 32'b00000000000000000010111110100010;
assign LUT_4[12631] = 32'b11111111111111111100001010011010;
assign LUT_4[12632] = 32'b11111111111111111111101111110111;
assign LUT_4[12633] = 32'b11111111111111111000111011101111;
assign LUT_4[12634] = 32'b11111111111111111111001010011011;
assign LUT_4[12635] = 32'b11111111111111111000010110010011;
assign LUT_4[12636] = 32'b11111111111111111100110000010011;
assign LUT_4[12637] = 32'b11111111111111110101111100001011;
assign LUT_4[12638] = 32'b11111111111111111100001010110111;
assign LUT_4[12639] = 32'b11111111111111110101010110101111;
assign LUT_4[12640] = 32'b00000000000000000111001100111011;
assign LUT_4[12641] = 32'b00000000000000000000011000110011;
assign LUT_4[12642] = 32'b00000000000000000110100111011111;
assign LUT_4[12643] = 32'b11111111111111111111110011010111;
assign LUT_4[12644] = 32'b00000000000000000100001101010111;
assign LUT_4[12645] = 32'b11111111111111111101011001001111;
assign LUT_4[12646] = 32'b00000000000000000011100111111011;
assign LUT_4[12647] = 32'b11111111111111111100110011110011;
assign LUT_4[12648] = 32'b00000000000000000000011001010000;
assign LUT_4[12649] = 32'b11111111111111111001100101001000;
assign LUT_4[12650] = 32'b11111111111111111111110011110100;
assign LUT_4[12651] = 32'b11111111111111111000111111101100;
assign LUT_4[12652] = 32'b11111111111111111101011001101100;
assign LUT_4[12653] = 32'b11111111111111110110100101100100;
assign LUT_4[12654] = 32'b11111111111111111100110100010000;
assign LUT_4[12655] = 32'b11111111111111110110000000001000;
assign LUT_4[12656] = 32'b00000000000000000100111110101001;
assign LUT_4[12657] = 32'b11111111111111111110001010100001;
assign LUT_4[12658] = 32'b00000000000000000100011001001101;
assign LUT_4[12659] = 32'b11111111111111111101100101000101;
assign LUT_4[12660] = 32'b00000000000000000001111111000101;
assign LUT_4[12661] = 32'b11111111111111111011001010111101;
assign LUT_4[12662] = 32'b00000000000000000001011001101001;
assign LUT_4[12663] = 32'b11111111111111111010100101100001;
assign LUT_4[12664] = 32'b11111111111111111110001010111110;
assign LUT_4[12665] = 32'b11111111111111110111010110110110;
assign LUT_4[12666] = 32'b11111111111111111101100101100010;
assign LUT_4[12667] = 32'b11111111111111110110110001011010;
assign LUT_4[12668] = 32'b11111111111111111011001011011010;
assign LUT_4[12669] = 32'b11111111111111110100010111010010;
assign LUT_4[12670] = 32'b11111111111111111010100101111110;
assign LUT_4[12671] = 32'b11111111111111110011110001110110;
assign LUT_4[12672] = 32'b00000000000000001010000000101000;
assign LUT_4[12673] = 32'b00000000000000000011001100100000;
assign LUT_4[12674] = 32'b00000000000000001001011011001100;
assign LUT_4[12675] = 32'b00000000000000000010100111000100;
assign LUT_4[12676] = 32'b00000000000000000111000001000100;
assign LUT_4[12677] = 32'b00000000000000000000001100111100;
assign LUT_4[12678] = 32'b00000000000000000110011011101000;
assign LUT_4[12679] = 32'b11111111111111111111100111100000;
assign LUT_4[12680] = 32'b00000000000000000011001100111101;
assign LUT_4[12681] = 32'b11111111111111111100011000110101;
assign LUT_4[12682] = 32'b00000000000000000010100111100001;
assign LUT_4[12683] = 32'b11111111111111111011110011011001;
assign LUT_4[12684] = 32'b00000000000000000000001101011001;
assign LUT_4[12685] = 32'b11111111111111111001011001010001;
assign LUT_4[12686] = 32'b11111111111111111111100111111101;
assign LUT_4[12687] = 32'b11111111111111111000110011110101;
assign LUT_4[12688] = 32'b00000000000000000111110010010110;
assign LUT_4[12689] = 32'b00000000000000000000111110001110;
assign LUT_4[12690] = 32'b00000000000000000111001100111010;
assign LUT_4[12691] = 32'b00000000000000000000011000110010;
assign LUT_4[12692] = 32'b00000000000000000100110010110010;
assign LUT_4[12693] = 32'b11111111111111111101111110101010;
assign LUT_4[12694] = 32'b00000000000000000100001101010110;
assign LUT_4[12695] = 32'b11111111111111111101011001001110;
assign LUT_4[12696] = 32'b00000000000000000000111110101011;
assign LUT_4[12697] = 32'b11111111111111111010001010100011;
assign LUT_4[12698] = 32'b00000000000000000000011001001111;
assign LUT_4[12699] = 32'b11111111111111111001100101000111;
assign LUT_4[12700] = 32'b11111111111111111101111111000111;
assign LUT_4[12701] = 32'b11111111111111110111001010111111;
assign LUT_4[12702] = 32'b11111111111111111101011001101011;
assign LUT_4[12703] = 32'b11111111111111110110100101100011;
assign LUT_4[12704] = 32'b00000000000000001000011011101111;
assign LUT_4[12705] = 32'b00000000000000000001100111100111;
assign LUT_4[12706] = 32'b00000000000000000111110110010011;
assign LUT_4[12707] = 32'b00000000000000000001000010001011;
assign LUT_4[12708] = 32'b00000000000000000101011100001011;
assign LUT_4[12709] = 32'b11111111111111111110101000000011;
assign LUT_4[12710] = 32'b00000000000000000100110110101111;
assign LUT_4[12711] = 32'b11111111111111111110000010100111;
assign LUT_4[12712] = 32'b00000000000000000001101000000100;
assign LUT_4[12713] = 32'b11111111111111111010110011111100;
assign LUT_4[12714] = 32'b00000000000000000001000010101000;
assign LUT_4[12715] = 32'b11111111111111111010001110100000;
assign LUT_4[12716] = 32'b11111111111111111110101000100000;
assign LUT_4[12717] = 32'b11111111111111110111110100011000;
assign LUT_4[12718] = 32'b11111111111111111110000011000100;
assign LUT_4[12719] = 32'b11111111111111110111001110111100;
assign LUT_4[12720] = 32'b00000000000000000110001101011101;
assign LUT_4[12721] = 32'b11111111111111111111011001010101;
assign LUT_4[12722] = 32'b00000000000000000101101000000001;
assign LUT_4[12723] = 32'b11111111111111111110110011111001;
assign LUT_4[12724] = 32'b00000000000000000011001101111001;
assign LUT_4[12725] = 32'b11111111111111111100011001110001;
assign LUT_4[12726] = 32'b00000000000000000010101000011101;
assign LUT_4[12727] = 32'b11111111111111111011110100010101;
assign LUT_4[12728] = 32'b11111111111111111111011001110010;
assign LUT_4[12729] = 32'b11111111111111111000100101101010;
assign LUT_4[12730] = 32'b11111111111111111110110100010110;
assign LUT_4[12731] = 32'b11111111111111111000000000001110;
assign LUT_4[12732] = 32'b11111111111111111100011010001110;
assign LUT_4[12733] = 32'b11111111111111110101100110000110;
assign LUT_4[12734] = 32'b11111111111111111011110100110010;
assign LUT_4[12735] = 32'b11111111111111110101000000101010;
assign LUT_4[12736] = 32'b00000000000000001011010111111100;
assign LUT_4[12737] = 32'b00000000000000000100100011110100;
assign LUT_4[12738] = 32'b00000000000000001010110010100000;
assign LUT_4[12739] = 32'b00000000000000000011111110011000;
assign LUT_4[12740] = 32'b00000000000000001000011000011000;
assign LUT_4[12741] = 32'b00000000000000000001100100010000;
assign LUT_4[12742] = 32'b00000000000000000111110010111100;
assign LUT_4[12743] = 32'b00000000000000000000111110110100;
assign LUT_4[12744] = 32'b00000000000000000100100100010001;
assign LUT_4[12745] = 32'b11111111111111111101110000001001;
assign LUT_4[12746] = 32'b00000000000000000011111110110101;
assign LUT_4[12747] = 32'b11111111111111111101001010101101;
assign LUT_4[12748] = 32'b00000000000000000001100100101101;
assign LUT_4[12749] = 32'b11111111111111111010110000100101;
assign LUT_4[12750] = 32'b00000000000000000000111111010001;
assign LUT_4[12751] = 32'b11111111111111111010001011001001;
assign LUT_4[12752] = 32'b00000000000000001001001001101010;
assign LUT_4[12753] = 32'b00000000000000000010010101100010;
assign LUT_4[12754] = 32'b00000000000000001000100100001110;
assign LUT_4[12755] = 32'b00000000000000000001110000000110;
assign LUT_4[12756] = 32'b00000000000000000110001010000110;
assign LUT_4[12757] = 32'b11111111111111111111010101111110;
assign LUT_4[12758] = 32'b00000000000000000101100100101010;
assign LUT_4[12759] = 32'b11111111111111111110110000100010;
assign LUT_4[12760] = 32'b00000000000000000010010101111111;
assign LUT_4[12761] = 32'b11111111111111111011100001110111;
assign LUT_4[12762] = 32'b00000000000000000001110000100011;
assign LUT_4[12763] = 32'b11111111111111111010111100011011;
assign LUT_4[12764] = 32'b11111111111111111111010110011011;
assign LUT_4[12765] = 32'b11111111111111111000100010010011;
assign LUT_4[12766] = 32'b11111111111111111110110000111111;
assign LUT_4[12767] = 32'b11111111111111110111111100110111;
assign LUT_4[12768] = 32'b00000000000000001001110011000011;
assign LUT_4[12769] = 32'b00000000000000000010111110111011;
assign LUT_4[12770] = 32'b00000000000000001001001101100111;
assign LUT_4[12771] = 32'b00000000000000000010011001011111;
assign LUT_4[12772] = 32'b00000000000000000110110011011111;
assign LUT_4[12773] = 32'b11111111111111111111111111010111;
assign LUT_4[12774] = 32'b00000000000000000110001110000011;
assign LUT_4[12775] = 32'b11111111111111111111011001111011;
assign LUT_4[12776] = 32'b00000000000000000010111111011000;
assign LUT_4[12777] = 32'b11111111111111111100001011010000;
assign LUT_4[12778] = 32'b00000000000000000010011001111100;
assign LUT_4[12779] = 32'b11111111111111111011100101110100;
assign LUT_4[12780] = 32'b11111111111111111111111111110100;
assign LUT_4[12781] = 32'b11111111111111111001001011101100;
assign LUT_4[12782] = 32'b11111111111111111111011010011000;
assign LUT_4[12783] = 32'b11111111111111111000100110010000;
assign LUT_4[12784] = 32'b00000000000000000111100100110001;
assign LUT_4[12785] = 32'b00000000000000000000110000101001;
assign LUT_4[12786] = 32'b00000000000000000110111111010101;
assign LUT_4[12787] = 32'b00000000000000000000001011001101;
assign LUT_4[12788] = 32'b00000000000000000100100101001101;
assign LUT_4[12789] = 32'b11111111111111111101110001000101;
assign LUT_4[12790] = 32'b00000000000000000011111111110001;
assign LUT_4[12791] = 32'b11111111111111111101001011101001;
assign LUT_4[12792] = 32'b00000000000000000000110001000110;
assign LUT_4[12793] = 32'b11111111111111111001111100111110;
assign LUT_4[12794] = 32'b00000000000000000000001011101010;
assign LUT_4[12795] = 32'b11111111111111111001010111100010;
assign LUT_4[12796] = 32'b11111111111111111101110001100010;
assign LUT_4[12797] = 32'b11111111111111110110111101011010;
assign LUT_4[12798] = 32'b11111111111111111101001100000110;
assign LUT_4[12799] = 32'b11111111111111110110010111111110;
assign LUT_4[12800] = 32'b00000000000000000001100011000101;
assign LUT_4[12801] = 32'b11111111111111111010101110111101;
assign LUT_4[12802] = 32'b00000000000000000000111101101001;
assign LUT_4[12803] = 32'b11111111111111111010001001100001;
assign LUT_4[12804] = 32'b11111111111111111110100011100001;
assign LUT_4[12805] = 32'b11111111111111110111101111011001;
assign LUT_4[12806] = 32'b11111111111111111101111110000101;
assign LUT_4[12807] = 32'b11111111111111110111001001111101;
assign LUT_4[12808] = 32'b11111111111111111010101111011010;
assign LUT_4[12809] = 32'b11111111111111110011111011010010;
assign LUT_4[12810] = 32'b11111111111111111010001001111110;
assign LUT_4[12811] = 32'b11111111111111110011010101110110;
assign LUT_4[12812] = 32'b11111111111111110111101111110110;
assign LUT_4[12813] = 32'b11111111111111110000111011101110;
assign LUT_4[12814] = 32'b11111111111111110111001010011010;
assign LUT_4[12815] = 32'b11111111111111110000010110010010;
assign LUT_4[12816] = 32'b11111111111111111111010100110011;
assign LUT_4[12817] = 32'b11111111111111111000100000101011;
assign LUT_4[12818] = 32'b11111111111111111110101111010111;
assign LUT_4[12819] = 32'b11111111111111110111111011001111;
assign LUT_4[12820] = 32'b11111111111111111100010101001111;
assign LUT_4[12821] = 32'b11111111111111110101100001000111;
assign LUT_4[12822] = 32'b11111111111111111011101111110011;
assign LUT_4[12823] = 32'b11111111111111110100111011101011;
assign LUT_4[12824] = 32'b11111111111111111000100001001000;
assign LUT_4[12825] = 32'b11111111111111110001101101000000;
assign LUT_4[12826] = 32'b11111111111111110111111011101100;
assign LUT_4[12827] = 32'b11111111111111110001000111100100;
assign LUT_4[12828] = 32'b11111111111111110101100001100100;
assign LUT_4[12829] = 32'b11111111111111101110101101011100;
assign LUT_4[12830] = 32'b11111111111111110100111100001000;
assign LUT_4[12831] = 32'b11111111111111101110001000000000;
assign LUT_4[12832] = 32'b11111111111111111111111110001100;
assign LUT_4[12833] = 32'b11111111111111111001001010000100;
assign LUT_4[12834] = 32'b11111111111111111111011000110000;
assign LUT_4[12835] = 32'b11111111111111111000100100101000;
assign LUT_4[12836] = 32'b11111111111111111100111110101000;
assign LUT_4[12837] = 32'b11111111111111110110001010100000;
assign LUT_4[12838] = 32'b11111111111111111100011001001100;
assign LUT_4[12839] = 32'b11111111111111110101100101000100;
assign LUT_4[12840] = 32'b11111111111111111001001010100001;
assign LUT_4[12841] = 32'b11111111111111110010010110011001;
assign LUT_4[12842] = 32'b11111111111111111000100101000101;
assign LUT_4[12843] = 32'b11111111111111110001110000111101;
assign LUT_4[12844] = 32'b11111111111111110110001010111101;
assign LUT_4[12845] = 32'b11111111111111101111010110110101;
assign LUT_4[12846] = 32'b11111111111111110101100101100001;
assign LUT_4[12847] = 32'b11111111111111101110110001011001;
assign LUT_4[12848] = 32'b11111111111111111101101111111010;
assign LUT_4[12849] = 32'b11111111111111110110111011110010;
assign LUT_4[12850] = 32'b11111111111111111101001010011110;
assign LUT_4[12851] = 32'b11111111111111110110010110010110;
assign LUT_4[12852] = 32'b11111111111111111010110000010110;
assign LUT_4[12853] = 32'b11111111111111110011111100001110;
assign LUT_4[12854] = 32'b11111111111111111010001010111010;
assign LUT_4[12855] = 32'b11111111111111110011010110110010;
assign LUT_4[12856] = 32'b11111111111111110110111100001111;
assign LUT_4[12857] = 32'b11111111111111110000001000000111;
assign LUT_4[12858] = 32'b11111111111111110110010110110011;
assign LUT_4[12859] = 32'b11111111111111101111100010101011;
assign LUT_4[12860] = 32'b11111111111111110011111100101011;
assign LUT_4[12861] = 32'b11111111111111101101001000100011;
assign LUT_4[12862] = 32'b11111111111111110011010111001111;
assign LUT_4[12863] = 32'b11111111111111101100100011000111;
assign LUT_4[12864] = 32'b00000000000000000010111010011001;
assign LUT_4[12865] = 32'b11111111111111111100000110010001;
assign LUT_4[12866] = 32'b00000000000000000010010100111101;
assign LUT_4[12867] = 32'b11111111111111111011100000110101;
assign LUT_4[12868] = 32'b11111111111111111111111010110101;
assign LUT_4[12869] = 32'b11111111111111111001000110101101;
assign LUT_4[12870] = 32'b11111111111111111111010101011001;
assign LUT_4[12871] = 32'b11111111111111111000100001010001;
assign LUT_4[12872] = 32'b11111111111111111100000110101110;
assign LUT_4[12873] = 32'b11111111111111110101010010100110;
assign LUT_4[12874] = 32'b11111111111111111011100001010010;
assign LUT_4[12875] = 32'b11111111111111110100101101001010;
assign LUT_4[12876] = 32'b11111111111111111001000111001010;
assign LUT_4[12877] = 32'b11111111111111110010010011000010;
assign LUT_4[12878] = 32'b11111111111111111000100001101110;
assign LUT_4[12879] = 32'b11111111111111110001101101100110;
assign LUT_4[12880] = 32'b00000000000000000000101100000111;
assign LUT_4[12881] = 32'b11111111111111111001110111111111;
assign LUT_4[12882] = 32'b00000000000000000000000110101011;
assign LUT_4[12883] = 32'b11111111111111111001010010100011;
assign LUT_4[12884] = 32'b11111111111111111101101100100011;
assign LUT_4[12885] = 32'b11111111111111110110111000011011;
assign LUT_4[12886] = 32'b11111111111111111101000111000111;
assign LUT_4[12887] = 32'b11111111111111110110010010111111;
assign LUT_4[12888] = 32'b11111111111111111001111000011100;
assign LUT_4[12889] = 32'b11111111111111110011000100010100;
assign LUT_4[12890] = 32'b11111111111111111001010011000000;
assign LUT_4[12891] = 32'b11111111111111110010011110111000;
assign LUT_4[12892] = 32'b11111111111111110110111000111000;
assign LUT_4[12893] = 32'b11111111111111110000000100110000;
assign LUT_4[12894] = 32'b11111111111111110110010011011100;
assign LUT_4[12895] = 32'b11111111111111101111011111010100;
assign LUT_4[12896] = 32'b00000000000000000001010101100000;
assign LUT_4[12897] = 32'b11111111111111111010100001011000;
assign LUT_4[12898] = 32'b00000000000000000000110000000100;
assign LUT_4[12899] = 32'b11111111111111111001111011111100;
assign LUT_4[12900] = 32'b11111111111111111110010101111100;
assign LUT_4[12901] = 32'b11111111111111110111100001110100;
assign LUT_4[12902] = 32'b11111111111111111101110000100000;
assign LUT_4[12903] = 32'b11111111111111110110111100011000;
assign LUT_4[12904] = 32'b11111111111111111010100001110101;
assign LUT_4[12905] = 32'b11111111111111110011101101101101;
assign LUT_4[12906] = 32'b11111111111111111001111100011001;
assign LUT_4[12907] = 32'b11111111111111110011001000010001;
assign LUT_4[12908] = 32'b11111111111111110111100010010001;
assign LUT_4[12909] = 32'b11111111111111110000101110001001;
assign LUT_4[12910] = 32'b11111111111111110110111100110101;
assign LUT_4[12911] = 32'b11111111111111110000001000101101;
assign LUT_4[12912] = 32'b11111111111111111111000111001110;
assign LUT_4[12913] = 32'b11111111111111111000010011000110;
assign LUT_4[12914] = 32'b11111111111111111110100001110010;
assign LUT_4[12915] = 32'b11111111111111110111101101101010;
assign LUT_4[12916] = 32'b11111111111111111100000111101010;
assign LUT_4[12917] = 32'b11111111111111110101010011100010;
assign LUT_4[12918] = 32'b11111111111111111011100010001110;
assign LUT_4[12919] = 32'b11111111111111110100101110000110;
assign LUT_4[12920] = 32'b11111111111111111000010011100011;
assign LUT_4[12921] = 32'b11111111111111110001011111011011;
assign LUT_4[12922] = 32'b11111111111111110111101110000111;
assign LUT_4[12923] = 32'b11111111111111110000111001111111;
assign LUT_4[12924] = 32'b11111111111111110101010011111111;
assign LUT_4[12925] = 32'b11111111111111101110011111110111;
assign LUT_4[12926] = 32'b11111111111111110100101110100011;
assign LUT_4[12927] = 32'b11111111111111101101111010011011;
assign LUT_4[12928] = 32'b00000000000000000100001001001101;
assign LUT_4[12929] = 32'b11111111111111111101010101000101;
assign LUT_4[12930] = 32'b00000000000000000011100011110001;
assign LUT_4[12931] = 32'b11111111111111111100101111101001;
assign LUT_4[12932] = 32'b00000000000000000001001001101001;
assign LUT_4[12933] = 32'b11111111111111111010010101100001;
assign LUT_4[12934] = 32'b00000000000000000000100100001101;
assign LUT_4[12935] = 32'b11111111111111111001110000000101;
assign LUT_4[12936] = 32'b11111111111111111101010101100010;
assign LUT_4[12937] = 32'b11111111111111110110100001011010;
assign LUT_4[12938] = 32'b11111111111111111100110000000110;
assign LUT_4[12939] = 32'b11111111111111110101111011111110;
assign LUT_4[12940] = 32'b11111111111111111010010101111110;
assign LUT_4[12941] = 32'b11111111111111110011100001110110;
assign LUT_4[12942] = 32'b11111111111111111001110000100010;
assign LUT_4[12943] = 32'b11111111111111110010111100011010;
assign LUT_4[12944] = 32'b00000000000000000001111010111011;
assign LUT_4[12945] = 32'b11111111111111111011000110110011;
assign LUT_4[12946] = 32'b00000000000000000001010101011111;
assign LUT_4[12947] = 32'b11111111111111111010100001010111;
assign LUT_4[12948] = 32'b11111111111111111110111011010111;
assign LUT_4[12949] = 32'b11111111111111111000000111001111;
assign LUT_4[12950] = 32'b11111111111111111110010101111011;
assign LUT_4[12951] = 32'b11111111111111110111100001110011;
assign LUT_4[12952] = 32'b11111111111111111011000111010000;
assign LUT_4[12953] = 32'b11111111111111110100010011001000;
assign LUT_4[12954] = 32'b11111111111111111010100001110100;
assign LUT_4[12955] = 32'b11111111111111110011101101101100;
assign LUT_4[12956] = 32'b11111111111111111000000111101100;
assign LUT_4[12957] = 32'b11111111111111110001010011100100;
assign LUT_4[12958] = 32'b11111111111111110111100010010000;
assign LUT_4[12959] = 32'b11111111111111110000101110001000;
assign LUT_4[12960] = 32'b00000000000000000010100100010100;
assign LUT_4[12961] = 32'b11111111111111111011110000001100;
assign LUT_4[12962] = 32'b00000000000000000001111110111000;
assign LUT_4[12963] = 32'b11111111111111111011001010110000;
assign LUT_4[12964] = 32'b11111111111111111111100100110000;
assign LUT_4[12965] = 32'b11111111111111111000110000101000;
assign LUT_4[12966] = 32'b11111111111111111110111111010100;
assign LUT_4[12967] = 32'b11111111111111111000001011001100;
assign LUT_4[12968] = 32'b11111111111111111011110000101001;
assign LUT_4[12969] = 32'b11111111111111110100111100100001;
assign LUT_4[12970] = 32'b11111111111111111011001011001101;
assign LUT_4[12971] = 32'b11111111111111110100010111000101;
assign LUT_4[12972] = 32'b11111111111111111000110001000101;
assign LUT_4[12973] = 32'b11111111111111110001111100111101;
assign LUT_4[12974] = 32'b11111111111111111000001011101001;
assign LUT_4[12975] = 32'b11111111111111110001010111100001;
assign LUT_4[12976] = 32'b00000000000000000000010110000010;
assign LUT_4[12977] = 32'b11111111111111111001100001111010;
assign LUT_4[12978] = 32'b11111111111111111111110000100110;
assign LUT_4[12979] = 32'b11111111111111111000111100011110;
assign LUT_4[12980] = 32'b11111111111111111101010110011110;
assign LUT_4[12981] = 32'b11111111111111110110100010010110;
assign LUT_4[12982] = 32'b11111111111111111100110001000010;
assign LUT_4[12983] = 32'b11111111111111110101111100111010;
assign LUT_4[12984] = 32'b11111111111111111001100010010111;
assign LUT_4[12985] = 32'b11111111111111110010101110001111;
assign LUT_4[12986] = 32'b11111111111111111000111100111011;
assign LUT_4[12987] = 32'b11111111111111110010001000110011;
assign LUT_4[12988] = 32'b11111111111111110110100010110011;
assign LUT_4[12989] = 32'b11111111111111101111101110101011;
assign LUT_4[12990] = 32'b11111111111111110101111101010111;
assign LUT_4[12991] = 32'b11111111111111101111001001001111;
assign LUT_4[12992] = 32'b00000000000000000101100000100001;
assign LUT_4[12993] = 32'b11111111111111111110101100011001;
assign LUT_4[12994] = 32'b00000000000000000100111011000101;
assign LUT_4[12995] = 32'b11111111111111111110000110111101;
assign LUT_4[12996] = 32'b00000000000000000010100000111101;
assign LUT_4[12997] = 32'b11111111111111111011101100110101;
assign LUT_4[12998] = 32'b00000000000000000001111011100001;
assign LUT_4[12999] = 32'b11111111111111111011000111011001;
assign LUT_4[13000] = 32'b11111111111111111110101100110110;
assign LUT_4[13001] = 32'b11111111111111110111111000101110;
assign LUT_4[13002] = 32'b11111111111111111110000111011010;
assign LUT_4[13003] = 32'b11111111111111110111010011010010;
assign LUT_4[13004] = 32'b11111111111111111011101101010010;
assign LUT_4[13005] = 32'b11111111111111110100111001001010;
assign LUT_4[13006] = 32'b11111111111111111011000111110110;
assign LUT_4[13007] = 32'b11111111111111110100010011101110;
assign LUT_4[13008] = 32'b00000000000000000011010010001111;
assign LUT_4[13009] = 32'b11111111111111111100011110000111;
assign LUT_4[13010] = 32'b00000000000000000010101100110011;
assign LUT_4[13011] = 32'b11111111111111111011111000101011;
assign LUT_4[13012] = 32'b00000000000000000000010010101011;
assign LUT_4[13013] = 32'b11111111111111111001011110100011;
assign LUT_4[13014] = 32'b11111111111111111111101101001111;
assign LUT_4[13015] = 32'b11111111111111111000111001000111;
assign LUT_4[13016] = 32'b11111111111111111100011110100100;
assign LUT_4[13017] = 32'b11111111111111110101101010011100;
assign LUT_4[13018] = 32'b11111111111111111011111001001000;
assign LUT_4[13019] = 32'b11111111111111110101000101000000;
assign LUT_4[13020] = 32'b11111111111111111001011111000000;
assign LUT_4[13021] = 32'b11111111111111110010101010111000;
assign LUT_4[13022] = 32'b11111111111111111000111001100100;
assign LUT_4[13023] = 32'b11111111111111110010000101011100;
assign LUT_4[13024] = 32'b00000000000000000011111011101000;
assign LUT_4[13025] = 32'b11111111111111111101000111100000;
assign LUT_4[13026] = 32'b00000000000000000011010110001100;
assign LUT_4[13027] = 32'b11111111111111111100100010000100;
assign LUT_4[13028] = 32'b00000000000000000000111100000100;
assign LUT_4[13029] = 32'b11111111111111111010000111111100;
assign LUT_4[13030] = 32'b00000000000000000000010110101000;
assign LUT_4[13031] = 32'b11111111111111111001100010100000;
assign LUT_4[13032] = 32'b11111111111111111101000111111101;
assign LUT_4[13033] = 32'b11111111111111110110010011110101;
assign LUT_4[13034] = 32'b11111111111111111100100010100001;
assign LUT_4[13035] = 32'b11111111111111110101101110011001;
assign LUT_4[13036] = 32'b11111111111111111010001000011001;
assign LUT_4[13037] = 32'b11111111111111110011010100010001;
assign LUT_4[13038] = 32'b11111111111111111001100010111101;
assign LUT_4[13039] = 32'b11111111111111110010101110110101;
assign LUT_4[13040] = 32'b00000000000000000001101101010110;
assign LUT_4[13041] = 32'b11111111111111111010111001001110;
assign LUT_4[13042] = 32'b00000000000000000001000111111010;
assign LUT_4[13043] = 32'b11111111111111111010010011110010;
assign LUT_4[13044] = 32'b11111111111111111110101101110010;
assign LUT_4[13045] = 32'b11111111111111110111111001101010;
assign LUT_4[13046] = 32'b11111111111111111110001000010110;
assign LUT_4[13047] = 32'b11111111111111110111010100001110;
assign LUT_4[13048] = 32'b11111111111111111010111001101011;
assign LUT_4[13049] = 32'b11111111111111110100000101100011;
assign LUT_4[13050] = 32'b11111111111111111010010100001111;
assign LUT_4[13051] = 32'b11111111111111110011100000000111;
assign LUT_4[13052] = 32'b11111111111111110111111010000111;
assign LUT_4[13053] = 32'b11111111111111110001000101111111;
assign LUT_4[13054] = 32'b11111111111111110111010100101011;
assign LUT_4[13055] = 32'b11111111111111110000100000100011;
assign LUT_4[13056] = 32'b00000000000000000110011110101000;
assign LUT_4[13057] = 32'b11111111111111111111101010100000;
assign LUT_4[13058] = 32'b00000000000000000101111001001100;
assign LUT_4[13059] = 32'b11111111111111111111000101000100;
assign LUT_4[13060] = 32'b00000000000000000011011111000100;
assign LUT_4[13061] = 32'b11111111111111111100101010111100;
assign LUT_4[13062] = 32'b00000000000000000010111001101000;
assign LUT_4[13063] = 32'b11111111111111111100000101100000;
assign LUT_4[13064] = 32'b11111111111111111111101010111101;
assign LUT_4[13065] = 32'b11111111111111111000110110110101;
assign LUT_4[13066] = 32'b11111111111111111111000101100001;
assign LUT_4[13067] = 32'b11111111111111111000010001011001;
assign LUT_4[13068] = 32'b11111111111111111100101011011001;
assign LUT_4[13069] = 32'b11111111111111110101110111010001;
assign LUT_4[13070] = 32'b11111111111111111100000101111101;
assign LUT_4[13071] = 32'b11111111111111110101010001110101;
assign LUT_4[13072] = 32'b00000000000000000100010000010110;
assign LUT_4[13073] = 32'b11111111111111111101011100001110;
assign LUT_4[13074] = 32'b00000000000000000011101010111010;
assign LUT_4[13075] = 32'b11111111111111111100110110110010;
assign LUT_4[13076] = 32'b00000000000000000001010000110010;
assign LUT_4[13077] = 32'b11111111111111111010011100101010;
assign LUT_4[13078] = 32'b00000000000000000000101011010110;
assign LUT_4[13079] = 32'b11111111111111111001110111001110;
assign LUT_4[13080] = 32'b11111111111111111101011100101011;
assign LUT_4[13081] = 32'b11111111111111110110101000100011;
assign LUT_4[13082] = 32'b11111111111111111100110111001111;
assign LUT_4[13083] = 32'b11111111111111110110000011000111;
assign LUT_4[13084] = 32'b11111111111111111010011101000111;
assign LUT_4[13085] = 32'b11111111111111110011101000111111;
assign LUT_4[13086] = 32'b11111111111111111001110111101011;
assign LUT_4[13087] = 32'b11111111111111110011000011100011;
assign LUT_4[13088] = 32'b00000000000000000100111001101111;
assign LUT_4[13089] = 32'b11111111111111111110000101100111;
assign LUT_4[13090] = 32'b00000000000000000100010100010011;
assign LUT_4[13091] = 32'b11111111111111111101100000001011;
assign LUT_4[13092] = 32'b00000000000000000001111010001011;
assign LUT_4[13093] = 32'b11111111111111111011000110000011;
assign LUT_4[13094] = 32'b00000000000000000001010100101111;
assign LUT_4[13095] = 32'b11111111111111111010100000100111;
assign LUT_4[13096] = 32'b11111111111111111110000110000100;
assign LUT_4[13097] = 32'b11111111111111110111010001111100;
assign LUT_4[13098] = 32'b11111111111111111101100000101000;
assign LUT_4[13099] = 32'b11111111111111110110101100100000;
assign LUT_4[13100] = 32'b11111111111111111011000110100000;
assign LUT_4[13101] = 32'b11111111111111110100010010011000;
assign LUT_4[13102] = 32'b11111111111111111010100001000100;
assign LUT_4[13103] = 32'b11111111111111110011101100111100;
assign LUT_4[13104] = 32'b00000000000000000010101011011101;
assign LUT_4[13105] = 32'b11111111111111111011110111010101;
assign LUT_4[13106] = 32'b00000000000000000010000110000001;
assign LUT_4[13107] = 32'b11111111111111111011010001111001;
assign LUT_4[13108] = 32'b11111111111111111111101011111001;
assign LUT_4[13109] = 32'b11111111111111111000110111110001;
assign LUT_4[13110] = 32'b11111111111111111111000110011101;
assign LUT_4[13111] = 32'b11111111111111111000010010010101;
assign LUT_4[13112] = 32'b11111111111111111011110111110010;
assign LUT_4[13113] = 32'b11111111111111110101000011101010;
assign LUT_4[13114] = 32'b11111111111111111011010010010110;
assign LUT_4[13115] = 32'b11111111111111110100011110001110;
assign LUT_4[13116] = 32'b11111111111111111000111000001110;
assign LUT_4[13117] = 32'b11111111111111110010000100000110;
assign LUT_4[13118] = 32'b11111111111111111000010010110010;
assign LUT_4[13119] = 32'b11111111111111110001011110101010;
assign LUT_4[13120] = 32'b00000000000000000111110101111100;
assign LUT_4[13121] = 32'b00000000000000000001000001110100;
assign LUT_4[13122] = 32'b00000000000000000111010000100000;
assign LUT_4[13123] = 32'b00000000000000000000011100011000;
assign LUT_4[13124] = 32'b00000000000000000100110110011000;
assign LUT_4[13125] = 32'b11111111111111111110000010010000;
assign LUT_4[13126] = 32'b00000000000000000100010000111100;
assign LUT_4[13127] = 32'b11111111111111111101011100110100;
assign LUT_4[13128] = 32'b00000000000000000001000010010001;
assign LUT_4[13129] = 32'b11111111111111111010001110001001;
assign LUT_4[13130] = 32'b00000000000000000000011100110101;
assign LUT_4[13131] = 32'b11111111111111111001101000101101;
assign LUT_4[13132] = 32'b11111111111111111110000010101101;
assign LUT_4[13133] = 32'b11111111111111110111001110100101;
assign LUT_4[13134] = 32'b11111111111111111101011101010001;
assign LUT_4[13135] = 32'b11111111111111110110101001001001;
assign LUT_4[13136] = 32'b00000000000000000101100111101010;
assign LUT_4[13137] = 32'b11111111111111111110110011100010;
assign LUT_4[13138] = 32'b00000000000000000101000010001110;
assign LUT_4[13139] = 32'b11111111111111111110001110000110;
assign LUT_4[13140] = 32'b00000000000000000010101000000110;
assign LUT_4[13141] = 32'b11111111111111111011110011111110;
assign LUT_4[13142] = 32'b00000000000000000010000010101010;
assign LUT_4[13143] = 32'b11111111111111111011001110100010;
assign LUT_4[13144] = 32'b11111111111111111110110011111111;
assign LUT_4[13145] = 32'b11111111111111110111111111110111;
assign LUT_4[13146] = 32'b11111111111111111110001110100011;
assign LUT_4[13147] = 32'b11111111111111110111011010011011;
assign LUT_4[13148] = 32'b11111111111111111011110100011011;
assign LUT_4[13149] = 32'b11111111111111110101000000010011;
assign LUT_4[13150] = 32'b11111111111111111011001110111111;
assign LUT_4[13151] = 32'b11111111111111110100011010110111;
assign LUT_4[13152] = 32'b00000000000000000110010001000011;
assign LUT_4[13153] = 32'b11111111111111111111011100111011;
assign LUT_4[13154] = 32'b00000000000000000101101011100111;
assign LUT_4[13155] = 32'b11111111111111111110110111011111;
assign LUT_4[13156] = 32'b00000000000000000011010001011111;
assign LUT_4[13157] = 32'b11111111111111111100011101010111;
assign LUT_4[13158] = 32'b00000000000000000010101100000011;
assign LUT_4[13159] = 32'b11111111111111111011110111111011;
assign LUT_4[13160] = 32'b11111111111111111111011101011000;
assign LUT_4[13161] = 32'b11111111111111111000101001010000;
assign LUT_4[13162] = 32'b11111111111111111110110111111100;
assign LUT_4[13163] = 32'b11111111111111111000000011110100;
assign LUT_4[13164] = 32'b11111111111111111100011101110100;
assign LUT_4[13165] = 32'b11111111111111110101101001101100;
assign LUT_4[13166] = 32'b11111111111111111011111000011000;
assign LUT_4[13167] = 32'b11111111111111110101000100010000;
assign LUT_4[13168] = 32'b00000000000000000100000010110001;
assign LUT_4[13169] = 32'b11111111111111111101001110101001;
assign LUT_4[13170] = 32'b00000000000000000011011101010101;
assign LUT_4[13171] = 32'b11111111111111111100101001001101;
assign LUT_4[13172] = 32'b00000000000000000001000011001101;
assign LUT_4[13173] = 32'b11111111111111111010001111000101;
assign LUT_4[13174] = 32'b00000000000000000000011101110001;
assign LUT_4[13175] = 32'b11111111111111111001101001101001;
assign LUT_4[13176] = 32'b11111111111111111101001111000110;
assign LUT_4[13177] = 32'b11111111111111110110011010111110;
assign LUT_4[13178] = 32'b11111111111111111100101001101010;
assign LUT_4[13179] = 32'b11111111111111110101110101100010;
assign LUT_4[13180] = 32'b11111111111111111010001111100010;
assign LUT_4[13181] = 32'b11111111111111110011011011011010;
assign LUT_4[13182] = 32'b11111111111111111001101010000110;
assign LUT_4[13183] = 32'b11111111111111110010110101111110;
assign LUT_4[13184] = 32'b00000000000000001001000100110000;
assign LUT_4[13185] = 32'b00000000000000000010010000101000;
assign LUT_4[13186] = 32'b00000000000000001000011111010100;
assign LUT_4[13187] = 32'b00000000000000000001101011001100;
assign LUT_4[13188] = 32'b00000000000000000110000101001100;
assign LUT_4[13189] = 32'b11111111111111111111010001000100;
assign LUT_4[13190] = 32'b00000000000000000101011111110000;
assign LUT_4[13191] = 32'b11111111111111111110101011101000;
assign LUT_4[13192] = 32'b00000000000000000010010001000101;
assign LUT_4[13193] = 32'b11111111111111111011011100111101;
assign LUT_4[13194] = 32'b00000000000000000001101011101001;
assign LUT_4[13195] = 32'b11111111111111111010110111100001;
assign LUT_4[13196] = 32'b11111111111111111111010001100001;
assign LUT_4[13197] = 32'b11111111111111111000011101011001;
assign LUT_4[13198] = 32'b11111111111111111110101100000101;
assign LUT_4[13199] = 32'b11111111111111110111110111111101;
assign LUT_4[13200] = 32'b00000000000000000110110110011110;
assign LUT_4[13201] = 32'b00000000000000000000000010010110;
assign LUT_4[13202] = 32'b00000000000000000110010001000010;
assign LUT_4[13203] = 32'b11111111111111111111011100111010;
assign LUT_4[13204] = 32'b00000000000000000011110110111010;
assign LUT_4[13205] = 32'b11111111111111111101000010110010;
assign LUT_4[13206] = 32'b00000000000000000011010001011110;
assign LUT_4[13207] = 32'b11111111111111111100011101010110;
assign LUT_4[13208] = 32'b00000000000000000000000010110011;
assign LUT_4[13209] = 32'b11111111111111111001001110101011;
assign LUT_4[13210] = 32'b11111111111111111111011101010111;
assign LUT_4[13211] = 32'b11111111111111111000101001001111;
assign LUT_4[13212] = 32'b11111111111111111101000011001111;
assign LUT_4[13213] = 32'b11111111111111110110001111000111;
assign LUT_4[13214] = 32'b11111111111111111100011101110011;
assign LUT_4[13215] = 32'b11111111111111110101101001101011;
assign LUT_4[13216] = 32'b00000000000000000111011111110111;
assign LUT_4[13217] = 32'b00000000000000000000101011101111;
assign LUT_4[13218] = 32'b00000000000000000110111010011011;
assign LUT_4[13219] = 32'b00000000000000000000000110010011;
assign LUT_4[13220] = 32'b00000000000000000100100000010011;
assign LUT_4[13221] = 32'b11111111111111111101101100001011;
assign LUT_4[13222] = 32'b00000000000000000011111010110111;
assign LUT_4[13223] = 32'b11111111111111111101000110101111;
assign LUT_4[13224] = 32'b00000000000000000000101100001100;
assign LUT_4[13225] = 32'b11111111111111111001111000000100;
assign LUT_4[13226] = 32'b00000000000000000000000110110000;
assign LUT_4[13227] = 32'b11111111111111111001010010101000;
assign LUT_4[13228] = 32'b11111111111111111101101100101000;
assign LUT_4[13229] = 32'b11111111111111110110111000100000;
assign LUT_4[13230] = 32'b11111111111111111101000111001100;
assign LUT_4[13231] = 32'b11111111111111110110010011000100;
assign LUT_4[13232] = 32'b00000000000000000101010001100101;
assign LUT_4[13233] = 32'b11111111111111111110011101011101;
assign LUT_4[13234] = 32'b00000000000000000100101100001001;
assign LUT_4[13235] = 32'b11111111111111111101111000000001;
assign LUT_4[13236] = 32'b00000000000000000010010010000001;
assign LUT_4[13237] = 32'b11111111111111111011011101111001;
assign LUT_4[13238] = 32'b00000000000000000001101100100101;
assign LUT_4[13239] = 32'b11111111111111111010111000011101;
assign LUT_4[13240] = 32'b11111111111111111110011101111010;
assign LUT_4[13241] = 32'b11111111111111110111101001110010;
assign LUT_4[13242] = 32'b11111111111111111101111000011110;
assign LUT_4[13243] = 32'b11111111111111110111000100010110;
assign LUT_4[13244] = 32'b11111111111111111011011110010110;
assign LUT_4[13245] = 32'b11111111111111110100101010001110;
assign LUT_4[13246] = 32'b11111111111111111010111000111010;
assign LUT_4[13247] = 32'b11111111111111110100000100110010;
assign LUT_4[13248] = 32'b00000000000000001010011100000100;
assign LUT_4[13249] = 32'b00000000000000000011100111111100;
assign LUT_4[13250] = 32'b00000000000000001001110110101000;
assign LUT_4[13251] = 32'b00000000000000000011000010100000;
assign LUT_4[13252] = 32'b00000000000000000111011100100000;
assign LUT_4[13253] = 32'b00000000000000000000101000011000;
assign LUT_4[13254] = 32'b00000000000000000110110111000100;
assign LUT_4[13255] = 32'b00000000000000000000000010111100;
assign LUT_4[13256] = 32'b00000000000000000011101000011001;
assign LUT_4[13257] = 32'b11111111111111111100110100010001;
assign LUT_4[13258] = 32'b00000000000000000011000010111101;
assign LUT_4[13259] = 32'b11111111111111111100001110110101;
assign LUT_4[13260] = 32'b00000000000000000000101000110101;
assign LUT_4[13261] = 32'b11111111111111111001110100101101;
assign LUT_4[13262] = 32'b00000000000000000000000011011001;
assign LUT_4[13263] = 32'b11111111111111111001001111010001;
assign LUT_4[13264] = 32'b00000000000000001000001101110010;
assign LUT_4[13265] = 32'b00000000000000000001011001101010;
assign LUT_4[13266] = 32'b00000000000000000111101000010110;
assign LUT_4[13267] = 32'b00000000000000000000110100001110;
assign LUT_4[13268] = 32'b00000000000000000101001110001110;
assign LUT_4[13269] = 32'b11111111111111111110011010000110;
assign LUT_4[13270] = 32'b00000000000000000100101000110010;
assign LUT_4[13271] = 32'b11111111111111111101110100101010;
assign LUT_4[13272] = 32'b00000000000000000001011010000111;
assign LUT_4[13273] = 32'b11111111111111111010100101111111;
assign LUT_4[13274] = 32'b00000000000000000000110100101011;
assign LUT_4[13275] = 32'b11111111111111111010000000100011;
assign LUT_4[13276] = 32'b11111111111111111110011010100011;
assign LUT_4[13277] = 32'b11111111111111110111100110011011;
assign LUT_4[13278] = 32'b11111111111111111101110101000111;
assign LUT_4[13279] = 32'b11111111111111110111000000111111;
assign LUT_4[13280] = 32'b00000000000000001000110111001011;
assign LUT_4[13281] = 32'b00000000000000000010000011000011;
assign LUT_4[13282] = 32'b00000000000000001000010001101111;
assign LUT_4[13283] = 32'b00000000000000000001011101100111;
assign LUT_4[13284] = 32'b00000000000000000101110111100111;
assign LUT_4[13285] = 32'b11111111111111111111000011011111;
assign LUT_4[13286] = 32'b00000000000000000101010010001011;
assign LUT_4[13287] = 32'b11111111111111111110011110000011;
assign LUT_4[13288] = 32'b00000000000000000010000011100000;
assign LUT_4[13289] = 32'b11111111111111111011001111011000;
assign LUT_4[13290] = 32'b00000000000000000001011110000100;
assign LUT_4[13291] = 32'b11111111111111111010101001111100;
assign LUT_4[13292] = 32'b11111111111111111111000011111100;
assign LUT_4[13293] = 32'b11111111111111111000001111110100;
assign LUT_4[13294] = 32'b11111111111111111110011110100000;
assign LUT_4[13295] = 32'b11111111111111110111101010011000;
assign LUT_4[13296] = 32'b00000000000000000110101000111001;
assign LUT_4[13297] = 32'b11111111111111111111110100110001;
assign LUT_4[13298] = 32'b00000000000000000110000011011101;
assign LUT_4[13299] = 32'b11111111111111111111001111010101;
assign LUT_4[13300] = 32'b00000000000000000011101001010101;
assign LUT_4[13301] = 32'b11111111111111111100110101001101;
assign LUT_4[13302] = 32'b00000000000000000011000011111001;
assign LUT_4[13303] = 32'b11111111111111111100001111110001;
assign LUT_4[13304] = 32'b11111111111111111111110101001110;
assign LUT_4[13305] = 32'b11111111111111111001000001000110;
assign LUT_4[13306] = 32'b11111111111111111111001111110010;
assign LUT_4[13307] = 32'b11111111111111111000011011101010;
assign LUT_4[13308] = 32'b11111111111111111100110101101010;
assign LUT_4[13309] = 32'b11111111111111110110000001100010;
assign LUT_4[13310] = 32'b11111111111111111100010000001110;
assign LUT_4[13311] = 32'b11111111111111110101011100000110;
assign LUT_4[13312] = 32'b00000000000000000100001001011100;
assign LUT_4[13313] = 32'b11111111111111111101010101010100;
assign LUT_4[13314] = 32'b00000000000000000011100100000000;
assign LUT_4[13315] = 32'b11111111111111111100101111111000;
assign LUT_4[13316] = 32'b00000000000000000001001001111000;
assign LUT_4[13317] = 32'b11111111111111111010010101110000;
assign LUT_4[13318] = 32'b00000000000000000000100100011100;
assign LUT_4[13319] = 32'b11111111111111111001110000010100;
assign LUT_4[13320] = 32'b11111111111111111101010101110001;
assign LUT_4[13321] = 32'b11111111111111110110100001101001;
assign LUT_4[13322] = 32'b11111111111111111100110000010101;
assign LUT_4[13323] = 32'b11111111111111110101111100001101;
assign LUT_4[13324] = 32'b11111111111111111010010110001101;
assign LUT_4[13325] = 32'b11111111111111110011100010000101;
assign LUT_4[13326] = 32'b11111111111111111001110000110001;
assign LUT_4[13327] = 32'b11111111111111110010111100101001;
assign LUT_4[13328] = 32'b00000000000000000001111011001010;
assign LUT_4[13329] = 32'b11111111111111111011000111000010;
assign LUT_4[13330] = 32'b00000000000000000001010101101110;
assign LUT_4[13331] = 32'b11111111111111111010100001100110;
assign LUT_4[13332] = 32'b11111111111111111110111011100110;
assign LUT_4[13333] = 32'b11111111111111111000000111011110;
assign LUT_4[13334] = 32'b11111111111111111110010110001010;
assign LUT_4[13335] = 32'b11111111111111110111100010000010;
assign LUT_4[13336] = 32'b11111111111111111011000111011111;
assign LUT_4[13337] = 32'b11111111111111110100010011010111;
assign LUT_4[13338] = 32'b11111111111111111010100010000011;
assign LUT_4[13339] = 32'b11111111111111110011101101111011;
assign LUT_4[13340] = 32'b11111111111111111000000111111011;
assign LUT_4[13341] = 32'b11111111111111110001010011110011;
assign LUT_4[13342] = 32'b11111111111111110111100010011111;
assign LUT_4[13343] = 32'b11111111111111110000101110010111;
assign LUT_4[13344] = 32'b00000000000000000010100100100011;
assign LUT_4[13345] = 32'b11111111111111111011110000011011;
assign LUT_4[13346] = 32'b00000000000000000001111111000111;
assign LUT_4[13347] = 32'b11111111111111111011001010111111;
assign LUT_4[13348] = 32'b11111111111111111111100100111111;
assign LUT_4[13349] = 32'b11111111111111111000110000110111;
assign LUT_4[13350] = 32'b11111111111111111110111111100011;
assign LUT_4[13351] = 32'b11111111111111111000001011011011;
assign LUT_4[13352] = 32'b11111111111111111011110000111000;
assign LUT_4[13353] = 32'b11111111111111110100111100110000;
assign LUT_4[13354] = 32'b11111111111111111011001011011100;
assign LUT_4[13355] = 32'b11111111111111110100010111010100;
assign LUT_4[13356] = 32'b11111111111111111000110001010100;
assign LUT_4[13357] = 32'b11111111111111110001111101001100;
assign LUT_4[13358] = 32'b11111111111111111000001011111000;
assign LUT_4[13359] = 32'b11111111111111110001010111110000;
assign LUT_4[13360] = 32'b00000000000000000000010110010001;
assign LUT_4[13361] = 32'b11111111111111111001100010001001;
assign LUT_4[13362] = 32'b11111111111111111111110000110101;
assign LUT_4[13363] = 32'b11111111111111111000111100101101;
assign LUT_4[13364] = 32'b11111111111111111101010110101101;
assign LUT_4[13365] = 32'b11111111111111110110100010100101;
assign LUT_4[13366] = 32'b11111111111111111100110001010001;
assign LUT_4[13367] = 32'b11111111111111110101111101001001;
assign LUT_4[13368] = 32'b11111111111111111001100010100110;
assign LUT_4[13369] = 32'b11111111111111110010101110011110;
assign LUT_4[13370] = 32'b11111111111111111000111101001010;
assign LUT_4[13371] = 32'b11111111111111110010001001000010;
assign LUT_4[13372] = 32'b11111111111111110110100011000010;
assign LUT_4[13373] = 32'b11111111111111101111101110111010;
assign LUT_4[13374] = 32'b11111111111111110101111101100110;
assign LUT_4[13375] = 32'b11111111111111101111001001011110;
assign LUT_4[13376] = 32'b00000000000000000101100000110000;
assign LUT_4[13377] = 32'b11111111111111111110101100101000;
assign LUT_4[13378] = 32'b00000000000000000100111011010100;
assign LUT_4[13379] = 32'b11111111111111111110000111001100;
assign LUT_4[13380] = 32'b00000000000000000010100001001100;
assign LUT_4[13381] = 32'b11111111111111111011101101000100;
assign LUT_4[13382] = 32'b00000000000000000001111011110000;
assign LUT_4[13383] = 32'b11111111111111111011000111101000;
assign LUT_4[13384] = 32'b11111111111111111110101101000101;
assign LUT_4[13385] = 32'b11111111111111110111111000111101;
assign LUT_4[13386] = 32'b11111111111111111110000111101001;
assign LUT_4[13387] = 32'b11111111111111110111010011100001;
assign LUT_4[13388] = 32'b11111111111111111011101101100001;
assign LUT_4[13389] = 32'b11111111111111110100111001011001;
assign LUT_4[13390] = 32'b11111111111111111011001000000101;
assign LUT_4[13391] = 32'b11111111111111110100010011111101;
assign LUT_4[13392] = 32'b00000000000000000011010010011110;
assign LUT_4[13393] = 32'b11111111111111111100011110010110;
assign LUT_4[13394] = 32'b00000000000000000010101101000010;
assign LUT_4[13395] = 32'b11111111111111111011111000111010;
assign LUT_4[13396] = 32'b00000000000000000000010010111010;
assign LUT_4[13397] = 32'b11111111111111111001011110110010;
assign LUT_4[13398] = 32'b11111111111111111111101101011110;
assign LUT_4[13399] = 32'b11111111111111111000111001010110;
assign LUT_4[13400] = 32'b11111111111111111100011110110011;
assign LUT_4[13401] = 32'b11111111111111110101101010101011;
assign LUT_4[13402] = 32'b11111111111111111011111001010111;
assign LUT_4[13403] = 32'b11111111111111110101000101001111;
assign LUT_4[13404] = 32'b11111111111111111001011111001111;
assign LUT_4[13405] = 32'b11111111111111110010101011000111;
assign LUT_4[13406] = 32'b11111111111111111000111001110011;
assign LUT_4[13407] = 32'b11111111111111110010000101101011;
assign LUT_4[13408] = 32'b00000000000000000011111011110111;
assign LUT_4[13409] = 32'b11111111111111111101000111101111;
assign LUT_4[13410] = 32'b00000000000000000011010110011011;
assign LUT_4[13411] = 32'b11111111111111111100100010010011;
assign LUT_4[13412] = 32'b00000000000000000000111100010011;
assign LUT_4[13413] = 32'b11111111111111111010001000001011;
assign LUT_4[13414] = 32'b00000000000000000000010110110111;
assign LUT_4[13415] = 32'b11111111111111111001100010101111;
assign LUT_4[13416] = 32'b11111111111111111101001000001100;
assign LUT_4[13417] = 32'b11111111111111110110010100000100;
assign LUT_4[13418] = 32'b11111111111111111100100010110000;
assign LUT_4[13419] = 32'b11111111111111110101101110101000;
assign LUT_4[13420] = 32'b11111111111111111010001000101000;
assign LUT_4[13421] = 32'b11111111111111110011010100100000;
assign LUT_4[13422] = 32'b11111111111111111001100011001100;
assign LUT_4[13423] = 32'b11111111111111110010101111000100;
assign LUT_4[13424] = 32'b00000000000000000001101101100101;
assign LUT_4[13425] = 32'b11111111111111111010111001011101;
assign LUT_4[13426] = 32'b00000000000000000001001000001001;
assign LUT_4[13427] = 32'b11111111111111111010010100000001;
assign LUT_4[13428] = 32'b11111111111111111110101110000001;
assign LUT_4[13429] = 32'b11111111111111110111111001111001;
assign LUT_4[13430] = 32'b11111111111111111110001000100101;
assign LUT_4[13431] = 32'b11111111111111110111010100011101;
assign LUT_4[13432] = 32'b11111111111111111010111001111010;
assign LUT_4[13433] = 32'b11111111111111110100000101110010;
assign LUT_4[13434] = 32'b11111111111111111010010100011110;
assign LUT_4[13435] = 32'b11111111111111110011100000010110;
assign LUT_4[13436] = 32'b11111111111111110111111010010110;
assign LUT_4[13437] = 32'b11111111111111110001000110001110;
assign LUT_4[13438] = 32'b11111111111111110111010100111010;
assign LUT_4[13439] = 32'b11111111111111110000100000110010;
assign LUT_4[13440] = 32'b00000000000000000110101111100100;
assign LUT_4[13441] = 32'b11111111111111111111111011011100;
assign LUT_4[13442] = 32'b00000000000000000110001010001000;
assign LUT_4[13443] = 32'b11111111111111111111010110000000;
assign LUT_4[13444] = 32'b00000000000000000011110000000000;
assign LUT_4[13445] = 32'b11111111111111111100111011111000;
assign LUT_4[13446] = 32'b00000000000000000011001010100100;
assign LUT_4[13447] = 32'b11111111111111111100010110011100;
assign LUT_4[13448] = 32'b11111111111111111111111011111001;
assign LUT_4[13449] = 32'b11111111111111111001000111110001;
assign LUT_4[13450] = 32'b11111111111111111111010110011101;
assign LUT_4[13451] = 32'b11111111111111111000100010010101;
assign LUT_4[13452] = 32'b11111111111111111100111100010101;
assign LUT_4[13453] = 32'b11111111111111110110001000001101;
assign LUT_4[13454] = 32'b11111111111111111100010110111001;
assign LUT_4[13455] = 32'b11111111111111110101100010110001;
assign LUT_4[13456] = 32'b00000000000000000100100001010010;
assign LUT_4[13457] = 32'b11111111111111111101101101001010;
assign LUT_4[13458] = 32'b00000000000000000011111011110110;
assign LUT_4[13459] = 32'b11111111111111111101000111101110;
assign LUT_4[13460] = 32'b00000000000000000001100001101110;
assign LUT_4[13461] = 32'b11111111111111111010101101100110;
assign LUT_4[13462] = 32'b00000000000000000000111100010010;
assign LUT_4[13463] = 32'b11111111111111111010001000001010;
assign LUT_4[13464] = 32'b11111111111111111101101101100111;
assign LUT_4[13465] = 32'b11111111111111110110111001011111;
assign LUT_4[13466] = 32'b11111111111111111101001000001011;
assign LUT_4[13467] = 32'b11111111111111110110010100000011;
assign LUT_4[13468] = 32'b11111111111111111010101110000011;
assign LUT_4[13469] = 32'b11111111111111110011111001111011;
assign LUT_4[13470] = 32'b11111111111111111010001000100111;
assign LUT_4[13471] = 32'b11111111111111110011010100011111;
assign LUT_4[13472] = 32'b00000000000000000101001010101011;
assign LUT_4[13473] = 32'b11111111111111111110010110100011;
assign LUT_4[13474] = 32'b00000000000000000100100101001111;
assign LUT_4[13475] = 32'b11111111111111111101110001000111;
assign LUT_4[13476] = 32'b00000000000000000010001011000111;
assign LUT_4[13477] = 32'b11111111111111111011010110111111;
assign LUT_4[13478] = 32'b00000000000000000001100101101011;
assign LUT_4[13479] = 32'b11111111111111111010110001100011;
assign LUT_4[13480] = 32'b11111111111111111110010111000000;
assign LUT_4[13481] = 32'b11111111111111110111100010111000;
assign LUT_4[13482] = 32'b11111111111111111101110001100100;
assign LUT_4[13483] = 32'b11111111111111110110111101011100;
assign LUT_4[13484] = 32'b11111111111111111011010111011100;
assign LUT_4[13485] = 32'b11111111111111110100100011010100;
assign LUT_4[13486] = 32'b11111111111111111010110010000000;
assign LUT_4[13487] = 32'b11111111111111110011111101111000;
assign LUT_4[13488] = 32'b00000000000000000010111100011001;
assign LUT_4[13489] = 32'b11111111111111111100001000010001;
assign LUT_4[13490] = 32'b00000000000000000010010110111101;
assign LUT_4[13491] = 32'b11111111111111111011100010110101;
assign LUT_4[13492] = 32'b11111111111111111111111100110101;
assign LUT_4[13493] = 32'b11111111111111111001001000101101;
assign LUT_4[13494] = 32'b11111111111111111111010111011001;
assign LUT_4[13495] = 32'b11111111111111111000100011010001;
assign LUT_4[13496] = 32'b11111111111111111100001000101110;
assign LUT_4[13497] = 32'b11111111111111110101010100100110;
assign LUT_4[13498] = 32'b11111111111111111011100011010010;
assign LUT_4[13499] = 32'b11111111111111110100101111001010;
assign LUT_4[13500] = 32'b11111111111111111001001001001010;
assign LUT_4[13501] = 32'b11111111111111110010010101000010;
assign LUT_4[13502] = 32'b11111111111111111000100011101110;
assign LUT_4[13503] = 32'b11111111111111110001101111100110;
assign LUT_4[13504] = 32'b00000000000000001000000110111000;
assign LUT_4[13505] = 32'b00000000000000000001010010110000;
assign LUT_4[13506] = 32'b00000000000000000111100001011100;
assign LUT_4[13507] = 32'b00000000000000000000101101010100;
assign LUT_4[13508] = 32'b00000000000000000101000111010100;
assign LUT_4[13509] = 32'b11111111111111111110010011001100;
assign LUT_4[13510] = 32'b00000000000000000100100001111000;
assign LUT_4[13511] = 32'b11111111111111111101101101110000;
assign LUT_4[13512] = 32'b00000000000000000001010011001101;
assign LUT_4[13513] = 32'b11111111111111111010011111000101;
assign LUT_4[13514] = 32'b00000000000000000000101101110001;
assign LUT_4[13515] = 32'b11111111111111111001111001101001;
assign LUT_4[13516] = 32'b11111111111111111110010011101001;
assign LUT_4[13517] = 32'b11111111111111110111011111100001;
assign LUT_4[13518] = 32'b11111111111111111101101110001101;
assign LUT_4[13519] = 32'b11111111111111110110111010000101;
assign LUT_4[13520] = 32'b00000000000000000101111000100110;
assign LUT_4[13521] = 32'b11111111111111111111000100011110;
assign LUT_4[13522] = 32'b00000000000000000101010011001010;
assign LUT_4[13523] = 32'b11111111111111111110011111000010;
assign LUT_4[13524] = 32'b00000000000000000010111001000010;
assign LUT_4[13525] = 32'b11111111111111111100000100111010;
assign LUT_4[13526] = 32'b00000000000000000010010011100110;
assign LUT_4[13527] = 32'b11111111111111111011011111011110;
assign LUT_4[13528] = 32'b11111111111111111111000100111011;
assign LUT_4[13529] = 32'b11111111111111111000010000110011;
assign LUT_4[13530] = 32'b11111111111111111110011111011111;
assign LUT_4[13531] = 32'b11111111111111110111101011010111;
assign LUT_4[13532] = 32'b11111111111111111100000101010111;
assign LUT_4[13533] = 32'b11111111111111110101010001001111;
assign LUT_4[13534] = 32'b11111111111111111011011111111011;
assign LUT_4[13535] = 32'b11111111111111110100101011110011;
assign LUT_4[13536] = 32'b00000000000000000110100001111111;
assign LUT_4[13537] = 32'b11111111111111111111101101110111;
assign LUT_4[13538] = 32'b00000000000000000101111100100011;
assign LUT_4[13539] = 32'b11111111111111111111001000011011;
assign LUT_4[13540] = 32'b00000000000000000011100010011011;
assign LUT_4[13541] = 32'b11111111111111111100101110010011;
assign LUT_4[13542] = 32'b00000000000000000010111100111111;
assign LUT_4[13543] = 32'b11111111111111111100001000110111;
assign LUT_4[13544] = 32'b11111111111111111111101110010100;
assign LUT_4[13545] = 32'b11111111111111111000111010001100;
assign LUT_4[13546] = 32'b11111111111111111111001000111000;
assign LUT_4[13547] = 32'b11111111111111111000010100110000;
assign LUT_4[13548] = 32'b11111111111111111100101110110000;
assign LUT_4[13549] = 32'b11111111111111110101111010101000;
assign LUT_4[13550] = 32'b11111111111111111100001001010100;
assign LUT_4[13551] = 32'b11111111111111110101010101001100;
assign LUT_4[13552] = 32'b00000000000000000100010011101101;
assign LUT_4[13553] = 32'b11111111111111111101011111100101;
assign LUT_4[13554] = 32'b00000000000000000011101110010001;
assign LUT_4[13555] = 32'b11111111111111111100111010001001;
assign LUT_4[13556] = 32'b00000000000000000001010100001001;
assign LUT_4[13557] = 32'b11111111111111111010100000000001;
assign LUT_4[13558] = 32'b00000000000000000000101110101101;
assign LUT_4[13559] = 32'b11111111111111111001111010100101;
assign LUT_4[13560] = 32'b11111111111111111101100000000010;
assign LUT_4[13561] = 32'b11111111111111110110101011111010;
assign LUT_4[13562] = 32'b11111111111111111100111010100110;
assign LUT_4[13563] = 32'b11111111111111110110000110011110;
assign LUT_4[13564] = 32'b11111111111111111010100000011110;
assign LUT_4[13565] = 32'b11111111111111110011101100010110;
assign LUT_4[13566] = 32'b11111111111111111001111011000010;
assign LUT_4[13567] = 32'b11111111111111110011000110111010;
assign LUT_4[13568] = 32'b00000000000000001001000100111111;
assign LUT_4[13569] = 32'b00000000000000000010010000110111;
assign LUT_4[13570] = 32'b00000000000000001000011111100011;
assign LUT_4[13571] = 32'b00000000000000000001101011011011;
assign LUT_4[13572] = 32'b00000000000000000110000101011011;
assign LUT_4[13573] = 32'b11111111111111111111010001010011;
assign LUT_4[13574] = 32'b00000000000000000101011111111111;
assign LUT_4[13575] = 32'b11111111111111111110101011110111;
assign LUT_4[13576] = 32'b00000000000000000010010001010100;
assign LUT_4[13577] = 32'b11111111111111111011011101001100;
assign LUT_4[13578] = 32'b00000000000000000001101011111000;
assign LUT_4[13579] = 32'b11111111111111111010110111110000;
assign LUT_4[13580] = 32'b11111111111111111111010001110000;
assign LUT_4[13581] = 32'b11111111111111111000011101101000;
assign LUT_4[13582] = 32'b11111111111111111110101100010100;
assign LUT_4[13583] = 32'b11111111111111110111111000001100;
assign LUT_4[13584] = 32'b00000000000000000110110110101101;
assign LUT_4[13585] = 32'b00000000000000000000000010100101;
assign LUT_4[13586] = 32'b00000000000000000110010001010001;
assign LUT_4[13587] = 32'b11111111111111111111011101001001;
assign LUT_4[13588] = 32'b00000000000000000011110111001001;
assign LUT_4[13589] = 32'b11111111111111111101000011000001;
assign LUT_4[13590] = 32'b00000000000000000011010001101101;
assign LUT_4[13591] = 32'b11111111111111111100011101100101;
assign LUT_4[13592] = 32'b00000000000000000000000011000010;
assign LUT_4[13593] = 32'b11111111111111111001001110111010;
assign LUT_4[13594] = 32'b11111111111111111111011101100110;
assign LUT_4[13595] = 32'b11111111111111111000101001011110;
assign LUT_4[13596] = 32'b11111111111111111101000011011110;
assign LUT_4[13597] = 32'b11111111111111110110001111010110;
assign LUT_4[13598] = 32'b11111111111111111100011110000010;
assign LUT_4[13599] = 32'b11111111111111110101101001111010;
assign LUT_4[13600] = 32'b00000000000000000111100000000110;
assign LUT_4[13601] = 32'b00000000000000000000101011111110;
assign LUT_4[13602] = 32'b00000000000000000110111010101010;
assign LUT_4[13603] = 32'b00000000000000000000000110100010;
assign LUT_4[13604] = 32'b00000000000000000100100000100010;
assign LUT_4[13605] = 32'b11111111111111111101101100011010;
assign LUT_4[13606] = 32'b00000000000000000011111011000110;
assign LUT_4[13607] = 32'b11111111111111111101000110111110;
assign LUT_4[13608] = 32'b00000000000000000000101100011011;
assign LUT_4[13609] = 32'b11111111111111111001111000010011;
assign LUT_4[13610] = 32'b00000000000000000000000110111111;
assign LUT_4[13611] = 32'b11111111111111111001010010110111;
assign LUT_4[13612] = 32'b11111111111111111101101100110111;
assign LUT_4[13613] = 32'b11111111111111110110111000101111;
assign LUT_4[13614] = 32'b11111111111111111101000111011011;
assign LUT_4[13615] = 32'b11111111111111110110010011010011;
assign LUT_4[13616] = 32'b00000000000000000101010001110100;
assign LUT_4[13617] = 32'b11111111111111111110011101101100;
assign LUT_4[13618] = 32'b00000000000000000100101100011000;
assign LUT_4[13619] = 32'b11111111111111111101111000010000;
assign LUT_4[13620] = 32'b00000000000000000010010010010000;
assign LUT_4[13621] = 32'b11111111111111111011011110001000;
assign LUT_4[13622] = 32'b00000000000000000001101100110100;
assign LUT_4[13623] = 32'b11111111111111111010111000101100;
assign LUT_4[13624] = 32'b11111111111111111110011110001001;
assign LUT_4[13625] = 32'b11111111111111110111101010000001;
assign LUT_4[13626] = 32'b11111111111111111101111000101101;
assign LUT_4[13627] = 32'b11111111111111110111000100100101;
assign LUT_4[13628] = 32'b11111111111111111011011110100101;
assign LUT_4[13629] = 32'b11111111111111110100101010011101;
assign LUT_4[13630] = 32'b11111111111111111010111001001001;
assign LUT_4[13631] = 32'b11111111111111110100000101000001;
assign LUT_4[13632] = 32'b00000000000000001010011100010011;
assign LUT_4[13633] = 32'b00000000000000000011101000001011;
assign LUT_4[13634] = 32'b00000000000000001001110110110111;
assign LUT_4[13635] = 32'b00000000000000000011000010101111;
assign LUT_4[13636] = 32'b00000000000000000111011100101111;
assign LUT_4[13637] = 32'b00000000000000000000101000100111;
assign LUT_4[13638] = 32'b00000000000000000110110111010011;
assign LUT_4[13639] = 32'b00000000000000000000000011001011;
assign LUT_4[13640] = 32'b00000000000000000011101000101000;
assign LUT_4[13641] = 32'b11111111111111111100110100100000;
assign LUT_4[13642] = 32'b00000000000000000011000011001100;
assign LUT_4[13643] = 32'b11111111111111111100001111000100;
assign LUT_4[13644] = 32'b00000000000000000000101001000100;
assign LUT_4[13645] = 32'b11111111111111111001110100111100;
assign LUT_4[13646] = 32'b00000000000000000000000011101000;
assign LUT_4[13647] = 32'b11111111111111111001001111100000;
assign LUT_4[13648] = 32'b00000000000000001000001110000001;
assign LUT_4[13649] = 32'b00000000000000000001011001111001;
assign LUT_4[13650] = 32'b00000000000000000111101000100101;
assign LUT_4[13651] = 32'b00000000000000000000110100011101;
assign LUT_4[13652] = 32'b00000000000000000101001110011101;
assign LUT_4[13653] = 32'b11111111111111111110011010010101;
assign LUT_4[13654] = 32'b00000000000000000100101001000001;
assign LUT_4[13655] = 32'b11111111111111111101110100111001;
assign LUT_4[13656] = 32'b00000000000000000001011010010110;
assign LUT_4[13657] = 32'b11111111111111111010100110001110;
assign LUT_4[13658] = 32'b00000000000000000000110100111010;
assign LUT_4[13659] = 32'b11111111111111111010000000110010;
assign LUT_4[13660] = 32'b11111111111111111110011010110010;
assign LUT_4[13661] = 32'b11111111111111110111100110101010;
assign LUT_4[13662] = 32'b11111111111111111101110101010110;
assign LUT_4[13663] = 32'b11111111111111110111000001001110;
assign LUT_4[13664] = 32'b00000000000000001000110111011010;
assign LUT_4[13665] = 32'b00000000000000000010000011010010;
assign LUT_4[13666] = 32'b00000000000000001000010001111110;
assign LUT_4[13667] = 32'b00000000000000000001011101110110;
assign LUT_4[13668] = 32'b00000000000000000101110111110110;
assign LUT_4[13669] = 32'b11111111111111111111000011101110;
assign LUT_4[13670] = 32'b00000000000000000101010010011010;
assign LUT_4[13671] = 32'b11111111111111111110011110010010;
assign LUT_4[13672] = 32'b00000000000000000010000011101111;
assign LUT_4[13673] = 32'b11111111111111111011001111100111;
assign LUT_4[13674] = 32'b00000000000000000001011110010011;
assign LUT_4[13675] = 32'b11111111111111111010101010001011;
assign LUT_4[13676] = 32'b11111111111111111111000100001011;
assign LUT_4[13677] = 32'b11111111111111111000010000000011;
assign LUT_4[13678] = 32'b11111111111111111110011110101111;
assign LUT_4[13679] = 32'b11111111111111110111101010100111;
assign LUT_4[13680] = 32'b00000000000000000110101001001000;
assign LUT_4[13681] = 32'b11111111111111111111110101000000;
assign LUT_4[13682] = 32'b00000000000000000110000011101100;
assign LUT_4[13683] = 32'b11111111111111111111001111100100;
assign LUT_4[13684] = 32'b00000000000000000011101001100100;
assign LUT_4[13685] = 32'b11111111111111111100110101011100;
assign LUT_4[13686] = 32'b00000000000000000011000100001000;
assign LUT_4[13687] = 32'b11111111111111111100010000000000;
assign LUT_4[13688] = 32'b11111111111111111111110101011101;
assign LUT_4[13689] = 32'b11111111111111111001000001010101;
assign LUT_4[13690] = 32'b11111111111111111111010000000001;
assign LUT_4[13691] = 32'b11111111111111111000011011111001;
assign LUT_4[13692] = 32'b11111111111111111100110101111001;
assign LUT_4[13693] = 32'b11111111111111110110000001110001;
assign LUT_4[13694] = 32'b11111111111111111100010000011101;
assign LUT_4[13695] = 32'b11111111111111110101011100010101;
assign LUT_4[13696] = 32'b00000000000000001011101011000111;
assign LUT_4[13697] = 32'b00000000000000000100110110111111;
assign LUT_4[13698] = 32'b00000000000000001011000101101011;
assign LUT_4[13699] = 32'b00000000000000000100010001100011;
assign LUT_4[13700] = 32'b00000000000000001000101011100011;
assign LUT_4[13701] = 32'b00000000000000000001110111011011;
assign LUT_4[13702] = 32'b00000000000000001000000110000111;
assign LUT_4[13703] = 32'b00000000000000000001010001111111;
assign LUT_4[13704] = 32'b00000000000000000100110111011100;
assign LUT_4[13705] = 32'b11111111111111111110000011010100;
assign LUT_4[13706] = 32'b00000000000000000100010010000000;
assign LUT_4[13707] = 32'b11111111111111111101011101111000;
assign LUT_4[13708] = 32'b00000000000000000001110111111000;
assign LUT_4[13709] = 32'b11111111111111111011000011110000;
assign LUT_4[13710] = 32'b00000000000000000001010010011100;
assign LUT_4[13711] = 32'b11111111111111111010011110010100;
assign LUT_4[13712] = 32'b00000000000000001001011100110101;
assign LUT_4[13713] = 32'b00000000000000000010101000101101;
assign LUT_4[13714] = 32'b00000000000000001000110111011001;
assign LUT_4[13715] = 32'b00000000000000000010000011010001;
assign LUT_4[13716] = 32'b00000000000000000110011101010001;
assign LUT_4[13717] = 32'b11111111111111111111101001001001;
assign LUT_4[13718] = 32'b00000000000000000101110111110101;
assign LUT_4[13719] = 32'b11111111111111111111000011101101;
assign LUT_4[13720] = 32'b00000000000000000010101001001010;
assign LUT_4[13721] = 32'b11111111111111111011110101000010;
assign LUT_4[13722] = 32'b00000000000000000010000011101110;
assign LUT_4[13723] = 32'b11111111111111111011001111100110;
assign LUT_4[13724] = 32'b11111111111111111111101001100110;
assign LUT_4[13725] = 32'b11111111111111111000110101011110;
assign LUT_4[13726] = 32'b11111111111111111111000100001010;
assign LUT_4[13727] = 32'b11111111111111111000010000000010;
assign LUT_4[13728] = 32'b00000000000000001010000110001110;
assign LUT_4[13729] = 32'b00000000000000000011010010000110;
assign LUT_4[13730] = 32'b00000000000000001001100000110010;
assign LUT_4[13731] = 32'b00000000000000000010101100101010;
assign LUT_4[13732] = 32'b00000000000000000111000110101010;
assign LUT_4[13733] = 32'b00000000000000000000010010100010;
assign LUT_4[13734] = 32'b00000000000000000110100001001110;
assign LUT_4[13735] = 32'b11111111111111111111101101000110;
assign LUT_4[13736] = 32'b00000000000000000011010010100011;
assign LUT_4[13737] = 32'b11111111111111111100011110011011;
assign LUT_4[13738] = 32'b00000000000000000010101101000111;
assign LUT_4[13739] = 32'b11111111111111111011111000111111;
assign LUT_4[13740] = 32'b00000000000000000000010010111111;
assign LUT_4[13741] = 32'b11111111111111111001011110110111;
assign LUT_4[13742] = 32'b11111111111111111111101101100011;
assign LUT_4[13743] = 32'b11111111111111111000111001011011;
assign LUT_4[13744] = 32'b00000000000000000111110111111100;
assign LUT_4[13745] = 32'b00000000000000000001000011110100;
assign LUT_4[13746] = 32'b00000000000000000111010010100000;
assign LUT_4[13747] = 32'b00000000000000000000011110011000;
assign LUT_4[13748] = 32'b00000000000000000100111000011000;
assign LUT_4[13749] = 32'b11111111111111111110000100010000;
assign LUT_4[13750] = 32'b00000000000000000100010010111100;
assign LUT_4[13751] = 32'b11111111111111111101011110110100;
assign LUT_4[13752] = 32'b00000000000000000001000100010001;
assign LUT_4[13753] = 32'b11111111111111111010010000001001;
assign LUT_4[13754] = 32'b00000000000000000000011110110101;
assign LUT_4[13755] = 32'b11111111111111111001101010101101;
assign LUT_4[13756] = 32'b11111111111111111110000100101101;
assign LUT_4[13757] = 32'b11111111111111110111010000100101;
assign LUT_4[13758] = 32'b11111111111111111101011111010001;
assign LUT_4[13759] = 32'b11111111111111110110101011001001;
assign LUT_4[13760] = 32'b00000000000000001101000010011011;
assign LUT_4[13761] = 32'b00000000000000000110001110010011;
assign LUT_4[13762] = 32'b00000000000000001100011100111111;
assign LUT_4[13763] = 32'b00000000000000000101101000110111;
assign LUT_4[13764] = 32'b00000000000000001010000010110111;
assign LUT_4[13765] = 32'b00000000000000000011001110101111;
assign LUT_4[13766] = 32'b00000000000000001001011101011011;
assign LUT_4[13767] = 32'b00000000000000000010101001010011;
assign LUT_4[13768] = 32'b00000000000000000110001110110000;
assign LUT_4[13769] = 32'b11111111111111111111011010101000;
assign LUT_4[13770] = 32'b00000000000000000101101001010100;
assign LUT_4[13771] = 32'b11111111111111111110110101001100;
assign LUT_4[13772] = 32'b00000000000000000011001111001100;
assign LUT_4[13773] = 32'b11111111111111111100011011000100;
assign LUT_4[13774] = 32'b00000000000000000010101001110000;
assign LUT_4[13775] = 32'b11111111111111111011110101101000;
assign LUT_4[13776] = 32'b00000000000000001010110100001001;
assign LUT_4[13777] = 32'b00000000000000000100000000000001;
assign LUT_4[13778] = 32'b00000000000000001010001110101101;
assign LUT_4[13779] = 32'b00000000000000000011011010100101;
assign LUT_4[13780] = 32'b00000000000000000111110100100101;
assign LUT_4[13781] = 32'b00000000000000000001000000011101;
assign LUT_4[13782] = 32'b00000000000000000111001111001001;
assign LUT_4[13783] = 32'b00000000000000000000011011000001;
assign LUT_4[13784] = 32'b00000000000000000100000000011110;
assign LUT_4[13785] = 32'b11111111111111111101001100010110;
assign LUT_4[13786] = 32'b00000000000000000011011011000010;
assign LUT_4[13787] = 32'b11111111111111111100100110111010;
assign LUT_4[13788] = 32'b00000000000000000001000000111010;
assign LUT_4[13789] = 32'b11111111111111111010001100110010;
assign LUT_4[13790] = 32'b00000000000000000000011011011110;
assign LUT_4[13791] = 32'b11111111111111111001100111010110;
assign LUT_4[13792] = 32'b00000000000000001011011101100010;
assign LUT_4[13793] = 32'b00000000000000000100101001011010;
assign LUT_4[13794] = 32'b00000000000000001010111000000110;
assign LUT_4[13795] = 32'b00000000000000000100000011111110;
assign LUT_4[13796] = 32'b00000000000000001000011101111110;
assign LUT_4[13797] = 32'b00000000000000000001101001110110;
assign LUT_4[13798] = 32'b00000000000000000111111000100010;
assign LUT_4[13799] = 32'b00000000000000000001000100011010;
assign LUT_4[13800] = 32'b00000000000000000100101001110111;
assign LUT_4[13801] = 32'b11111111111111111101110101101111;
assign LUT_4[13802] = 32'b00000000000000000100000100011011;
assign LUT_4[13803] = 32'b11111111111111111101010000010011;
assign LUT_4[13804] = 32'b00000000000000000001101010010011;
assign LUT_4[13805] = 32'b11111111111111111010110110001011;
assign LUT_4[13806] = 32'b00000000000000000001000100110111;
assign LUT_4[13807] = 32'b11111111111111111010010000101111;
assign LUT_4[13808] = 32'b00000000000000001001001111010000;
assign LUT_4[13809] = 32'b00000000000000000010011011001000;
assign LUT_4[13810] = 32'b00000000000000001000101001110100;
assign LUT_4[13811] = 32'b00000000000000000001110101101100;
assign LUT_4[13812] = 32'b00000000000000000110001111101100;
assign LUT_4[13813] = 32'b11111111111111111111011011100100;
assign LUT_4[13814] = 32'b00000000000000000101101010010000;
assign LUT_4[13815] = 32'b11111111111111111110110110001000;
assign LUT_4[13816] = 32'b00000000000000000010011011100101;
assign LUT_4[13817] = 32'b11111111111111111011100111011101;
assign LUT_4[13818] = 32'b00000000000000000001110110001001;
assign LUT_4[13819] = 32'b11111111111111111011000010000001;
assign LUT_4[13820] = 32'b11111111111111111111011100000001;
assign LUT_4[13821] = 32'b11111111111111111000100111111001;
assign LUT_4[13822] = 32'b11111111111111111110110110100101;
assign LUT_4[13823] = 32'b11111111111111111000000010011101;
assign LUT_4[13824] = 32'b00000000000000000011001101100100;
assign LUT_4[13825] = 32'b11111111111111111100011001011100;
assign LUT_4[13826] = 32'b00000000000000000010101000001000;
assign LUT_4[13827] = 32'b11111111111111111011110100000000;
assign LUT_4[13828] = 32'b00000000000000000000001110000000;
assign LUT_4[13829] = 32'b11111111111111111001011001111000;
assign LUT_4[13830] = 32'b11111111111111111111101000100100;
assign LUT_4[13831] = 32'b11111111111111111000110100011100;
assign LUT_4[13832] = 32'b11111111111111111100011001111001;
assign LUT_4[13833] = 32'b11111111111111110101100101110001;
assign LUT_4[13834] = 32'b11111111111111111011110100011101;
assign LUT_4[13835] = 32'b11111111111111110101000000010101;
assign LUT_4[13836] = 32'b11111111111111111001011010010101;
assign LUT_4[13837] = 32'b11111111111111110010100110001101;
assign LUT_4[13838] = 32'b11111111111111111000110100111001;
assign LUT_4[13839] = 32'b11111111111111110010000000110001;
assign LUT_4[13840] = 32'b00000000000000000000111111010010;
assign LUT_4[13841] = 32'b11111111111111111010001011001010;
assign LUT_4[13842] = 32'b00000000000000000000011001110110;
assign LUT_4[13843] = 32'b11111111111111111001100101101110;
assign LUT_4[13844] = 32'b11111111111111111101111111101110;
assign LUT_4[13845] = 32'b11111111111111110111001011100110;
assign LUT_4[13846] = 32'b11111111111111111101011010010010;
assign LUT_4[13847] = 32'b11111111111111110110100110001010;
assign LUT_4[13848] = 32'b11111111111111111010001011100111;
assign LUT_4[13849] = 32'b11111111111111110011010111011111;
assign LUT_4[13850] = 32'b11111111111111111001100110001011;
assign LUT_4[13851] = 32'b11111111111111110010110010000011;
assign LUT_4[13852] = 32'b11111111111111110111001100000011;
assign LUT_4[13853] = 32'b11111111111111110000010111111011;
assign LUT_4[13854] = 32'b11111111111111110110100110100111;
assign LUT_4[13855] = 32'b11111111111111101111110010011111;
assign LUT_4[13856] = 32'b00000000000000000001101000101011;
assign LUT_4[13857] = 32'b11111111111111111010110100100011;
assign LUT_4[13858] = 32'b00000000000000000001000011001111;
assign LUT_4[13859] = 32'b11111111111111111010001111000111;
assign LUT_4[13860] = 32'b11111111111111111110101001000111;
assign LUT_4[13861] = 32'b11111111111111110111110100111111;
assign LUT_4[13862] = 32'b11111111111111111110000011101011;
assign LUT_4[13863] = 32'b11111111111111110111001111100011;
assign LUT_4[13864] = 32'b11111111111111111010110101000000;
assign LUT_4[13865] = 32'b11111111111111110100000000111000;
assign LUT_4[13866] = 32'b11111111111111111010001111100100;
assign LUT_4[13867] = 32'b11111111111111110011011011011100;
assign LUT_4[13868] = 32'b11111111111111110111110101011100;
assign LUT_4[13869] = 32'b11111111111111110001000001010100;
assign LUT_4[13870] = 32'b11111111111111110111010000000000;
assign LUT_4[13871] = 32'b11111111111111110000011011111000;
assign LUT_4[13872] = 32'b11111111111111111111011010011001;
assign LUT_4[13873] = 32'b11111111111111111000100110010001;
assign LUT_4[13874] = 32'b11111111111111111110110100111101;
assign LUT_4[13875] = 32'b11111111111111111000000000110101;
assign LUT_4[13876] = 32'b11111111111111111100011010110101;
assign LUT_4[13877] = 32'b11111111111111110101100110101101;
assign LUT_4[13878] = 32'b11111111111111111011110101011001;
assign LUT_4[13879] = 32'b11111111111111110101000001010001;
assign LUT_4[13880] = 32'b11111111111111111000100110101110;
assign LUT_4[13881] = 32'b11111111111111110001110010100110;
assign LUT_4[13882] = 32'b11111111111111111000000001010010;
assign LUT_4[13883] = 32'b11111111111111110001001101001010;
assign LUT_4[13884] = 32'b11111111111111110101100111001010;
assign LUT_4[13885] = 32'b11111111111111101110110011000010;
assign LUT_4[13886] = 32'b11111111111111110101000001101110;
assign LUT_4[13887] = 32'b11111111111111101110001101100110;
assign LUT_4[13888] = 32'b00000000000000000100100100111000;
assign LUT_4[13889] = 32'b11111111111111111101110000110000;
assign LUT_4[13890] = 32'b00000000000000000011111111011100;
assign LUT_4[13891] = 32'b11111111111111111101001011010100;
assign LUT_4[13892] = 32'b00000000000000000001100101010100;
assign LUT_4[13893] = 32'b11111111111111111010110001001100;
assign LUT_4[13894] = 32'b00000000000000000000111111111000;
assign LUT_4[13895] = 32'b11111111111111111010001011110000;
assign LUT_4[13896] = 32'b11111111111111111101110001001101;
assign LUT_4[13897] = 32'b11111111111111110110111101000101;
assign LUT_4[13898] = 32'b11111111111111111101001011110001;
assign LUT_4[13899] = 32'b11111111111111110110010111101001;
assign LUT_4[13900] = 32'b11111111111111111010110001101001;
assign LUT_4[13901] = 32'b11111111111111110011111101100001;
assign LUT_4[13902] = 32'b11111111111111111010001100001101;
assign LUT_4[13903] = 32'b11111111111111110011011000000101;
assign LUT_4[13904] = 32'b00000000000000000010010110100110;
assign LUT_4[13905] = 32'b11111111111111111011100010011110;
assign LUT_4[13906] = 32'b00000000000000000001110001001010;
assign LUT_4[13907] = 32'b11111111111111111010111101000010;
assign LUT_4[13908] = 32'b11111111111111111111010111000010;
assign LUT_4[13909] = 32'b11111111111111111000100010111010;
assign LUT_4[13910] = 32'b11111111111111111110110001100110;
assign LUT_4[13911] = 32'b11111111111111110111111101011110;
assign LUT_4[13912] = 32'b11111111111111111011100010111011;
assign LUT_4[13913] = 32'b11111111111111110100101110110011;
assign LUT_4[13914] = 32'b11111111111111111010111101011111;
assign LUT_4[13915] = 32'b11111111111111110100001001010111;
assign LUT_4[13916] = 32'b11111111111111111000100011010111;
assign LUT_4[13917] = 32'b11111111111111110001101111001111;
assign LUT_4[13918] = 32'b11111111111111110111111101111011;
assign LUT_4[13919] = 32'b11111111111111110001001001110011;
assign LUT_4[13920] = 32'b00000000000000000010111111111111;
assign LUT_4[13921] = 32'b11111111111111111100001011110111;
assign LUT_4[13922] = 32'b00000000000000000010011010100011;
assign LUT_4[13923] = 32'b11111111111111111011100110011011;
assign LUT_4[13924] = 32'b00000000000000000000000000011011;
assign LUT_4[13925] = 32'b11111111111111111001001100010011;
assign LUT_4[13926] = 32'b11111111111111111111011010111111;
assign LUT_4[13927] = 32'b11111111111111111000100110110111;
assign LUT_4[13928] = 32'b11111111111111111100001100010100;
assign LUT_4[13929] = 32'b11111111111111110101011000001100;
assign LUT_4[13930] = 32'b11111111111111111011100110111000;
assign LUT_4[13931] = 32'b11111111111111110100110010110000;
assign LUT_4[13932] = 32'b11111111111111111001001100110000;
assign LUT_4[13933] = 32'b11111111111111110010011000101000;
assign LUT_4[13934] = 32'b11111111111111111000100111010100;
assign LUT_4[13935] = 32'b11111111111111110001110011001100;
assign LUT_4[13936] = 32'b00000000000000000000110001101101;
assign LUT_4[13937] = 32'b11111111111111111001111101100101;
assign LUT_4[13938] = 32'b00000000000000000000001100010001;
assign LUT_4[13939] = 32'b11111111111111111001011000001001;
assign LUT_4[13940] = 32'b11111111111111111101110010001001;
assign LUT_4[13941] = 32'b11111111111111110110111110000001;
assign LUT_4[13942] = 32'b11111111111111111101001100101101;
assign LUT_4[13943] = 32'b11111111111111110110011000100101;
assign LUT_4[13944] = 32'b11111111111111111001111110000010;
assign LUT_4[13945] = 32'b11111111111111110011001001111010;
assign LUT_4[13946] = 32'b11111111111111111001011000100110;
assign LUT_4[13947] = 32'b11111111111111110010100100011110;
assign LUT_4[13948] = 32'b11111111111111110110111110011110;
assign LUT_4[13949] = 32'b11111111111111110000001010010110;
assign LUT_4[13950] = 32'b11111111111111110110011001000010;
assign LUT_4[13951] = 32'b11111111111111101111100100111010;
assign LUT_4[13952] = 32'b00000000000000000101110011101100;
assign LUT_4[13953] = 32'b11111111111111111110111111100100;
assign LUT_4[13954] = 32'b00000000000000000101001110010000;
assign LUT_4[13955] = 32'b11111111111111111110011010001000;
assign LUT_4[13956] = 32'b00000000000000000010110100001000;
assign LUT_4[13957] = 32'b11111111111111111100000000000000;
assign LUT_4[13958] = 32'b00000000000000000010001110101100;
assign LUT_4[13959] = 32'b11111111111111111011011010100100;
assign LUT_4[13960] = 32'b11111111111111111111000000000001;
assign LUT_4[13961] = 32'b11111111111111111000001011111001;
assign LUT_4[13962] = 32'b11111111111111111110011010100101;
assign LUT_4[13963] = 32'b11111111111111110111100110011101;
assign LUT_4[13964] = 32'b11111111111111111100000000011101;
assign LUT_4[13965] = 32'b11111111111111110101001100010101;
assign LUT_4[13966] = 32'b11111111111111111011011011000001;
assign LUT_4[13967] = 32'b11111111111111110100100110111001;
assign LUT_4[13968] = 32'b00000000000000000011100101011010;
assign LUT_4[13969] = 32'b11111111111111111100110001010010;
assign LUT_4[13970] = 32'b00000000000000000010111111111110;
assign LUT_4[13971] = 32'b11111111111111111100001011110110;
assign LUT_4[13972] = 32'b00000000000000000000100101110110;
assign LUT_4[13973] = 32'b11111111111111111001110001101110;
assign LUT_4[13974] = 32'b00000000000000000000000000011010;
assign LUT_4[13975] = 32'b11111111111111111001001100010010;
assign LUT_4[13976] = 32'b11111111111111111100110001101111;
assign LUT_4[13977] = 32'b11111111111111110101111101100111;
assign LUT_4[13978] = 32'b11111111111111111100001100010011;
assign LUT_4[13979] = 32'b11111111111111110101011000001011;
assign LUT_4[13980] = 32'b11111111111111111001110010001011;
assign LUT_4[13981] = 32'b11111111111111110010111110000011;
assign LUT_4[13982] = 32'b11111111111111111001001100101111;
assign LUT_4[13983] = 32'b11111111111111110010011000100111;
assign LUT_4[13984] = 32'b00000000000000000100001110110011;
assign LUT_4[13985] = 32'b11111111111111111101011010101011;
assign LUT_4[13986] = 32'b00000000000000000011101001010111;
assign LUT_4[13987] = 32'b11111111111111111100110101001111;
assign LUT_4[13988] = 32'b00000000000000000001001111001111;
assign LUT_4[13989] = 32'b11111111111111111010011011000111;
assign LUT_4[13990] = 32'b00000000000000000000101001110011;
assign LUT_4[13991] = 32'b11111111111111111001110101101011;
assign LUT_4[13992] = 32'b11111111111111111101011011001000;
assign LUT_4[13993] = 32'b11111111111111110110100111000000;
assign LUT_4[13994] = 32'b11111111111111111100110101101100;
assign LUT_4[13995] = 32'b11111111111111110110000001100100;
assign LUT_4[13996] = 32'b11111111111111111010011011100100;
assign LUT_4[13997] = 32'b11111111111111110011100111011100;
assign LUT_4[13998] = 32'b11111111111111111001110110001000;
assign LUT_4[13999] = 32'b11111111111111110011000010000000;
assign LUT_4[14000] = 32'b00000000000000000010000000100001;
assign LUT_4[14001] = 32'b11111111111111111011001100011001;
assign LUT_4[14002] = 32'b00000000000000000001011011000101;
assign LUT_4[14003] = 32'b11111111111111111010100110111101;
assign LUT_4[14004] = 32'b11111111111111111111000000111101;
assign LUT_4[14005] = 32'b11111111111111111000001100110101;
assign LUT_4[14006] = 32'b11111111111111111110011011100001;
assign LUT_4[14007] = 32'b11111111111111110111100111011001;
assign LUT_4[14008] = 32'b11111111111111111011001100110110;
assign LUT_4[14009] = 32'b11111111111111110100011000101110;
assign LUT_4[14010] = 32'b11111111111111111010100111011010;
assign LUT_4[14011] = 32'b11111111111111110011110011010010;
assign LUT_4[14012] = 32'b11111111111111111000001101010010;
assign LUT_4[14013] = 32'b11111111111111110001011001001010;
assign LUT_4[14014] = 32'b11111111111111110111100111110110;
assign LUT_4[14015] = 32'b11111111111111110000110011101110;
assign LUT_4[14016] = 32'b00000000000000000111001011000000;
assign LUT_4[14017] = 32'b00000000000000000000010110111000;
assign LUT_4[14018] = 32'b00000000000000000110100101100100;
assign LUT_4[14019] = 32'b11111111111111111111110001011100;
assign LUT_4[14020] = 32'b00000000000000000100001011011100;
assign LUT_4[14021] = 32'b11111111111111111101010111010100;
assign LUT_4[14022] = 32'b00000000000000000011100110000000;
assign LUT_4[14023] = 32'b11111111111111111100110001111000;
assign LUT_4[14024] = 32'b00000000000000000000010111010101;
assign LUT_4[14025] = 32'b11111111111111111001100011001101;
assign LUT_4[14026] = 32'b11111111111111111111110001111001;
assign LUT_4[14027] = 32'b11111111111111111000111101110001;
assign LUT_4[14028] = 32'b11111111111111111101010111110001;
assign LUT_4[14029] = 32'b11111111111111110110100011101001;
assign LUT_4[14030] = 32'b11111111111111111100110010010101;
assign LUT_4[14031] = 32'b11111111111111110101111110001101;
assign LUT_4[14032] = 32'b00000000000000000100111100101110;
assign LUT_4[14033] = 32'b11111111111111111110001000100110;
assign LUT_4[14034] = 32'b00000000000000000100010111010010;
assign LUT_4[14035] = 32'b11111111111111111101100011001010;
assign LUT_4[14036] = 32'b00000000000000000001111101001010;
assign LUT_4[14037] = 32'b11111111111111111011001001000010;
assign LUT_4[14038] = 32'b00000000000000000001010111101110;
assign LUT_4[14039] = 32'b11111111111111111010100011100110;
assign LUT_4[14040] = 32'b11111111111111111110001001000011;
assign LUT_4[14041] = 32'b11111111111111110111010100111011;
assign LUT_4[14042] = 32'b11111111111111111101100011100111;
assign LUT_4[14043] = 32'b11111111111111110110101111011111;
assign LUT_4[14044] = 32'b11111111111111111011001001011111;
assign LUT_4[14045] = 32'b11111111111111110100010101010111;
assign LUT_4[14046] = 32'b11111111111111111010100100000011;
assign LUT_4[14047] = 32'b11111111111111110011101111111011;
assign LUT_4[14048] = 32'b00000000000000000101100110000111;
assign LUT_4[14049] = 32'b11111111111111111110110001111111;
assign LUT_4[14050] = 32'b00000000000000000101000000101011;
assign LUT_4[14051] = 32'b11111111111111111110001100100011;
assign LUT_4[14052] = 32'b00000000000000000010100110100011;
assign LUT_4[14053] = 32'b11111111111111111011110010011011;
assign LUT_4[14054] = 32'b00000000000000000010000001000111;
assign LUT_4[14055] = 32'b11111111111111111011001100111111;
assign LUT_4[14056] = 32'b11111111111111111110110010011100;
assign LUT_4[14057] = 32'b11111111111111110111111110010100;
assign LUT_4[14058] = 32'b11111111111111111110001101000000;
assign LUT_4[14059] = 32'b11111111111111110111011000111000;
assign LUT_4[14060] = 32'b11111111111111111011110010111000;
assign LUT_4[14061] = 32'b11111111111111110100111110110000;
assign LUT_4[14062] = 32'b11111111111111111011001101011100;
assign LUT_4[14063] = 32'b11111111111111110100011001010100;
assign LUT_4[14064] = 32'b00000000000000000011010111110101;
assign LUT_4[14065] = 32'b11111111111111111100100011101101;
assign LUT_4[14066] = 32'b00000000000000000010110010011001;
assign LUT_4[14067] = 32'b11111111111111111011111110010001;
assign LUT_4[14068] = 32'b00000000000000000000011000010001;
assign LUT_4[14069] = 32'b11111111111111111001100100001001;
assign LUT_4[14070] = 32'b11111111111111111111110010110101;
assign LUT_4[14071] = 32'b11111111111111111000111110101101;
assign LUT_4[14072] = 32'b11111111111111111100100100001010;
assign LUT_4[14073] = 32'b11111111111111110101110000000010;
assign LUT_4[14074] = 32'b11111111111111111011111110101110;
assign LUT_4[14075] = 32'b11111111111111110101001010100110;
assign LUT_4[14076] = 32'b11111111111111111001100100100110;
assign LUT_4[14077] = 32'b11111111111111110010110000011110;
assign LUT_4[14078] = 32'b11111111111111111000111111001010;
assign LUT_4[14079] = 32'b11111111111111110010001011000010;
assign LUT_4[14080] = 32'b00000000000000001000001001000111;
assign LUT_4[14081] = 32'b00000000000000000001010100111111;
assign LUT_4[14082] = 32'b00000000000000000111100011101011;
assign LUT_4[14083] = 32'b00000000000000000000101111100011;
assign LUT_4[14084] = 32'b00000000000000000101001001100011;
assign LUT_4[14085] = 32'b11111111111111111110010101011011;
assign LUT_4[14086] = 32'b00000000000000000100100100000111;
assign LUT_4[14087] = 32'b11111111111111111101101111111111;
assign LUT_4[14088] = 32'b00000000000000000001010101011100;
assign LUT_4[14089] = 32'b11111111111111111010100001010100;
assign LUT_4[14090] = 32'b00000000000000000000110000000000;
assign LUT_4[14091] = 32'b11111111111111111001111011111000;
assign LUT_4[14092] = 32'b11111111111111111110010101111000;
assign LUT_4[14093] = 32'b11111111111111110111100001110000;
assign LUT_4[14094] = 32'b11111111111111111101110000011100;
assign LUT_4[14095] = 32'b11111111111111110110111100010100;
assign LUT_4[14096] = 32'b00000000000000000101111010110101;
assign LUT_4[14097] = 32'b11111111111111111111000110101101;
assign LUT_4[14098] = 32'b00000000000000000101010101011001;
assign LUT_4[14099] = 32'b11111111111111111110100001010001;
assign LUT_4[14100] = 32'b00000000000000000010111011010001;
assign LUT_4[14101] = 32'b11111111111111111100000111001001;
assign LUT_4[14102] = 32'b00000000000000000010010101110101;
assign LUT_4[14103] = 32'b11111111111111111011100001101101;
assign LUT_4[14104] = 32'b11111111111111111111000111001010;
assign LUT_4[14105] = 32'b11111111111111111000010011000010;
assign LUT_4[14106] = 32'b11111111111111111110100001101110;
assign LUT_4[14107] = 32'b11111111111111110111101101100110;
assign LUT_4[14108] = 32'b11111111111111111100000111100110;
assign LUT_4[14109] = 32'b11111111111111110101010011011110;
assign LUT_4[14110] = 32'b11111111111111111011100010001010;
assign LUT_4[14111] = 32'b11111111111111110100101110000010;
assign LUT_4[14112] = 32'b00000000000000000110100100001110;
assign LUT_4[14113] = 32'b11111111111111111111110000000110;
assign LUT_4[14114] = 32'b00000000000000000101111110110010;
assign LUT_4[14115] = 32'b11111111111111111111001010101010;
assign LUT_4[14116] = 32'b00000000000000000011100100101010;
assign LUT_4[14117] = 32'b11111111111111111100110000100010;
assign LUT_4[14118] = 32'b00000000000000000010111111001110;
assign LUT_4[14119] = 32'b11111111111111111100001011000110;
assign LUT_4[14120] = 32'b11111111111111111111110000100011;
assign LUT_4[14121] = 32'b11111111111111111000111100011011;
assign LUT_4[14122] = 32'b11111111111111111111001011000111;
assign LUT_4[14123] = 32'b11111111111111111000010110111111;
assign LUT_4[14124] = 32'b11111111111111111100110000111111;
assign LUT_4[14125] = 32'b11111111111111110101111100110111;
assign LUT_4[14126] = 32'b11111111111111111100001011100011;
assign LUT_4[14127] = 32'b11111111111111110101010111011011;
assign LUT_4[14128] = 32'b00000000000000000100010101111100;
assign LUT_4[14129] = 32'b11111111111111111101100001110100;
assign LUT_4[14130] = 32'b00000000000000000011110000100000;
assign LUT_4[14131] = 32'b11111111111111111100111100011000;
assign LUT_4[14132] = 32'b00000000000000000001010110011000;
assign LUT_4[14133] = 32'b11111111111111111010100010010000;
assign LUT_4[14134] = 32'b00000000000000000000110000111100;
assign LUT_4[14135] = 32'b11111111111111111001111100110100;
assign LUT_4[14136] = 32'b11111111111111111101100010010001;
assign LUT_4[14137] = 32'b11111111111111110110101110001001;
assign LUT_4[14138] = 32'b11111111111111111100111100110101;
assign LUT_4[14139] = 32'b11111111111111110110001000101101;
assign LUT_4[14140] = 32'b11111111111111111010100010101101;
assign LUT_4[14141] = 32'b11111111111111110011101110100101;
assign LUT_4[14142] = 32'b11111111111111111001111101010001;
assign LUT_4[14143] = 32'b11111111111111110011001001001001;
assign LUT_4[14144] = 32'b00000000000000001001100000011011;
assign LUT_4[14145] = 32'b00000000000000000010101100010011;
assign LUT_4[14146] = 32'b00000000000000001000111010111111;
assign LUT_4[14147] = 32'b00000000000000000010000110110111;
assign LUT_4[14148] = 32'b00000000000000000110100000110111;
assign LUT_4[14149] = 32'b11111111111111111111101100101111;
assign LUT_4[14150] = 32'b00000000000000000101111011011011;
assign LUT_4[14151] = 32'b11111111111111111111000111010011;
assign LUT_4[14152] = 32'b00000000000000000010101100110000;
assign LUT_4[14153] = 32'b11111111111111111011111000101000;
assign LUT_4[14154] = 32'b00000000000000000010000111010100;
assign LUT_4[14155] = 32'b11111111111111111011010011001100;
assign LUT_4[14156] = 32'b11111111111111111111101101001100;
assign LUT_4[14157] = 32'b11111111111111111000111001000100;
assign LUT_4[14158] = 32'b11111111111111111111000111110000;
assign LUT_4[14159] = 32'b11111111111111111000010011101000;
assign LUT_4[14160] = 32'b00000000000000000111010010001001;
assign LUT_4[14161] = 32'b00000000000000000000011110000001;
assign LUT_4[14162] = 32'b00000000000000000110101100101101;
assign LUT_4[14163] = 32'b11111111111111111111111000100101;
assign LUT_4[14164] = 32'b00000000000000000100010010100101;
assign LUT_4[14165] = 32'b11111111111111111101011110011101;
assign LUT_4[14166] = 32'b00000000000000000011101101001001;
assign LUT_4[14167] = 32'b11111111111111111100111001000001;
assign LUT_4[14168] = 32'b00000000000000000000011110011110;
assign LUT_4[14169] = 32'b11111111111111111001101010010110;
assign LUT_4[14170] = 32'b11111111111111111111111001000010;
assign LUT_4[14171] = 32'b11111111111111111001000100111010;
assign LUT_4[14172] = 32'b11111111111111111101011110111010;
assign LUT_4[14173] = 32'b11111111111111110110101010110010;
assign LUT_4[14174] = 32'b11111111111111111100111001011110;
assign LUT_4[14175] = 32'b11111111111111110110000101010110;
assign LUT_4[14176] = 32'b00000000000000000111111011100010;
assign LUT_4[14177] = 32'b00000000000000000001000111011010;
assign LUT_4[14178] = 32'b00000000000000000111010110000110;
assign LUT_4[14179] = 32'b00000000000000000000100001111110;
assign LUT_4[14180] = 32'b00000000000000000100111011111110;
assign LUT_4[14181] = 32'b11111111111111111110000111110110;
assign LUT_4[14182] = 32'b00000000000000000100010110100010;
assign LUT_4[14183] = 32'b11111111111111111101100010011010;
assign LUT_4[14184] = 32'b00000000000000000001000111110111;
assign LUT_4[14185] = 32'b11111111111111111010010011101111;
assign LUT_4[14186] = 32'b00000000000000000000100010011011;
assign LUT_4[14187] = 32'b11111111111111111001101110010011;
assign LUT_4[14188] = 32'b11111111111111111110001000010011;
assign LUT_4[14189] = 32'b11111111111111110111010100001011;
assign LUT_4[14190] = 32'b11111111111111111101100010110111;
assign LUT_4[14191] = 32'b11111111111111110110101110101111;
assign LUT_4[14192] = 32'b00000000000000000101101101010000;
assign LUT_4[14193] = 32'b11111111111111111110111001001000;
assign LUT_4[14194] = 32'b00000000000000000101000111110100;
assign LUT_4[14195] = 32'b11111111111111111110010011101100;
assign LUT_4[14196] = 32'b00000000000000000010101101101100;
assign LUT_4[14197] = 32'b11111111111111111011111001100100;
assign LUT_4[14198] = 32'b00000000000000000010001000010000;
assign LUT_4[14199] = 32'b11111111111111111011010100001000;
assign LUT_4[14200] = 32'b11111111111111111110111001100101;
assign LUT_4[14201] = 32'b11111111111111111000000101011101;
assign LUT_4[14202] = 32'b11111111111111111110010100001001;
assign LUT_4[14203] = 32'b11111111111111110111100000000001;
assign LUT_4[14204] = 32'b11111111111111111011111010000001;
assign LUT_4[14205] = 32'b11111111111111110101000101111001;
assign LUT_4[14206] = 32'b11111111111111111011010100100101;
assign LUT_4[14207] = 32'b11111111111111110100100000011101;
assign LUT_4[14208] = 32'b00000000000000001010101111001111;
assign LUT_4[14209] = 32'b00000000000000000011111011000111;
assign LUT_4[14210] = 32'b00000000000000001010001001110011;
assign LUT_4[14211] = 32'b00000000000000000011010101101011;
assign LUT_4[14212] = 32'b00000000000000000111101111101011;
assign LUT_4[14213] = 32'b00000000000000000000111011100011;
assign LUT_4[14214] = 32'b00000000000000000111001010001111;
assign LUT_4[14215] = 32'b00000000000000000000010110000111;
assign LUT_4[14216] = 32'b00000000000000000011111011100100;
assign LUT_4[14217] = 32'b11111111111111111101000111011100;
assign LUT_4[14218] = 32'b00000000000000000011010110001000;
assign LUT_4[14219] = 32'b11111111111111111100100010000000;
assign LUT_4[14220] = 32'b00000000000000000000111100000000;
assign LUT_4[14221] = 32'b11111111111111111010000111111000;
assign LUT_4[14222] = 32'b00000000000000000000010110100100;
assign LUT_4[14223] = 32'b11111111111111111001100010011100;
assign LUT_4[14224] = 32'b00000000000000001000100000111101;
assign LUT_4[14225] = 32'b00000000000000000001101100110101;
assign LUT_4[14226] = 32'b00000000000000000111111011100001;
assign LUT_4[14227] = 32'b00000000000000000001000111011001;
assign LUT_4[14228] = 32'b00000000000000000101100001011001;
assign LUT_4[14229] = 32'b11111111111111111110101101010001;
assign LUT_4[14230] = 32'b00000000000000000100111011111101;
assign LUT_4[14231] = 32'b11111111111111111110000111110101;
assign LUT_4[14232] = 32'b00000000000000000001101101010010;
assign LUT_4[14233] = 32'b11111111111111111010111001001010;
assign LUT_4[14234] = 32'b00000000000000000001000111110110;
assign LUT_4[14235] = 32'b11111111111111111010010011101110;
assign LUT_4[14236] = 32'b11111111111111111110101101101110;
assign LUT_4[14237] = 32'b11111111111111110111111001100110;
assign LUT_4[14238] = 32'b11111111111111111110001000010010;
assign LUT_4[14239] = 32'b11111111111111110111010100001010;
assign LUT_4[14240] = 32'b00000000000000001001001010010110;
assign LUT_4[14241] = 32'b00000000000000000010010110001110;
assign LUT_4[14242] = 32'b00000000000000001000100100111010;
assign LUT_4[14243] = 32'b00000000000000000001110000110010;
assign LUT_4[14244] = 32'b00000000000000000110001010110010;
assign LUT_4[14245] = 32'b11111111111111111111010110101010;
assign LUT_4[14246] = 32'b00000000000000000101100101010110;
assign LUT_4[14247] = 32'b11111111111111111110110001001110;
assign LUT_4[14248] = 32'b00000000000000000010010110101011;
assign LUT_4[14249] = 32'b11111111111111111011100010100011;
assign LUT_4[14250] = 32'b00000000000000000001110001001111;
assign LUT_4[14251] = 32'b11111111111111111010111101000111;
assign LUT_4[14252] = 32'b11111111111111111111010111000111;
assign LUT_4[14253] = 32'b11111111111111111000100010111111;
assign LUT_4[14254] = 32'b11111111111111111110110001101011;
assign LUT_4[14255] = 32'b11111111111111110111111101100011;
assign LUT_4[14256] = 32'b00000000000000000110111100000100;
assign LUT_4[14257] = 32'b00000000000000000000000111111100;
assign LUT_4[14258] = 32'b00000000000000000110010110101000;
assign LUT_4[14259] = 32'b11111111111111111111100010100000;
assign LUT_4[14260] = 32'b00000000000000000011111100100000;
assign LUT_4[14261] = 32'b11111111111111111101001000011000;
assign LUT_4[14262] = 32'b00000000000000000011010111000100;
assign LUT_4[14263] = 32'b11111111111111111100100010111100;
assign LUT_4[14264] = 32'b00000000000000000000001000011001;
assign LUT_4[14265] = 32'b11111111111111111001010100010001;
assign LUT_4[14266] = 32'b11111111111111111111100010111101;
assign LUT_4[14267] = 32'b11111111111111111000101110110101;
assign LUT_4[14268] = 32'b11111111111111111101001000110101;
assign LUT_4[14269] = 32'b11111111111111110110010100101101;
assign LUT_4[14270] = 32'b11111111111111111100100011011001;
assign LUT_4[14271] = 32'b11111111111111110101101111010001;
assign LUT_4[14272] = 32'b00000000000000001100000110100011;
assign LUT_4[14273] = 32'b00000000000000000101010010011011;
assign LUT_4[14274] = 32'b00000000000000001011100001000111;
assign LUT_4[14275] = 32'b00000000000000000100101100111111;
assign LUT_4[14276] = 32'b00000000000000001001000110111111;
assign LUT_4[14277] = 32'b00000000000000000010010010110111;
assign LUT_4[14278] = 32'b00000000000000001000100001100011;
assign LUT_4[14279] = 32'b00000000000000000001101101011011;
assign LUT_4[14280] = 32'b00000000000000000101010010111000;
assign LUT_4[14281] = 32'b11111111111111111110011110110000;
assign LUT_4[14282] = 32'b00000000000000000100101101011100;
assign LUT_4[14283] = 32'b11111111111111111101111001010100;
assign LUT_4[14284] = 32'b00000000000000000010010011010100;
assign LUT_4[14285] = 32'b11111111111111111011011111001100;
assign LUT_4[14286] = 32'b00000000000000000001101101111000;
assign LUT_4[14287] = 32'b11111111111111111010111001110000;
assign LUT_4[14288] = 32'b00000000000000001001111000010001;
assign LUT_4[14289] = 32'b00000000000000000011000100001001;
assign LUT_4[14290] = 32'b00000000000000001001010010110101;
assign LUT_4[14291] = 32'b00000000000000000010011110101101;
assign LUT_4[14292] = 32'b00000000000000000110111000101101;
assign LUT_4[14293] = 32'b00000000000000000000000100100101;
assign LUT_4[14294] = 32'b00000000000000000110010011010001;
assign LUT_4[14295] = 32'b11111111111111111111011111001001;
assign LUT_4[14296] = 32'b00000000000000000011000100100110;
assign LUT_4[14297] = 32'b11111111111111111100010000011110;
assign LUT_4[14298] = 32'b00000000000000000010011111001010;
assign LUT_4[14299] = 32'b11111111111111111011101011000010;
assign LUT_4[14300] = 32'b00000000000000000000000101000010;
assign LUT_4[14301] = 32'b11111111111111111001010000111010;
assign LUT_4[14302] = 32'b11111111111111111111011111100110;
assign LUT_4[14303] = 32'b11111111111111111000101011011110;
assign LUT_4[14304] = 32'b00000000000000001010100001101010;
assign LUT_4[14305] = 32'b00000000000000000011101101100010;
assign LUT_4[14306] = 32'b00000000000000001001111100001110;
assign LUT_4[14307] = 32'b00000000000000000011001000000110;
assign LUT_4[14308] = 32'b00000000000000000111100010000110;
assign LUT_4[14309] = 32'b00000000000000000000101101111110;
assign LUT_4[14310] = 32'b00000000000000000110111100101010;
assign LUT_4[14311] = 32'b00000000000000000000001000100010;
assign LUT_4[14312] = 32'b00000000000000000011101101111111;
assign LUT_4[14313] = 32'b11111111111111111100111001110111;
assign LUT_4[14314] = 32'b00000000000000000011001000100011;
assign LUT_4[14315] = 32'b11111111111111111100010100011011;
assign LUT_4[14316] = 32'b00000000000000000000101110011011;
assign LUT_4[14317] = 32'b11111111111111111001111010010011;
assign LUT_4[14318] = 32'b00000000000000000000001000111111;
assign LUT_4[14319] = 32'b11111111111111111001010100110111;
assign LUT_4[14320] = 32'b00000000000000001000010011011000;
assign LUT_4[14321] = 32'b00000000000000000001011111010000;
assign LUT_4[14322] = 32'b00000000000000000111101101111100;
assign LUT_4[14323] = 32'b00000000000000000000111001110100;
assign LUT_4[14324] = 32'b00000000000000000101010011110100;
assign LUT_4[14325] = 32'b11111111111111111110011111101100;
assign LUT_4[14326] = 32'b00000000000000000100101110011000;
assign LUT_4[14327] = 32'b11111111111111111101111010010000;
assign LUT_4[14328] = 32'b00000000000000000001011111101101;
assign LUT_4[14329] = 32'b11111111111111111010101011100101;
assign LUT_4[14330] = 32'b00000000000000000000111010010001;
assign LUT_4[14331] = 32'b11111111111111111010000110001001;
assign LUT_4[14332] = 32'b11111111111111111110100000001001;
assign LUT_4[14333] = 32'b11111111111111110111101100000001;
assign LUT_4[14334] = 32'b11111111111111111101111010101101;
assign LUT_4[14335] = 32'b11111111111111110111000110100101;
assign LUT_4[14336] = 32'b11111111111111111101111110000111;
assign LUT_4[14337] = 32'b11111111111111110111001001111111;
assign LUT_4[14338] = 32'b11111111111111111101011000101011;
assign LUT_4[14339] = 32'b11111111111111110110100100100011;
assign LUT_4[14340] = 32'b11111111111111111010111110100011;
assign LUT_4[14341] = 32'b11111111111111110100001010011011;
assign LUT_4[14342] = 32'b11111111111111111010011001000111;
assign LUT_4[14343] = 32'b11111111111111110011100100111111;
assign LUT_4[14344] = 32'b11111111111111110111001010011100;
assign LUT_4[14345] = 32'b11111111111111110000010110010100;
assign LUT_4[14346] = 32'b11111111111111110110100101000000;
assign LUT_4[14347] = 32'b11111111111111101111110000111000;
assign LUT_4[14348] = 32'b11111111111111110100001010111000;
assign LUT_4[14349] = 32'b11111111111111101101010110110000;
assign LUT_4[14350] = 32'b11111111111111110011100101011100;
assign LUT_4[14351] = 32'b11111111111111101100110001010100;
assign LUT_4[14352] = 32'b11111111111111111011101111110101;
assign LUT_4[14353] = 32'b11111111111111110100111011101101;
assign LUT_4[14354] = 32'b11111111111111111011001010011001;
assign LUT_4[14355] = 32'b11111111111111110100010110010001;
assign LUT_4[14356] = 32'b11111111111111111000110000010001;
assign LUT_4[14357] = 32'b11111111111111110001111100001001;
assign LUT_4[14358] = 32'b11111111111111111000001010110101;
assign LUT_4[14359] = 32'b11111111111111110001010110101101;
assign LUT_4[14360] = 32'b11111111111111110100111100001010;
assign LUT_4[14361] = 32'b11111111111111101110001000000010;
assign LUT_4[14362] = 32'b11111111111111110100010110101110;
assign LUT_4[14363] = 32'b11111111111111101101100010100110;
assign LUT_4[14364] = 32'b11111111111111110001111100100110;
assign LUT_4[14365] = 32'b11111111111111101011001000011110;
assign LUT_4[14366] = 32'b11111111111111110001010111001010;
assign LUT_4[14367] = 32'b11111111111111101010100011000010;
assign LUT_4[14368] = 32'b11111111111111111100011001001110;
assign LUT_4[14369] = 32'b11111111111111110101100101000110;
assign LUT_4[14370] = 32'b11111111111111111011110011110010;
assign LUT_4[14371] = 32'b11111111111111110100111111101010;
assign LUT_4[14372] = 32'b11111111111111111001011001101010;
assign LUT_4[14373] = 32'b11111111111111110010100101100010;
assign LUT_4[14374] = 32'b11111111111111111000110100001110;
assign LUT_4[14375] = 32'b11111111111111110010000000000110;
assign LUT_4[14376] = 32'b11111111111111110101100101100011;
assign LUT_4[14377] = 32'b11111111111111101110110001011011;
assign LUT_4[14378] = 32'b11111111111111110101000000000111;
assign LUT_4[14379] = 32'b11111111111111101110001011111111;
assign LUT_4[14380] = 32'b11111111111111110010100101111111;
assign LUT_4[14381] = 32'b11111111111111101011110001110111;
assign LUT_4[14382] = 32'b11111111111111110010000000100011;
assign LUT_4[14383] = 32'b11111111111111101011001100011011;
assign LUT_4[14384] = 32'b11111111111111111010001010111100;
assign LUT_4[14385] = 32'b11111111111111110011010110110100;
assign LUT_4[14386] = 32'b11111111111111111001100101100000;
assign LUT_4[14387] = 32'b11111111111111110010110001011000;
assign LUT_4[14388] = 32'b11111111111111110111001011011000;
assign LUT_4[14389] = 32'b11111111111111110000010111010000;
assign LUT_4[14390] = 32'b11111111111111110110100101111100;
assign LUT_4[14391] = 32'b11111111111111101111110001110100;
assign LUT_4[14392] = 32'b11111111111111110011010111010001;
assign LUT_4[14393] = 32'b11111111111111101100100011001001;
assign LUT_4[14394] = 32'b11111111111111110010110001110101;
assign LUT_4[14395] = 32'b11111111111111101011111101101101;
assign LUT_4[14396] = 32'b11111111111111110000010111101101;
assign LUT_4[14397] = 32'b11111111111111101001100011100101;
assign LUT_4[14398] = 32'b11111111111111101111110010010001;
assign LUT_4[14399] = 32'b11111111111111101000111110001001;
assign LUT_4[14400] = 32'b11111111111111111111010101011011;
assign LUT_4[14401] = 32'b11111111111111111000100001010011;
assign LUT_4[14402] = 32'b11111111111111111110101111111111;
assign LUT_4[14403] = 32'b11111111111111110111111011110111;
assign LUT_4[14404] = 32'b11111111111111111100010101110111;
assign LUT_4[14405] = 32'b11111111111111110101100001101111;
assign LUT_4[14406] = 32'b11111111111111111011110000011011;
assign LUT_4[14407] = 32'b11111111111111110100111100010011;
assign LUT_4[14408] = 32'b11111111111111111000100001110000;
assign LUT_4[14409] = 32'b11111111111111110001101101101000;
assign LUT_4[14410] = 32'b11111111111111110111111100010100;
assign LUT_4[14411] = 32'b11111111111111110001001000001100;
assign LUT_4[14412] = 32'b11111111111111110101100010001100;
assign LUT_4[14413] = 32'b11111111111111101110101110000100;
assign LUT_4[14414] = 32'b11111111111111110100111100110000;
assign LUT_4[14415] = 32'b11111111111111101110001000101000;
assign LUT_4[14416] = 32'b11111111111111111101000111001001;
assign LUT_4[14417] = 32'b11111111111111110110010011000001;
assign LUT_4[14418] = 32'b11111111111111111100100001101101;
assign LUT_4[14419] = 32'b11111111111111110101101101100101;
assign LUT_4[14420] = 32'b11111111111111111010000111100101;
assign LUT_4[14421] = 32'b11111111111111110011010011011101;
assign LUT_4[14422] = 32'b11111111111111111001100010001001;
assign LUT_4[14423] = 32'b11111111111111110010101110000001;
assign LUT_4[14424] = 32'b11111111111111110110010011011110;
assign LUT_4[14425] = 32'b11111111111111101111011111010110;
assign LUT_4[14426] = 32'b11111111111111110101101110000010;
assign LUT_4[14427] = 32'b11111111111111101110111001111010;
assign LUT_4[14428] = 32'b11111111111111110011010011111010;
assign LUT_4[14429] = 32'b11111111111111101100011111110010;
assign LUT_4[14430] = 32'b11111111111111110010101110011110;
assign LUT_4[14431] = 32'b11111111111111101011111010010110;
assign LUT_4[14432] = 32'b11111111111111111101110000100010;
assign LUT_4[14433] = 32'b11111111111111110110111100011010;
assign LUT_4[14434] = 32'b11111111111111111101001011000110;
assign LUT_4[14435] = 32'b11111111111111110110010110111110;
assign LUT_4[14436] = 32'b11111111111111111010110000111110;
assign LUT_4[14437] = 32'b11111111111111110011111100110110;
assign LUT_4[14438] = 32'b11111111111111111010001011100010;
assign LUT_4[14439] = 32'b11111111111111110011010111011010;
assign LUT_4[14440] = 32'b11111111111111110110111100110111;
assign LUT_4[14441] = 32'b11111111111111110000001000101111;
assign LUT_4[14442] = 32'b11111111111111110110010111011011;
assign LUT_4[14443] = 32'b11111111111111101111100011010011;
assign LUT_4[14444] = 32'b11111111111111110011111101010011;
assign LUT_4[14445] = 32'b11111111111111101101001001001011;
assign LUT_4[14446] = 32'b11111111111111110011010111110111;
assign LUT_4[14447] = 32'b11111111111111101100100011101111;
assign LUT_4[14448] = 32'b11111111111111111011100010010000;
assign LUT_4[14449] = 32'b11111111111111110100101110001000;
assign LUT_4[14450] = 32'b11111111111111111010111100110100;
assign LUT_4[14451] = 32'b11111111111111110100001000101100;
assign LUT_4[14452] = 32'b11111111111111111000100010101100;
assign LUT_4[14453] = 32'b11111111111111110001101110100100;
assign LUT_4[14454] = 32'b11111111111111110111111101010000;
assign LUT_4[14455] = 32'b11111111111111110001001001001000;
assign LUT_4[14456] = 32'b11111111111111110100101110100101;
assign LUT_4[14457] = 32'b11111111111111101101111010011101;
assign LUT_4[14458] = 32'b11111111111111110100001001001001;
assign LUT_4[14459] = 32'b11111111111111101101010101000001;
assign LUT_4[14460] = 32'b11111111111111110001101111000001;
assign LUT_4[14461] = 32'b11111111111111101010111010111001;
assign LUT_4[14462] = 32'b11111111111111110001001001100101;
assign LUT_4[14463] = 32'b11111111111111101010010101011101;
assign LUT_4[14464] = 32'b00000000000000000000100100001111;
assign LUT_4[14465] = 32'b11111111111111111001110000000111;
assign LUT_4[14466] = 32'b11111111111111111111111110110011;
assign LUT_4[14467] = 32'b11111111111111111001001010101011;
assign LUT_4[14468] = 32'b11111111111111111101100100101011;
assign LUT_4[14469] = 32'b11111111111111110110110000100011;
assign LUT_4[14470] = 32'b11111111111111111100111111001111;
assign LUT_4[14471] = 32'b11111111111111110110001011000111;
assign LUT_4[14472] = 32'b11111111111111111001110000100100;
assign LUT_4[14473] = 32'b11111111111111110010111100011100;
assign LUT_4[14474] = 32'b11111111111111111001001011001000;
assign LUT_4[14475] = 32'b11111111111111110010010111000000;
assign LUT_4[14476] = 32'b11111111111111110110110001000000;
assign LUT_4[14477] = 32'b11111111111111101111111100111000;
assign LUT_4[14478] = 32'b11111111111111110110001011100100;
assign LUT_4[14479] = 32'b11111111111111101111010111011100;
assign LUT_4[14480] = 32'b11111111111111111110010101111101;
assign LUT_4[14481] = 32'b11111111111111110111100001110101;
assign LUT_4[14482] = 32'b11111111111111111101110000100001;
assign LUT_4[14483] = 32'b11111111111111110110111100011001;
assign LUT_4[14484] = 32'b11111111111111111011010110011001;
assign LUT_4[14485] = 32'b11111111111111110100100010010001;
assign LUT_4[14486] = 32'b11111111111111111010110000111101;
assign LUT_4[14487] = 32'b11111111111111110011111100110101;
assign LUT_4[14488] = 32'b11111111111111110111100010010010;
assign LUT_4[14489] = 32'b11111111111111110000101110001010;
assign LUT_4[14490] = 32'b11111111111111110110111100110110;
assign LUT_4[14491] = 32'b11111111111111110000001000101110;
assign LUT_4[14492] = 32'b11111111111111110100100010101110;
assign LUT_4[14493] = 32'b11111111111111101101101110100110;
assign LUT_4[14494] = 32'b11111111111111110011111101010010;
assign LUT_4[14495] = 32'b11111111111111101101001001001010;
assign LUT_4[14496] = 32'b11111111111111111110111111010110;
assign LUT_4[14497] = 32'b11111111111111111000001011001110;
assign LUT_4[14498] = 32'b11111111111111111110011001111010;
assign LUT_4[14499] = 32'b11111111111111110111100101110010;
assign LUT_4[14500] = 32'b11111111111111111011111111110010;
assign LUT_4[14501] = 32'b11111111111111110101001011101010;
assign LUT_4[14502] = 32'b11111111111111111011011010010110;
assign LUT_4[14503] = 32'b11111111111111110100100110001110;
assign LUT_4[14504] = 32'b11111111111111111000001011101011;
assign LUT_4[14505] = 32'b11111111111111110001010111100011;
assign LUT_4[14506] = 32'b11111111111111110111100110001111;
assign LUT_4[14507] = 32'b11111111111111110000110010000111;
assign LUT_4[14508] = 32'b11111111111111110101001100000111;
assign LUT_4[14509] = 32'b11111111111111101110010111111111;
assign LUT_4[14510] = 32'b11111111111111110100100110101011;
assign LUT_4[14511] = 32'b11111111111111101101110010100011;
assign LUT_4[14512] = 32'b11111111111111111100110001000100;
assign LUT_4[14513] = 32'b11111111111111110101111100111100;
assign LUT_4[14514] = 32'b11111111111111111100001011101000;
assign LUT_4[14515] = 32'b11111111111111110101010111100000;
assign LUT_4[14516] = 32'b11111111111111111001110001100000;
assign LUT_4[14517] = 32'b11111111111111110010111101011000;
assign LUT_4[14518] = 32'b11111111111111111001001100000100;
assign LUT_4[14519] = 32'b11111111111111110010010111111100;
assign LUT_4[14520] = 32'b11111111111111110101111101011001;
assign LUT_4[14521] = 32'b11111111111111101111001001010001;
assign LUT_4[14522] = 32'b11111111111111110101010111111101;
assign LUT_4[14523] = 32'b11111111111111101110100011110101;
assign LUT_4[14524] = 32'b11111111111111110010111101110101;
assign LUT_4[14525] = 32'b11111111111111101100001001101101;
assign LUT_4[14526] = 32'b11111111111111110010011000011001;
assign LUT_4[14527] = 32'b11111111111111101011100100010001;
assign LUT_4[14528] = 32'b00000000000000000001111011100011;
assign LUT_4[14529] = 32'b11111111111111111011000111011011;
assign LUT_4[14530] = 32'b00000000000000000001010110000111;
assign LUT_4[14531] = 32'b11111111111111111010100001111111;
assign LUT_4[14532] = 32'b11111111111111111110111011111111;
assign LUT_4[14533] = 32'b11111111111111111000000111110111;
assign LUT_4[14534] = 32'b11111111111111111110010110100011;
assign LUT_4[14535] = 32'b11111111111111110111100010011011;
assign LUT_4[14536] = 32'b11111111111111111011000111111000;
assign LUT_4[14537] = 32'b11111111111111110100010011110000;
assign LUT_4[14538] = 32'b11111111111111111010100010011100;
assign LUT_4[14539] = 32'b11111111111111110011101110010100;
assign LUT_4[14540] = 32'b11111111111111111000001000010100;
assign LUT_4[14541] = 32'b11111111111111110001010100001100;
assign LUT_4[14542] = 32'b11111111111111110111100010111000;
assign LUT_4[14543] = 32'b11111111111111110000101110110000;
assign LUT_4[14544] = 32'b11111111111111111111101101010001;
assign LUT_4[14545] = 32'b11111111111111111000111001001001;
assign LUT_4[14546] = 32'b11111111111111111111000111110101;
assign LUT_4[14547] = 32'b11111111111111111000010011101101;
assign LUT_4[14548] = 32'b11111111111111111100101101101101;
assign LUT_4[14549] = 32'b11111111111111110101111001100101;
assign LUT_4[14550] = 32'b11111111111111111100001000010001;
assign LUT_4[14551] = 32'b11111111111111110101010100001001;
assign LUT_4[14552] = 32'b11111111111111111000111001100110;
assign LUT_4[14553] = 32'b11111111111111110010000101011110;
assign LUT_4[14554] = 32'b11111111111111111000010100001010;
assign LUT_4[14555] = 32'b11111111111111110001100000000010;
assign LUT_4[14556] = 32'b11111111111111110101111010000010;
assign LUT_4[14557] = 32'b11111111111111101111000101111010;
assign LUT_4[14558] = 32'b11111111111111110101010100100110;
assign LUT_4[14559] = 32'b11111111111111101110100000011110;
assign LUT_4[14560] = 32'b00000000000000000000010110101010;
assign LUT_4[14561] = 32'b11111111111111111001100010100010;
assign LUT_4[14562] = 32'b11111111111111111111110001001110;
assign LUT_4[14563] = 32'b11111111111111111000111101000110;
assign LUT_4[14564] = 32'b11111111111111111101010111000110;
assign LUT_4[14565] = 32'b11111111111111110110100010111110;
assign LUT_4[14566] = 32'b11111111111111111100110001101010;
assign LUT_4[14567] = 32'b11111111111111110101111101100010;
assign LUT_4[14568] = 32'b11111111111111111001100010111111;
assign LUT_4[14569] = 32'b11111111111111110010101110110111;
assign LUT_4[14570] = 32'b11111111111111111000111101100011;
assign LUT_4[14571] = 32'b11111111111111110010001001011011;
assign LUT_4[14572] = 32'b11111111111111110110100011011011;
assign LUT_4[14573] = 32'b11111111111111101111101111010011;
assign LUT_4[14574] = 32'b11111111111111110101111101111111;
assign LUT_4[14575] = 32'b11111111111111101111001001110111;
assign LUT_4[14576] = 32'b11111111111111111110001000011000;
assign LUT_4[14577] = 32'b11111111111111110111010100010000;
assign LUT_4[14578] = 32'b11111111111111111101100010111100;
assign LUT_4[14579] = 32'b11111111111111110110101110110100;
assign LUT_4[14580] = 32'b11111111111111111011001000110100;
assign LUT_4[14581] = 32'b11111111111111110100010100101100;
assign LUT_4[14582] = 32'b11111111111111111010100011011000;
assign LUT_4[14583] = 32'b11111111111111110011101111010000;
assign LUT_4[14584] = 32'b11111111111111110111010100101101;
assign LUT_4[14585] = 32'b11111111111111110000100000100101;
assign LUT_4[14586] = 32'b11111111111111110110101111010001;
assign LUT_4[14587] = 32'b11111111111111101111111011001001;
assign LUT_4[14588] = 32'b11111111111111110100010101001001;
assign LUT_4[14589] = 32'b11111111111111101101100001000001;
assign LUT_4[14590] = 32'b11111111111111110011101111101101;
assign LUT_4[14591] = 32'b11111111111111101100111011100101;
assign LUT_4[14592] = 32'b00000000000000000010111001101010;
assign LUT_4[14593] = 32'b11111111111111111100000101100010;
assign LUT_4[14594] = 32'b00000000000000000010010100001110;
assign LUT_4[14595] = 32'b11111111111111111011100000000110;
assign LUT_4[14596] = 32'b11111111111111111111111010000110;
assign LUT_4[14597] = 32'b11111111111111111001000101111110;
assign LUT_4[14598] = 32'b11111111111111111111010100101010;
assign LUT_4[14599] = 32'b11111111111111111000100000100010;
assign LUT_4[14600] = 32'b11111111111111111100000101111111;
assign LUT_4[14601] = 32'b11111111111111110101010001110111;
assign LUT_4[14602] = 32'b11111111111111111011100000100011;
assign LUT_4[14603] = 32'b11111111111111110100101100011011;
assign LUT_4[14604] = 32'b11111111111111111001000110011011;
assign LUT_4[14605] = 32'b11111111111111110010010010010011;
assign LUT_4[14606] = 32'b11111111111111111000100000111111;
assign LUT_4[14607] = 32'b11111111111111110001101100110111;
assign LUT_4[14608] = 32'b00000000000000000000101011011000;
assign LUT_4[14609] = 32'b11111111111111111001110111010000;
assign LUT_4[14610] = 32'b00000000000000000000000101111100;
assign LUT_4[14611] = 32'b11111111111111111001010001110100;
assign LUT_4[14612] = 32'b11111111111111111101101011110100;
assign LUT_4[14613] = 32'b11111111111111110110110111101100;
assign LUT_4[14614] = 32'b11111111111111111101000110011000;
assign LUT_4[14615] = 32'b11111111111111110110010010010000;
assign LUT_4[14616] = 32'b11111111111111111001110111101101;
assign LUT_4[14617] = 32'b11111111111111110011000011100101;
assign LUT_4[14618] = 32'b11111111111111111001010010010001;
assign LUT_4[14619] = 32'b11111111111111110010011110001001;
assign LUT_4[14620] = 32'b11111111111111110110111000001001;
assign LUT_4[14621] = 32'b11111111111111110000000100000001;
assign LUT_4[14622] = 32'b11111111111111110110010010101101;
assign LUT_4[14623] = 32'b11111111111111101111011110100101;
assign LUT_4[14624] = 32'b00000000000000000001010100110001;
assign LUT_4[14625] = 32'b11111111111111111010100000101001;
assign LUT_4[14626] = 32'b00000000000000000000101111010101;
assign LUT_4[14627] = 32'b11111111111111111001111011001101;
assign LUT_4[14628] = 32'b11111111111111111110010101001101;
assign LUT_4[14629] = 32'b11111111111111110111100001000101;
assign LUT_4[14630] = 32'b11111111111111111101101111110001;
assign LUT_4[14631] = 32'b11111111111111110110111011101001;
assign LUT_4[14632] = 32'b11111111111111111010100001000110;
assign LUT_4[14633] = 32'b11111111111111110011101100111110;
assign LUT_4[14634] = 32'b11111111111111111001111011101010;
assign LUT_4[14635] = 32'b11111111111111110011000111100010;
assign LUT_4[14636] = 32'b11111111111111110111100001100010;
assign LUT_4[14637] = 32'b11111111111111110000101101011010;
assign LUT_4[14638] = 32'b11111111111111110110111100000110;
assign LUT_4[14639] = 32'b11111111111111110000000111111110;
assign LUT_4[14640] = 32'b11111111111111111111000110011111;
assign LUT_4[14641] = 32'b11111111111111111000010010010111;
assign LUT_4[14642] = 32'b11111111111111111110100001000011;
assign LUT_4[14643] = 32'b11111111111111110111101100111011;
assign LUT_4[14644] = 32'b11111111111111111100000110111011;
assign LUT_4[14645] = 32'b11111111111111110101010010110011;
assign LUT_4[14646] = 32'b11111111111111111011100001011111;
assign LUT_4[14647] = 32'b11111111111111110100101101010111;
assign LUT_4[14648] = 32'b11111111111111111000010010110100;
assign LUT_4[14649] = 32'b11111111111111110001011110101100;
assign LUT_4[14650] = 32'b11111111111111110111101101011000;
assign LUT_4[14651] = 32'b11111111111111110000111001010000;
assign LUT_4[14652] = 32'b11111111111111110101010011010000;
assign LUT_4[14653] = 32'b11111111111111101110011111001000;
assign LUT_4[14654] = 32'b11111111111111110100101101110100;
assign LUT_4[14655] = 32'b11111111111111101101111001101100;
assign LUT_4[14656] = 32'b00000000000000000100010000111110;
assign LUT_4[14657] = 32'b11111111111111111101011100110110;
assign LUT_4[14658] = 32'b00000000000000000011101011100010;
assign LUT_4[14659] = 32'b11111111111111111100110111011010;
assign LUT_4[14660] = 32'b00000000000000000001010001011010;
assign LUT_4[14661] = 32'b11111111111111111010011101010010;
assign LUT_4[14662] = 32'b00000000000000000000101011111110;
assign LUT_4[14663] = 32'b11111111111111111001110111110110;
assign LUT_4[14664] = 32'b11111111111111111101011101010011;
assign LUT_4[14665] = 32'b11111111111111110110101001001011;
assign LUT_4[14666] = 32'b11111111111111111100110111110111;
assign LUT_4[14667] = 32'b11111111111111110110000011101111;
assign LUT_4[14668] = 32'b11111111111111111010011101101111;
assign LUT_4[14669] = 32'b11111111111111110011101001100111;
assign LUT_4[14670] = 32'b11111111111111111001111000010011;
assign LUT_4[14671] = 32'b11111111111111110011000100001011;
assign LUT_4[14672] = 32'b00000000000000000010000010101100;
assign LUT_4[14673] = 32'b11111111111111111011001110100100;
assign LUT_4[14674] = 32'b00000000000000000001011101010000;
assign LUT_4[14675] = 32'b11111111111111111010101001001000;
assign LUT_4[14676] = 32'b11111111111111111111000011001000;
assign LUT_4[14677] = 32'b11111111111111111000001111000000;
assign LUT_4[14678] = 32'b11111111111111111110011101101100;
assign LUT_4[14679] = 32'b11111111111111110111101001100100;
assign LUT_4[14680] = 32'b11111111111111111011001111000001;
assign LUT_4[14681] = 32'b11111111111111110100011010111001;
assign LUT_4[14682] = 32'b11111111111111111010101001100101;
assign LUT_4[14683] = 32'b11111111111111110011110101011101;
assign LUT_4[14684] = 32'b11111111111111111000001111011101;
assign LUT_4[14685] = 32'b11111111111111110001011011010101;
assign LUT_4[14686] = 32'b11111111111111110111101010000001;
assign LUT_4[14687] = 32'b11111111111111110000110101111001;
assign LUT_4[14688] = 32'b00000000000000000010101100000101;
assign LUT_4[14689] = 32'b11111111111111111011110111111101;
assign LUT_4[14690] = 32'b00000000000000000010000110101001;
assign LUT_4[14691] = 32'b11111111111111111011010010100001;
assign LUT_4[14692] = 32'b11111111111111111111101100100001;
assign LUT_4[14693] = 32'b11111111111111111000111000011001;
assign LUT_4[14694] = 32'b11111111111111111111000111000101;
assign LUT_4[14695] = 32'b11111111111111111000010010111101;
assign LUT_4[14696] = 32'b11111111111111111011111000011010;
assign LUT_4[14697] = 32'b11111111111111110101000100010010;
assign LUT_4[14698] = 32'b11111111111111111011010010111110;
assign LUT_4[14699] = 32'b11111111111111110100011110110110;
assign LUT_4[14700] = 32'b11111111111111111000111000110110;
assign LUT_4[14701] = 32'b11111111111111110010000100101110;
assign LUT_4[14702] = 32'b11111111111111111000010011011010;
assign LUT_4[14703] = 32'b11111111111111110001011111010010;
assign LUT_4[14704] = 32'b00000000000000000000011101110011;
assign LUT_4[14705] = 32'b11111111111111111001101001101011;
assign LUT_4[14706] = 32'b11111111111111111111111000010111;
assign LUT_4[14707] = 32'b11111111111111111001000100001111;
assign LUT_4[14708] = 32'b11111111111111111101011110001111;
assign LUT_4[14709] = 32'b11111111111111110110101010000111;
assign LUT_4[14710] = 32'b11111111111111111100111000110011;
assign LUT_4[14711] = 32'b11111111111111110110000100101011;
assign LUT_4[14712] = 32'b11111111111111111001101010001000;
assign LUT_4[14713] = 32'b11111111111111110010110110000000;
assign LUT_4[14714] = 32'b11111111111111111001000100101100;
assign LUT_4[14715] = 32'b11111111111111110010010000100100;
assign LUT_4[14716] = 32'b11111111111111110110101010100100;
assign LUT_4[14717] = 32'b11111111111111101111110110011100;
assign LUT_4[14718] = 32'b11111111111111110110000101001000;
assign LUT_4[14719] = 32'b11111111111111101111010001000000;
assign LUT_4[14720] = 32'b00000000000000000101011111110010;
assign LUT_4[14721] = 32'b11111111111111111110101011101010;
assign LUT_4[14722] = 32'b00000000000000000100111010010110;
assign LUT_4[14723] = 32'b11111111111111111110000110001110;
assign LUT_4[14724] = 32'b00000000000000000010100000001110;
assign LUT_4[14725] = 32'b11111111111111111011101100000110;
assign LUT_4[14726] = 32'b00000000000000000001111010110010;
assign LUT_4[14727] = 32'b11111111111111111011000110101010;
assign LUT_4[14728] = 32'b11111111111111111110101100000111;
assign LUT_4[14729] = 32'b11111111111111110111110111111111;
assign LUT_4[14730] = 32'b11111111111111111110000110101011;
assign LUT_4[14731] = 32'b11111111111111110111010010100011;
assign LUT_4[14732] = 32'b11111111111111111011101100100011;
assign LUT_4[14733] = 32'b11111111111111110100111000011011;
assign LUT_4[14734] = 32'b11111111111111111011000111000111;
assign LUT_4[14735] = 32'b11111111111111110100010010111111;
assign LUT_4[14736] = 32'b00000000000000000011010001100000;
assign LUT_4[14737] = 32'b11111111111111111100011101011000;
assign LUT_4[14738] = 32'b00000000000000000010101100000100;
assign LUT_4[14739] = 32'b11111111111111111011110111111100;
assign LUT_4[14740] = 32'b00000000000000000000010001111100;
assign LUT_4[14741] = 32'b11111111111111111001011101110100;
assign LUT_4[14742] = 32'b11111111111111111111101100100000;
assign LUT_4[14743] = 32'b11111111111111111000111000011000;
assign LUT_4[14744] = 32'b11111111111111111100011101110101;
assign LUT_4[14745] = 32'b11111111111111110101101001101101;
assign LUT_4[14746] = 32'b11111111111111111011111000011001;
assign LUT_4[14747] = 32'b11111111111111110101000100010001;
assign LUT_4[14748] = 32'b11111111111111111001011110010001;
assign LUT_4[14749] = 32'b11111111111111110010101010001001;
assign LUT_4[14750] = 32'b11111111111111111000111000110101;
assign LUT_4[14751] = 32'b11111111111111110010000100101101;
assign LUT_4[14752] = 32'b00000000000000000011111010111001;
assign LUT_4[14753] = 32'b11111111111111111101000110110001;
assign LUT_4[14754] = 32'b00000000000000000011010101011101;
assign LUT_4[14755] = 32'b11111111111111111100100001010101;
assign LUT_4[14756] = 32'b00000000000000000000111011010101;
assign LUT_4[14757] = 32'b11111111111111111010000111001101;
assign LUT_4[14758] = 32'b00000000000000000000010101111001;
assign LUT_4[14759] = 32'b11111111111111111001100001110001;
assign LUT_4[14760] = 32'b11111111111111111101000111001110;
assign LUT_4[14761] = 32'b11111111111111110110010011000110;
assign LUT_4[14762] = 32'b11111111111111111100100001110010;
assign LUT_4[14763] = 32'b11111111111111110101101101101010;
assign LUT_4[14764] = 32'b11111111111111111010000111101010;
assign LUT_4[14765] = 32'b11111111111111110011010011100010;
assign LUT_4[14766] = 32'b11111111111111111001100010001110;
assign LUT_4[14767] = 32'b11111111111111110010101110000110;
assign LUT_4[14768] = 32'b00000000000000000001101100100111;
assign LUT_4[14769] = 32'b11111111111111111010111000011111;
assign LUT_4[14770] = 32'b00000000000000000001000111001011;
assign LUT_4[14771] = 32'b11111111111111111010010011000011;
assign LUT_4[14772] = 32'b11111111111111111110101101000011;
assign LUT_4[14773] = 32'b11111111111111110111111000111011;
assign LUT_4[14774] = 32'b11111111111111111110000111100111;
assign LUT_4[14775] = 32'b11111111111111110111010011011111;
assign LUT_4[14776] = 32'b11111111111111111010111000111100;
assign LUT_4[14777] = 32'b11111111111111110100000100110100;
assign LUT_4[14778] = 32'b11111111111111111010010011100000;
assign LUT_4[14779] = 32'b11111111111111110011011111011000;
assign LUT_4[14780] = 32'b11111111111111110111111001011000;
assign LUT_4[14781] = 32'b11111111111111110001000101010000;
assign LUT_4[14782] = 32'b11111111111111110111010011111100;
assign LUT_4[14783] = 32'b11111111111111110000011111110100;
assign LUT_4[14784] = 32'b00000000000000000110110111000110;
assign LUT_4[14785] = 32'b00000000000000000000000010111110;
assign LUT_4[14786] = 32'b00000000000000000110010001101010;
assign LUT_4[14787] = 32'b11111111111111111111011101100010;
assign LUT_4[14788] = 32'b00000000000000000011110111100010;
assign LUT_4[14789] = 32'b11111111111111111101000011011010;
assign LUT_4[14790] = 32'b00000000000000000011010010000110;
assign LUT_4[14791] = 32'b11111111111111111100011101111110;
assign LUT_4[14792] = 32'b00000000000000000000000011011011;
assign LUT_4[14793] = 32'b11111111111111111001001111010011;
assign LUT_4[14794] = 32'b11111111111111111111011101111111;
assign LUT_4[14795] = 32'b11111111111111111000101001110111;
assign LUT_4[14796] = 32'b11111111111111111101000011110111;
assign LUT_4[14797] = 32'b11111111111111110110001111101111;
assign LUT_4[14798] = 32'b11111111111111111100011110011011;
assign LUT_4[14799] = 32'b11111111111111110101101010010011;
assign LUT_4[14800] = 32'b00000000000000000100101000110100;
assign LUT_4[14801] = 32'b11111111111111111101110100101100;
assign LUT_4[14802] = 32'b00000000000000000100000011011000;
assign LUT_4[14803] = 32'b11111111111111111101001111010000;
assign LUT_4[14804] = 32'b00000000000000000001101001010000;
assign LUT_4[14805] = 32'b11111111111111111010110101001000;
assign LUT_4[14806] = 32'b00000000000000000001000011110100;
assign LUT_4[14807] = 32'b11111111111111111010001111101100;
assign LUT_4[14808] = 32'b11111111111111111101110101001001;
assign LUT_4[14809] = 32'b11111111111111110111000001000001;
assign LUT_4[14810] = 32'b11111111111111111101001111101101;
assign LUT_4[14811] = 32'b11111111111111110110011011100101;
assign LUT_4[14812] = 32'b11111111111111111010110101100101;
assign LUT_4[14813] = 32'b11111111111111110100000001011101;
assign LUT_4[14814] = 32'b11111111111111111010010000001001;
assign LUT_4[14815] = 32'b11111111111111110011011100000001;
assign LUT_4[14816] = 32'b00000000000000000101010010001101;
assign LUT_4[14817] = 32'b11111111111111111110011110000101;
assign LUT_4[14818] = 32'b00000000000000000100101100110001;
assign LUT_4[14819] = 32'b11111111111111111101111000101001;
assign LUT_4[14820] = 32'b00000000000000000010010010101001;
assign LUT_4[14821] = 32'b11111111111111111011011110100001;
assign LUT_4[14822] = 32'b00000000000000000001101101001101;
assign LUT_4[14823] = 32'b11111111111111111010111001000101;
assign LUT_4[14824] = 32'b11111111111111111110011110100010;
assign LUT_4[14825] = 32'b11111111111111110111101010011010;
assign LUT_4[14826] = 32'b11111111111111111101111001000110;
assign LUT_4[14827] = 32'b11111111111111110111000100111110;
assign LUT_4[14828] = 32'b11111111111111111011011110111110;
assign LUT_4[14829] = 32'b11111111111111110100101010110110;
assign LUT_4[14830] = 32'b11111111111111111010111001100010;
assign LUT_4[14831] = 32'b11111111111111110100000101011010;
assign LUT_4[14832] = 32'b00000000000000000011000011111011;
assign LUT_4[14833] = 32'b11111111111111111100001111110011;
assign LUT_4[14834] = 32'b00000000000000000010011110011111;
assign LUT_4[14835] = 32'b11111111111111111011101010010111;
assign LUT_4[14836] = 32'b00000000000000000000000100010111;
assign LUT_4[14837] = 32'b11111111111111111001010000001111;
assign LUT_4[14838] = 32'b11111111111111111111011110111011;
assign LUT_4[14839] = 32'b11111111111111111000101010110011;
assign LUT_4[14840] = 32'b11111111111111111100010000010000;
assign LUT_4[14841] = 32'b11111111111111110101011100001000;
assign LUT_4[14842] = 32'b11111111111111111011101010110100;
assign LUT_4[14843] = 32'b11111111111111110100110110101100;
assign LUT_4[14844] = 32'b11111111111111111001010000101100;
assign LUT_4[14845] = 32'b11111111111111110010011100100100;
assign LUT_4[14846] = 32'b11111111111111111000101011010000;
assign LUT_4[14847] = 32'b11111111111111110001110111001000;
assign LUT_4[14848] = 32'b11111111111111111101000010001111;
assign LUT_4[14849] = 32'b11111111111111110110001110000111;
assign LUT_4[14850] = 32'b11111111111111111100011100110011;
assign LUT_4[14851] = 32'b11111111111111110101101000101011;
assign LUT_4[14852] = 32'b11111111111111111010000010101011;
assign LUT_4[14853] = 32'b11111111111111110011001110100011;
assign LUT_4[14854] = 32'b11111111111111111001011101001111;
assign LUT_4[14855] = 32'b11111111111111110010101001000111;
assign LUT_4[14856] = 32'b11111111111111110110001110100100;
assign LUT_4[14857] = 32'b11111111111111101111011010011100;
assign LUT_4[14858] = 32'b11111111111111110101101001001000;
assign LUT_4[14859] = 32'b11111111111111101110110101000000;
assign LUT_4[14860] = 32'b11111111111111110011001111000000;
assign LUT_4[14861] = 32'b11111111111111101100011010111000;
assign LUT_4[14862] = 32'b11111111111111110010101001100100;
assign LUT_4[14863] = 32'b11111111111111101011110101011100;
assign LUT_4[14864] = 32'b11111111111111111010110011111101;
assign LUT_4[14865] = 32'b11111111111111110011111111110101;
assign LUT_4[14866] = 32'b11111111111111111010001110100001;
assign LUT_4[14867] = 32'b11111111111111110011011010011001;
assign LUT_4[14868] = 32'b11111111111111110111110100011001;
assign LUT_4[14869] = 32'b11111111111111110001000000010001;
assign LUT_4[14870] = 32'b11111111111111110111001110111101;
assign LUT_4[14871] = 32'b11111111111111110000011010110101;
assign LUT_4[14872] = 32'b11111111111111110100000000010010;
assign LUT_4[14873] = 32'b11111111111111101101001100001010;
assign LUT_4[14874] = 32'b11111111111111110011011010110110;
assign LUT_4[14875] = 32'b11111111111111101100100110101110;
assign LUT_4[14876] = 32'b11111111111111110001000000101110;
assign LUT_4[14877] = 32'b11111111111111101010001100100110;
assign LUT_4[14878] = 32'b11111111111111110000011011010010;
assign LUT_4[14879] = 32'b11111111111111101001100111001010;
assign LUT_4[14880] = 32'b11111111111111111011011101010110;
assign LUT_4[14881] = 32'b11111111111111110100101001001110;
assign LUT_4[14882] = 32'b11111111111111111010110111111010;
assign LUT_4[14883] = 32'b11111111111111110100000011110010;
assign LUT_4[14884] = 32'b11111111111111111000011101110010;
assign LUT_4[14885] = 32'b11111111111111110001101001101010;
assign LUT_4[14886] = 32'b11111111111111110111111000010110;
assign LUT_4[14887] = 32'b11111111111111110001000100001110;
assign LUT_4[14888] = 32'b11111111111111110100101001101011;
assign LUT_4[14889] = 32'b11111111111111101101110101100011;
assign LUT_4[14890] = 32'b11111111111111110100000100001111;
assign LUT_4[14891] = 32'b11111111111111101101010000000111;
assign LUT_4[14892] = 32'b11111111111111110001101010000111;
assign LUT_4[14893] = 32'b11111111111111101010110101111111;
assign LUT_4[14894] = 32'b11111111111111110001000100101011;
assign LUT_4[14895] = 32'b11111111111111101010010000100011;
assign LUT_4[14896] = 32'b11111111111111111001001111000100;
assign LUT_4[14897] = 32'b11111111111111110010011010111100;
assign LUT_4[14898] = 32'b11111111111111111000101001101000;
assign LUT_4[14899] = 32'b11111111111111110001110101100000;
assign LUT_4[14900] = 32'b11111111111111110110001111100000;
assign LUT_4[14901] = 32'b11111111111111101111011011011000;
assign LUT_4[14902] = 32'b11111111111111110101101010000100;
assign LUT_4[14903] = 32'b11111111111111101110110101111100;
assign LUT_4[14904] = 32'b11111111111111110010011011011001;
assign LUT_4[14905] = 32'b11111111111111101011100111010001;
assign LUT_4[14906] = 32'b11111111111111110001110101111101;
assign LUT_4[14907] = 32'b11111111111111101011000001110101;
assign LUT_4[14908] = 32'b11111111111111101111011011110101;
assign LUT_4[14909] = 32'b11111111111111101000100111101101;
assign LUT_4[14910] = 32'b11111111111111101110110110011001;
assign LUT_4[14911] = 32'b11111111111111101000000010010001;
assign LUT_4[14912] = 32'b11111111111111111110011001100011;
assign LUT_4[14913] = 32'b11111111111111110111100101011011;
assign LUT_4[14914] = 32'b11111111111111111101110100000111;
assign LUT_4[14915] = 32'b11111111111111110110111111111111;
assign LUT_4[14916] = 32'b11111111111111111011011001111111;
assign LUT_4[14917] = 32'b11111111111111110100100101110111;
assign LUT_4[14918] = 32'b11111111111111111010110100100011;
assign LUT_4[14919] = 32'b11111111111111110100000000011011;
assign LUT_4[14920] = 32'b11111111111111110111100101111000;
assign LUT_4[14921] = 32'b11111111111111110000110001110000;
assign LUT_4[14922] = 32'b11111111111111110111000000011100;
assign LUT_4[14923] = 32'b11111111111111110000001100010100;
assign LUT_4[14924] = 32'b11111111111111110100100110010100;
assign LUT_4[14925] = 32'b11111111111111101101110010001100;
assign LUT_4[14926] = 32'b11111111111111110100000000111000;
assign LUT_4[14927] = 32'b11111111111111101101001100110000;
assign LUT_4[14928] = 32'b11111111111111111100001011010001;
assign LUT_4[14929] = 32'b11111111111111110101010111001001;
assign LUT_4[14930] = 32'b11111111111111111011100101110101;
assign LUT_4[14931] = 32'b11111111111111110100110001101101;
assign LUT_4[14932] = 32'b11111111111111111001001011101101;
assign LUT_4[14933] = 32'b11111111111111110010010111100101;
assign LUT_4[14934] = 32'b11111111111111111000100110010001;
assign LUT_4[14935] = 32'b11111111111111110001110010001001;
assign LUT_4[14936] = 32'b11111111111111110101010111100110;
assign LUT_4[14937] = 32'b11111111111111101110100011011110;
assign LUT_4[14938] = 32'b11111111111111110100110010001010;
assign LUT_4[14939] = 32'b11111111111111101101111110000010;
assign LUT_4[14940] = 32'b11111111111111110010011000000010;
assign LUT_4[14941] = 32'b11111111111111101011100011111010;
assign LUT_4[14942] = 32'b11111111111111110001110010100110;
assign LUT_4[14943] = 32'b11111111111111101010111110011110;
assign LUT_4[14944] = 32'b11111111111111111100110100101010;
assign LUT_4[14945] = 32'b11111111111111110110000000100010;
assign LUT_4[14946] = 32'b11111111111111111100001111001110;
assign LUT_4[14947] = 32'b11111111111111110101011011000110;
assign LUT_4[14948] = 32'b11111111111111111001110101000110;
assign LUT_4[14949] = 32'b11111111111111110011000000111110;
assign LUT_4[14950] = 32'b11111111111111111001001111101010;
assign LUT_4[14951] = 32'b11111111111111110010011011100010;
assign LUT_4[14952] = 32'b11111111111111110110000000111111;
assign LUT_4[14953] = 32'b11111111111111101111001100110111;
assign LUT_4[14954] = 32'b11111111111111110101011011100011;
assign LUT_4[14955] = 32'b11111111111111101110100111011011;
assign LUT_4[14956] = 32'b11111111111111110011000001011011;
assign LUT_4[14957] = 32'b11111111111111101100001101010011;
assign LUT_4[14958] = 32'b11111111111111110010011011111111;
assign LUT_4[14959] = 32'b11111111111111101011100111110111;
assign LUT_4[14960] = 32'b11111111111111111010100110011000;
assign LUT_4[14961] = 32'b11111111111111110011110010010000;
assign LUT_4[14962] = 32'b11111111111111111010000000111100;
assign LUT_4[14963] = 32'b11111111111111110011001100110100;
assign LUT_4[14964] = 32'b11111111111111110111100110110100;
assign LUT_4[14965] = 32'b11111111111111110000110010101100;
assign LUT_4[14966] = 32'b11111111111111110111000001011000;
assign LUT_4[14967] = 32'b11111111111111110000001101010000;
assign LUT_4[14968] = 32'b11111111111111110011110010101101;
assign LUT_4[14969] = 32'b11111111111111101100111110100101;
assign LUT_4[14970] = 32'b11111111111111110011001101010001;
assign LUT_4[14971] = 32'b11111111111111101100011001001001;
assign LUT_4[14972] = 32'b11111111111111110000110011001001;
assign LUT_4[14973] = 32'b11111111111111101001111111000001;
assign LUT_4[14974] = 32'b11111111111111110000001101101101;
assign LUT_4[14975] = 32'b11111111111111101001011001100101;
assign LUT_4[14976] = 32'b11111111111111111111101000010111;
assign LUT_4[14977] = 32'b11111111111111111000110100001111;
assign LUT_4[14978] = 32'b11111111111111111111000010111011;
assign LUT_4[14979] = 32'b11111111111111111000001110110011;
assign LUT_4[14980] = 32'b11111111111111111100101000110011;
assign LUT_4[14981] = 32'b11111111111111110101110100101011;
assign LUT_4[14982] = 32'b11111111111111111100000011010111;
assign LUT_4[14983] = 32'b11111111111111110101001111001111;
assign LUT_4[14984] = 32'b11111111111111111000110100101100;
assign LUT_4[14985] = 32'b11111111111111110010000000100100;
assign LUT_4[14986] = 32'b11111111111111111000001111010000;
assign LUT_4[14987] = 32'b11111111111111110001011011001000;
assign LUT_4[14988] = 32'b11111111111111110101110101001000;
assign LUT_4[14989] = 32'b11111111111111101111000001000000;
assign LUT_4[14990] = 32'b11111111111111110101001111101100;
assign LUT_4[14991] = 32'b11111111111111101110011011100100;
assign LUT_4[14992] = 32'b11111111111111111101011010000101;
assign LUT_4[14993] = 32'b11111111111111110110100101111101;
assign LUT_4[14994] = 32'b11111111111111111100110100101001;
assign LUT_4[14995] = 32'b11111111111111110110000000100001;
assign LUT_4[14996] = 32'b11111111111111111010011010100001;
assign LUT_4[14997] = 32'b11111111111111110011100110011001;
assign LUT_4[14998] = 32'b11111111111111111001110101000101;
assign LUT_4[14999] = 32'b11111111111111110011000000111101;
assign LUT_4[15000] = 32'b11111111111111110110100110011010;
assign LUT_4[15001] = 32'b11111111111111101111110010010010;
assign LUT_4[15002] = 32'b11111111111111110110000000111110;
assign LUT_4[15003] = 32'b11111111111111101111001100110110;
assign LUT_4[15004] = 32'b11111111111111110011100110110110;
assign LUT_4[15005] = 32'b11111111111111101100110010101110;
assign LUT_4[15006] = 32'b11111111111111110011000001011010;
assign LUT_4[15007] = 32'b11111111111111101100001101010010;
assign LUT_4[15008] = 32'b11111111111111111110000011011110;
assign LUT_4[15009] = 32'b11111111111111110111001111010110;
assign LUT_4[15010] = 32'b11111111111111111101011110000010;
assign LUT_4[15011] = 32'b11111111111111110110101001111010;
assign LUT_4[15012] = 32'b11111111111111111011000011111010;
assign LUT_4[15013] = 32'b11111111111111110100001111110010;
assign LUT_4[15014] = 32'b11111111111111111010011110011110;
assign LUT_4[15015] = 32'b11111111111111110011101010010110;
assign LUT_4[15016] = 32'b11111111111111110111001111110011;
assign LUT_4[15017] = 32'b11111111111111110000011011101011;
assign LUT_4[15018] = 32'b11111111111111110110101010010111;
assign LUT_4[15019] = 32'b11111111111111101111110110001111;
assign LUT_4[15020] = 32'b11111111111111110100010000001111;
assign LUT_4[15021] = 32'b11111111111111101101011100000111;
assign LUT_4[15022] = 32'b11111111111111110011101010110011;
assign LUT_4[15023] = 32'b11111111111111101100110110101011;
assign LUT_4[15024] = 32'b11111111111111111011110101001100;
assign LUT_4[15025] = 32'b11111111111111110101000001000100;
assign LUT_4[15026] = 32'b11111111111111111011001111110000;
assign LUT_4[15027] = 32'b11111111111111110100011011101000;
assign LUT_4[15028] = 32'b11111111111111111000110101101000;
assign LUT_4[15029] = 32'b11111111111111110010000001100000;
assign LUT_4[15030] = 32'b11111111111111111000010000001100;
assign LUT_4[15031] = 32'b11111111111111110001011100000100;
assign LUT_4[15032] = 32'b11111111111111110101000001100001;
assign LUT_4[15033] = 32'b11111111111111101110001101011001;
assign LUT_4[15034] = 32'b11111111111111110100011100000101;
assign LUT_4[15035] = 32'b11111111111111101101100111111101;
assign LUT_4[15036] = 32'b11111111111111110010000001111101;
assign LUT_4[15037] = 32'b11111111111111101011001101110101;
assign LUT_4[15038] = 32'b11111111111111110001011100100001;
assign LUT_4[15039] = 32'b11111111111111101010101000011001;
assign LUT_4[15040] = 32'b00000000000000000000111111101011;
assign LUT_4[15041] = 32'b11111111111111111010001011100011;
assign LUT_4[15042] = 32'b00000000000000000000011010001111;
assign LUT_4[15043] = 32'b11111111111111111001100110000111;
assign LUT_4[15044] = 32'b11111111111111111110000000000111;
assign LUT_4[15045] = 32'b11111111111111110111001011111111;
assign LUT_4[15046] = 32'b11111111111111111101011010101011;
assign LUT_4[15047] = 32'b11111111111111110110100110100011;
assign LUT_4[15048] = 32'b11111111111111111010001100000000;
assign LUT_4[15049] = 32'b11111111111111110011010111111000;
assign LUT_4[15050] = 32'b11111111111111111001100110100100;
assign LUT_4[15051] = 32'b11111111111111110010110010011100;
assign LUT_4[15052] = 32'b11111111111111110111001100011100;
assign LUT_4[15053] = 32'b11111111111111110000011000010100;
assign LUT_4[15054] = 32'b11111111111111110110100111000000;
assign LUT_4[15055] = 32'b11111111111111101111110010111000;
assign LUT_4[15056] = 32'b11111111111111111110110001011001;
assign LUT_4[15057] = 32'b11111111111111110111111101010001;
assign LUT_4[15058] = 32'b11111111111111111110001011111101;
assign LUT_4[15059] = 32'b11111111111111110111010111110101;
assign LUT_4[15060] = 32'b11111111111111111011110001110101;
assign LUT_4[15061] = 32'b11111111111111110100111101101101;
assign LUT_4[15062] = 32'b11111111111111111011001100011001;
assign LUT_4[15063] = 32'b11111111111111110100011000010001;
assign LUT_4[15064] = 32'b11111111111111110111111101101110;
assign LUT_4[15065] = 32'b11111111111111110001001001100110;
assign LUT_4[15066] = 32'b11111111111111110111011000010010;
assign LUT_4[15067] = 32'b11111111111111110000100100001010;
assign LUT_4[15068] = 32'b11111111111111110100111110001010;
assign LUT_4[15069] = 32'b11111111111111101110001010000010;
assign LUT_4[15070] = 32'b11111111111111110100011000101110;
assign LUT_4[15071] = 32'b11111111111111101101100100100110;
assign LUT_4[15072] = 32'b11111111111111111111011010110010;
assign LUT_4[15073] = 32'b11111111111111111000100110101010;
assign LUT_4[15074] = 32'b11111111111111111110110101010110;
assign LUT_4[15075] = 32'b11111111111111111000000001001110;
assign LUT_4[15076] = 32'b11111111111111111100011011001110;
assign LUT_4[15077] = 32'b11111111111111110101100111000110;
assign LUT_4[15078] = 32'b11111111111111111011110101110010;
assign LUT_4[15079] = 32'b11111111111111110101000001101010;
assign LUT_4[15080] = 32'b11111111111111111000100111000111;
assign LUT_4[15081] = 32'b11111111111111110001110010111111;
assign LUT_4[15082] = 32'b11111111111111111000000001101011;
assign LUT_4[15083] = 32'b11111111111111110001001101100011;
assign LUT_4[15084] = 32'b11111111111111110101100111100011;
assign LUT_4[15085] = 32'b11111111111111101110110011011011;
assign LUT_4[15086] = 32'b11111111111111110101000010000111;
assign LUT_4[15087] = 32'b11111111111111101110001101111111;
assign LUT_4[15088] = 32'b11111111111111111101001100100000;
assign LUT_4[15089] = 32'b11111111111111110110011000011000;
assign LUT_4[15090] = 32'b11111111111111111100100111000100;
assign LUT_4[15091] = 32'b11111111111111110101110010111100;
assign LUT_4[15092] = 32'b11111111111111111010001100111100;
assign LUT_4[15093] = 32'b11111111111111110011011000110100;
assign LUT_4[15094] = 32'b11111111111111111001100111100000;
assign LUT_4[15095] = 32'b11111111111111110010110011011000;
assign LUT_4[15096] = 32'b11111111111111110110011000110101;
assign LUT_4[15097] = 32'b11111111111111101111100100101101;
assign LUT_4[15098] = 32'b11111111111111110101110011011001;
assign LUT_4[15099] = 32'b11111111111111101110111111010001;
assign LUT_4[15100] = 32'b11111111111111110011011001010001;
assign LUT_4[15101] = 32'b11111111111111101100100101001001;
assign LUT_4[15102] = 32'b11111111111111110010110011110101;
assign LUT_4[15103] = 32'b11111111111111101011111111101101;
assign LUT_4[15104] = 32'b00000000000000000001111101110010;
assign LUT_4[15105] = 32'b11111111111111111011001001101010;
assign LUT_4[15106] = 32'b00000000000000000001011000010110;
assign LUT_4[15107] = 32'b11111111111111111010100100001110;
assign LUT_4[15108] = 32'b11111111111111111110111110001110;
assign LUT_4[15109] = 32'b11111111111111111000001010000110;
assign LUT_4[15110] = 32'b11111111111111111110011000110010;
assign LUT_4[15111] = 32'b11111111111111110111100100101010;
assign LUT_4[15112] = 32'b11111111111111111011001010000111;
assign LUT_4[15113] = 32'b11111111111111110100010101111111;
assign LUT_4[15114] = 32'b11111111111111111010100100101011;
assign LUT_4[15115] = 32'b11111111111111110011110000100011;
assign LUT_4[15116] = 32'b11111111111111111000001010100011;
assign LUT_4[15117] = 32'b11111111111111110001010110011011;
assign LUT_4[15118] = 32'b11111111111111110111100101000111;
assign LUT_4[15119] = 32'b11111111111111110000110000111111;
assign LUT_4[15120] = 32'b11111111111111111111101111100000;
assign LUT_4[15121] = 32'b11111111111111111000111011011000;
assign LUT_4[15122] = 32'b11111111111111111111001010000100;
assign LUT_4[15123] = 32'b11111111111111111000010101111100;
assign LUT_4[15124] = 32'b11111111111111111100101111111100;
assign LUT_4[15125] = 32'b11111111111111110101111011110100;
assign LUT_4[15126] = 32'b11111111111111111100001010100000;
assign LUT_4[15127] = 32'b11111111111111110101010110011000;
assign LUT_4[15128] = 32'b11111111111111111000111011110101;
assign LUT_4[15129] = 32'b11111111111111110010000111101101;
assign LUT_4[15130] = 32'b11111111111111111000010110011001;
assign LUT_4[15131] = 32'b11111111111111110001100010010001;
assign LUT_4[15132] = 32'b11111111111111110101111100010001;
assign LUT_4[15133] = 32'b11111111111111101111001000001001;
assign LUT_4[15134] = 32'b11111111111111110101010110110101;
assign LUT_4[15135] = 32'b11111111111111101110100010101101;
assign LUT_4[15136] = 32'b00000000000000000000011000111001;
assign LUT_4[15137] = 32'b11111111111111111001100100110001;
assign LUT_4[15138] = 32'b11111111111111111111110011011101;
assign LUT_4[15139] = 32'b11111111111111111000111111010101;
assign LUT_4[15140] = 32'b11111111111111111101011001010101;
assign LUT_4[15141] = 32'b11111111111111110110100101001101;
assign LUT_4[15142] = 32'b11111111111111111100110011111001;
assign LUT_4[15143] = 32'b11111111111111110101111111110001;
assign LUT_4[15144] = 32'b11111111111111111001100101001110;
assign LUT_4[15145] = 32'b11111111111111110010110001000110;
assign LUT_4[15146] = 32'b11111111111111111000111111110010;
assign LUT_4[15147] = 32'b11111111111111110010001011101010;
assign LUT_4[15148] = 32'b11111111111111110110100101101010;
assign LUT_4[15149] = 32'b11111111111111101111110001100010;
assign LUT_4[15150] = 32'b11111111111111110110000000001110;
assign LUT_4[15151] = 32'b11111111111111101111001100000110;
assign LUT_4[15152] = 32'b11111111111111111110001010100111;
assign LUT_4[15153] = 32'b11111111111111110111010110011111;
assign LUT_4[15154] = 32'b11111111111111111101100101001011;
assign LUT_4[15155] = 32'b11111111111111110110110001000011;
assign LUT_4[15156] = 32'b11111111111111111011001011000011;
assign LUT_4[15157] = 32'b11111111111111110100010110111011;
assign LUT_4[15158] = 32'b11111111111111111010100101100111;
assign LUT_4[15159] = 32'b11111111111111110011110001011111;
assign LUT_4[15160] = 32'b11111111111111110111010110111100;
assign LUT_4[15161] = 32'b11111111111111110000100010110100;
assign LUT_4[15162] = 32'b11111111111111110110110001100000;
assign LUT_4[15163] = 32'b11111111111111101111111101011000;
assign LUT_4[15164] = 32'b11111111111111110100010111011000;
assign LUT_4[15165] = 32'b11111111111111101101100011010000;
assign LUT_4[15166] = 32'b11111111111111110011110001111100;
assign LUT_4[15167] = 32'b11111111111111101100111101110100;
assign LUT_4[15168] = 32'b00000000000000000011010101000110;
assign LUT_4[15169] = 32'b11111111111111111100100000111110;
assign LUT_4[15170] = 32'b00000000000000000010101111101010;
assign LUT_4[15171] = 32'b11111111111111111011111011100010;
assign LUT_4[15172] = 32'b00000000000000000000010101100010;
assign LUT_4[15173] = 32'b11111111111111111001100001011010;
assign LUT_4[15174] = 32'b11111111111111111111110000000110;
assign LUT_4[15175] = 32'b11111111111111111000111011111110;
assign LUT_4[15176] = 32'b11111111111111111100100001011011;
assign LUT_4[15177] = 32'b11111111111111110101101101010011;
assign LUT_4[15178] = 32'b11111111111111111011111011111111;
assign LUT_4[15179] = 32'b11111111111111110101000111110111;
assign LUT_4[15180] = 32'b11111111111111111001100001110111;
assign LUT_4[15181] = 32'b11111111111111110010101101101111;
assign LUT_4[15182] = 32'b11111111111111111000111100011011;
assign LUT_4[15183] = 32'b11111111111111110010001000010011;
assign LUT_4[15184] = 32'b00000000000000000001000110110100;
assign LUT_4[15185] = 32'b11111111111111111010010010101100;
assign LUT_4[15186] = 32'b00000000000000000000100001011000;
assign LUT_4[15187] = 32'b11111111111111111001101101010000;
assign LUT_4[15188] = 32'b11111111111111111110000111010000;
assign LUT_4[15189] = 32'b11111111111111110111010011001000;
assign LUT_4[15190] = 32'b11111111111111111101100001110100;
assign LUT_4[15191] = 32'b11111111111111110110101101101100;
assign LUT_4[15192] = 32'b11111111111111111010010011001001;
assign LUT_4[15193] = 32'b11111111111111110011011111000001;
assign LUT_4[15194] = 32'b11111111111111111001101101101101;
assign LUT_4[15195] = 32'b11111111111111110010111001100101;
assign LUT_4[15196] = 32'b11111111111111110111010011100101;
assign LUT_4[15197] = 32'b11111111111111110000011111011101;
assign LUT_4[15198] = 32'b11111111111111110110101110001001;
assign LUT_4[15199] = 32'b11111111111111101111111010000001;
assign LUT_4[15200] = 32'b00000000000000000001110000001101;
assign LUT_4[15201] = 32'b11111111111111111010111100000101;
assign LUT_4[15202] = 32'b00000000000000000001001010110001;
assign LUT_4[15203] = 32'b11111111111111111010010110101001;
assign LUT_4[15204] = 32'b11111111111111111110110000101001;
assign LUT_4[15205] = 32'b11111111111111110111111100100001;
assign LUT_4[15206] = 32'b11111111111111111110001011001101;
assign LUT_4[15207] = 32'b11111111111111110111010111000101;
assign LUT_4[15208] = 32'b11111111111111111010111100100010;
assign LUT_4[15209] = 32'b11111111111111110100001000011010;
assign LUT_4[15210] = 32'b11111111111111111010010111000110;
assign LUT_4[15211] = 32'b11111111111111110011100010111110;
assign LUT_4[15212] = 32'b11111111111111110111111100111110;
assign LUT_4[15213] = 32'b11111111111111110001001000110110;
assign LUT_4[15214] = 32'b11111111111111110111010111100010;
assign LUT_4[15215] = 32'b11111111111111110000100011011010;
assign LUT_4[15216] = 32'b11111111111111111111100001111011;
assign LUT_4[15217] = 32'b11111111111111111000101101110011;
assign LUT_4[15218] = 32'b11111111111111111110111100011111;
assign LUT_4[15219] = 32'b11111111111111111000001000010111;
assign LUT_4[15220] = 32'b11111111111111111100100010010111;
assign LUT_4[15221] = 32'b11111111111111110101101110001111;
assign LUT_4[15222] = 32'b11111111111111111011111100111011;
assign LUT_4[15223] = 32'b11111111111111110101001000110011;
assign LUT_4[15224] = 32'b11111111111111111000101110010000;
assign LUT_4[15225] = 32'b11111111111111110001111010001000;
assign LUT_4[15226] = 32'b11111111111111111000001000110100;
assign LUT_4[15227] = 32'b11111111111111110001010100101100;
assign LUT_4[15228] = 32'b11111111111111110101101110101100;
assign LUT_4[15229] = 32'b11111111111111101110111010100100;
assign LUT_4[15230] = 32'b11111111111111110101001001010000;
assign LUT_4[15231] = 32'b11111111111111101110010101001000;
assign LUT_4[15232] = 32'b00000000000000000100100011111010;
assign LUT_4[15233] = 32'b11111111111111111101101111110010;
assign LUT_4[15234] = 32'b00000000000000000011111110011110;
assign LUT_4[15235] = 32'b11111111111111111101001010010110;
assign LUT_4[15236] = 32'b00000000000000000001100100010110;
assign LUT_4[15237] = 32'b11111111111111111010110000001110;
assign LUT_4[15238] = 32'b00000000000000000000111110111010;
assign LUT_4[15239] = 32'b11111111111111111010001010110010;
assign LUT_4[15240] = 32'b11111111111111111101110000001111;
assign LUT_4[15241] = 32'b11111111111111110110111100000111;
assign LUT_4[15242] = 32'b11111111111111111101001010110011;
assign LUT_4[15243] = 32'b11111111111111110110010110101011;
assign LUT_4[15244] = 32'b11111111111111111010110000101011;
assign LUT_4[15245] = 32'b11111111111111110011111100100011;
assign LUT_4[15246] = 32'b11111111111111111010001011001111;
assign LUT_4[15247] = 32'b11111111111111110011010111000111;
assign LUT_4[15248] = 32'b00000000000000000010010101101000;
assign LUT_4[15249] = 32'b11111111111111111011100001100000;
assign LUT_4[15250] = 32'b00000000000000000001110000001100;
assign LUT_4[15251] = 32'b11111111111111111010111100000100;
assign LUT_4[15252] = 32'b11111111111111111111010110000100;
assign LUT_4[15253] = 32'b11111111111111111000100001111100;
assign LUT_4[15254] = 32'b11111111111111111110110000101000;
assign LUT_4[15255] = 32'b11111111111111110111111100100000;
assign LUT_4[15256] = 32'b11111111111111111011100001111101;
assign LUT_4[15257] = 32'b11111111111111110100101101110101;
assign LUT_4[15258] = 32'b11111111111111111010111100100001;
assign LUT_4[15259] = 32'b11111111111111110100001000011001;
assign LUT_4[15260] = 32'b11111111111111111000100010011001;
assign LUT_4[15261] = 32'b11111111111111110001101110010001;
assign LUT_4[15262] = 32'b11111111111111110111111100111101;
assign LUT_4[15263] = 32'b11111111111111110001001000110101;
assign LUT_4[15264] = 32'b00000000000000000010111111000001;
assign LUT_4[15265] = 32'b11111111111111111100001010111001;
assign LUT_4[15266] = 32'b00000000000000000010011001100101;
assign LUT_4[15267] = 32'b11111111111111111011100101011101;
assign LUT_4[15268] = 32'b11111111111111111111111111011101;
assign LUT_4[15269] = 32'b11111111111111111001001011010101;
assign LUT_4[15270] = 32'b11111111111111111111011010000001;
assign LUT_4[15271] = 32'b11111111111111111000100101111001;
assign LUT_4[15272] = 32'b11111111111111111100001011010110;
assign LUT_4[15273] = 32'b11111111111111110101010111001110;
assign LUT_4[15274] = 32'b11111111111111111011100101111010;
assign LUT_4[15275] = 32'b11111111111111110100110001110010;
assign LUT_4[15276] = 32'b11111111111111111001001011110010;
assign LUT_4[15277] = 32'b11111111111111110010010111101010;
assign LUT_4[15278] = 32'b11111111111111111000100110010110;
assign LUT_4[15279] = 32'b11111111111111110001110010001110;
assign LUT_4[15280] = 32'b00000000000000000000110000101111;
assign LUT_4[15281] = 32'b11111111111111111001111100100111;
assign LUT_4[15282] = 32'b00000000000000000000001011010011;
assign LUT_4[15283] = 32'b11111111111111111001010111001011;
assign LUT_4[15284] = 32'b11111111111111111101110001001011;
assign LUT_4[15285] = 32'b11111111111111110110111101000011;
assign LUT_4[15286] = 32'b11111111111111111101001011101111;
assign LUT_4[15287] = 32'b11111111111111110110010111100111;
assign LUT_4[15288] = 32'b11111111111111111001111101000100;
assign LUT_4[15289] = 32'b11111111111111110011001000111100;
assign LUT_4[15290] = 32'b11111111111111111001010111101000;
assign LUT_4[15291] = 32'b11111111111111110010100011100000;
assign LUT_4[15292] = 32'b11111111111111110110111101100000;
assign LUT_4[15293] = 32'b11111111111111110000001001011000;
assign LUT_4[15294] = 32'b11111111111111110110011000000100;
assign LUT_4[15295] = 32'b11111111111111101111100011111100;
assign LUT_4[15296] = 32'b00000000000000000101111011001110;
assign LUT_4[15297] = 32'b11111111111111111111000111000110;
assign LUT_4[15298] = 32'b00000000000000000101010101110010;
assign LUT_4[15299] = 32'b11111111111111111110100001101010;
assign LUT_4[15300] = 32'b00000000000000000010111011101010;
assign LUT_4[15301] = 32'b11111111111111111100000111100010;
assign LUT_4[15302] = 32'b00000000000000000010010110001110;
assign LUT_4[15303] = 32'b11111111111111111011100010000110;
assign LUT_4[15304] = 32'b11111111111111111111000111100011;
assign LUT_4[15305] = 32'b11111111111111111000010011011011;
assign LUT_4[15306] = 32'b11111111111111111110100010000111;
assign LUT_4[15307] = 32'b11111111111111110111101101111111;
assign LUT_4[15308] = 32'b11111111111111111100000111111111;
assign LUT_4[15309] = 32'b11111111111111110101010011110111;
assign LUT_4[15310] = 32'b11111111111111111011100010100011;
assign LUT_4[15311] = 32'b11111111111111110100101110011011;
assign LUT_4[15312] = 32'b00000000000000000011101100111100;
assign LUT_4[15313] = 32'b11111111111111111100111000110100;
assign LUT_4[15314] = 32'b00000000000000000011000111100000;
assign LUT_4[15315] = 32'b11111111111111111100010011011000;
assign LUT_4[15316] = 32'b00000000000000000000101101011000;
assign LUT_4[15317] = 32'b11111111111111111001111001010000;
assign LUT_4[15318] = 32'b00000000000000000000000111111100;
assign LUT_4[15319] = 32'b11111111111111111001010011110100;
assign LUT_4[15320] = 32'b11111111111111111100111001010001;
assign LUT_4[15321] = 32'b11111111111111110110000101001001;
assign LUT_4[15322] = 32'b11111111111111111100010011110101;
assign LUT_4[15323] = 32'b11111111111111110101011111101101;
assign LUT_4[15324] = 32'b11111111111111111001111001101101;
assign LUT_4[15325] = 32'b11111111111111110011000101100101;
assign LUT_4[15326] = 32'b11111111111111111001010100010001;
assign LUT_4[15327] = 32'b11111111111111110010100000001001;
assign LUT_4[15328] = 32'b00000000000000000100010110010101;
assign LUT_4[15329] = 32'b11111111111111111101100010001101;
assign LUT_4[15330] = 32'b00000000000000000011110000111001;
assign LUT_4[15331] = 32'b11111111111111111100111100110001;
assign LUT_4[15332] = 32'b00000000000000000001010110110001;
assign LUT_4[15333] = 32'b11111111111111111010100010101001;
assign LUT_4[15334] = 32'b00000000000000000000110001010101;
assign LUT_4[15335] = 32'b11111111111111111001111101001101;
assign LUT_4[15336] = 32'b11111111111111111101100010101010;
assign LUT_4[15337] = 32'b11111111111111110110101110100010;
assign LUT_4[15338] = 32'b11111111111111111100111101001110;
assign LUT_4[15339] = 32'b11111111111111110110001001000110;
assign LUT_4[15340] = 32'b11111111111111111010100011000110;
assign LUT_4[15341] = 32'b11111111111111110011101110111110;
assign LUT_4[15342] = 32'b11111111111111111001111101101010;
assign LUT_4[15343] = 32'b11111111111111110011001001100010;
assign LUT_4[15344] = 32'b00000000000000000010001000000011;
assign LUT_4[15345] = 32'b11111111111111111011010011111011;
assign LUT_4[15346] = 32'b00000000000000000001100010100111;
assign LUT_4[15347] = 32'b11111111111111111010101110011111;
assign LUT_4[15348] = 32'b11111111111111111111001000011111;
assign LUT_4[15349] = 32'b11111111111111111000010100010111;
assign LUT_4[15350] = 32'b11111111111111111110100011000011;
assign LUT_4[15351] = 32'b11111111111111110111101110111011;
assign LUT_4[15352] = 32'b11111111111111111011010100011000;
assign LUT_4[15353] = 32'b11111111111111110100100000010000;
assign LUT_4[15354] = 32'b11111111111111111010101110111100;
assign LUT_4[15355] = 32'b11111111111111110011111010110100;
assign LUT_4[15356] = 32'b11111111111111111000010100110100;
assign LUT_4[15357] = 32'b11111111111111110001100000101100;
assign LUT_4[15358] = 32'b11111111111111110111101111011000;
assign LUT_4[15359] = 32'b11111111111111110000111011010000;
assign LUT_4[15360] = 32'b11111111111111111111101000100110;
assign LUT_4[15361] = 32'b11111111111111111000110100011110;
assign LUT_4[15362] = 32'b11111111111111111111000011001010;
assign LUT_4[15363] = 32'b11111111111111111000001111000010;
assign LUT_4[15364] = 32'b11111111111111111100101001000010;
assign LUT_4[15365] = 32'b11111111111111110101110100111010;
assign LUT_4[15366] = 32'b11111111111111111100000011100110;
assign LUT_4[15367] = 32'b11111111111111110101001111011110;
assign LUT_4[15368] = 32'b11111111111111111000110100111011;
assign LUT_4[15369] = 32'b11111111111111110010000000110011;
assign LUT_4[15370] = 32'b11111111111111111000001111011111;
assign LUT_4[15371] = 32'b11111111111111110001011011010111;
assign LUT_4[15372] = 32'b11111111111111110101110101010111;
assign LUT_4[15373] = 32'b11111111111111101111000001001111;
assign LUT_4[15374] = 32'b11111111111111110101001111111011;
assign LUT_4[15375] = 32'b11111111111111101110011011110011;
assign LUT_4[15376] = 32'b11111111111111111101011010010100;
assign LUT_4[15377] = 32'b11111111111111110110100110001100;
assign LUT_4[15378] = 32'b11111111111111111100110100111000;
assign LUT_4[15379] = 32'b11111111111111110110000000110000;
assign LUT_4[15380] = 32'b11111111111111111010011010110000;
assign LUT_4[15381] = 32'b11111111111111110011100110101000;
assign LUT_4[15382] = 32'b11111111111111111001110101010100;
assign LUT_4[15383] = 32'b11111111111111110011000001001100;
assign LUT_4[15384] = 32'b11111111111111110110100110101001;
assign LUT_4[15385] = 32'b11111111111111101111110010100001;
assign LUT_4[15386] = 32'b11111111111111110110000001001101;
assign LUT_4[15387] = 32'b11111111111111101111001101000101;
assign LUT_4[15388] = 32'b11111111111111110011100111000101;
assign LUT_4[15389] = 32'b11111111111111101100110010111101;
assign LUT_4[15390] = 32'b11111111111111110011000001101001;
assign LUT_4[15391] = 32'b11111111111111101100001101100001;
assign LUT_4[15392] = 32'b11111111111111111110000011101101;
assign LUT_4[15393] = 32'b11111111111111110111001111100101;
assign LUT_4[15394] = 32'b11111111111111111101011110010001;
assign LUT_4[15395] = 32'b11111111111111110110101010001001;
assign LUT_4[15396] = 32'b11111111111111111011000100001001;
assign LUT_4[15397] = 32'b11111111111111110100010000000001;
assign LUT_4[15398] = 32'b11111111111111111010011110101101;
assign LUT_4[15399] = 32'b11111111111111110011101010100101;
assign LUT_4[15400] = 32'b11111111111111110111010000000010;
assign LUT_4[15401] = 32'b11111111111111110000011011111010;
assign LUT_4[15402] = 32'b11111111111111110110101010100110;
assign LUT_4[15403] = 32'b11111111111111101111110110011110;
assign LUT_4[15404] = 32'b11111111111111110100010000011110;
assign LUT_4[15405] = 32'b11111111111111101101011100010110;
assign LUT_4[15406] = 32'b11111111111111110011101011000010;
assign LUT_4[15407] = 32'b11111111111111101100110110111010;
assign LUT_4[15408] = 32'b11111111111111111011110101011011;
assign LUT_4[15409] = 32'b11111111111111110101000001010011;
assign LUT_4[15410] = 32'b11111111111111111011001111111111;
assign LUT_4[15411] = 32'b11111111111111110100011011110111;
assign LUT_4[15412] = 32'b11111111111111111000110101110111;
assign LUT_4[15413] = 32'b11111111111111110010000001101111;
assign LUT_4[15414] = 32'b11111111111111111000010000011011;
assign LUT_4[15415] = 32'b11111111111111110001011100010011;
assign LUT_4[15416] = 32'b11111111111111110101000001110000;
assign LUT_4[15417] = 32'b11111111111111101110001101101000;
assign LUT_4[15418] = 32'b11111111111111110100011100010100;
assign LUT_4[15419] = 32'b11111111111111101101101000001100;
assign LUT_4[15420] = 32'b11111111111111110010000010001100;
assign LUT_4[15421] = 32'b11111111111111101011001110000100;
assign LUT_4[15422] = 32'b11111111111111110001011100110000;
assign LUT_4[15423] = 32'b11111111111111101010101000101000;
assign LUT_4[15424] = 32'b00000000000000000000111111111010;
assign LUT_4[15425] = 32'b11111111111111111010001011110010;
assign LUT_4[15426] = 32'b00000000000000000000011010011110;
assign LUT_4[15427] = 32'b11111111111111111001100110010110;
assign LUT_4[15428] = 32'b11111111111111111110000000010110;
assign LUT_4[15429] = 32'b11111111111111110111001100001110;
assign LUT_4[15430] = 32'b11111111111111111101011010111010;
assign LUT_4[15431] = 32'b11111111111111110110100110110010;
assign LUT_4[15432] = 32'b11111111111111111010001100001111;
assign LUT_4[15433] = 32'b11111111111111110011011000000111;
assign LUT_4[15434] = 32'b11111111111111111001100110110011;
assign LUT_4[15435] = 32'b11111111111111110010110010101011;
assign LUT_4[15436] = 32'b11111111111111110111001100101011;
assign LUT_4[15437] = 32'b11111111111111110000011000100011;
assign LUT_4[15438] = 32'b11111111111111110110100111001111;
assign LUT_4[15439] = 32'b11111111111111101111110011000111;
assign LUT_4[15440] = 32'b11111111111111111110110001101000;
assign LUT_4[15441] = 32'b11111111111111110111111101100000;
assign LUT_4[15442] = 32'b11111111111111111110001100001100;
assign LUT_4[15443] = 32'b11111111111111110111011000000100;
assign LUT_4[15444] = 32'b11111111111111111011110010000100;
assign LUT_4[15445] = 32'b11111111111111110100111101111100;
assign LUT_4[15446] = 32'b11111111111111111011001100101000;
assign LUT_4[15447] = 32'b11111111111111110100011000100000;
assign LUT_4[15448] = 32'b11111111111111110111111101111101;
assign LUT_4[15449] = 32'b11111111111111110001001001110101;
assign LUT_4[15450] = 32'b11111111111111110111011000100001;
assign LUT_4[15451] = 32'b11111111111111110000100100011001;
assign LUT_4[15452] = 32'b11111111111111110100111110011001;
assign LUT_4[15453] = 32'b11111111111111101110001010010001;
assign LUT_4[15454] = 32'b11111111111111110100011000111101;
assign LUT_4[15455] = 32'b11111111111111101101100100110101;
assign LUT_4[15456] = 32'b11111111111111111111011011000001;
assign LUT_4[15457] = 32'b11111111111111111000100110111001;
assign LUT_4[15458] = 32'b11111111111111111110110101100101;
assign LUT_4[15459] = 32'b11111111111111111000000001011101;
assign LUT_4[15460] = 32'b11111111111111111100011011011101;
assign LUT_4[15461] = 32'b11111111111111110101100111010101;
assign LUT_4[15462] = 32'b11111111111111111011110110000001;
assign LUT_4[15463] = 32'b11111111111111110101000001111001;
assign LUT_4[15464] = 32'b11111111111111111000100111010110;
assign LUT_4[15465] = 32'b11111111111111110001110011001110;
assign LUT_4[15466] = 32'b11111111111111111000000001111010;
assign LUT_4[15467] = 32'b11111111111111110001001101110010;
assign LUT_4[15468] = 32'b11111111111111110101100111110010;
assign LUT_4[15469] = 32'b11111111111111101110110011101010;
assign LUT_4[15470] = 32'b11111111111111110101000010010110;
assign LUT_4[15471] = 32'b11111111111111101110001110001110;
assign LUT_4[15472] = 32'b11111111111111111101001100101111;
assign LUT_4[15473] = 32'b11111111111111110110011000100111;
assign LUT_4[15474] = 32'b11111111111111111100100111010011;
assign LUT_4[15475] = 32'b11111111111111110101110011001011;
assign LUT_4[15476] = 32'b11111111111111111010001101001011;
assign LUT_4[15477] = 32'b11111111111111110011011001000011;
assign LUT_4[15478] = 32'b11111111111111111001100111101111;
assign LUT_4[15479] = 32'b11111111111111110010110011100111;
assign LUT_4[15480] = 32'b11111111111111110110011001000100;
assign LUT_4[15481] = 32'b11111111111111101111100100111100;
assign LUT_4[15482] = 32'b11111111111111110101110011101000;
assign LUT_4[15483] = 32'b11111111111111101110111111100000;
assign LUT_4[15484] = 32'b11111111111111110011011001100000;
assign LUT_4[15485] = 32'b11111111111111101100100101011000;
assign LUT_4[15486] = 32'b11111111111111110010110100000100;
assign LUT_4[15487] = 32'b11111111111111101011111111111100;
assign LUT_4[15488] = 32'b00000000000000000010001110101110;
assign LUT_4[15489] = 32'b11111111111111111011011010100110;
assign LUT_4[15490] = 32'b00000000000000000001101001010010;
assign LUT_4[15491] = 32'b11111111111111111010110101001010;
assign LUT_4[15492] = 32'b11111111111111111111001111001010;
assign LUT_4[15493] = 32'b11111111111111111000011011000010;
assign LUT_4[15494] = 32'b11111111111111111110101001101110;
assign LUT_4[15495] = 32'b11111111111111110111110101100110;
assign LUT_4[15496] = 32'b11111111111111111011011011000011;
assign LUT_4[15497] = 32'b11111111111111110100100110111011;
assign LUT_4[15498] = 32'b11111111111111111010110101100111;
assign LUT_4[15499] = 32'b11111111111111110100000001011111;
assign LUT_4[15500] = 32'b11111111111111111000011011011111;
assign LUT_4[15501] = 32'b11111111111111110001100111010111;
assign LUT_4[15502] = 32'b11111111111111110111110110000011;
assign LUT_4[15503] = 32'b11111111111111110001000001111011;
assign LUT_4[15504] = 32'b00000000000000000000000000011100;
assign LUT_4[15505] = 32'b11111111111111111001001100010100;
assign LUT_4[15506] = 32'b11111111111111111111011011000000;
assign LUT_4[15507] = 32'b11111111111111111000100110111000;
assign LUT_4[15508] = 32'b11111111111111111101000000111000;
assign LUT_4[15509] = 32'b11111111111111110110001100110000;
assign LUT_4[15510] = 32'b11111111111111111100011011011100;
assign LUT_4[15511] = 32'b11111111111111110101100111010100;
assign LUT_4[15512] = 32'b11111111111111111001001100110001;
assign LUT_4[15513] = 32'b11111111111111110010011000101001;
assign LUT_4[15514] = 32'b11111111111111111000100111010101;
assign LUT_4[15515] = 32'b11111111111111110001110011001101;
assign LUT_4[15516] = 32'b11111111111111110110001101001101;
assign LUT_4[15517] = 32'b11111111111111101111011001000101;
assign LUT_4[15518] = 32'b11111111111111110101100111110001;
assign LUT_4[15519] = 32'b11111111111111101110110011101001;
assign LUT_4[15520] = 32'b00000000000000000000101001110101;
assign LUT_4[15521] = 32'b11111111111111111001110101101101;
assign LUT_4[15522] = 32'b00000000000000000000000100011001;
assign LUT_4[15523] = 32'b11111111111111111001010000010001;
assign LUT_4[15524] = 32'b11111111111111111101101010010001;
assign LUT_4[15525] = 32'b11111111111111110110110110001001;
assign LUT_4[15526] = 32'b11111111111111111101000100110101;
assign LUT_4[15527] = 32'b11111111111111110110010000101101;
assign LUT_4[15528] = 32'b11111111111111111001110110001010;
assign LUT_4[15529] = 32'b11111111111111110011000010000010;
assign LUT_4[15530] = 32'b11111111111111111001010000101110;
assign LUT_4[15531] = 32'b11111111111111110010011100100110;
assign LUT_4[15532] = 32'b11111111111111110110110110100110;
assign LUT_4[15533] = 32'b11111111111111110000000010011110;
assign LUT_4[15534] = 32'b11111111111111110110010001001010;
assign LUT_4[15535] = 32'b11111111111111101111011101000010;
assign LUT_4[15536] = 32'b11111111111111111110011011100011;
assign LUT_4[15537] = 32'b11111111111111110111100111011011;
assign LUT_4[15538] = 32'b11111111111111111101110110000111;
assign LUT_4[15539] = 32'b11111111111111110111000001111111;
assign LUT_4[15540] = 32'b11111111111111111011011011111111;
assign LUT_4[15541] = 32'b11111111111111110100100111110111;
assign LUT_4[15542] = 32'b11111111111111111010110110100011;
assign LUT_4[15543] = 32'b11111111111111110100000010011011;
assign LUT_4[15544] = 32'b11111111111111110111100111111000;
assign LUT_4[15545] = 32'b11111111111111110000110011110000;
assign LUT_4[15546] = 32'b11111111111111110111000010011100;
assign LUT_4[15547] = 32'b11111111111111110000001110010100;
assign LUT_4[15548] = 32'b11111111111111110100101000010100;
assign LUT_4[15549] = 32'b11111111111111101101110100001100;
assign LUT_4[15550] = 32'b11111111111111110100000010111000;
assign LUT_4[15551] = 32'b11111111111111101101001110110000;
assign LUT_4[15552] = 32'b00000000000000000011100110000010;
assign LUT_4[15553] = 32'b11111111111111111100110001111010;
assign LUT_4[15554] = 32'b00000000000000000011000000100110;
assign LUT_4[15555] = 32'b11111111111111111100001100011110;
assign LUT_4[15556] = 32'b00000000000000000000100110011110;
assign LUT_4[15557] = 32'b11111111111111111001110010010110;
assign LUT_4[15558] = 32'b00000000000000000000000001000010;
assign LUT_4[15559] = 32'b11111111111111111001001100111010;
assign LUT_4[15560] = 32'b11111111111111111100110010010111;
assign LUT_4[15561] = 32'b11111111111111110101111110001111;
assign LUT_4[15562] = 32'b11111111111111111100001100111011;
assign LUT_4[15563] = 32'b11111111111111110101011000110011;
assign LUT_4[15564] = 32'b11111111111111111001110010110011;
assign LUT_4[15565] = 32'b11111111111111110010111110101011;
assign LUT_4[15566] = 32'b11111111111111111001001101010111;
assign LUT_4[15567] = 32'b11111111111111110010011001001111;
assign LUT_4[15568] = 32'b00000000000000000001010111110000;
assign LUT_4[15569] = 32'b11111111111111111010100011101000;
assign LUT_4[15570] = 32'b00000000000000000000110010010100;
assign LUT_4[15571] = 32'b11111111111111111001111110001100;
assign LUT_4[15572] = 32'b11111111111111111110011000001100;
assign LUT_4[15573] = 32'b11111111111111110111100100000100;
assign LUT_4[15574] = 32'b11111111111111111101110010110000;
assign LUT_4[15575] = 32'b11111111111111110110111110101000;
assign LUT_4[15576] = 32'b11111111111111111010100100000101;
assign LUT_4[15577] = 32'b11111111111111110011101111111101;
assign LUT_4[15578] = 32'b11111111111111111001111110101001;
assign LUT_4[15579] = 32'b11111111111111110011001010100001;
assign LUT_4[15580] = 32'b11111111111111110111100100100001;
assign LUT_4[15581] = 32'b11111111111111110000110000011001;
assign LUT_4[15582] = 32'b11111111111111110110111111000101;
assign LUT_4[15583] = 32'b11111111111111110000001010111101;
assign LUT_4[15584] = 32'b00000000000000000010000001001001;
assign LUT_4[15585] = 32'b11111111111111111011001101000001;
assign LUT_4[15586] = 32'b00000000000000000001011011101101;
assign LUT_4[15587] = 32'b11111111111111111010100111100101;
assign LUT_4[15588] = 32'b11111111111111111111000001100101;
assign LUT_4[15589] = 32'b11111111111111111000001101011101;
assign LUT_4[15590] = 32'b11111111111111111110011100001001;
assign LUT_4[15591] = 32'b11111111111111110111101000000001;
assign LUT_4[15592] = 32'b11111111111111111011001101011110;
assign LUT_4[15593] = 32'b11111111111111110100011001010110;
assign LUT_4[15594] = 32'b11111111111111111010101000000010;
assign LUT_4[15595] = 32'b11111111111111110011110011111010;
assign LUT_4[15596] = 32'b11111111111111111000001101111010;
assign LUT_4[15597] = 32'b11111111111111110001011001110010;
assign LUT_4[15598] = 32'b11111111111111110111101000011110;
assign LUT_4[15599] = 32'b11111111111111110000110100010110;
assign LUT_4[15600] = 32'b11111111111111111111110010110111;
assign LUT_4[15601] = 32'b11111111111111111000111110101111;
assign LUT_4[15602] = 32'b11111111111111111111001101011011;
assign LUT_4[15603] = 32'b11111111111111111000011001010011;
assign LUT_4[15604] = 32'b11111111111111111100110011010011;
assign LUT_4[15605] = 32'b11111111111111110101111111001011;
assign LUT_4[15606] = 32'b11111111111111111100001101110111;
assign LUT_4[15607] = 32'b11111111111111110101011001101111;
assign LUT_4[15608] = 32'b11111111111111111000111111001100;
assign LUT_4[15609] = 32'b11111111111111110010001011000100;
assign LUT_4[15610] = 32'b11111111111111111000011001110000;
assign LUT_4[15611] = 32'b11111111111111110001100101101000;
assign LUT_4[15612] = 32'b11111111111111110101111111101000;
assign LUT_4[15613] = 32'b11111111111111101111001011100000;
assign LUT_4[15614] = 32'b11111111111111110101011010001100;
assign LUT_4[15615] = 32'b11111111111111101110100110000100;
assign LUT_4[15616] = 32'b00000000000000000100100100001001;
assign LUT_4[15617] = 32'b11111111111111111101110000000001;
assign LUT_4[15618] = 32'b00000000000000000011111110101101;
assign LUT_4[15619] = 32'b11111111111111111101001010100101;
assign LUT_4[15620] = 32'b00000000000000000001100100100101;
assign LUT_4[15621] = 32'b11111111111111111010110000011101;
assign LUT_4[15622] = 32'b00000000000000000000111111001001;
assign LUT_4[15623] = 32'b11111111111111111010001011000001;
assign LUT_4[15624] = 32'b11111111111111111101110000011110;
assign LUT_4[15625] = 32'b11111111111111110110111100010110;
assign LUT_4[15626] = 32'b11111111111111111101001011000010;
assign LUT_4[15627] = 32'b11111111111111110110010110111010;
assign LUT_4[15628] = 32'b11111111111111111010110000111010;
assign LUT_4[15629] = 32'b11111111111111110011111100110010;
assign LUT_4[15630] = 32'b11111111111111111010001011011110;
assign LUT_4[15631] = 32'b11111111111111110011010111010110;
assign LUT_4[15632] = 32'b00000000000000000010010101110111;
assign LUT_4[15633] = 32'b11111111111111111011100001101111;
assign LUT_4[15634] = 32'b00000000000000000001110000011011;
assign LUT_4[15635] = 32'b11111111111111111010111100010011;
assign LUT_4[15636] = 32'b11111111111111111111010110010011;
assign LUT_4[15637] = 32'b11111111111111111000100010001011;
assign LUT_4[15638] = 32'b11111111111111111110110000110111;
assign LUT_4[15639] = 32'b11111111111111110111111100101111;
assign LUT_4[15640] = 32'b11111111111111111011100010001100;
assign LUT_4[15641] = 32'b11111111111111110100101110000100;
assign LUT_4[15642] = 32'b11111111111111111010111100110000;
assign LUT_4[15643] = 32'b11111111111111110100001000101000;
assign LUT_4[15644] = 32'b11111111111111111000100010101000;
assign LUT_4[15645] = 32'b11111111111111110001101110100000;
assign LUT_4[15646] = 32'b11111111111111110111111101001100;
assign LUT_4[15647] = 32'b11111111111111110001001001000100;
assign LUT_4[15648] = 32'b00000000000000000010111111010000;
assign LUT_4[15649] = 32'b11111111111111111100001011001000;
assign LUT_4[15650] = 32'b00000000000000000010011001110100;
assign LUT_4[15651] = 32'b11111111111111111011100101101100;
assign LUT_4[15652] = 32'b11111111111111111111111111101100;
assign LUT_4[15653] = 32'b11111111111111111001001011100100;
assign LUT_4[15654] = 32'b11111111111111111111011010010000;
assign LUT_4[15655] = 32'b11111111111111111000100110001000;
assign LUT_4[15656] = 32'b11111111111111111100001011100101;
assign LUT_4[15657] = 32'b11111111111111110101010111011101;
assign LUT_4[15658] = 32'b11111111111111111011100110001001;
assign LUT_4[15659] = 32'b11111111111111110100110010000001;
assign LUT_4[15660] = 32'b11111111111111111001001100000001;
assign LUT_4[15661] = 32'b11111111111111110010010111111001;
assign LUT_4[15662] = 32'b11111111111111111000100110100101;
assign LUT_4[15663] = 32'b11111111111111110001110010011101;
assign LUT_4[15664] = 32'b00000000000000000000110000111110;
assign LUT_4[15665] = 32'b11111111111111111001111100110110;
assign LUT_4[15666] = 32'b00000000000000000000001011100010;
assign LUT_4[15667] = 32'b11111111111111111001010111011010;
assign LUT_4[15668] = 32'b11111111111111111101110001011010;
assign LUT_4[15669] = 32'b11111111111111110110111101010010;
assign LUT_4[15670] = 32'b11111111111111111101001011111110;
assign LUT_4[15671] = 32'b11111111111111110110010111110110;
assign LUT_4[15672] = 32'b11111111111111111001111101010011;
assign LUT_4[15673] = 32'b11111111111111110011001001001011;
assign LUT_4[15674] = 32'b11111111111111111001010111110111;
assign LUT_4[15675] = 32'b11111111111111110010100011101111;
assign LUT_4[15676] = 32'b11111111111111110110111101101111;
assign LUT_4[15677] = 32'b11111111111111110000001001100111;
assign LUT_4[15678] = 32'b11111111111111110110011000010011;
assign LUT_4[15679] = 32'b11111111111111101111100100001011;
assign LUT_4[15680] = 32'b00000000000000000101111011011101;
assign LUT_4[15681] = 32'b11111111111111111111000111010101;
assign LUT_4[15682] = 32'b00000000000000000101010110000001;
assign LUT_4[15683] = 32'b11111111111111111110100001111001;
assign LUT_4[15684] = 32'b00000000000000000010111011111001;
assign LUT_4[15685] = 32'b11111111111111111100000111110001;
assign LUT_4[15686] = 32'b00000000000000000010010110011101;
assign LUT_4[15687] = 32'b11111111111111111011100010010101;
assign LUT_4[15688] = 32'b11111111111111111111000111110010;
assign LUT_4[15689] = 32'b11111111111111111000010011101010;
assign LUT_4[15690] = 32'b11111111111111111110100010010110;
assign LUT_4[15691] = 32'b11111111111111110111101110001110;
assign LUT_4[15692] = 32'b11111111111111111100001000001110;
assign LUT_4[15693] = 32'b11111111111111110101010100000110;
assign LUT_4[15694] = 32'b11111111111111111011100010110010;
assign LUT_4[15695] = 32'b11111111111111110100101110101010;
assign LUT_4[15696] = 32'b00000000000000000011101101001011;
assign LUT_4[15697] = 32'b11111111111111111100111001000011;
assign LUT_4[15698] = 32'b00000000000000000011000111101111;
assign LUT_4[15699] = 32'b11111111111111111100010011100111;
assign LUT_4[15700] = 32'b00000000000000000000101101100111;
assign LUT_4[15701] = 32'b11111111111111111001111001011111;
assign LUT_4[15702] = 32'b00000000000000000000001000001011;
assign LUT_4[15703] = 32'b11111111111111111001010100000011;
assign LUT_4[15704] = 32'b11111111111111111100111001100000;
assign LUT_4[15705] = 32'b11111111111111110110000101011000;
assign LUT_4[15706] = 32'b11111111111111111100010100000100;
assign LUT_4[15707] = 32'b11111111111111110101011111111100;
assign LUT_4[15708] = 32'b11111111111111111001111001111100;
assign LUT_4[15709] = 32'b11111111111111110011000101110100;
assign LUT_4[15710] = 32'b11111111111111111001010100100000;
assign LUT_4[15711] = 32'b11111111111111110010100000011000;
assign LUT_4[15712] = 32'b00000000000000000100010110100100;
assign LUT_4[15713] = 32'b11111111111111111101100010011100;
assign LUT_4[15714] = 32'b00000000000000000011110001001000;
assign LUT_4[15715] = 32'b11111111111111111100111101000000;
assign LUT_4[15716] = 32'b00000000000000000001010111000000;
assign LUT_4[15717] = 32'b11111111111111111010100010111000;
assign LUT_4[15718] = 32'b00000000000000000000110001100100;
assign LUT_4[15719] = 32'b11111111111111111001111101011100;
assign LUT_4[15720] = 32'b11111111111111111101100010111001;
assign LUT_4[15721] = 32'b11111111111111110110101110110001;
assign LUT_4[15722] = 32'b11111111111111111100111101011101;
assign LUT_4[15723] = 32'b11111111111111110110001001010101;
assign LUT_4[15724] = 32'b11111111111111111010100011010101;
assign LUT_4[15725] = 32'b11111111111111110011101111001101;
assign LUT_4[15726] = 32'b11111111111111111001111101111001;
assign LUT_4[15727] = 32'b11111111111111110011001001110001;
assign LUT_4[15728] = 32'b00000000000000000010001000010010;
assign LUT_4[15729] = 32'b11111111111111111011010100001010;
assign LUT_4[15730] = 32'b00000000000000000001100010110110;
assign LUT_4[15731] = 32'b11111111111111111010101110101110;
assign LUT_4[15732] = 32'b11111111111111111111001000101110;
assign LUT_4[15733] = 32'b11111111111111111000010100100110;
assign LUT_4[15734] = 32'b11111111111111111110100011010010;
assign LUT_4[15735] = 32'b11111111111111110111101111001010;
assign LUT_4[15736] = 32'b11111111111111111011010100100111;
assign LUT_4[15737] = 32'b11111111111111110100100000011111;
assign LUT_4[15738] = 32'b11111111111111111010101111001011;
assign LUT_4[15739] = 32'b11111111111111110011111011000011;
assign LUT_4[15740] = 32'b11111111111111111000010101000011;
assign LUT_4[15741] = 32'b11111111111111110001100000111011;
assign LUT_4[15742] = 32'b11111111111111110111101111100111;
assign LUT_4[15743] = 32'b11111111111111110000111011011111;
assign LUT_4[15744] = 32'b00000000000000000111001010010001;
assign LUT_4[15745] = 32'b00000000000000000000010110001001;
assign LUT_4[15746] = 32'b00000000000000000110100100110101;
assign LUT_4[15747] = 32'b11111111111111111111110000101101;
assign LUT_4[15748] = 32'b00000000000000000100001010101101;
assign LUT_4[15749] = 32'b11111111111111111101010110100101;
assign LUT_4[15750] = 32'b00000000000000000011100101010001;
assign LUT_4[15751] = 32'b11111111111111111100110001001001;
assign LUT_4[15752] = 32'b00000000000000000000010110100110;
assign LUT_4[15753] = 32'b11111111111111111001100010011110;
assign LUT_4[15754] = 32'b11111111111111111111110001001010;
assign LUT_4[15755] = 32'b11111111111111111000111101000010;
assign LUT_4[15756] = 32'b11111111111111111101010111000010;
assign LUT_4[15757] = 32'b11111111111111110110100010111010;
assign LUT_4[15758] = 32'b11111111111111111100110001100110;
assign LUT_4[15759] = 32'b11111111111111110101111101011110;
assign LUT_4[15760] = 32'b00000000000000000100111011111111;
assign LUT_4[15761] = 32'b11111111111111111110000111110111;
assign LUT_4[15762] = 32'b00000000000000000100010110100011;
assign LUT_4[15763] = 32'b11111111111111111101100010011011;
assign LUT_4[15764] = 32'b00000000000000000001111100011011;
assign LUT_4[15765] = 32'b11111111111111111011001000010011;
assign LUT_4[15766] = 32'b00000000000000000001010110111111;
assign LUT_4[15767] = 32'b11111111111111111010100010110111;
assign LUT_4[15768] = 32'b11111111111111111110001000010100;
assign LUT_4[15769] = 32'b11111111111111110111010100001100;
assign LUT_4[15770] = 32'b11111111111111111101100010111000;
assign LUT_4[15771] = 32'b11111111111111110110101110110000;
assign LUT_4[15772] = 32'b11111111111111111011001000110000;
assign LUT_4[15773] = 32'b11111111111111110100010100101000;
assign LUT_4[15774] = 32'b11111111111111111010100011010100;
assign LUT_4[15775] = 32'b11111111111111110011101111001100;
assign LUT_4[15776] = 32'b00000000000000000101100101011000;
assign LUT_4[15777] = 32'b11111111111111111110110001010000;
assign LUT_4[15778] = 32'b00000000000000000100111111111100;
assign LUT_4[15779] = 32'b11111111111111111110001011110100;
assign LUT_4[15780] = 32'b00000000000000000010100101110100;
assign LUT_4[15781] = 32'b11111111111111111011110001101100;
assign LUT_4[15782] = 32'b00000000000000000010000000011000;
assign LUT_4[15783] = 32'b11111111111111111011001100010000;
assign LUT_4[15784] = 32'b11111111111111111110110001101101;
assign LUT_4[15785] = 32'b11111111111111110111111101100101;
assign LUT_4[15786] = 32'b11111111111111111110001100010001;
assign LUT_4[15787] = 32'b11111111111111110111011000001001;
assign LUT_4[15788] = 32'b11111111111111111011110010001001;
assign LUT_4[15789] = 32'b11111111111111110100111110000001;
assign LUT_4[15790] = 32'b11111111111111111011001100101101;
assign LUT_4[15791] = 32'b11111111111111110100011000100101;
assign LUT_4[15792] = 32'b00000000000000000011010111000110;
assign LUT_4[15793] = 32'b11111111111111111100100010111110;
assign LUT_4[15794] = 32'b00000000000000000010110001101010;
assign LUT_4[15795] = 32'b11111111111111111011111101100010;
assign LUT_4[15796] = 32'b00000000000000000000010111100010;
assign LUT_4[15797] = 32'b11111111111111111001100011011010;
assign LUT_4[15798] = 32'b11111111111111111111110010000110;
assign LUT_4[15799] = 32'b11111111111111111000111101111110;
assign LUT_4[15800] = 32'b11111111111111111100100011011011;
assign LUT_4[15801] = 32'b11111111111111110101101111010011;
assign LUT_4[15802] = 32'b11111111111111111011111101111111;
assign LUT_4[15803] = 32'b11111111111111110101001001110111;
assign LUT_4[15804] = 32'b11111111111111111001100011110111;
assign LUT_4[15805] = 32'b11111111111111110010101111101111;
assign LUT_4[15806] = 32'b11111111111111111000111110011011;
assign LUT_4[15807] = 32'b11111111111111110010001010010011;
assign LUT_4[15808] = 32'b00000000000000001000100001100101;
assign LUT_4[15809] = 32'b00000000000000000001101101011101;
assign LUT_4[15810] = 32'b00000000000000000111111100001001;
assign LUT_4[15811] = 32'b00000000000000000001001000000001;
assign LUT_4[15812] = 32'b00000000000000000101100010000001;
assign LUT_4[15813] = 32'b11111111111111111110101101111001;
assign LUT_4[15814] = 32'b00000000000000000100111100100101;
assign LUT_4[15815] = 32'b11111111111111111110001000011101;
assign LUT_4[15816] = 32'b00000000000000000001101101111010;
assign LUT_4[15817] = 32'b11111111111111111010111001110010;
assign LUT_4[15818] = 32'b00000000000000000001001000011110;
assign LUT_4[15819] = 32'b11111111111111111010010100010110;
assign LUT_4[15820] = 32'b11111111111111111110101110010110;
assign LUT_4[15821] = 32'b11111111111111110111111010001110;
assign LUT_4[15822] = 32'b11111111111111111110001000111010;
assign LUT_4[15823] = 32'b11111111111111110111010100110010;
assign LUT_4[15824] = 32'b00000000000000000110010011010011;
assign LUT_4[15825] = 32'b11111111111111111111011111001011;
assign LUT_4[15826] = 32'b00000000000000000101101101110111;
assign LUT_4[15827] = 32'b11111111111111111110111001101111;
assign LUT_4[15828] = 32'b00000000000000000011010011101111;
assign LUT_4[15829] = 32'b11111111111111111100011111100111;
assign LUT_4[15830] = 32'b00000000000000000010101110010011;
assign LUT_4[15831] = 32'b11111111111111111011111010001011;
assign LUT_4[15832] = 32'b11111111111111111111011111101000;
assign LUT_4[15833] = 32'b11111111111111111000101011100000;
assign LUT_4[15834] = 32'b11111111111111111110111010001100;
assign LUT_4[15835] = 32'b11111111111111111000000110000100;
assign LUT_4[15836] = 32'b11111111111111111100100000000100;
assign LUT_4[15837] = 32'b11111111111111110101101011111100;
assign LUT_4[15838] = 32'b11111111111111111011111010101000;
assign LUT_4[15839] = 32'b11111111111111110101000110100000;
assign LUT_4[15840] = 32'b00000000000000000110111100101100;
assign LUT_4[15841] = 32'b00000000000000000000001000100100;
assign LUT_4[15842] = 32'b00000000000000000110010111010000;
assign LUT_4[15843] = 32'b11111111111111111111100011001000;
assign LUT_4[15844] = 32'b00000000000000000011111101001000;
assign LUT_4[15845] = 32'b11111111111111111101001001000000;
assign LUT_4[15846] = 32'b00000000000000000011010111101100;
assign LUT_4[15847] = 32'b11111111111111111100100011100100;
assign LUT_4[15848] = 32'b00000000000000000000001001000001;
assign LUT_4[15849] = 32'b11111111111111111001010100111001;
assign LUT_4[15850] = 32'b11111111111111111111100011100101;
assign LUT_4[15851] = 32'b11111111111111111000101111011101;
assign LUT_4[15852] = 32'b11111111111111111101001001011101;
assign LUT_4[15853] = 32'b11111111111111110110010101010101;
assign LUT_4[15854] = 32'b11111111111111111100100100000001;
assign LUT_4[15855] = 32'b11111111111111110101101111111001;
assign LUT_4[15856] = 32'b00000000000000000100101110011010;
assign LUT_4[15857] = 32'b11111111111111111101111010010010;
assign LUT_4[15858] = 32'b00000000000000000100001000111110;
assign LUT_4[15859] = 32'b11111111111111111101010100110110;
assign LUT_4[15860] = 32'b00000000000000000001101110110110;
assign LUT_4[15861] = 32'b11111111111111111010111010101110;
assign LUT_4[15862] = 32'b00000000000000000001001001011010;
assign LUT_4[15863] = 32'b11111111111111111010010101010010;
assign LUT_4[15864] = 32'b11111111111111111101111010101111;
assign LUT_4[15865] = 32'b11111111111111110111000110100111;
assign LUT_4[15866] = 32'b11111111111111111101010101010011;
assign LUT_4[15867] = 32'b11111111111111110110100001001011;
assign LUT_4[15868] = 32'b11111111111111111010111011001011;
assign LUT_4[15869] = 32'b11111111111111110100000111000011;
assign LUT_4[15870] = 32'b11111111111111111010010101101111;
assign LUT_4[15871] = 32'b11111111111111110011100001100111;
assign LUT_4[15872] = 32'b11111111111111111110101100101110;
assign LUT_4[15873] = 32'b11111111111111110111111000100110;
assign LUT_4[15874] = 32'b11111111111111111110000111010010;
assign LUT_4[15875] = 32'b11111111111111110111010011001010;
assign LUT_4[15876] = 32'b11111111111111111011101101001010;
assign LUT_4[15877] = 32'b11111111111111110100111001000010;
assign LUT_4[15878] = 32'b11111111111111111011000111101110;
assign LUT_4[15879] = 32'b11111111111111110100010011100110;
assign LUT_4[15880] = 32'b11111111111111110111111001000011;
assign LUT_4[15881] = 32'b11111111111111110001000100111011;
assign LUT_4[15882] = 32'b11111111111111110111010011100111;
assign LUT_4[15883] = 32'b11111111111111110000011111011111;
assign LUT_4[15884] = 32'b11111111111111110100111001011111;
assign LUT_4[15885] = 32'b11111111111111101110000101010111;
assign LUT_4[15886] = 32'b11111111111111110100010100000011;
assign LUT_4[15887] = 32'b11111111111111101101011111111011;
assign LUT_4[15888] = 32'b11111111111111111100011110011100;
assign LUT_4[15889] = 32'b11111111111111110101101010010100;
assign LUT_4[15890] = 32'b11111111111111111011111001000000;
assign LUT_4[15891] = 32'b11111111111111110101000100111000;
assign LUT_4[15892] = 32'b11111111111111111001011110111000;
assign LUT_4[15893] = 32'b11111111111111110010101010110000;
assign LUT_4[15894] = 32'b11111111111111111000111001011100;
assign LUT_4[15895] = 32'b11111111111111110010000101010100;
assign LUT_4[15896] = 32'b11111111111111110101101010110001;
assign LUT_4[15897] = 32'b11111111111111101110110110101001;
assign LUT_4[15898] = 32'b11111111111111110101000101010101;
assign LUT_4[15899] = 32'b11111111111111101110010001001101;
assign LUT_4[15900] = 32'b11111111111111110010101011001101;
assign LUT_4[15901] = 32'b11111111111111101011110111000101;
assign LUT_4[15902] = 32'b11111111111111110010000101110001;
assign LUT_4[15903] = 32'b11111111111111101011010001101001;
assign LUT_4[15904] = 32'b11111111111111111101000111110101;
assign LUT_4[15905] = 32'b11111111111111110110010011101101;
assign LUT_4[15906] = 32'b11111111111111111100100010011001;
assign LUT_4[15907] = 32'b11111111111111110101101110010001;
assign LUT_4[15908] = 32'b11111111111111111010001000010001;
assign LUT_4[15909] = 32'b11111111111111110011010100001001;
assign LUT_4[15910] = 32'b11111111111111111001100010110101;
assign LUT_4[15911] = 32'b11111111111111110010101110101101;
assign LUT_4[15912] = 32'b11111111111111110110010100001010;
assign LUT_4[15913] = 32'b11111111111111101111100000000010;
assign LUT_4[15914] = 32'b11111111111111110101101110101110;
assign LUT_4[15915] = 32'b11111111111111101110111010100110;
assign LUT_4[15916] = 32'b11111111111111110011010100100110;
assign LUT_4[15917] = 32'b11111111111111101100100000011110;
assign LUT_4[15918] = 32'b11111111111111110010101111001010;
assign LUT_4[15919] = 32'b11111111111111101011111011000010;
assign LUT_4[15920] = 32'b11111111111111111010111001100011;
assign LUT_4[15921] = 32'b11111111111111110100000101011011;
assign LUT_4[15922] = 32'b11111111111111111010010100000111;
assign LUT_4[15923] = 32'b11111111111111110011011111111111;
assign LUT_4[15924] = 32'b11111111111111110111111001111111;
assign LUT_4[15925] = 32'b11111111111111110001000101110111;
assign LUT_4[15926] = 32'b11111111111111110111010100100011;
assign LUT_4[15927] = 32'b11111111111111110000100000011011;
assign LUT_4[15928] = 32'b11111111111111110100000101111000;
assign LUT_4[15929] = 32'b11111111111111101101010001110000;
assign LUT_4[15930] = 32'b11111111111111110011100000011100;
assign LUT_4[15931] = 32'b11111111111111101100101100010100;
assign LUT_4[15932] = 32'b11111111111111110001000110010100;
assign LUT_4[15933] = 32'b11111111111111101010010010001100;
assign LUT_4[15934] = 32'b11111111111111110000100000111000;
assign LUT_4[15935] = 32'b11111111111111101001101100110000;
assign LUT_4[15936] = 32'b00000000000000000000000100000010;
assign LUT_4[15937] = 32'b11111111111111111001001111111010;
assign LUT_4[15938] = 32'b11111111111111111111011110100110;
assign LUT_4[15939] = 32'b11111111111111111000101010011110;
assign LUT_4[15940] = 32'b11111111111111111101000100011110;
assign LUT_4[15941] = 32'b11111111111111110110010000010110;
assign LUT_4[15942] = 32'b11111111111111111100011111000010;
assign LUT_4[15943] = 32'b11111111111111110101101010111010;
assign LUT_4[15944] = 32'b11111111111111111001010000010111;
assign LUT_4[15945] = 32'b11111111111111110010011100001111;
assign LUT_4[15946] = 32'b11111111111111111000101010111011;
assign LUT_4[15947] = 32'b11111111111111110001110110110011;
assign LUT_4[15948] = 32'b11111111111111110110010000110011;
assign LUT_4[15949] = 32'b11111111111111101111011100101011;
assign LUT_4[15950] = 32'b11111111111111110101101011010111;
assign LUT_4[15951] = 32'b11111111111111101110110111001111;
assign LUT_4[15952] = 32'b11111111111111111101110101110000;
assign LUT_4[15953] = 32'b11111111111111110111000001101000;
assign LUT_4[15954] = 32'b11111111111111111101010000010100;
assign LUT_4[15955] = 32'b11111111111111110110011100001100;
assign LUT_4[15956] = 32'b11111111111111111010110110001100;
assign LUT_4[15957] = 32'b11111111111111110100000010000100;
assign LUT_4[15958] = 32'b11111111111111111010010000110000;
assign LUT_4[15959] = 32'b11111111111111110011011100101000;
assign LUT_4[15960] = 32'b11111111111111110111000010000101;
assign LUT_4[15961] = 32'b11111111111111110000001101111101;
assign LUT_4[15962] = 32'b11111111111111110110011100101001;
assign LUT_4[15963] = 32'b11111111111111101111101000100001;
assign LUT_4[15964] = 32'b11111111111111110100000010100001;
assign LUT_4[15965] = 32'b11111111111111101101001110011001;
assign LUT_4[15966] = 32'b11111111111111110011011101000101;
assign LUT_4[15967] = 32'b11111111111111101100101000111101;
assign LUT_4[15968] = 32'b11111111111111111110011111001001;
assign LUT_4[15969] = 32'b11111111111111110111101011000001;
assign LUT_4[15970] = 32'b11111111111111111101111001101101;
assign LUT_4[15971] = 32'b11111111111111110111000101100101;
assign LUT_4[15972] = 32'b11111111111111111011011111100101;
assign LUT_4[15973] = 32'b11111111111111110100101011011101;
assign LUT_4[15974] = 32'b11111111111111111010111010001001;
assign LUT_4[15975] = 32'b11111111111111110100000110000001;
assign LUT_4[15976] = 32'b11111111111111110111101011011110;
assign LUT_4[15977] = 32'b11111111111111110000110111010110;
assign LUT_4[15978] = 32'b11111111111111110111000110000010;
assign LUT_4[15979] = 32'b11111111111111110000010001111010;
assign LUT_4[15980] = 32'b11111111111111110100101011111010;
assign LUT_4[15981] = 32'b11111111111111101101110111110010;
assign LUT_4[15982] = 32'b11111111111111110100000110011110;
assign LUT_4[15983] = 32'b11111111111111101101010010010110;
assign LUT_4[15984] = 32'b11111111111111111100010000110111;
assign LUT_4[15985] = 32'b11111111111111110101011100101111;
assign LUT_4[15986] = 32'b11111111111111111011101011011011;
assign LUT_4[15987] = 32'b11111111111111110100110111010011;
assign LUT_4[15988] = 32'b11111111111111111001010001010011;
assign LUT_4[15989] = 32'b11111111111111110010011101001011;
assign LUT_4[15990] = 32'b11111111111111111000101011110111;
assign LUT_4[15991] = 32'b11111111111111110001110111101111;
assign LUT_4[15992] = 32'b11111111111111110101011101001100;
assign LUT_4[15993] = 32'b11111111111111101110101001000100;
assign LUT_4[15994] = 32'b11111111111111110100110111110000;
assign LUT_4[15995] = 32'b11111111111111101110000011101000;
assign LUT_4[15996] = 32'b11111111111111110010011101101000;
assign LUT_4[15997] = 32'b11111111111111101011101001100000;
assign LUT_4[15998] = 32'b11111111111111110001111000001100;
assign LUT_4[15999] = 32'b11111111111111101011000100000100;
assign LUT_4[16000] = 32'b00000000000000000001010010110110;
assign LUT_4[16001] = 32'b11111111111111111010011110101110;
assign LUT_4[16002] = 32'b00000000000000000000101101011010;
assign LUT_4[16003] = 32'b11111111111111111001111001010010;
assign LUT_4[16004] = 32'b11111111111111111110010011010010;
assign LUT_4[16005] = 32'b11111111111111110111011111001010;
assign LUT_4[16006] = 32'b11111111111111111101101101110110;
assign LUT_4[16007] = 32'b11111111111111110110111001101110;
assign LUT_4[16008] = 32'b11111111111111111010011111001011;
assign LUT_4[16009] = 32'b11111111111111110011101011000011;
assign LUT_4[16010] = 32'b11111111111111111001111001101111;
assign LUT_4[16011] = 32'b11111111111111110011000101100111;
assign LUT_4[16012] = 32'b11111111111111110111011111100111;
assign LUT_4[16013] = 32'b11111111111111110000101011011111;
assign LUT_4[16014] = 32'b11111111111111110110111010001011;
assign LUT_4[16015] = 32'b11111111111111110000000110000011;
assign LUT_4[16016] = 32'b11111111111111111111000100100100;
assign LUT_4[16017] = 32'b11111111111111111000010000011100;
assign LUT_4[16018] = 32'b11111111111111111110011111001000;
assign LUT_4[16019] = 32'b11111111111111110111101011000000;
assign LUT_4[16020] = 32'b11111111111111111100000101000000;
assign LUT_4[16021] = 32'b11111111111111110101010000111000;
assign LUT_4[16022] = 32'b11111111111111111011011111100100;
assign LUT_4[16023] = 32'b11111111111111110100101011011100;
assign LUT_4[16024] = 32'b11111111111111111000010000111001;
assign LUT_4[16025] = 32'b11111111111111110001011100110001;
assign LUT_4[16026] = 32'b11111111111111110111101011011101;
assign LUT_4[16027] = 32'b11111111111111110000110111010101;
assign LUT_4[16028] = 32'b11111111111111110101010001010101;
assign LUT_4[16029] = 32'b11111111111111101110011101001101;
assign LUT_4[16030] = 32'b11111111111111110100101011111001;
assign LUT_4[16031] = 32'b11111111111111101101110111110001;
assign LUT_4[16032] = 32'b11111111111111111111101101111101;
assign LUT_4[16033] = 32'b11111111111111111000111001110101;
assign LUT_4[16034] = 32'b11111111111111111111001000100001;
assign LUT_4[16035] = 32'b11111111111111111000010100011001;
assign LUT_4[16036] = 32'b11111111111111111100101110011001;
assign LUT_4[16037] = 32'b11111111111111110101111010010001;
assign LUT_4[16038] = 32'b11111111111111111100001000111101;
assign LUT_4[16039] = 32'b11111111111111110101010100110101;
assign LUT_4[16040] = 32'b11111111111111111000111010010010;
assign LUT_4[16041] = 32'b11111111111111110010000110001010;
assign LUT_4[16042] = 32'b11111111111111111000010100110110;
assign LUT_4[16043] = 32'b11111111111111110001100000101110;
assign LUT_4[16044] = 32'b11111111111111110101111010101110;
assign LUT_4[16045] = 32'b11111111111111101111000110100110;
assign LUT_4[16046] = 32'b11111111111111110101010101010010;
assign LUT_4[16047] = 32'b11111111111111101110100001001010;
assign LUT_4[16048] = 32'b11111111111111111101011111101011;
assign LUT_4[16049] = 32'b11111111111111110110101011100011;
assign LUT_4[16050] = 32'b11111111111111111100111010001111;
assign LUT_4[16051] = 32'b11111111111111110110000110000111;
assign LUT_4[16052] = 32'b11111111111111111010100000000111;
assign LUT_4[16053] = 32'b11111111111111110011101011111111;
assign LUT_4[16054] = 32'b11111111111111111001111010101011;
assign LUT_4[16055] = 32'b11111111111111110011000110100011;
assign LUT_4[16056] = 32'b11111111111111110110101100000000;
assign LUT_4[16057] = 32'b11111111111111101111110111111000;
assign LUT_4[16058] = 32'b11111111111111110110000110100100;
assign LUT_4[16059] = 32'b11111111111111101111010010011100;
assign LUT_4[16060] = 32'b11111111111111110011101100011100;
assign LUT_4[16061] = 32'b11111111111111101100111000010100;
assign LUT_4[16062] = 32'b11111111111111110011000111000000;
assign LUT_4[16063] = 32'b11111111111111101100010010111000;
assign LUT_4[16064] = 32'b00000000000000000010101010001010;
assign LUT_4[16065] = 32'b11111111111111111011110110000010;
assign LUT_4[16066] = 32'b00000000000000000010000100101110;
assign LUT_4[16067] = 32'b11111111111111111011010000100110;
assign LUT_4[16068] = 32'b11111111111111111111101010100110;
assign LUT_4[16069] = 32'b11111111111111111000110110011110;
assign LUT_4[16070] = 32'b11111111111111111111000101001010;
assign LUT_4[16071] = 32'b11111111111111111000010001000010;
assign LUT_4[16072] = 32'b11111111111111111011110110011111;
assign LUT_4[16073] = 32'b11111111111111110101000010010111;
assign LUT_4[16074] = 32'b11111111111111111011010001000011;
assign LUT_4[16075] = 32'b11111111111111110100011100111011;
assign LUT_4[16076] = 32'b11111111111111111000110110111011;
assign LUT_4[16077] = 32'b11111111111111110010000010110011;
assign LUT_4[16078] = 32'b11111111111111111000010001011111;
assign LUT_4[16079] = 32'b11111111111111110001011101010111;
assign LUT_4[16080] = 32'b00000000000000000000011011111000;
assign LUT_4[16081] = 32'b11111111111111111001100111110000;
assign LUT_4[16082] = 32'b11111111111111111111110110011100;
assign LUT_4[16083] = 32'b11111111111111111001000010010100;
assign LUT_4[16084] = 32'b11111111111111111101011100010100;
assign LUT_4[16085] = 32'b11111111111111110110101000001100;
assign LUT_4[16086] = 32'b11111111111111111100110110111000;
assign LUT_4[16087] = 32'b11111111111111110110000010110000;
assign LUT_4[16088] = 32'b11111111111111111001101000001101;
assign LUT_4[16089] = 32'b11111111111111110010110100000101;
assign LUT_4[16090] = 32'b11111111111111111001000010110001;
assign LUT_4[16091] = 32'b11111111111111110010001110101001;
assign LUT_4[16092] = 32'b11111111111111110110101000101001;
assign LUT_4[16093] = 32'b11111111111111101111110100100001;
assign LUT_4[16094] = 32'b11111111111111110110000011001101;
assign LUT_4[16095] = 32'b11111111111111101111001111000101;
assign LUT_4[16096] = 32'b00000000000000000001000101010001;
assign LUT_4[16097] = 32'b11111111111111111010010001001001;
assign LUT_4[16098] = 32'b00000000000000000000011111110101;
assign LUT_4[16099] = 32'b11111111111111111001101011101101;
assign LUT_4[16100] = 32'b11111111111111111110000101101101;
assign LUT_4[16101] = 32'b11111111111111110111010001100101;
assign LUT_4[16102] = 32'b11111111111111111101100000010001;
assign LUT_4[16103] = 32'b11111111111111110110101100001001;
assign LUT_4[16104] = 32'b11111111111111111010010001100110;
assign LUT_4[16105] = 32'b11111111111111110011011101011110;
assign LUT_4[16106] = 32'b11111111111111111001101100001010;
assign LUT_4[16107] = 32'b11111111111111110010111000000010;
assign LUT_4[16108] = 32'b11111111111111110111010010000010;
assign LUT_4[16109] = 32'b11111111111111110000011101111010;
assign LUT_4[16110] = 32'b11111111111111110110101100100110;
assign LUT_4[16111] = 32'b11111111111111101111111000011110;
assign LUT_4[16112] = 32'b11111111111111111110110110111111;
assign LUT_4[16113] = 32'b11111111111111111000000010110111;
assign LUT_4[16114] = 32'b11111111111111111110010001100011;
assign LUT_4[16115] = 32'b11111111111111110111011101011011;
assign LUT_4[16116] = 32'b11111111111111111011110111011011;
assign LUT_4[16117] = 32'b11111111111111110101000011010011;
assign LUT_4[16118] = 32'b11111111111111111011010001111111;
assign LUT_4[16119] = 32'b11111111111111110100011101110111;
assign LUT_4[16120] = 32'b11111111111111111000000011010100;
assign LUT_4[16121] = 32'b11111111111111110001001111001100;
assign LUT_4[16122] = 32'b11111111111111110111011101111000;
assign LUT_4[16123] = 32'b11111111111111110000101001110000;
assign LUT_4[16124] = 32'b11111111111111110101000011110000;
assign LUT_4[16125] = 32'b11111111111111101110001111101000;
assign LUT_4[16126] = 32'b11111111111111110100011110010100;
assign LUT_4[16127] = 32'b11111111111111101101101010001100;
assign LUT_4[16128] = 32'b00000000000000000011101000010001;
assign LUT_4[16129] = 32'b11111111111111111100110100001001;
assign LUT_4[16130] = 32'b00000000000000000011000010110101;
assign LUT_4[16131] = 32'b11111111111111111100001110101101;
assign LUT_4[16132] = 32'b00000000000000000000101000101101;
assign LUT_4[16133] = 32'b11111111111111111001110100100101;
assign LUT_4[16134] = 32'b00000000000000000000000011010001;
assign LUT_4[16135] = 32'b11111111111111111001001111001001;
assign LUT_4[16136] = 32'b11111111111111111100110100100110;
assign LUT_4[16137] = 32'b11111111111111110110000000011110;
assign LUT_4[16138] = 32'b11111111111111111100001111001010;
assign LUT_4[16139] = 32'b11111111111111110101011011000010;
assign LUT_4[16140] = 32'b11111111111111111001110101000010;
assign LUT_4[16141] = 32'b11111111111111110011000000111010;
assign LUT_4[16142] = 32'b11111111111111111001001111100110;
assign LUT_4[16143] = 32'b11111111111111110010011011011110;
assign LUT_4[16144] = 32'b00000000000000000001011001111111;
assign LUT_4[16145] = 32'b11111111111111111010100101110111;
assign LUT_4[16146] = 32'b00000000000000000000110100100011;
assign LUT_4[16147] = 32'b11111111111111111010000000011011;
assign LUT_4[16148] = 32'b11111111111111111110011010011011;
assign LUT_4[16149] = 32'b11111111111111110111100110010011;
assign LUT_4[16150] = 32'b11111111111111111101110100111111;
assign LUT_4[16151] = 32'b11111111111111110111000000110111;
assign LUT_4[16152] = 32'b11111111111111111010100110010100;
assign LUT_4[16153] = 32'b11111111111111110011110010001100;
assign LUT_4[16154] = 32'b11111111111111111010000000111000;
assign LUT_4[16155] = 32'b11111111111111110011001100110000;
assign LUT_4[16156] = 32'b11111111111111110111100110110000;
assign LUT_4[16157] = 32'b11111111111111110000110010101000;
assign LUT_4[16158] = 32'b11111111111111110111000001010100;
assign LUT_4[16159] = 32'b11111111111111110000001101001100;
assign LUT_4[16160] = 32'b00000000000000000010000011011000;
assign LUT_4[16161] = 32'b11111111111111111011001111010000;
assign LUT_4[16162] = 32'b00000000000000000001011101111100;
assign LUT_4[16163] = 32'b11111111111111111010101001110100;
assign LUT_4[16164] = 32'b11111111111111111111000011110100;
assign LUT_4[16165] = 32'b11111111111111111000001111101100;
assign LUT_4[16166] = 32'b11111111111111111110011110011000;
assign LUT_4[16167] = 32'b11111111111111110111101010010000;
assign LUT_4[16168] = 32'b11111111111111111011001111101101;
assign LUT_4[16169] = 32'b11111111111111110100011011100101;
assign LUT_4[16170] = 32'b11111111111111111010101010010001;
assign LUT_4[16171] = 32'b11111111111111110011110110001001;
assign LUT_4[16172] = 32'b11111111111111111000010000001001;
assign LUT_4[16173] = 32'b11111111111111110001011100000001;
assign LUT_4[16174] = 32'b11111111111111110111101010101101;
assign LUT_4[16175] = 32'b11111111111111110000110110100101;
assign LUT_4[16176] = 32'b11111111111111111111110101000110;
assign LUT_4[16177] = 32'b11111111111111111001000000111110;
assign LUT_4[16178] = 32'b11111111111111111111001111101010;
assign LUT_4[16179] = 32'b11111111111111111000011011100010;
assign LUT_4[16180] = 32'b11111111111111111100110101100010;
assign LUT_4[16181] = 32'b11111111111111110110000001011010;
assign LUT_4[16182] = 32'b11111111111111111100010000000110;
assign LUT_4[16183] = 32'b11111111111111110101011011111110;
assign LUT_4[16184] = 32'b11111111111111111001000001011011;
assign LUT_4[16185] = 32'b11111111111111110010001101010011;
assign LUT_4[16186] = 32'b11111111111111111000011011111111;
assign LUT_4[16187] = 32'b11111111111111110001100111110111;
assign LUT_4[16188] = 32'b11111111111111110110000001110111;
assign LUT_4[16189] = 32'b11111111111111101111001101101111;
assign LUT_4[16190] = 32'b11111111111111110101011100011011;
assign LUT_4[16191] = 32'b11111111111111101110101000010011;
assign LUT_4[16192] = 32'b00000000000000000100111111100101;
assign LUT_4[16193] = 32'b11111111111111111110001011011101;
assign LUT_4[16194] = 32'b00000000000000000100011010001001;
assign LUT_4[16195] = 32'b11111111111111111101100110000001;
assign LUT_4[16196] = 32'b00000000000000000010000000000001;
assign LUT_4[16197] = 32'b11111111111111111011001011111001;
assign LUT_4[16198] = 32'b00000000000000000001011010100101;
assign LUT_4[16199] = 32'b11111111111111111010100110011101;
assign LUT_4[16200] = 32'b11111111111111111110001011111010;
assign LUT_4[16201] = 32'b11111111111111110111010111110010;
assign LUT_4[16202] = 32'b11111111111111111101100110011110;
assign LUT_4[16203] = 32'b11111111111111110110110010010110;
assign LUT_4[16204] = 32'b11111111111111111011001100010110;
assign LUT_4[16205] = 32'b11111111111111110100011000001110;
assign LUT_4[16206] = 32'b11111111111111111010100110111010;
assign LUT_4[16207] = 32'b11111111111111110011110010110010;
assign LUT_4[16208] = 32'b00000000000000000010110001010011;
assign LUT_4[16209] = 32'b11111111111111111011111101001011;
assign LUT_4[16210] = 32'b00000000000000000010001011110111;
assign LUT_4[16211] = 32'b11111111111111111011010111101111;
assign LUT_4[16212] = 32'b11111111111111111111110001101111;
assign LUT_4[16213] = 32'b11111111111111111000111101100111;
assign LUT_4[16214] = 32'b11111111111111111111001100010011;
assign LUT_4[16215] = 32'b11111111111111111000011000001011;
assign LUT_4[16216] = 32'b11111111111111111011111101101000;
assign LUT_4[16217] = 32'b11111111111111110101001001100000;
assign LUT_4[16218] = 32'b11111111111111111011011000001100;
assign LUT_4[16219] = 32'b11111111111111110100100100000100;
assign LUT_4[16220] = 32'b11111111111111111000111110000100;
assign LUT_4[16221] = 32'b11111111111111110010001001111100;
assign LUT_4[16222] = 32'b11111111111111111000011000101000;
assign LUT_4[16223] = 32'b11111111111111110001100100100000;
assign LUT_4[16224] = 32'b00000000000000000011011010101100;
assign LUT_4[16225] = 32'b11111111111111111100100110100100;
assign LUT_4[16226] = 32'b00000000000000000010110101010000;
assign LUT_4[16227] = 32'b11111111111111111100000001001000;
assign LUT_4[16228] = 32'b00000000000000000000011011001000;
assign LUT_4[16229] = 32'b11111111111111111001100111000000;
assign LUT_4[16230] = 32'b11111111111111111111110101101100;
assign LUT_4[16231] = 32'b11111111111111111001000001100100;
assign LUT_4[16232] = 32'b11111111111111111100100111000001;
assign LUT_4[16233] = 32'b11111111111111110101110010111001;
assign LUT_4[16234] = 32'b11111111111111111100000001100101;
assign LUT_4[16235] = 32'b11111111111111110101001101011101;
assign LUT_4[16236] = 32'b11111111111111111001100111011101;
assign LUT_4[16237] = 32'b11111111111111110010110011010101;
assign LUT_4[16238] = 32'b11111111111111111001000010000001;
assign LUT_4[16239] = 32'b11111111111111110010001101111001;
assign LUT_4[16240] = 32'b00000000000000000001001100011010;
assign LUT_4[16241] = 32'b11111111111111111010011000010010;
assign LUT_4[16242] = 32'b00000000000000000000100110111110;
assign LUT_4[16243] = 32'b11111111111111111001110010110110;
assign LUT_4[16244] = 32'b11111111111111111110001100110110;
assign LUT_4[16245] = 32'b11111111111111110111011000101110;
assign LUT_4[16246] = 32'b11111111111111111101100111011010;
assign LUT_4[16247] = 32'b11111111111111110110110011010010;
assign LUT_4[16248] = 32'b11111111111111111010011000101111;
assign LUT_4[16249] = 32'b11111111111111110011100100100111;
assign LUT_4[16250] = 32'b11111111111111111001110011010011;
assign LUT_4[16251] = 32'b11111111111111110010111111001011;
assign LUT_4[16252] = 32'b11111111111111110111011001001011;
assign LUT_4[16253] = 32'b11111111111111110000100101000011;
assign LUT_4[16254] = 32'b11111111111111110110110011101111;
assign LUT_4[16255] = 32'b11111111111111101111111111100111;
assign LUT_4[16256] = 32'b00000000000000000110001110011001;
assign LUT_4[16257] = 32'b11111111111111111111011010010001;
assign LUT_4[16258] = 32'b00000000000000000101101000111101;
assign LUT_4[16259] = 32'b11111111111111111110110100110101;
assign LUT_4[16260] = 32'b00000000000000000011001110110101;
assign LUT_4[16261] = 32'b11111111111111111100011010101101;
assign LUT_4[16262] = 32'b00000000000000000010101001011001;
assign LUT_4[16263] = 32'b11111111111111111011110101010001;
assign LUT_4[16264] = 32'b11111111111111111111011010101110;
assign LUT_4[16265] = 32'b11111111111111111000100110100110;
assign LUT_4[16266] = 32'b11111111111111111110110101010010;
assign LUT_4[16267] = 32'b11111111111111111000000001001010;
assign LUT_4[16268] = 32'b11111111111111111100011011001010;
assign LUT_4[16269] = 32'b11111111111111110101100111000010;
assign LUT_4[16270] = 32'b11111111111111111011110101101110;
assign LUT_4[16271] = 32'b11111111111111110101000001100110;
assign LUT_4[16272] = 32'b00000000000000000100000000000111;
assign LUT_4[16273] = 32'b11111111111111111101001011111111;
assign LUT_4[16274] = 32'b00000000000000000011011010101011;
assign LUT_4[16275] = 32'b11111111111111111100100110100011;
assign LUT_4[16276] = 32'b00000000000000000001000000100011;
assign LUT_4[16277] = 32'b11111111111111111010001100011011;
assign LUT_4[16278] = 32'b00000000000000000000011011000111;
assign LUT_4[16279] = 32'b11111111111111111001100110111111;
assign LUT_4[16280] = 32'b11111111111111111101001100011100;
assign LUT_4[16281] = 32'b11111111111111110110011000010100;
assign LUT_4[16282] = 32'b11111111111111111100100111000000;
assign LUT_4[16283] = 32'b11111111111111110101110010111000;
assign LUT_4[16284] = 32'b11111111111111111010001100111000;
assign LUT_4[16285] = 32'b11111111111111110011011000110000;
assign LUT_4[16286] = 32'b11111111111111111001100111011100;
assign LUT_4[16287] = 32'b11111111111111110010110011010100;
assign LUT_4[16288] = 32'b00000000000000000100101001100000;
assign LUT_4[16289] = 32'b11111111111111111101110101011000;
assign LUT_4[16290] = 32'b00000000000000000100000100000100;
assign LUT_4[16291] = 32'b11111111111111111101001111111100;
assign LUT_4[16292] = 32'b00000000000000000001101001111100;
assign LUT_4[16293] = 32'b11111111111111111010110101110100;
assign LUT_4[16294] = 32'b00000000000000000001000100100000;
assign LUT_4[16295] = 32'b11111111111111111010010000011000;
assign LUT_4[16296] = 32'b11111111111111111101110101110101;
assign LUT_4[16297] = 32'b11111111111111110111000001101101;
assign LUT_4[16298] = 32'b11111111111111111101010000011001;
assign LUT_4[16299] = 32'b11111111111111110110011100010001;
assign LUT_4[16300] = 32'b11111111111111111010110110010001;
assign LUT_4[16301] = 32'b11111111111111110100000010001001;
assign LUT_4[16302] = 32'b11111111111111111010010000110101;
assign LUT_4[16303] = 32'b11111111111111110011011100101101;
assign LUT_4[16304] = 32'b00000000000000000010011011001110;
assign LUT_4[16305] = 32'b11111111111111111011100111000110;
assign LUT_4[16306] = 32'b00000000000000000001110101110010;
assign LUT_4[16307] = 32'b11111111111111111011000001101010;
assign LUT_4[16308] = 32'b11111111111111111111011011101010;
assign LUT_4[16309] = 32'b11111111111111111000100111100010;
assign LUT_4[16310] = 32'b11111111111111111110110110001110;
assign LUT_4[16311] = 32'b11111111111111111000000010000110;
assign LUT_4[16312] = 32'b11111111111111111011100111100011;
assign LUT_4[16313] = 32'b11111111111111110100110011011011;
assign LUT_4[16314] = 32'b11111111111111111011000010000111;
assign LUT_4[16315] = 32'b11111111111111110100001101111111;
assign LUT_4[16316] = 32'b11111111111111111000100111111111;
assign LUT_4[16317] = 32'b11111111111111110001110011110111;
assign LUT_4[16318] = 32'b11111111111111111000000010100011;
assign LUT_4[16319] = 32'b11111111111111110001001110011011;
assign LUT_4[16320] = 32'b00000000000000000111100101101101;
assign LUT_4[16321] = 32'b00000000000000000000110001100101;
assign LUT_4[16322] = 32'b00000000000000000111000000010001;
assign LUT_4[16323] = 32'b00000000000000000000001100001001;
assign LUT_4[16324] = 32'b00000000000000000100100110001001;
assign LUT_4[16325] = 32'b11111111111111111101110010000001;
assign LUT_4[16326] = 32'b00000000000000000100000000101101;
assign LUT_4[16327] = 32'b11111111111111111101001100100101;
assign LUT_4[16328] = 32'b00000000000000000000110010000010;
assign LUT_4[16329] = 32'b11111111111111111001111101111010;
assign LUT_4[16330] = 32'b00000000000000000000001100100110;
assign LUT_4[16331] = 32'b11111111111111111001011000011110;
assign LUT_4[16332] = 32'b11111111111111111101110010011110;
assign LUT_4[16333] = 32'b11111111111111110110111110010110;
assign LUT_4[16334] = 32'b11111111111111111101001101000010;
assign LUT_4[16335] = 32'b11111111111111110110011000111010;
assign LUT_4[16336] = 32'b00000000000000000101010111011011;
assign LUT_4[16337] = 32'b11111111111111111110100011010011;
assign LUT_4[16338] = 32'b00000000000000000100110001111111;
assign LUT_4[16339] = 32'b11111111111111111101111101110111;
assign LUT_4[16340] = 32'b00000000000000000010010111110111;
assign LUT_4[16341] = 32'b11111111111111111011100011101111;
assign LUT_4[16342] = 32'b00000000000000000001110010011011;
assign LUT_4[16343] = 32'b11111111111111111010111110010011;
assign LUT_4[16344] = 32'b11111111111111111110100011110000;
assign LUT_4[16345] = 32'b11111111111111110111101111101000;
assign LUT_4[16346] = 32'b11111111111111111101111110010100;
assign LUT_4[16347] = 32'b11111111111111110111001010001100;
assign LUT_4[16348] = 32'b11111111111111111011100100001100;
assign LUT_4[16349] = 32'b11111111111111110100110000000100;
assign LUT_4[16350] = 32'b11111111111111111010111110110000;
assign LUT_4[16351] = 32'b11111111111111110100001010101000;
assign LUT_4[16352] = 32'b00000000000000000110000000110100;
assign LUT_4[16353] = 32'b11111111111111111111001100101100;
assign LUT_4[16354] = 32'b00000000000000000101011011011000;
assign LUT_4[16355] = 32'b11111111111111111110100111010000;
assign LUT_4[16356] = 32'b00000000000000000011000001010000;
assign LUT_4[16357] = 32'b11111111111111111100001101001000;
assign LUT_4[16358] = 32'b00000000000000000010011011110100;
assign LUT_4[16359] = 32'b11111111111111111011100111101100;
assign LUT_4[16360] = 32'b11111111111111111111001101001001;
assign LUT_4[16361] = 32'b11111111111111111000011001000001;
assign LUT_4[16362] = 32'b11111111111111111110100111101101;
assign LUT_4[16363] = 32'b11111111111111110111110011100101;
assign LUT_4[16364] = 32'b11111111111111111100001101100101;
assign LUT_4[16365] = 32'b11111111111111110101011001011101;
assign LUT_4[16366] = 32'b11111111111111111011101000001001;
assign LUT_4[16367] = 32'b11111111111111110100110100000001;
assign LUT_4[16368] = 32'b00000000000000000011110010100010;
assign LUT_4[16369] = 32'b11111111111111111100111110011010;
assign LUT_4[16370] = 32'b00000000000000000011001101000110;
assign LUT_4[16371] = 32'b11111111111111111100011000111110;
assign LUT_4[16372] = 32'b00000000000000000000110010111110;
assign LUT_4[16373] = 32'b11111111111111111001111110110110;
assign LUT_4[16374] = 32'b00000000000000000000001101100010;
assign LUT_4[16375] = 32'b11111111111111111001011001011010;
assign LUT_4[16376] = 32'b11111111111111111100111110110111;
assign LUT_4[16377] = 32'b11111111111111110110001010101111;
assign LUT_4[16378] = 32'b11111111111111111100011001011011;
assign LUT_4[16379] = 32'b11111111111111110101100101010011;
assign LUT_4[16380] = 32'b11111111111111111001111111010011;
assign LUT_4[16381] = 32'b11111111111111110011001011001011;
assign LUT_4[16382] = 32'b11111111111111111001011001110111;
assign LUT_4[16383] = 32'b11111111111111110010100101101111;
assign LUT_4[16384] = 32'b00000000000000000101011101001100;
assign LUT_4[16385] = 32'b11111111111111111110101001000100;
assign LUT_4[16386] = 32'b00000000000000000100110111110000;
assign LUT_4[16387] = 32'b11111111111111111110000011101000;
assign LUT_4[16388] = 32'b00000000000000000010011101101000;
assign LUT_4[16389] = 32'b11111111111111111011101001100000;
assign LUT_4[16390] = 32'b00000000000000000001111000001100;
assign LUT_4[16391] = 32'b11111111111111111011000100000100;
assign LUT_4[16392] = 32'b11111111111111111110101001100001;
assign LUT_4[16393] = 32'b11111111111111110111110101011001;
assign LUT_4[16394] = 32'b11111111111111111110000100000101;
assign LUT_4[16395] = 32'b11111111111111110111001111111101;
assign LUT_4[16396] = 32'b11111111111111111011101001111101;
assign LUT_4[16397] = 32'b11111111111111110100110101110101;
assign LUT_4[16398] = 32'b11111111111111111011000100100001;
assign LUT_4[16399] = 32'b11111111111111110100010000011001;
assign LUT_4[16400] = 32'b00000000000000000011001110111010;
assign LUT_4[16401] = 32'b11111111111111111100011010110010;
assign LUT_4[16402] = 32'b00000000000000000010101001011110;
assign LUT_4[16403] = 32'b11111111111111111011110101010110;
assign LUT_4[16404] = 32'b00000000000000000000001111010110;
assign LUT_4[16405] = 32'b11111111111111111001011011001110;
assign LUT_4[16406] = 32'b11111111111111111111101001111010;
assign LUT_4[16407] = 32'b11111111111111111000110101110010;
assign LUT_4[16408] = 32'b11111111111111111100011011001111;
assign LUT_4[16409] = 32'b11111111111111110101100111000111;
assign LUT_4[16410] = 32'b11111111111111111011110101110011;
assign LUT_4[16411] = 32'b11111111111111110101000001101011;
assign LUT_4[16412] = 32'b11111111111111111001011011101011;
assign LUT_4[16413] = 32'b11111111111111110010100111100011;
assign LUT_4[16414] = 32'b11111111111111111000110110001111;
assign LUT_4[16415] = 32'b11111111111111110010000010000111;
assign LUT_4[16416] = 32'b00000000000000000011111000010011;
assign LUT_4[16417] = 32'b11111111111111111101000100001011;
assign LUT_4[16418] = 32'b00000000000000000011010010110111;
assign LUT_4[16419] = 32'b11111111111111111100011110101111;
assign LUT_4[16420] = 32'b00000000000000000000111000101111;
assign LUT_4[16421] = 32'b11111111111111111010000100100111;
assign LUT_4[16422] = 32'b00000000000000000000010011010011;
assign LUT_4[16423] = 32'b11111111111111111001011111001011;
assign LUT_4[16424] = 32'b11111111111111111101000100101000;
assign LUT_4[16425] = 32'b11111111111111110110010000100000;
assign LUT_4[16426] = 32'b11111111111111111100011111001100;
assign LUT_4[16427] = 32'b11111111111111110101101011000100;
assign LUT_4[16428] = 32'b11111111111111111010000101000100;
assign LUT_4[16429] = 32'b11111111111111110011010000111100;
assign LUT_4[16430] = 32'b11111111111111111001011111101000;
assign LUT_4[16431] = 32'b11111111111111110010101011100000;
assign LUT_4[16432] = 32'b00000000000000000001101010000001;
assign LUT_4[16433] = 32'b11111111111111111010110101111001;
assign LUT_4[16434] = 32'b00000000000000000001000100100101;
assign LUT_4[16435] = 32'b11111111111111111010010000011101;
assign LUT_4[16436] = 32'b11111111111111111110101010011101;
assign LUT_4[16437] = 32'b11111111111111110111110110010101;
assign LUT_4[16438] = 32'b11111111111111111110000101000001;
assign LUT_4[16439] = 32'b11111111111111110111010000111001;
assign LUT_4[16440] = 32'b11111111111111111010110110010110;
assign LUT_4[16441] = 32'b11111111111111110100000010001110;
assign LUT_4[16442] = 32'b11111111111111111010010000111010;
assign LUT_4[16443] = 32'b11111111111111110011011100110010;
assign LUT_4[16444] = 32'b11111111111111110111110110110010;
assign LUT_4[16445] = 32'b11111111111111110001000010101010;
assign LUT_4[16446] = 32'b11111111111111110111010001010110;
assign LUT_4[16447] = 32'b11111111111111110000011101001110;
assign LUT_4[16448] = 32'b00000000000000000110110100100000;
assign LUT_4[16449] = 32'b00000000000000000000000000011000;
assign LUT_4[16450] = 32'b00000000000000000110001111000100;
assign LUT_4[16451] = 32'b11111111111111111111011010111100;
assign LUT_4[16452] = 32'b00000000000000000011110100111100;
assign LUT_4[16453] = 32'b11111111111111111101000000110100;
assign LUT_4[16454] = 32'b00000000000000000011001111100000;
assign LUT_4[16455] = 32'b11111111111111111100011011011000;
assign LUT_4[16456] = 32'b00000000000000000000000000110101;
assign LUT_4[16457] = 32'b11111111111111111001001100101101;
assign LUT_4[16458] = 32'b11111111111111111111011011011001;
assign LUT_4[16459] = 32'b11111111111111111000100111010001;
assign LUT_4[16460] = 32'b11111111111111111101000001010001;
assign LUT_4[16461] = 32'b11111111111111110110001101001001;
assign LUT_4[16462] = 32'b11111111111111111100011011110101;
assign LUT_4[16463] = 32'b11111111111111110101100111101101;
assign LUT_4[16464] = 32'b00000000000000000100100110001110;
assign LUT_4[16465] = 32'b11111111111111111101110010000110;
assign LUT_4[16466] = 32'b00000000000000000100000000110010;
assign LUT_4[16467] = 32'b11111111111111111101001100101010;
assign LUT_4[16468] = 32'b00000000000000000001100110101010;
assign LUT_4[16469] = 32'b11111111111111111010110010100010;
assign LUT_4[16470] = 32'b00000000000000000001000001001110;
assign LUT_4[16471] = 32'b11111111111111111010001101000110;
assign LUT_4[16472] = 32'b11111111111111111101110010100011;
assign LUT_4[16473] = 32'b11111111111111110110111110011011;
assign LUT_4[16474] = 32'b11111111111111111101001101000111;
assign LUT_4[16475] = 32'b11111111111111110110011000111111;
assign LUT_4[16476] = 32'b11111111111111111010110010111111;
assign LUT_4[16477] = 32'b11111111111111110011111110110111;
assign LUT_4[16478] = 32'b11111111111111111010001101100011;
assign LUT_4[16479] = 32'b11111111111111110011011001011011;
assign LUT_4[16480] = 32'b00000000000000000101001111100111;
assign LUT_4[16481] = 32'b11111111111111111110011011011111;
assign LUT_4[16482] = 32'b00000000000000000100101010001011;
assign LUT_4[16483] = 32'b11111111111111111101110110000011;
assign LUT_4[16484] = 32'b00000000000000000010010000000011;
assign LUT_4[16485] = 32'b11111111111111111011011011111011;
assign LUT_4[16486] = 32'b00000000000000000001101010100111;
assign LUT_4[16487] = 32'b11111111111111111010110110011111;
assign LUT_4[16488] = 32'b11111111111111111110011011111100;
assign LUT_4[16489] = 32'b11111111111111110111100111110100;
assign LUT_4[16490] = 32'b11111111111111111101110110100000;
assign LUT_4[16491] = 32'b11111111111111110111000010011000;
assign LUT_4[16492] = 32'b11111111111111111011011100011000;
assign LUT_4[16493] = 32'b11111111111111110100101000010000;
assign LUT_4[16494] = 32'b11111111111111111010110110111100;
assign LUT_4[16495] = 32'b11111111111111110100000010110100;
assign LUT_4[16496] = 32'b00000000000000000011000001010101;
assign LUT_4[16497] = 32'b11111111111111111100001101001101;
assign LUT_4[16498] = 32'b00000000000000000010011011111001;
assign LUT_4[16499] = 32'b11111111111111111011100111110001;
assign LUT_4[16500] = 32'b00000000000000000000000001110001;
assign LUT_4[16501] = 32'b11111111111111111001001101101001;
assign LUT_4[16502] = 32'b11111111111111111111011100010101;
assign LUT_4[16503] = 32'b11111111111111111000101000001101;
assign LUT_4[16504] = 32'b11111111111111111100001101101010;
assign LUT_4[16505] = 32'b11111111111111110101011001100010;
assign LUT_4[16506] = 32'b11111111111111111011101000001110;
assign LUT_4[16507] = 32'b11111111111111110100110100000110;
assign LUT_4[16508] = 32'b11111111111111111001001110000110;
assign LUT_4[16509] = 32'b11111111111111110010011001111110;
assign LUT_4[16510] = 32'b11111111111111111000101000101010;
assign LUT_4[16511] = 32'b11111111111111110001110100100010;
assign LUT_4[16512] = 32'b00000000000000001000000011010100;
assign LUT_4[16513] = 32'b00000000000000000001001111001100;
assign LUT_4[16514] = 32'b00000000000000000111011101111000;
assign LUT_4[16515] = 32'b00000000000000000000101001110000;
assign LUT_4[16516] = 32'b00000000000000000101000011110000;
assign LUT_4[16517] = 32'b11111111111111111110001111101000;
assign LUT_4[16518] = 32'b00000000000000000100011110010100;
assign LUT_4[16519] = 32'b11111111111111111101101010001100;
assign LUT_4[16520] = 32'b00000000000000000001001111101001;
assign LUT_4[16521] = 32'b11111111111111111010011011100001;
assign LUT_4[16522] = 32'b00000000000000000000101010001101;
assign LUT_4[16523] = 32'b11111111111111111001110110000101;
assign LUT_4[16524] = 32'b11111111111111111110010000000101;
assign LUT_4[16525] = 32'b11111111111111110111011011111101;
assign LUT_4[16526] = 32'b11111111111111111101101010101001;
assign LUT_4[16527] = 32'b11111111111111110110110110100001;
assign LUT_4[16528] = 32'b00000000000000000101110101000010;
assign LUT_4[16529] = 32'b11111111111111111111000000111010;
assign LUT_4[16530] = 32'b00000000000000000101001111100110;
assign LUT_4[16531] = 32'b11111111111111111110011011011110;
assign LUT_4[16532] = 32'b00000000000000000010110101011110;
assign LUT_4[16533] = 32'b11111111111111111100000001010110;
assign LUT_4[16534] = 32'b00000000000000000010010000000010;
assign LUT_4[16535] = 32'b11111111111111111011011011111010;
assign LUT_4[16536] = 32'b11111111111111111111000001010111;
assign LUT_4[16537] = 32'b11111111111111111000001101001111;
assign LUT_4[16538] = 32'b11111111111111111110011011111011;
assign LUT_4[16539] = 32'b11111111111111110111100111110011;
assign LUT_4[16540] = 32'b11111111111111111100000001110011;
assign LUT_4[16541] = 32'b11111111111111110101001101101011;
assign LUT_4[16542] = 32'b11111111111111111011011100010111;
assign LUT_4[16543] = 32'b11111111111111110100101000001111;
assign LUT_4[16544] = 32'b00000000000000000110011110011011;
assign LUT_4[16545] = 32'b11111111111111111111101010010011;
assign LUT_4[16546] = 32'b00000000000000000101111000111111;
assign LUT_4[16547] = 32'b11111111111111111111000100110111;
assign LUT_4[16548] = 32'b00000000000000000011011110110111;
assign LUT_4[16549] = 32'b11111111111111111100101010101111;
assign LUT_4[16550] = 32'b00000000000000000010111001011011;
assign LUT_4[16551] = 32'b11111111111111111100000101010011;
assign LUT_4[16552] = 32'b11111111111111111111101010110000;
assign LUT_4[16553] = 32'b11111111111111111000110110101000;
assign LUT_4[16554] = 32'b11111111111111111111000101010100;
assign LUT_4[16555] = 32'b11111111111111111000010001001100;
assign LUT_4[16556] = 32'b11111111111111111100101011001100;
assign LUT_4[16557] = 32'b11111111111111110101110111000100;
assign LUT_4[16558] = 32'b11111111111111111100000101110000;
assign LUT_4[16559] = 32'b11111111111111110101010001101000;
assign LUT_4[16560] = 32'b00000000000000000100010000001001;
assign LUT_4[16561] = 32'b11111111111111111101011100000001;
assign LUT_4[16562] = 32'b00000000000000000011101010101101;
assign LUT_4[16563] = 32'b11111111111111111100110110100101;
assign LUT_4[16564] = 32'b00000000000000000001010000100101;
assign LUT_4[16565] = 32'b11111111111111111010011100011101;
assign LUT_4[16566] = 32'b00000000000000000000101011001001;
assign LUT_4[16567] = 32'b11111111111111111001110111000001;
assign LUT_4[16568] = 32'b11111111111111111101011100011110;
assign LUT_4[16569] = 32'b11111111111111110110101000010110;
assign LUT_4[16570] = 32'b11111111111111111100110111000010;
assign LUT_4[16571] = 32'b11111111111111110110000010111010;
assign LUT_4[16572] = 32'b11111111111111111010011100111010;
assign LUT_4[16573] = 32'b11111111111111110011101000110010;
assign LUT_4[16574] = 32'b11111111111111111001110111011110;
assign LUT_4[16575] = 32'b11111111111111110011000011010110;
assign LUT_4[16576] = 32'b00000000000000001001011010101000;
assign LUT_4[16577] = 32'b00000000000000000010100110100000;
assign LUT_4[16578] = 32'b00000000000000001000110101001100;
assign LUT_4[16579] = 32'b00000000000000000010000001000100;
assign LUT_4[16580] = 32'b00000000000000000110011011000100;
assign LUT_4[16581] = 32'b11111111111111111111100110111100;
assign LUT_4[16582] = 32'b00000000000000000101110101101000;
assign LUT_4[16583] = 32'b11111111111111111111000001100000;
assign LUT_4[16584] = 32'b00000000000000000010100110111101;
assign LUT_4[16585] = 32'b11111111111111111011110010110101;
assign LUT_4[16586] = 32'b00000000000000000010000001100001;
assign LUT_4[16587] = 32'b11111111111111111011001101011001;
assign LUT_4[16588] = 32'b11111111111111111111100111011001;
assign LUT_4[16589] = 32'b11111111111111111000110011010001;
assign LUT_4[16590] = 32'b11111111111111111111000001111101;
assign LUT_4[16591] = 32'b11111111111111111000001101110101;
assign LUT_4[16592] = 32'b00000000000000000111001100010110;
assign LUT_4[16593] = 32'b00000000000000000000011000001110;
assign LUT_4[16594] = 32'b00000000000000000110100110111010;
assign LUT_4[16595] = 32'b11111111111111111111110010110010;
assign LUT_4[16596] = 32'b00000000000000000100001100110010;
assign LUT_4[16597] = 32'b11111111111111111101011000101010;
assign LUT_4[16598] = 32'b00000000000000000011100111010110;
assign LUT_4[16599] = 32'b11111111111111111100110011001110;
assign LUT_4[16600] = 32'b00000000000000000000011000101011;
assign LUT_4[16601] = 32'b11111111111111111001100100100011;
assign LUT_4[16602] = 32'b11111111111111111111110011001111;
assign LUT_4[16603] = 32'b11111111111111111000111111000111;
assign LUT_4[16604] = 32'b11111111111111111101011001000111;
assign LUT_4[16605] = 32'b11111111111111110110100100111111;
assign LUT_4[16606] = 32'b11111111111111111100110011101011;
assign LUT_4[16607] = 32'b11111111111111110101111111100011;
assign LUT_4[16608] = 32'b00000000000000000111110101101111;
assign LUT_4[16609] = 32'b00000000000000000001000001100111;
assign LUT_4[16610] = 32'b00000000000000000111010000010011;
assign LUT_4[16611] = 32'b00000000000000000000011100001011;
assign LUT_4[16612] = 32'b00000000000000000100110110001011;
assign LUT_4[16613] = 32'b11111111111111111110000010000011;
assign LUT_4[16614] = 32'b00000000000000000100010000101111;
assign LUT_4[16615] = 32'b11111111111111111101011100100111;
assign LUT_4[16616] = 32'b00000000000000000001000010000100;
assign LUT_4[16617] = 32'b11111111111111111010001101111100;
assign LUT_4[16618] = 32'b00000000000000000000011100101000;
assign LUT_4[16619] = 32'b11111111111111111001101000100000;
assign LUT_4[16620] = 32'b11111111111111111110000010100000;
assign LUT_4[16621] = 32'b11111111111111110111001110011000;
assign LUT_4[16622] = 32'b11111111111111111101011101000100;
assign LUT_4[16623] = 32'b11111111111111110110101000111100;
assign LUT_4[16624] = 32'b00000000000000000101100111011101;
assign LUT_4[16625] = 32'b11111111111111111110110011010101;
assign LUT_4[16626] = 32'b00000000000000000101000010000001;
assign LUT_4[16627] = 32'b11111111111111111110001101111001;
assign LUT_4[16628] = 32'b00000000000000000010100111111001;
assign LUT_4[16629] = 32'b11111111111111111011110011110001;
assign LUT_4[16630] = 32'b00000000000000000010000010011101;
assign LUT_4[16631] = 32'b11111111111111111011001110010101;
assign LUT_4[16632] = 32'b11111111111111111110110011110010;
assign LUT_4[16633] = 32'b11111111111111110111111111101010;
assign LUT_4[16634] = 32'b11111111111111111110001110010110;
assign LUT_4[16635] = 32'b11111111111111110111011010001110;
assign LUT_4[16636] = 32'b11111111111111111011110100001110;
assign LUT_4[16637] = 32'b11111111111111110101000000000110;
assign LUT_4[16638] = 32'b11111111111111111011001110110010;
assign LUT_4[16639] = 32'b11111111111111110100011010101010;
assign LUT_4[16640] = 32'b00000000000000001010011000101111;
assign LUT_4[16641] = 32'b00000000000000000011100100100111;
assign LUT_4[16642] = 32'b00000000000000001001110011010011;
assign LUT_4[16643] = 32'b00000000000000000010111111001011;
assign LUT_4[16644] = 32'b00000000000000000111011001001011;
assign LUT_4[16645] = 32'b00000000000000000000100101000011;
assign LUT_4[16646] = 32'b00000000000000000110110011101111;
assign LUT_4[16647] = 32'b11111111111111111111111111100111;
assign LUT_4[16648] = 32'b00000000000000000011100101000100;
assign LUT_4[16649] = 32'b11111111111111111100110000111100;
assign LUT_4[16650] = 32'b00000000000000000010111111101000;
assign LUT_4[16651] = 32'b11111111111111111100001011100000;
assign LUT_4[16652] = 32'b00000000000000000000100101100000;
assign LUT_4[16653] = 32'b11111111111111111001110001011000;
assign LUT_4[16654] = 32'b00000000000000000000000000000100;
assign LUT_4[16655] = 32'b11111111111111111001001011111100;
assign LUT_4[16656] = 32'b00000000000000001000001010011101;
assign LUT_4[16657] = 32'b00000000000000000001010110010101;
assign LUT_4[16658] = 32'b00000000000000000111100101000001;
assign LUT_4[16659] = 32'b00000000000000000000110000111001;
assign LUT_4[16660] = 32'b00000000000000000101001010111001;
assign LUT_4[16661] = 32'b11111111111111111110010110110001;
assign LUT_4[16662] = 32'b00000000000000000100100101011101;
assign LUT_4[16663] = 32'b11111111111111111101110001010101;
assign LUT_4[16664] = 32'b00000000000000000001010110110010;
assign LUT_4[16665] = 32'b11111111111111111010100010101010;
assign LUT_4[16666] = 32'b00000000000000000000110001010110;
assign LUT_4[16667] = 32'b11111111111111111001111101001110;
assign LUT_4[16668] = 32'b11111111111111111110010111001110;
assign LUT_4[16669] = 32'b11111111111111110111100011000110;
assign LUT_4[16670] = 32'b11111111111111111101110001110010;
assign LUT_4[16671] = 32'b11111111111111110110111101101010;
assign LUT_4[16672] = 32'b00000000000000001000110011110110;
assign LUT_4[16673] = 32'b00000000000000000001111111101110;
assign LUT_4[16674] = 32'b00000000000000001000001110011010;
assign LUT_4[16675] = 32'b00000000000000000001011010010010;
assign LUT_4[16676] = 32'b00000000000000000101110100010010;
assign LUT_4[16677] = 32'b11111111111111111111000000001010;
assign LUT_4[16678] = 32'b00000000000000000101001110110110;
assign LUT_4[16679] = 32'b11111111111111111110011010101110;
assign LUT_4[16680] = 32'b00000000000000000010000000001011;
assign LUT_4[16681] = 32'b11111111111111111011001100000011;
assign LUT_4[16682] = 32'b00000000000000000001011010101111;
assign LUT_4[16683] = 32'b11111111111111111010100110100111;
assign LUT_4[16684] = 32'b11111111111111111111000000100111;
assign LUT_4[16685] = 32'b11111111111111111000001100011111;
assign LUT_4[16686] = 32'b11111111111111111110011011001011;
assign LUT_4[16687] = 32'b11111111111111110111100111000011;
assign LUT_4[16688] = 32'b00000000000000000110100101100100;
assign LUT_4[16689] = 32'b11111111111111111111110001011100;
assign LUT_4[16690] = 32'b00000000000000000110000000001000;
assign LUT_4[16691] = 32'b11111111111111111111001100000000;
assign LUT_4[16692] = 32'b00000000000000000011100110000000;
assign LUT_4[16693] = 32'b11111111111111111100110001111000;
assign LUT_4[16694] = 32'b00000000000000000011000000100100;
assign LUT_4[16695] = 32'b11111111111111111100001100011100;
assign LUT_4[16696] = 32'b11111111111111111111110001111001;
assign LUT_4[16697] = 32'b11111111111111111000111101110001;
assign LUT_4[16698] = 32'b11111111111111111111001100011101;
assign LUT_4[16699] = 32'b11111111111111111000011000010101;
assign LUT_4[16700] = 32'b11111111111111111100110010010101;
assign LUT_4[16701] = 32'b11111111111111110101111110001101;
assign LUT_4[16702] = 32'b11111111111111111100001100111001;
assign LUT_4[16703] = 32'b11111111111111110101011000110001;
assign LUT_4[16704] = 32'b00000000000000001011110000000011;
assign LUT_4[16705] = 32'b00000000000000000100111011111011;
assign LUT_4[16706] = 32'b00000000000000001011001010100111;
assign LUT_4[16707] = 32'b00000000000000000100010110011111;
assign LUT_4[16708] = 32'b00000000000000001000110000011111;
assign LUT_4[16709] = 32'b00000000000000000001111100010111;
assign LUT_4[16710] = 32'b00000000000000001000001011000011;
assign LUT_4[16711] = 32'b00000000000000000001010110111011;
assign LUT_4[16712] = 32'b00000000000000000100111100011000;
assign LUT_4[16713] = 32'b11111111111111111110001000010000;
assign LUT_4[16714] = 32'b00000000000000000100010110111100;
assign LUT_4[16715] = 32'b11111111111111111101100010110100;
assign LUT_4[16716] = 32'b00000000000000000001111100110100;
assign LUT_4[16717] = 32'b11111111111111111011001000101100;
assign LUT_4[16718] = 32'b00000000000000000001010111011000;
assign LUT_4[16719] = 32'b11111111111111111010100011010000;
assign LUT_4[16720] = 32'b00000000000000001001100001110001;
assign LUT_4[16721] = 32'b00000000000000000010101101101001;
assign LUT_4[16722] = 32'b00000000000000001000111100010101;
assign LUT_4[16723] = 32'b00000000000000000010001000001101;
assign LUT_4[16724] = 32'b00000000000000000110100010001101;
assign LUT_4[16725] = 32'b11111111111111111111101110000101;
assign LUT_4[16726] = 32'b00000000000000000101111100110001;
assign LUT_4[16727] = 32'b11111111111111111111001000101001;
assign LUT_4[16728] = 32'b00000000000000000010101110000110;
assign LUT_4[16729] = 32'b11111111111111111011111001111110;
assign LUT_4[16730] = 32'b00000000000000000010001000101010;
assign LUT_4[16731] = 32'b11111111111111111011010100100010;
assign LUT_4[16732] = 32'b11111111111111111111101110100010;
assign LUT_4[16733] = 32'b11111111111111111000111010011010;
assign LUT_4[16734] = 32'b11111111111111111111001001000110;
assign LUT_4[16735] = 32'b11111111111111111000010100111110;
assign LUT_4[16736] = 32'b00000000000000001010001011001010;
assign LUT_4[16737] = 32'b00000000000000000011010111000010;
assign LUT_4[16738] = 32'b00000000000000001001100101101110;
assign LUT_4[16739] = 32'b00000000000000000010110001100110;
assign LUT_4[16740] = 32'b00000000000000000111001011100110;
assign LUT_4[16741] = 32'b00000000000000000000010111011110;
assign LUT_4[16742] = 32'b00000000000000000110100110001010;
assign LUT_4[16743] = 32'b11111111111111111111110010000010;
assign LUT_4[16744] = 32'b00000000000000000011010111011111;
assign LUT_4[16745] = 32'b11111111111111111100100011010111;
assign LUT_4[16746] = 32'b00000000000000000010110010000011;
assign LUT_4[16747] = 32'b11111111111111111011111101111011;
assign LUT_4[16748] = 32'b00000000000000000000010111111011;
assign LUT_4[16749] = 32'b11111111111111111001100011110011;
assign LUT_4[16750] = 32'b11111111111111111111110010011111;
assign LUT_4[16751] = 32'b11111111111111111000111110010111;
assign LUT_4[16752] = 32'b00000000000000000111111100111000;
assign LUT_4[16753] = 32'b00000000000000000001001000110000;
assign LUT_4[16754] = 32'b00000000000000000111010111011100;
assign LUT_4[16755] = 32'b00000000000000000000100011010100;
assign LUT_4[16756] = 32'b00000000000000000100111101010100;
assign LUT_4[16757] = 32'b11111111111111111110001001001100;
assign LUT_4[16758] = 32'b00000000000000000100010111111000;
assign LUT_4[16759] = 32'b11111111111111111101100011110000;
assign LUT_4[16760] = 32'b00000000000000000001001001001101;
assign LUT_4[16761] = 32'b11111111111111111010010101000101;
assign LUT_4[16762] = 32'b00000000000000000000100011110001;
assign LUT_4[16763] = 32'b11111111111111111001101111101001;
assign LUT_4[16764] = 32'b11111111111111111110001001101001;
assign LUT_4[16765] = 32'b11111111111111110111010101100001;
assign LUT_4[16766] = 32'b11111111111111111101100100001101;
assign LUT_4[16767] = 32'b11111111111111110110110000000101;
assign LUT_4[16768] = 32'b00000000000000001100111110110111;
assign LUT_4[16769] = 32'b00000000000000000110001010101111;
assign LUT_4[16770] = 32'b00000000000000001100011001011011;
assign LUT_4[16771] = 32'b00000000000000000101100101010011;
assign LUT_4[16772] = 32'b00000000000000001001111111010011;
assign LUT_4[16773] = 32'b00000000000000000011001011001011;
assign LUT_4[16774] = 32'b00000000000000001001011001110111;
assign LUT_4[16775] = 32'b00000000000000000010100101101111;
assign LUT_4[16776] = 32'b00000000000000000110001011001100;
assign LUT_4[16777] = 32'b11111111111111111111010111000100;
assign LUT_4[16778] = 32'b00000000000000000101100101110000;
assign LUT_4[16779] = 32'b11111111111111111110110001101000;
assign LUT_4[16780] = 32'b00000000000000000011001011101000;
assign LUT_4[16781] = 32'b11111111111111111100010111100000;
assign LUT_4[16782] = 32'b00000000000000000010100110001100;
assign LUT_4[16783] = 32'b11111111111111111011110010000100;
assign LUT_4[16784] = 32'b00000000000000001010110000100101;
assign LUT_4[16785] = 32'b00000000000000000011111100011101;
assign LUT_4[16786] = 32'b00000000000000001010001011001001;
assign LUT_4[16787] = 32'b00000000000000000011010111000001;
assign LUT_4[16788] = 32'b00000000000000000111110001000001;
assign LUT_4[16789] = 32'b00000000000000000000111100111001;
assign LUT_4[16790] = 32'b00000000000000000111001011100101;
assign LUT_4[16791] = 32'b00000000000000000000010111011101;
assign LUT_4[16792] = 32'b00000000000000000011111100111010;
assign LUT_4[16793] = 32'b11111111111111111101001000110010;
assign LUT_4[16794] = 32'b00000000000000000011010111011110;
assign LUT_4[16795] = 32'b11111111111111111100100011010110;
assign LUT_4[16796] = 32'b00000000000000000000111101010110;
assign LUT_4[16797] = 32'b11111111111111111010001001001110;
assign LUT_4[16798] = 32'b00000000000000000000010111111010;
assign LUT_4[16799] = 32'b11111111111111111001100011110010;
assign LUT_4[16800] = 32'b00000000000000001011011001111110;
assign LUT_4[16801] = 32'b00000000000000000100100101110110;
assign LUT_4[16802] = 32'b00000000000000001010110100100010;
assign LUT_4[16803] = 32'b00000000000000000100000000011010;
assign LUT_4[16804] = 32'b00000000000000001000011010011010;
assign LUT_4[16805] = 32'b00000000000000000001100110010010;
assign LUT_4[16806] = 32'b00000000000000000111110100111110;
assign LUT_4[16807] = 32'b00000000000000000001000000110110;
assign LUT_4[16808] = 32'b00000000000000000100100110010011;
assign LUT_4[16809] = 32'b11111111111111111101110010001011;
assign LUT_4[16810] = 32'b00000000000000000100000000110111;
assign LUT_4[16811] = 32'b11111111111111111101001100101111;
assign LUT_4[16812] = 32'b00000000000000000001100110101111;
assign LUT_4[16813] = 32'b11111111111111111010110010100111;
assign LUT_4[16814] = 32'b00000000000000000001000001010011;
assign LUT_4[16815] = 32'b11111111111111111010001101001011;
assign LUT_4[16816] = 32'b00000000000000001001001011101100;
assign LUT_4[16817] = 32'b00000000000000000010010111100100;
assign LUT_4[16818] = 32'b00000000000000001000100110010000;
assign LUT_4[16819] = 32'b00000000000000000001110010001000;
assign LUT_4[16820] = 32'b00000000000000000110001100001000;
assign LUT_4[16821] = 32'b11111111111111111111011000000000;
assign LUT_4[16822] = 32'b00000000000000000101100110101100;
assign LUT_4[16823] = 32'b11111111111111111110110010100100;
assign LUT_4[16824] = 32'b00000000000000000010011000000001;
assign LUT_4[16825] = 32'b11111111111111111011100011111001;
assign LUT_4[16826] = 32'b00000000000000000001110010100101;
assign LUT_4[16827] = 32'b11111111111111111010111110011101;
assign LUT_4[16828] = 32'b11111111111111111111011000011101;
assign LUT_4[16829] = 32'b11111111111111111000100100010101;
assign LUT_4[16830] = 32'b11111111111111111110110011000001;
assign LUT_4[16831] = 32'b11111111111111110111111110111001;
assign LUT_4[16832] = 32'b00000000000000001110010110001011;
assign LUT_4[16833] = 32'b00000000000000000111100010000011;
assign LUT_4[16834] = 32'b00000000000000001101110000101111;
assign LUT_4[16835] = 32'b00000000000000000110111100100111;
assign LUT_4[16836] = 32'b00000000000000001011010110100111;
assign LUT_4[16837] = 32'b00000000000000000100100010011111;
assign LUT_4[16838] = 32'b00000000000000001010110001001011;
assign LUT_4[16839] = 32'b00000000000000000011111101000011;
assign LUT_4[16840] = 32'b00000000000000000111100010100000;
assign LUT_4[16841] = 32'b00000000000000000000101110011000;
assign LUT_4[16842] = 32'b00000000000000000110111101000100;
assign LUT_4[16843] = 32'b00000000000000000000001000111100;
assign LUT_4[16844] = 32'b00000000000000000100100010111100;
assign LUT_4[16845] = 32'b11111111111111111101101110110100;
assign LUT_4[16846] = 32'b00000000000000000011111101100000;
assign LUT_4[16847] = 32'b11111111111111111101001001011000;
assign LUT_4[16848] = 32'b00000000000000001100000111111001;
assign LUT_4[16849] = 32'b00000000000000000101010011110001;
assign LUT_4[16850] = 32'b00000000000000001011100010011101;
assign LUT_4[16851] = 32'b00000000000000000100101110010101;
assign LUT_4[16852] = 32'b00000000000000001001001000010101;
assign LUT_4[16853] = 32'b00000000000000000010010100001101;
assign LUT_4[16854] = 32'b00000000000000001000100010111001;
assign LUT_4[16855] = 32'b00000000000000000001101110110001;
assign LUT_4[16856] = 32'b00000000000000000101010100001110;
assign LUT_4[16857] = 32'b11111111111111111110100000000110;
assign LUT_4[16858] = 32'b00000000000000000100101110110010;
assign LUT_4[16859] = 32'b11111111111111111101111010101010;
assign LUT_4[16860] = 32'b00000000000000000010010100101010;
assign LUT_4[16861] = 32'b11111111111111111011100000100010;
assign LUT_4[16862] = 32'b00000000000000000001101111001110;
assign LUT_4[16863] = 32'b11111111111111111010111011000110;
assign LUT_4[16864] = 32'b00000000000000001100110001010010;
assign LUT_4[16865] = 32'b00000000000000000101111101001010;
assign LUT_4[16866] = 32'b00000000000000001100001011110110;
assign LUT_4[16867] = 32'b00000000000000000101010111101110;
assign LUT_4[16868] = 32'b00000000000000001001110001101110;
assign LUT_4[16869] = 32'b00000000000000000010111101100110;
assign LUT_4[16870] = 32'b00000000000000001001001100010010;
assign LUT_4[16871] = 32'b00000000000000000010011000001010;
assign LUT_4[16872] = 32'b00000000000000000101111101100111;
assign LUT_4[16873] = 32'b11111111111111111111001001011111;
assign LUT_4[16874] = 32'b00000000000000000101011000001011;
assign LUT_4[16875] = 32'b11111111111111111110100100000011;
assign LUT_4[16876] = 32'b00000000000000000010111110000011;
assign LUT_4[16877] = 32'b11111111111111111100001001111011;
assign LUT_4[16878] = 32'b00000000000000000010011000100111;
assign LUT_4[16879] = 32'b11111111111111111011100100011111;
assign LUT_4[16880] = 32'b00000000000000001010100011000000;
assign LUT_4[16881] = 32'b00000000000000000011101110111000;
assign LUT_4[16882] = 32'b00000000000000001001111101100100;
assign LUT_4[16883] = 32'b00000000000000000011001001011100;
assign LUT_4[16884] = 32'b00000000000000000111100011011100;
assign LUT_4[16885] = 32'b00000000000000000000101111010100;
assign LUT_4[16886] = 32'b00000000000000000110111110000000;
assign LUT_4[16887] = 32'b00000000000000000000001001111000;
assign LUT_4[16888] = 32'b00000000000000000011101111010101;
assign LUT_4[16889] = 32'b11111111111111111100111011001101;
assign LUT_4[16890] = 32'b00000000000000000011001001111001;
assign LUT_4[16891] = 32'b11111111111111111100010101110001;
assign LUT_4[16892] = 32'b00000000000000000000101111110001;
assign LUT_4[16893] = 32'b11111111111111111001111011101001;
assign LUT_4[16894] = 32'b00000000000000000000001010010101;
assign LUT_4[16895] = 32'b11111111111111111001010110001101;
assign LUT_4[16896] = 32'b00000000000000000100100001010100;
assign LUT_4[16897] = 32'b11111111111111111101101101001100;
assign LUT_4[16898] = 32'b00000000000000000011111011111000;
assign LUT_4[16899] = 32'b11111111111111111101000111110000;
assign LUT_4[16900] = 32'b00000000000000000001100001110000;
assign LUT_4[16901] = 32'b11111111111111111010101101101000;
assign LUT_4[16902] = 32'b00000000000000000000111100010100;
assign LUT_4[16903] = 32'b11111111111111111010001000001100;
assign LUT_4[16904] = 32'b11111111111111111101101101101001;
assign LUT_4[16905] = 32'b11111111111111110110111001100001;
assign LUT_4[16906] = 32'b11111111111111111101001000001101;
assign LUT_4[16907] = 32'b11111111111111110110010100000101;
assign LUT_4[16908] = 32'b11111111111111111010101110000101;
assign LUT_4[16909] = 32'b11111111111111110011111001111101;
assign LUT_4[16910] = 32'b11111111111111111010001000101001;
assign LUT_4[16911] = 32'b11111111111111110011010100100001;
assign LUT_4[16912] = 32'b00000000000000000010010011000010;
assign LUT_4[16913] = 32'b11111111111111111011011110111010;
assign LUT_4[16914] = 32'b00000000000000000001101101100110;
assign LUT_4[16915] = 32'b11111111111111111010111001011110;
assign LUT_4[16916] = 32'b11111111111111111111010011011110;
assign LUT_4[16917] = 32'b11111111111111111000011111010110;
assign LUT_4[16918] = 32'b11111111111111111110101110000010;
assign LUT_4[16919] = 32'b11111111111111110111111001111010;
assign LUT_4[16920] = 32'b11111111111111111011011111010111;
assign LUT_4[16921] = 32'b11111111111111110100101011001111;
assign LUT_4[16922] = 32'b11111111111111111010111001111011;
assign LUT_4[16923] = 32'b11111111111111110100000101110011;
assign LUT_4[16924] = 32'b11111111111111111000011111110011;
assign LUT_4[16925] = 32'b11111111111111110001101011101011;
assign LUT_4[16926] = 32'b11111111111111110111111010010111;
assign LUT_4[16927] = 32'b11111111111111110001000110001111;
assign LUT_4[16928] = 32'b00000000000000000010111100011011;
assign LUT_4[16929] = 32'b11111111111111111100001000010011;
assign LUT_4[16930] = 32'b00000000000000000010010110111111;
assign LUT_4[16931] = 32'b11111111111111111011100010110111;
assign LUT_4[16932] = 32'b11111111111111111111111100110111;
assign LUT_4[16933] = 32'b11111111111111111001001000101111;
assign LUT_4[16934] = 32'b11111111111111111111010111011011;
assign LUT_4[16935] = 32'b11111111111111111000100011010011;
assign LUT_4[16936] = 32'b11111111111111111100001000110000;
assign LUT_4[16937] = 32'b11111111111111110101010100101000;
assign LUT_4[16938] = 32'b11111111111111111011100011010100;
assign LUT_4[16939] = 32'b11111111111111110100101111001100;
assign LUT_4[16940] = 32'b11111111111111111001001001001100;
assign LUT_4[16941] = 32'b11111111111111110010010101000100;
assign LUT_4[16942] = 32'b11111111111111111000100011110000;
assign LUT_4[16943] = 32'b11111111111111110001101111101000;
assign LUT_4[16944] = 32'b00000000000000000000101110001001;
assign LUT_4[16945] = 32'b11111111111111111001111010000001;
assign LUT_4[16946] = 32'b00000000000000000000001000101101;
assign LUT_4[16947] = 32'b11111111111111111001010100100101;
assign LUT_4[16948] = 32'b11111111111111111101101110100101;
assign LUT_4[16949] = 32'b11111111111111110110111010011101;
assign LUT_4[16950] = 32'b11111111111111111101001001001001;
assign LUT_4[16951] = 32'b11111111111111110110010101000001;
assign LUT_4[16952] = 32'b11111111111111111001111010011110;
assign LUT_4[16953] = 32'b11111111111111110011000110010110;
assign LUT_4[16954] = 32'b11111111111111111001010101000010;
assign LUT_4[16955] = 32'b11111111111111110010100000111010;
assign LUT_4[16956] = 32'b11111111111111110110111010111010;
assign LUT_4[16957] = 32'b11111111111111110000000110110010;
assign LUT_4[16958] = 32'b11111111111111110110010101011110;
assign LUT_4[16959] = 32'b11111111111111101111100001010110;
assign LUT_4[16960] = 32'b00000000000000000101111000101000;
assign LUT_4[16961] = 32'b11111111111111111111000100100000;
assign LUT_4[16962] = 32'b00000000000000000101010011001100;
assign LUT_4[16963] = 32'b11111111111111111110011111000100;
assign LUT_4[16964] = 32'b00000000000000000010111001000100;
assign LUT_4[16965] = 32'b11111111111111111100000100111100;
assign LUT_4[16966] = 32'b00000000000000000010010011101000;
assign LUT_4[16967] = 32'b11111111111111111011011111100000;
assign LUT_4[16968] = 32'b11111111111111111111000100111101;
assign LUT_4[16969] = 32'b11111111111111111000010000110101;
assign LUT_4[16970] = 32'b11111111111111111110011111100001;
assign LUT_4[16971] = 32'b11111111111111110111101011011001;
assign LUT_4[16972] = 32'b11111111111111111100000101011001;
assign LUT_4[16973] = 32'b11111111111111110101010001010001;
assign LUT_4[16974] = 32'b11111111111111111011011111111101;
assign LUT_4[16975] = 32'b11111111111111110100101011110101;
assign LUT_4[16976] = 32'b00000000000000000011101010010110;
assign LUT_4[16977] = 32'b11111111111111111100110110001110;
assign LUT_4[16978] = 32'b00000000000000000011000100111010;
assign LUT_4[16979] = 32'b11111111111111111100010000110010;
assign LUT_4[16980] = 32'b00000000000000000000101010110010;
assign LUT_4[16981] = 32'b11111111111111111001110110101010;
assign LUT_4[16982] = 32'b00000000000000000000000101010110;
assign LUT_4[16983] = 32'b11111111111111111001010001001110;
assign LUT_4[16984] = 32'b11111111111111111100110110101011;
assign LUT_4[16985] = 32'b11111111111111110110000010100011;
assign LUT_4[16986] = 32'b11111111111111111100010001001111;
assign LUT_4[16987] = 32'b11111111111111110101011101000111;
assign LUT_4[16988] = 32'b11111111111111111001110111000111;
assign LUT_4[16989] = 32'b11111111111111110011000010111111;
assign LUT_4[16990] = 32'b11111111111111111001010001101011;
assign LUT_4[16991] = 32'b11111111111111110010011101100011;
assign LUT_4[16992] = 32'b00000000000000000100010011101111;
assign LUT_4[16993] = 32'b11111111111111111101011111100111;
assign LUT_4[16994] = 32'b00000000000000000011101110010011;
assign LUT_4[16995] = 32'b11111111111111111100111010001011;
assign LUT_4[16996] = 32'b00000000000000000001010100001011;
assign LUT_4[16997] = 32'b11111111111111111010100000000011;
assign LUT_4[16998] = 32'b00000000000000000000101110101111;
assign LUT_4[16999] = 32'b11111111111111111001111010100111;
assign LUT_4[17000] = 32'b11111111111111111101100000000100;
assign LUT_4[17001] = 32'b11111111111111110110101011111100;
assign LUT_4[17002] = 32'b11111111111111111100111010101000;
assign LUT_4[17003] = 32'b11111111111111110110000110100000;
assign LUT_4[17004] = 32'b11111111111111111010100000100000;
assign LUT_4[17005] = 32'b11111111111111110011101100011000;
assign LUT_4[17006] = 32'b11111111111111111001111011000100;
assign LUT_4[17007] = 32'b11111111111111110011000110111100;
assign LUT_4[17008] = 32'b00000000000000000010000101011101;
assign LUT_4[17009] = 32'b11111111111111111011010001010101;
assign LUT_4[17010] = 32'b00000000000000000001100000000001;
assign LUT_4[17011] = 32'b11111111111111111010101011111001;
assign LUT_4[17012] = 32'b11111111111111111111000101111001;
assign LUT_4[17013] = 32'b11111111111111111000010001110001;
assign LUT_4[17014] = 32'b11111111111111111110100000011101;
assign LUT_4[17015] = 32'b11111111111111110111101100010101;
assign LUT_4[17016] = 32'b11111111111111111011010001110010;
assign LUT_4[17017] = 32'b11111111111111110100011101101010;
assign LUT_4[17018] = 32'b11111111111111111010101100010110;
assign LUT_4[17019] = 32'b11111111111111110011111000001110;
assign LUT_4[17020] = 32'b11111111111111111000010010001110;
assign LUT_4[17021] = 32'b11111111111111110001011110000110;
assign LUT_4[17022] = 32'b11111111111111110111101100110010;
assign LUT_4[17023] = 32'b11111111111111110000111000101010;
assign LUT_4[17024] = 32'b00000000000000000111000111011100;
assign LUT_4[17025] = 32'b00000000000000000000010011010100;
assign LUT_4[17026] = 32'b00000000000000000110100010000000;
assign LUT_4[17027] = 32'b11111111111111111111101101111000;
assign LUT_4[17028] = 32'b00000000000000000100000111111000;
assign LUT_4[17029] = 32'b11111111111111111101010011110000;
assign LUT_4[17030] = 32'b00000000000000000011100010011100;
assign LUT_4[17031] = 32'b11111111111111111100101110010100;
assign LUT_4[17032] = 32'b00000000000000000000010011110001;
assign LUT_4[17033] = 32'b11111111111111111001011111101001;
assign LUT_4[17034] = 32'b11111111111111111111101110010101;
assign LUT_4[17035] = 32'b11111111111111111000111010001101;
assign LUT_4[17036] = 32'b11111111111111111101010100001101;
assign LUT_4[17037] = 32'b11111111111111110110100000000101;
assign LUT_4[17038] = 32'b11111111111111111100101110110001;
assign LUT_4[17039] = 32'b11111111111111110101111010101001;
assign LUT_4[17040] = 32'b00000000000000000100111001001010;
assign LUT_4[17041] = 32'b11111111111111111110000101000010;
assign LUT_4[17042] = 32'b00000000000000000100010011101110;
assign LUT_4[17043] = 32'b11111111111111111101011111100110;
assign LUT_4[17044] = 32'b00000000000000000001111001100110;
assign LUT_4[17045] = 32'b11111111111111111011000101011110;
assign LUT_4[17046] = 32'b00000000000000000001010100001010;
assign LUT_4[17047] = 32'b11111111111111111010100000000010;
assign LUT_4[17048] = 32'b11111111111111111110000101011111;
assign LUT_4[17049] = 32'b11111111111111110111010001010111;
assign LUT_4[17050] = 32'b11111111111111111101100000000011;
assign LUT_4[17051] = 32'b11111111111111110110101011111011;
assign LUT_4[17052] = 32'b11111111111111111011000101111011;
assign LUT_4[17053] = 32'b11111111111111110100010001110011;
assign LUT_4[17054] = 32'b11111111111111111010100000011111;
assign LUT_4[17055] = 32'b11111111111111110011101100010111;
assign LUT_4[17056] = 32'b00000000000000000101100010100011;
assign LUT_4[17057] = 32'b11111111111111111110101110011011;
assign LUT_4[17058] = 32'b00000000000000000100111101000111;
assign LUT_4[17059] = 32'b11111111111111111110001000111111;
assign LUT_4[17060] = 32'b00000000000000000010100010111111;
assign LUT_4[17061] = 32'b11111111111111111011101110110111;
assign LUT_4[17062] = 32'b00000000000000000001111101100011;
assign LUT_4[17063] = 32'b11111111111111111011001001011011;
assign LUT_4[17064] = 32'b11111111111111111110101110111000;
assign LUT_4[17065] = 32'b11111111111111110111111010110000;
assign LUT_4[17066] = 32'b11111111111111111110001001011100;
assign LUT_4[17067] = 32'b11111111111111110111010101010100;
assign LUT_4[17068] = 32'b11111111111111111011101111010100;
assign LUT_4[17069] = 32'b11111111111111110100111011001100;
assign LUT_4[17070] = 32'b11111111111111111011001001111000;
assign LUT_4[17071] = 32'b11111111111111110100010101110000;
assign LUT_4[17072] = 32'b00000000000000000011010100010001;
assign LUT_4[17073] = 32'b11111111111111111100100000001001;
assign LUT_4[17074] = 32'b00000000000000000010101110110101;
assign LUT_4[17075] = 32'b11111111111111111011111010101101;
assign LUT_4[17076] = 32'b00000000000000000000010100101101;
assign LUT_4[17077] = 32'b11111111111111111001100000100101;
assign LUT_4[17078] = 32'b11111111111111111111101111010001;
assign LUT_4[17079] = 32'b11111111111111111000111011001001;
assign LUT_4[17080] = 32'b11111111111111111100100000100110;
assign LUT_4[17081] = 32'b11111111111111110101101100011110;
assign LUT_4[17082] = 32'b11111111111111111011111011001010;
assign LUT_4[17083] = 32'b11111111111111110101000111000010;
assign LUT_4[17084] = 32'b11111111111111111001100001000010;
assign LUT_4[17085] = 32'b11111111111111110010101100111010;
assign LUT_4[17086] = 32'b11111111111111111000111011100110;
assign LUT_4[17087] = 32'b11111111111111110010000111011110;
assign LUT_4[17088] = 32'b00000000000000001000011110110000;
assign LUT_4[17089] = 32'b00000000000000000001101010101000;
assign LUT_4[17090] = 32'b00000000000000000111111001010100;
assign LUT_4[17091] = 32'b00000000000000000001000101001100;
assign LUT_4[17092] = 32'b00000000000000000101011111001100;
assign LUT_4[17093] = 32'b11111111111111111110101011000100;
assign LUT_4[17094] = 32'b00000000000000000100111001110000;
assign LUT_4[17095] = 32'b11111111111111111110000101101000;
assign LUT_4[17096] = 32'b00000000000000000001101011000101;
assign LUT_4[17097] = 32'b11111111111111111010110110111101;
assign LUT_4[17098] = 32'b00000000000000000001000101101001;
assign LUT_4[17099] = 32'b11111111111111111010010001100001;
assign LUT_4[17100] = 32'b11111111111111111110101011100001;
assign LUT_4[17101] = 32'b11111111111111110111110111011001;
assign LUT_4[17102] = 32'b11111111111111111110000110000101;
assign LUT_4[17103] = 32'b11111111111111110111010001111101;
assign LUT_4[17104] = 32'b00000000000000000110010000011110;
assign LUT_4[17105] = 32'b11111111111111111111011100010110;
assign LUT_4[17106] = 32'b00000000000000000101101011000010;
assign LUT_4[17107] = 32'b11111111111111111110110110111010;
assign LUT_4[17108] = 32'b00000000000000000011010000111010;
assign LUT_4[17109] = 32'b11111111111111111100011100110010;
assign LUT_4[17110] = 32'b00000000000000000010101011011110;
assign LUT_4[17111] = 32'b11111111111111111011110111010110;
assign LUT_4[17112] = 32'b11111111111111111111011100110011;
assign LUT_4[17113] = 32'b11111111111111111000101000101011;
assign LUT_4[17114] = 32'b11111111111111111110110111010111;
assign LUT_4[17115] = 32'b11111111111111111000000011001111;
assign LUT_4[17116] = 32'b11111111111111111100011101001111;
assign LUT_4[17117] = 32'b11111111111111110101101001000111;
assign LUT_4[17118] = 32'b11111111111111111011110111110011;
assign LUT_4[17119] = 32'b11111111111111110101000011101011;
assign LUT_4[17120] = 32'b00000000000000000110111001110111;
assign LUT_4[17121] = 32'b00000000000000000000000101101111;
assign LUT_4[17122] = 32'b00000000000000000110010100011011;
assign LUT_4[17123] = 32'b11111111111111111111100000010011;
assign LUT_4[17124] = 32'b00000000000000000011111010010011;
assign LUT_4[17125] = 32'b11111111111111111101000110001011;
assign LUT_4[17126] = 32'b00000000000000000011010100110111;
assign LUT_4[17127] = 32'b11111111111111111100100000101111;
assign LUT_4[17128] = 32'b00000000000000000000000110001100;
assign LUT_4[17129] = 32'b11111111111111111001010010000100;
assign LUT_4[17130] = 32'b11111111111111111111100000110000;
assign LUT_4[17131] = 32'b11111111111111111000101100101000;
assign LUT_4[17132] = 32'b11111111111111111101000110101000;
assign LUT_4[17133] = 32'b11111111111111110110010010100000;
assign LUT_4[17134] = 32'b11111111111111111100100001001100;
assign LUT_4[17135] = 32'b11111111111111110101101101000100;
assign LUT_4[17136] = 32'b00000000000000000100101011100101;
assign LUT_4[17137] = 32'b11111111111111111101110111011101;
assign LUT_4[17138] = 32'b00000000000000000100000110001001;
assign LUT_4[17139] = 32'b11111111111111111101010010000001;
assign LUT_4[17140] = 32'b00000000000000000001101100000001;
assign LUT_4[17141] = 32'b11111111111111111010110111111001;
assign LUT_4[17142] = 32'b00000000000000000001000110100101;
assign LUT_4[17143] = 32'b11111111111111111010010010011101;
assign LUT_4[17144] = 32'b11111111111111111101110111111010;
assign LUT_4[17145] = 32'b11111111111111110111000011110010;
assign LUT_4[17146] = 32'b11111111111111111101010010011110;
assign LUT_4[17147] = 32'b11111111111111110110011110010110;
assign LUT_4[17148] = 32'b11111111111111111010111000010110;
assign LUT_4[17149] = 32'b11111111111111110100000100001110;
assign LUT_4[17150] = 32'b11111111111111111010010010111010;
assign LUT_4[17151] = 32'b11111111111111110011011110110010;
assign LUT_4[17152] = 32'b00000000000000001001011100110111;
assign LUT_4[17153] = 32'b00000000000000000010101000101111;
assign LUT_4[17154] = 32'b00000000000000001000110111011011;
assign LUT_4[17155] = 32'b00000000000000000010000011010011;
assign LUT_4[17156] = 32'b00000000000000000110011101010011;
assign LUT_4[17157] = 32'b11111111111111111111101001001011;
assign LUT_4[17158] = 32'b00000000000000000101110111110111;
assign LUT_4[17159] = 32'b11111111111111111111000011101111;
assign LUT_4[17160] = 32'b00000000000000000010101001001100;
assign LUT_4[17161] = 32'b11111111111111111011110101000100;
assign LUT_4[17162] = 32'b00000000000000000010000011110000;
assign LUT_4[17163] = 32'b11111111111111111011001111101000;
assign LUT_4[17164] = 32'b11111111111111111111101001101000;
assign LUT_4[17165] = 32'b11111111111111111000110101100000;
assign LUT_4[17166] = 32'b11111111111111111111000100001100;
assign LUT_4[17167] = 32'b11111111111111111000010000000100;
assign LUT_4[17168] = 32'b00000000000000000111001110100101;
assign LUT_4[17169] = 32'b00000000000000000000011010011101;
assign LUT_4[17170] = 32'b00000000000000000110101001001001;
assign LUT_4[17171] = 32'b11111111111111111111110101000001;
assign LUT_4[17172] = 32'b00000000000000000100001111000001;
assign LUT_4[17173] = 32'b11111111111111111101011010111001;
assign LUT_4[17174] = 32'b00000000000000000011101001100101;
assign LUT_4[17175] = 32'b11111111111111111100110101011101;
assign LUT_4[17176] = 32'b00000000000000000000011010111010;
assign LUT_4[17177] = 32'b11111111111111111001100110110010;
assign LUT_4[17178] = 32'b11111111111111111111110101011110;
assign LUT_4[17179] = 32'b11111111111111111001000001010110;
assign LUT_4[17180] = 32'b11111111111111111101011011010110;
assign LUT_4[17181] = 32'b11111111111111110110100111001110;
assign LUT_4[17182] = 32'b11111111111111111100110101111010;
assign LUT_4[17183] = 32'b11111111111111110110000001110010;
assign LUT_4[17184] = 32'b00000000000000000111110111111110;
assign LUT_4[17185] = 32'b00000000000000000001000011110110;
assign LUT_4[17186] = 32'b00000000000000000111010010100010;
assign LUT_4[17187] = 32'b00000000000000000000011110011010;
assign LUT_4[17188] = 32'b00000000000000000100111000011010;
assign LUT_4[17189] = 32'b11111111111111111110000100010010;
assign LUT_4[17190] = 32'b00000000000000000100010010111110;
assign LUT_4[17191] = 32'b11111111111111111101011110110110;
assign LUT_4[17192] = 32'b00000000000000000001000100010011;
assign LUT_4[17193] = 32'b11111111111111111010010000001011;
assign LUT_4[17194] = 32'b00000000000000000000011110110111;
assign LUT_4[17195] = 32'b11111111111111111001101010101111;
assign LUT_4[17196] = 32'b11111111111111111110000100101111;
assign LUT_4[17197] = 32'b11111111111111110111010000100111;
assign LUT_4[17198] = 32'b11111111111111111101011111010011;
assign LUT_4[17199] = 32'b11111111111111110110101011001011;
assign LUT_4[17200] = 32'b00000000000000000101101001101100;
assign LUT_4[17201] = 32'b11111111111111111110110101100100;
assign LUT_4[17202] = 32'b00000000000000000101000100010000;
assign LUT_4[17203] = 32'b11111111111111111110010000001000;
assign LUT_4[17204] = 32'b00000000000000000010101010001000;
assign LUT_4[17205] = 32'b11111111111111111011110110000000;
assign LUT_4[17206] = 32'b00000000000000000010000100101100;
assign LUT_4[17207] = 32'b11111111111111111011010000100100;
assign LUT_4[17208] = 32'b11111111111111111110110110000001;
assign LUT_4[17209] = 32'b11111111111111111000000001111001;
assign LUT_4[17210] = 32'b11111111111111111110010000100101;
assign LUT_4[17211] = 32'b11111111111111110111011100011101;
assign LUT_4[17212] = 32'b11111111111111111011110110011101;
assign LUT_4[17213] = 32'b11111111111111110101000010010101;
assign LUT_4[17214] = 32'b11111111111111111011010001000001;
assign LUT_4[17215] = 32'b11111111111111110100011100111001;
assign LUT_4[17216] = 32'b00000000000000001010110100001011;
assign LUT_4[17217] = 32'b00000000000000000100000000000011;
assign LUT_4[17218] = 32'b00000000000000001010001110101111;
assign LUT_4[17219] = 32'b00000000000000000011011010100111;
assign LUT_4[17220] = 32'b00000000000000000111110100100111;
assign LUT_4[17221] = 32'b00000000000000000001000000011111;
assign LUT_4[17222] = 32'b00000000000000000111001111001011;
assign LUT_4[17223] = 32'b00000000000000000000011011000011;
assign LUT_4[17224] = 32'b00000000000000000100000000100000;
assign LUT_4[17225] = 32'b11111111111111111101001100011000;
assign LUT_4[17226] = 32'b00000000000000000011011011000100;
assign LUT_4[17227] = 32'b11111111111111111100100110111100;
assign LUT_4[17228] = 32'b00000000000000000001000000111100;
assign LUT_4[17229] = 32'b11111111111111111010001100110100;
assign LUT_4[17230] = 32'b00000000000000000000011011100000;
assign LUT_4[17231] = 32'b11111111111111111001100111011000;
assign LUT_4[17232] = 32'b00000000000000001000100101111001;
assign LUT_4[17233] = 32'b00000000000000000001110001110001;
assign LUT_4[17234] = 32'b00000000000000001000000000011101;
assign LUT_4[17235] = 32'b00000000000000000001001100010101;
assign LUT_4[17236] = 32'b00000000000000000101100110010101;
assign LUT_4[17237] = 32'b11111111111111111110110010001101;
assign LUT_4[17238] = 32'b00000000000000000101000000111001;
assign LUT_4[17239] = 32'b11111111111111111110001100110001;
assign LUT_4[17240] = 32'b00000000000000000001110010001110;
assign LUT_4[17241] = 32'b11111111111111111010111110000110;
assign LUT_4[17242] = 32'b00000000000000000001001100110010;
assign LUT_4[17243] = 32'b11111111111111111010011000101010;
assign LUT_4[17244] = 32'b11111111111111111110110010101010;
assign LUT_4[17245] = 32'b11111111111111110111111110100010;
assign LUT_4[17246] = 32'b11111111111111111110001101001110;
assign LUT_4[17247] = 32'b11111111111111110111011001000110;
assign LUT_4[17248] = 32'b00000000000000001001001111010010;
assign LUT_4[17249] = 32'b00000000000000000010011011001010;
assign LUT_4[17250] = 32'b00000000000000001000101001110110;
assign LUT_4[17251] = 32'b00000000000000000001110101101110;
assign LUT_4[17252] = 32'b00000000000000000110001111101110;
assign LUT_4[17253] = 32'b11111111111111111111011011100110;
assign LUT_4[17254] = 32'b00000000000000000101101010010010;
assign LUT_4[17255] = 32'b11111111111111111110110110001010;
assign LUT_4[17256] = 32'b00000000000000000010011011100111;
assign LUT_4[17257] = 32'b11111111111111111011100111011111;
assign LUT_4[17258] = 32'b00000000000000000001110110001011;
assign LUT_4[17259] = 32'b11111111111111111011000010000011;
assign LUT_4[17260] = 32'b11111111111111111111011100000011;
assign LUT_4[17261] = 32'b11111111111111111000100111111011;
assign LUT_4[17262] = 32'b11111111111111111110110110100111;
assign LUT_4[17263] = 32'b11111111111111111000000010011111;
assign LUT_4[17264] = 32'b00000000000000000111000001000000;
assign LUT_4[17265] = 32'b00000000000000000000001100111000;
assign LUT_4[17266] = 32'b00000000000000000110011011100100;
assign LUT_4[17267] = 32'b11111111111111111111100111011100;
assign LUT_4[17268] = 32'b00000000000000000100000001011100;
assign LUT_4[17269] = 32'b11111111111111111101001101010100;
assign LUT_4[17270] = 32'b00000000000000000011011100000000;
assign LUT_4[17271] = 32'b11111111111111111100100111111000;
assign LUT_4[17272] = 32'b00000000000000000000001101010101;
assign LUT_4[17273] = 32'b11111111111111111001011001001101;
assign LUT_4[17274] = 32'b11111111111111111111100111111001;
assign LUT_4[17275] = 32'b11111111111111111000110011110001;
assign LUT_4[17276] = 32'b11111111111111111101001101110001;
assign LUT_4[17277] = 32'b11111111111111110110011001101001;
assign LUT_4[17278] = 32'b11111111111111111100101000010101;
assign LUT_4[17279] = 32'b11111111111111110101110100001101;
assign LUT_4[17280] = 32'b00000000000000001100000010111111;
assign LUT_4[17281] = 32'b00000000000000000101001110110111;
assign LUT_4[17282] = 32'b00000000000000001011011101100011;
assign LUT_4[17283] = 32'b00000000000000000100101001011011;
assign LUT_4[17284] = 32'b00000000000000001001000011011011;
assign LUT_4[17285] = 32'b00000000000000000010001111010011;
assign LUT_4[17286] = 32'b00000000000000001000011101111111;
assign LUT_4[17287] = 32'b00000000000000000001101001110111;
assign LUT_4[17288] = 32'b00000000000000000101001111010100;
assign LUT_4[17289] = 32'b11111111111111111110011011001100;
assign LUT_4[17290] = 32'b00000000000000000100101001111000;
assign LUT_4[17291] = 32'b11111111111111111101110101110000;
assign LUT_4[17292] = 32'b00000000000000000010001111110000;
assign LUT_4[17293] = 32'b11111111111111111011011011101000;
assign LUT_4[17294] = 32'b00000000000000000001101010010100;
assign LUT_4[17295] = 32'b11111111111111111010110110001100;
assign LUT_4[17296] = 32'b00000000000000001001110100101101;
assign LUT_4[17297] = 32'b00000000000000000011000000100101;
assign LUT_4[17298] = 32'b00000000000000001001001111010001;
assign LUT_4[17299] = 32'b00000000000000000010011011001001;
assign LUT_4[17300] = 32'b00000000000000000110110101001001;
assign LUT_4[17301] = 32'b00000000000000000000000001000001;
assign LUT_4[17302] = 32'b00000000000000000110001111101101;
assign LUT_4[17303] = 32'b11111111111111111111011011100101;
assign LUT_4[17304] = 32'b00000000000000000011000001000010;
assign LUT_4[17305] = 32'b11111111111111111100001100111010;
assign LUT_4[17306] = 32'b00000000000000000010011011100110;
assign LUT_4[17307] = 32'b11111111111111111011100111011110;
assign LUT_4[17308] = 32'b00000000000000000000000001011110;
assign LUT_4[17309] = 32'b11111111111111111001001101010110;
assign LUT_4[17310] = 32'b11111111111111111111011100000010;
assign LUT_4[17311] = 32'b11111111111111111000100111111010;
assign LUT_4[17312] = 32'b00000000000000001010011110000110;
assign LUT_4[17313] = 32'b00000000000000000011101001111110;
assign LUT_4[17314] = 32'b00000000000000001001111000101010;
assign LUT_4[17315] = 32'b00000000000000000011000100100010;
assign LUT_4[17316] = 32'b00000000000000000111011110100010;
assign LUT_4[17317] = 32'b00000000000000000000101010011010;
assign LUT_4[17318] = 32'b00000000000000000110111001000110;
assign LUT_4[17319] = 32'b00000000000000000000000100111110;
assign LUT_4[17320] = 32'b00000000000000000011101010011011;
assign LUT_4[17321] = 32'b11111111111111111100110110010011;
assign LUT_4[17322] = 32'b00000000000000000011000100111111;
assign LUT_4[17323] = 32'b11111111111111111100010000110111;
assign LUT_4[17324] = 32'b00000000000000000000101010110111;
assign LUT_4[17325] = 32'b11111111111111111001110110101111;
assign LUT_4[17326] = 32'b00000000000000000000000101011011;
assign LUT_4[17327] = 32'b11111111111111111001010001010011;
assign LUT_4[17328] = 32'b00000000000000001000001111110100;
assign LUT_4[17329] = 32'b00000000000000000001011011101100;
assign LUT_4[17330] = 32'b00000000000000000111101010011000;
assign LUT_4[17331] = 32'b00000000000000000000110110010000;
assign LUT_4[17332] = 32'b00000000000000000101010000010000;
assign LUT_4[17333] = 32'b11111111111111111110011100001000;
assign LUT_4[17334] = 32'b00000000000000000100101010110100;
assign LUT_4[17335] = 32'b11111111111111111101110110101100;
assign LUT_4[17336] = 32'b00000000000000000001011100001001;
assign LUT_4[17337] = 32'b11111111111111111010101000000001;
assign LUT_4[17338] = 32'b00000000000000000000110110101101;
assign LUT_4[17339] = 32'b11111111111111111010000010100101;
assign LUT_4[17340] = 32'b11111111111111111110011100100101;
assign LUT_4[17341] = 32'b11111111111111110111101000011101;
assign LUT_4[17342] = 32'b11111111111111111101110111001001;
assign LUT_4[17343] = 32'b11111111111111110111000011000001;
assign LUT_4[17344] = 32'b00000000000000001101011010010011;
assign LUT_4[17345] = 32'b00000000000000000110100110001011;
assign LUT_4[17346] = 32'b00000000000000001100110100110111;
assign LUT_4[17347] = 32'b00000000000000000110000000101111;
assign LUT_4[17348] = 32'b00000000000000001010011010101111;
assign LUT_4[17349] = 32'b00000000000000000011100110100111;
assign LUT_4[17350] = 32'b00000000000000001001110101010011;
assign LUT_4[17351] = 32'b00000000000000000011000001001011;
assign LUT_4[17352] = 32'b00000000000000000110100110101000;
assign LUT_4[17353] = 32'b11111111111111111111110010100000;
assign LUT_4[17354] = 32'b00000000000000000110000001001100;
assign LUT_4[17355] = 32'b11111111111111111111001101000100;
assign LUT_4[17356] = 32'b00000000000000000011100111000100;
assign LUT_4[17357] = 32'b11111111111111111100110010111100;
assign LUT_4[17358] = 32'b00000000000000000011000001101000;
assign LUT_4[17359] = 32'b11111111111111111100001101100000;
assign LUT_4[17360] = 32'b00000000000000001011001100000001;
assign LUT_4[17361] = 32'b00000000000000000100010111111001;
assign LUT_4[17362] = 32'b00000000000000001010100110100101;
assign LUT_4[17363] = 32'b00000000000000000011110010011101;
assign LUT_4[17364] = 32'b00000000000000001000001100011101;
assign LUT_4[17365] = 32'b00000000000000000001011000010101;
assign LUT_4[17366] = 32'b00000000000000000111100111000001;
assign LUT_4[17367] = 32'b00000000000000000000110010111001;
assign LUT_4[17368] = 32'b00000000000000000100011000010110;
assign LUT_4[17369] = 32'b11111111111111111101100100001110;
assign LUT_4[17370] = 32'b00000000000000000011110010111010;
assign LUT_4[17371] = 32'b11111111111111111100111110110010;
assign LUT_4[17372] = 32'b00000000000000000001011000110010;
assign LUT_4[17373] = 32'b11111111111111111010100100101010;
assign LUT_4[17374] = 32'b00000000000000000000110011010110;
assign LUT_4[17375] = 32'b11111111111111111001111111001110;
assign LUT_4[17376] = 32'b00000000000000001011110101011010;
assign LUT_4[17377] = 32'b00000000000000000101000001010010;
assign LUT_4[17378] = 32'b00000000000000001011001111111110;
assign LUT_4[17379] = 32'b00000000000000000100011011110110;
assign LUT_4[17380] = 32'b00000000000000001000110101110110;
assign LUT_4[17381] = 32'b00000000000000000010000001101110;
assign LUT_4[17382] = 32'b00000000000000001000010000011010;
assign LUT_4[17383] = 32'b00000000000000000001011100010010;
assign LUT_4[17384] = 32'b00000000000000000101000001101111;
assign LUT_4[17385] = 32'b11111111111111111110001101100111;
assign LUT_4[17386] = 32'b00000000000000000100011100010011;
assign LUT_4[17387] = 32'b11111111111111111101101000001011;
assign LUT_4[17388] = 32'b00000000000000000010000010001011;
assign LUT_4[17389] = 32'b11111111111111111011001110000011;
assign LUT_4[17390] = 32'b00000000000000000001011100101111;
assign LUT_4[17391] = 32'b11111111111111111010101000100111;
assign LUT_4[17392] = 32'b00000000000000001001100111001000;
assign LUT_4[17393] = 32'b00000000000000000010110011000000;
assign LUT_4[17394] = 32'b00000000000000001001000001101100;
assign LUT_4[17395] = 32'b00000000000000000010001101100100;
assign LUT_4[17396] = 32'b00000000000000000110100111100100;
assign LUT_4[17397] = 32'b11111111111111111111110011011100;
assign LUT_4[17398] = 32'b00000000000000000110000010001000;
assign LUT_4[17399] = 32'b11111111111111111111001110000000;
assign LUT_4[17400] = 32'b00000000000000000010110011011101;
assign LUT_4[17401] = 32'b11111111111111111011111111010101;
assign LUT_4[17402] = 32'b00000000000000000010001110000001;
assign LUT_4[17403] = 32'b11111111111111111011011001111001;
assign LUT_4[17404] = 32'b11111111111111111111110011111001;
assign LUT_4[17405] = 32'b11111111111111111000111111110001;
assign LUT_4[17406] = 32'b11111111111111111111001110011101;
assign LUT_4[17407] = 32'b11111111111111111000011010010101;
assign LUT_4[17408] = 32'b00000000000000000111000111101011;
assign LUT_4[17409] = 32'b00000000000000000000010011100011;
assign LUT_4[17410] = 32'b00000000000000000110100010001111;
assign LUT_4[17411] = 32'b11111111111111111111101110000111;
assign LUT_4[17412] = 32'b00000000000000000100001000000111;
assign LUT_4[17413] = 32'b11111111111111111101010011111111;
assign LUT_4[17414] = 32'b00000000000000000011100010101011;
assign LUT_4[17415] = 32'b11111111111111111100101110100011;
assign LUT_4[17416] = 32'b00000000000000000000010100000000;
assign LUT_4[17417] = 32'b11111111111111111001011111111000;
assign LUT_4[17418] = 32'b11111111111111111111101110100100;
assign LUT_4[17419] = 32'b11111111111111111000111010011100;
assign LUT_4[17420] = 32'b11111111111111111101010100011100;
assign LUT_4[17421] = 32'b11111111111111110110100000010100;
assign LUT_4[17422] = 32'b11111111111111111100101111000000;
assign LUT_4[17423] = 32'b11111111111111110101111010111000;
assign LUT_4[17424] = 32'b00000000000000000100111001011001;
assign LUT_4[17425] = 32'b11111111111111111110000101010001;
assign LUT_4[17426] = 32'b00000000000000000100010011111101;
assign LUT_4[17427] = 32'b11111111111111111101011111110101;
assign LUT_4[17428] = 32'b00000000000000000001111001110101;
assign LUT_4[17429] = 32'b11111111111111111011000101101101;
assign LUT_4[17430] = 32'b00000000000000000001010100011001;
assign LUT_4[17431] = 32'b11111111111111111010100000010001;
assign LUT_4[17432] = 32'b11111111111111111110000101101110;
assign LUT_4[17433] = 32'b11111111111111110111010001100110;
assign LUT_4[17434] = 32'b11111111111111111101100000010010;
assign LUT_4[17435] = 32'b11111111111111110110101100001010;
assign LUT_4[17436] = 32'b11111111111111111011000110001010;
assign LUT_4[17437] = 32'b11111111111111110100010010000010;
assign LUT_4[17438] = 32'b11111111111111111010100000101110;
assign LUT_4[17439] = 32'b11111111111111110011101100100110;
assign LUT_4[17440] = 32'b00000000000000000101100010110010;
assign LUT_4[17441] = 32'b11111111111111111110101110101010;
assign LUT_4[17442] = 32'b00000000000000000100111101010110;
assign LUT_4[17443] = 32'b11111111111111111110001001001110;
assign LUT_4[17444] = 32'b00000000000000000010100011001110;
assign LUT_4[17445] = 32'b11111111111111111011101111000110;
assign LUT_4[17446] = 32'b00000000000000000001111101110010;
assign LUT_4[17447] = 32'b11111111111111111011001001101010;
assign LUT_4[17448] = 32'b11111111111111111110101111000111;
assign LUT_4[17449] = 32'b11111111111111110111111010111111;
assign LUT_4[17450] = 32'b11111111111111111110001001101011;
assign LUT_4[17451] = 32'b11111111111111110111010101100011;
assign LUT_4[17452] = 32'b11111111111111111011101111100011;
assign LUT_4[17453] = 32'b11111111111111110100111011011011;
assign LUT_4[17454] = 32'b11111111111111111011001010000111;
assign LUT_4[17455] = 32'b11111111111111110100010101111111;
assign LUT_4[17456] = 32'b00000000000000000011010100100000;
assign LUT_4[17457] = 32'b11111111111111111100100000011000;
assign LUT_4[17458] = 32'b00000000000000000010101111000100;
assign LUT_4[17459] = 32'b11111111111111111011111010111100;
assign LUT_4[17460] = 32'b00000000000000000000010100111100;
assign LUT_4[17461] = 32'b11111111111111111001100000110100;
assign LUT_4[17462] = 32'b11111111111111111111101111100000;
assign LUT_4[17463] = 32'b11111111111111111000111011011000;
assign LUT_4[17464] = 32'b11111111111111111100100000110101;
assign LUT_4[17465] = 32'b11111111111111110101101100101101;
assign LUT_4[17466] = 32'b11111111111111111011111011011001;
assign LUT_4[17467] = 32'b11111111111111110101000111010001;
assign LUT_4[17468] = 32'b11111111111111111001100001010001;
assign LUT_4[17469] = 32'b11111111111111110010101101001001;
assign LUT_4[17470] = 32'b11111111111111111000111011110101;
assign LUT_4[17471] = 32'b11111111111111110010000111101101;
assign LUT_4[17472] = 32'b00000000000000001000011110111111;
assign LUT_4[17473] = 32'b00000000000000000001101010110111;
assign LUT_4[17474] = 32'b00000000000000000111111001100011;
assign LUT_4[17475] = 32'b00000000000000000001000101011011;
assign LUT_4[17476] = 32'b00000000000000000101011111011011;
assign LUT_4[17477] = 32'b11111111111111111110101011010011;
assign LUT_4[17478] = 32'b00000000000000000100111001111111;
assign LUT_4[17479] = 32'b11111111111111111110000101110111;
assign LUT_4[17480] = 32'b00000000000000000001101011010100;
assign LUT_4[17481] = 32'b11111111111111111010110111001100;
assign LUT_4[17482] = 32'b00000000000000000001000101111000;
assign LUT_4[17483] = 32'b11111111111111111010010001110000;
assign LUT_4[17484] = 32'b11111111111111111110101011110000;
assign LUT_4[17485] = 32'b11111111111111110111110111101000;
assign LUT_4[17486] = 32'b11111111111111111110000110010100;
assign LUT_4[17487] = 32'b11111111111111110111010010001100;
assign LUT_4[17488] = 32'b00000000000000000110010000101101;
assign LUT_4[17489] = 32'b11111111111111111111011100100101;
assign LUT_4[17490] = 32'b00000000000000000101101011010001;
assign LUT_4[17491] = 32'b11111111111111111110110111001001;
assign LUT_4[17492] = 32'b00000000000000000011010001001001;
assign LUT_4[17493] = 32'b11111111111111111100011101000001;
assign LUT_4[17494] = 32'b00000000000000000010101011101101;
assign LUT_4[17495] = 32'b11111111111111111011110111100101;
assign LUT_4[17496] = 32'b11111111111111111111011101000010;
assign LUT_4[17497] = 32'b11111111111111111000101000111010;
assign LUT_4[17498] = 32'b11111111111111111110110111100110;
assign LUT_4[17499] = 32'b11111111111111111000000011011110;
assign LUT_4[17500] = 32'b11111111111111111100011101011110;
assign LUT_4[17501] = 32'b11111111111111110101101001010110;
assign LUT_4[17502] = 32'b11111111111111111011111000000010;
assign LUT_4[17503] = 32'b11111111111111110101000011111010;
assign LUT_4[17504] = 32'b00000000000000000110111010000110;
assign LUT_4[17505] = 32'b00000000000000000000000101111110;
assign LUT_4[17506] = 32'b00000000000000000110010100101010;
assign LUT_4[17507] = 32'b11111111111111111111100000100010;
assign LUT_4[17508] = 32'b00000000000000000011111010100010;
assign LUT_4[17509] = 32'b11111111111111111101000110011010;
assign LUT_4[17510] = 32'b00000000000000000011010101000110;
assign LUT_4[17511] = 32'b11111111111111111100100000111110;
assign LUT_4[17512] = 32'b00000000000000000000000110011011;
assign LUT_4[17513] = 32'b11111111111111111001010010010011;
assign LUT_4[17514] = 32'b11111111111111111111100000111111;
assign LUT_4[17515] = 32'b11111111111111111000101100110111;
assign LUT_4[17516] = 32'b11111111111111111101000110110111;
assign LUT_4[17517] = 32'b11111111111111110110010010101111;
assign LUT_4[17518] = 32'b11111111111111111100100001011011;
assign LUT_4[17519] = 32'b11111111111111110101101101010011;
assign LUT_4[17520] = 32'b00000000000000000100101011110100;
assign LUT_4[17521] = 32'b11111111111111111101110111101100;
assign LUT_4[17522] = 32'b00000000000000000100000110011000;
assign LUT_4[17523] = 32'b11111111111111111101010010010000;
assign LUT_4[17524] = 32'b00000000000000000001101100010000;
assign LUT_4[17525] = 32'b11111111111111111010111000001000;
assign LUT_4[17526] = 32'b00000000000000000001000110110100;
assign LUT_4[17527] = 32'b11111111111111111010010010101100;
assign LUT_4[17528] = 32'b11111111111111111101111000001001;
assign LUT_4[17529] = 32'b11111111111111110111000100000001;
assign LUT_4[17530] = 32'b11111111111111111101010010101101;
assign LUT_4[17531] = 32'b11111111111111110110011110100101;
assign LUT_4[17532] = 32'b11111111111111111010111000100101;
assign LUT_4[17533] = 32'b11111111111111110100000100011101;
assign LUT_4[17534] = 32'b11111111111111111010010011001001;
assign LUT_4[17535] = 32'b11111111111111110011011111000001;
assign LUT_4[17536] = 32'b00000000000000001001101101110011;
assign LUT_4[17537] = 32'b00000000000000000010111001101011;
assign LUT_4[17538] = 32'b00000000000000001001001000010111;
assign LUT_4[17539] = 32'b00000000000000000010010100001111;
assign LUT_4[17540] = 32'b00000000000000000110101110001111;
assign LUT_4[17541] = 32'b11111111111111111111111010000111;
assign LUT_4[17542] = 32'b00000000000000000110001000110011;
assign LUT_4[17543] = 32'b11111111111111111111010100101011;
assign LUT_4[17544] = 32'b00000000000000000010111010001000;
assign LUT_4[17545] = 32'b11111111111111111100000110000000;
assign LUT_4[17546] = 32'b00000000000000000010010100101100;
assign LUT_4[17547] = 32'b11111111111111111011100000100100;
assign LUT_4[17548] = 32'b11111111111111111111111010100100;
assign LUT_4[17549] = 32'b11111111111111111001000110011100;
assign LUT_4[17550] = 32'b11111111111111111111010101001000;
assign LUT_4[17551] = 32'b11111111111111111000100001000000;
assign LUT_4[17552] = 32'b00000000000000000111011111100001;
assign LUT_4[17553] = 32'b00000000000000000000101011011001;
assign LUT_4[17554] = 32'b00000000000000000110111010000101;
assign LUT_4[17555] = 32'b00000000000000000000000101111101;
assign LUT_4[17556] = 32'b00000000000000000100011111111101;
assign LUT_4[17557] = 32'b11111111111111111101101011110101;
assign LUT_4[17558] = 32'b00000000000000000011111010100001;
assign LUT_4[17559] = 32'b11111111111111111101000110011001;
assign LUT_4[17560] = 32'b00000000000000000000101011110110;
assign LUT_4[17561] = 32'b11111111111111111001110111101110;
assign LUT_4[17562] = 32'b00000000000000000000000110011010;
assign LUT_4[17563] = 32'b11111111111111111001010010010010;
assign LUT_4[17564] = 32'b11111111111111111101101100010010;
assign LUT_4[17565] = 32'b11111111111111110110111000001010;
assign LUT_4[17566] = 32'b11111111111111111101000110110110;
assign LUT_4[17567] = 32'b11111111111111110110010010101110;
assign LUT_4[17568] = 32'b00000000000000001000001000111010;
assign LUT_4[17569] = 32'b00000000000000000001010100110010;
assign LUT_4[17570] = 32'b00000000000000000111100011011110;
assign LUT_4[17571] = 32'b00000000000000000000101111010110;
assign LUT_4[17572] = 32'b00000000000000000101001001010110;
assign LUT_4[17573] = 32'b11111111111111111110010101001110;
assign LUT_4[17574] = 32'b00000000000000000100100011111010;
assign LUT_4[17575] = 32'b11111111111111111101101111110010;
assign LUT_4[17576] = 32'b00000000000000000001010101001111;
assign LUT_4[17577] = 32'b11111111111111111010100001000111;
assign LUT_4[17578] = 32'b00000000000000000000101111110011;
assign LUT_4[17579] = 32'b11111111111111111001111011101011;
assign LUT_4[17580] = 32'b11111111111111111110010101101011;
assign LUT_4[17581] = 32'b11111111111111110111100001100011;
assign LUT_4[17582] = 32'b11111111111111111101110000001111;
assign LUT_4[17583] = 32'b11111111111111110110111100000111;
assign LUT_4[17584] = 32'b00000000000000000101111010101000;
assign LUT_4[17585] = 32'b11111111111111111111000110100000;
assign LUT_4[17586] = 32'b00000000000000000101010101001100;
assign LUT_4[17587] = 32'b11111111111111111110100001000100;
assign LUT_4[17588] = 32'b00000000000000000010111011000100;
assign LUT_4[17589] = 32'b11111111111111111100000110111100;
assign LUT_4[17590] = 32'b00000000000000000010010101101000;
assign LUT_4[17591] = 32'b11111111111111111011100001100000;
assign LUT_4[17592] = 32'b11111111111111111111000110111101;
assign LUT_4[17593] = 32'b11111111111111111000010010110101;
assign LUT_4[17594] = 32'b11111111111111111110100001100001;
assign LUT_4[17595] = 32'b11111111111111110111101101011001;
assign LUT_4[17596] = 32'b11111111111111111100000111011001;
assign LUT_4[17597] = 32'b11111111111111110101010011010001;
assign LUT_4[17598] = 32'b11111111111111111011100001111101;
assign LUT_4[17599] = 32'b11111111111111110100101101110101;
assign LUT_4[17600] = 32'b00000000000000001011000101000111;
assign LUT_4[17601] = 32'b00000000000000000100010000111111;
assign LUT_4[17602] = 32'b00000000000000001010011111101011;
assign LUT_4[17603] = 32'b00000000000000000011101011100011;
assign LUT_4[17604] = 32'b00000000000000001000000101100011;
assign LUT_4[17605] = 32'b00000000000000000001010001011011;
assign LUT_4[17606] = 32'b00000000000000000111100000000111;
assign LUT_4[17607] = 32'b00000000000000000000101011111111;
assign LUT_4[17608] = 32'b00000000000000000100010001011100;
assign LUT_4[17609] = 32'b11111111111111111101011101010100;
assign LUT_4[17610] = 32'b00000000000000000011101100000000;
assign LUT_4[17611] = 32'b11111111111111111100110111111000;
assign LUT_4[17612] = 32'b00000000000000000001010001111000;
assign LUT_4[17613] = 32'b11111111111111111010011101110000;
assign LUT_4[17614] = 32'b00000000000000000000101100011100;
assign LUT_4[17615] = 32'b11111111111111111001111000010100;
assign LUT_4[17616] = 32'b00000000000000001000110110110101;
assign LUT_4[17617] = 32'b00000000000000000010000010101101;
assign LUT_4[17618] = 32'b00000000000000001000010001011001;
assign LUT_4[17619] = 32'b00000000000000000001011101010001;
assign LUT_4[17620] = 32'b00000000000000000101110111010001;
assign LUT_4[17621] = 32'b11111111111111111111000011001001;
assign LUT_4[17622] = 32'b00000000000000000101010001110101;
assign LUT_4[17623] = 32'b11111111111111111110011101101101;
assign LUT_4[17624] = 32'b00000000000000000010000011001010;
assign LUT_4[17625] = 32'b11111111111111111011001111000010;
assign LUT_4[17626] = 32'b00000000000000000001011101101110;
assign LUT_4[17627] = 32'b11111111111111111010101001100110;
assign LUT_4[17628] = 32'b11111111111111111111000011100110;
assign LUT_4[17629] = 32'b11111111111111111000001111011110;
assign LUT_4[17630] = 32'b11111111111111111110011110001010;
assign LUT_4[17631] = 32'b11111111111111110111101010000010;
assign LUT_4[17632] = 32'b00000000000000001001100000001110;
assign LUT_4[17633] = 32'b00000000000000000010101100000110;
assign LUT_4[17634] = 32'b00000000000000001000111010110010;
assign LUT_4[17635] = 32'b00000000000000000010000110101010;
assign LUT_4[17636] = 32'b00000000000000000110100000101010;
assign LUT_4[17637] = 32'b11111111111111111111101100100010;
assign LUT_4[17638] = 32'b00000000000000000101111011001110;
assign LUT_4[17639] = 32'b11111111111111111111000111000110;
assign LUT_4[17640] = 32'b00000000000000000010101100100011;
assign LUT_4[17641] = 32'b11111111111111111011111000011011;
assign LUT_4[17642] = 32'b00000000000000000010000111000111;
assign LUT_4[17643] = 32'b11111111111111111011010010111111;
assign LUT_4[17644] = 32'b11111111111111111111101100111111;
assign LUT_4[17645] = 32'b11111111111111111000111000110111;
assign LUT_4[17646] = 32'b11111111111111111111000111100011;
assign LUT_4[17647] = 32'b11111111111111111000010011011011;
assign LUT_4[17648] = 32'b00000000000000000111010001111100;
assign LUT_4[17649] = 32'b00000000000000000000011101110100;
assign LUT_4[17650] = 32'b00000000000000000110101100100000;
assign LUT_4[17651] = 32'b11111111111111111111111000011000;
assign LUT_4[17652] = 32'b00000000000000000100010010011000;
assign LUT_4[17653] = 32'b11111111111111111101011110010000;
assign LUT_4[17654] = 32'b00000000000000000011101100111100;
assign LUT_4[17655] = 32'b11111111111111111100111000110100;
assign LUT_4[17656] = 32'b00000000000000000000011110010001;
assign LUT_4[17657] = 32'b11111111111111111001101010001001;
assign LUT_4[17658] = 32'b11111111111111111111111000110101;
assign LUT_4[17659] = 32'b11111111111111111001000100101101;
assign LUT_4[17660] = 32'b11111111111111111101011110101101;
assign LUT_4[17661] = 32'b11111111111111110110101010100101;
assign LUT_4[17662] = 32'b11111111111111111100111001010001;
assign LUT_4[17663] = 32'b11111111111111110110000101001001;
assign LUT_4[17664] = 32'b00000000000000001100000011001110;
assign LUT_4[17665] = 32'b00000000000000000101001111000110;
assign LUT_4[17666] = 32'b00000000000000001011011101110010;
assign LUT_4[17667] = 32'b00000000000000000100101001101010;
assign LUT_4[17668] = 32'b00000000000000001001000011101010;
assign LUT_4[17669] = 32'b00000000000000000010001111100010;
assign LUT_4[17670] = 32'b00000000000000001000011110001110;
assign LUT_4[17671] = 32'b00000000000000000001101010000110;
assign LUT_4[17672] = 32'b00000000000000000101001111100011;
assign LUT_4[17673] = 32'b11111111111111111110011011011011;
assign LUT_4[17674] = 32'b00000000000000000100101010000111;
assign LUT_4[17675] = 32'b11111111111111111101110101111111;
assign LUT_4[17676] = 32'b00000000000000000010001111111111;
assign LUT_4[17677] = 32'b11111111111111111011011011110111;
assign LUT_4[17678] = 32'b00000000000000000001101010100011;
assign LUT_4[17679] = 32'b11111111111111111010110110011011;
assign LUT_4[17680] = 32'b00000000000000001001110100111100;
assign LUT_4[17681] = 32'b00000000000000000011000000110100;
assign LUT_4[17682] = 32'b00000000000000001001001111100000;
assign LUT_4[17683] = 32'b00000000000000000010011011011000;
assign LUT_4[17684] = 32'b00000000000000000110110101011000;
assign LUT_4[17685] = 32'b00000000000000000000000001010000;
assign LUT_4[17686] = 32'b00000000000000000110001111111100;
assign LUT_4[17687] = 32'b11111111111111111111011011110100;
assign LUT_4[17688] = 32'b00000000000000000011000001010001;
assign LUT_4[17689] = 32'b11111111111111111100001101001001;
assign LUT_4[17690] = 32'b00000000000000000010011011110101;
assign LUT_4[17691] = 32'b11111111111111111011100111101101;
assign LUT_4[17692] = 32'b00000000000000000000000001101101;
assign LUT_4[17693] = 32'b11111111111111111001001101100101;
assign LUT_4[17694] = 32'b11111111111111111111011100010001;
assign LUT_4[17695] = 32'b11111111111111111000101000001001;
assign LUT_4[17696] = 32'b00000000000000001010011110010101;
assign LUT_4[17697] = 32'b00000000000000000011101010001101;
assign LUT_4[17698] = 32'b00000000000000001001111000111001;
assign LUT_4[17699] = 32'b00000000000000000011000100110001;
assign LUT_4[17700] = 32'b00000000000000000111011110110001;
assign LUT_4[17701] = 32'b00000000000000000000101010101001;
assign LUT_4[17702] = 32'b00000000000000000110111001010101;
assign LUT_4[17703] = 32'b00000000000000000000000101001101;
assign LUT_4[17704] = 32'b00000000000000000011101010101010;
assign LUT_4[17705] = 32'b11111111111111111100110110100010;
assign LUT_4[17706] = 32'b00000000000000000011000101001110;
assign LUT_4[17707] = 32'b11111111111111111100010001000110;
assign LUT_4[17708] = 32'b00000000000000000000101011000110;
assign LUT_4[17709] = 32'b11111111111111111001110110111110;
assign LUT_4[17710] = 32'b00000000000000000000000101101010;
assign LUT_4[17711] = 32'b11111111111111111001010001100010;
assign LUT_4[17712] = 32'b00000000000000001000010000000011;
assign LUT_4[17713] = 32'b00000000000000000001011011111011;
assign LUT_4[17714] = 32'b00000000000000000111101010100111;
assign LUT_4[17715] = 32'b00000000000000000000110110011111;
assign LUT_4[17716] = 32'b00000000000000000101010000011111;
assign LUT_4[17717] = 32'b11111111111111111110011100010111;
assign LUT_4[17718] = 32'b00000000000000000100101011000011;
assign LUT_4[17719] = 32'b11111111111111111101110110111011;
assign LUT_4[17720] = 32'b00000000000000000001011100011000;
assign LUT_4[17721] = 32'b11111111111111111010101000010000;
assign LUT_4[17722] = 32'b00000000000000000000110110111100;
assign LUT_4[17723] = 32'b11111111111111111010000010110100;
assign LUT_4[17724] = 32'b11111111111111111110011100110100;
assign LUT_4[17725] = 32'b11111111111111110111101000101100;
assign LUT_4[17726] = 32'b11111111111111111101110111011000;
assign LUT_4[17727] = 32'b11111111111111110111000011010000;
assign LUT_4[17728] = 32'b00000000000000001101011010100010;
assign LUT_4[17729] = 32'b00000000000000000110100110011010;
assign LUT_4[17730] = 32'b00000000000000001100110101000110;
assign LUT_4[17731] = 32'b00000000000000000110000000111110;
assign LUT_4[17732] = 32'b00000000000000001010011010111110;
assign LUT_4[17733] = 32'b00000000000000000011100110110110;
assign LUT_4[17734] = 32'b00000000000000001001110101100010;
assign LUT_4[17735] = 32'b00000000000000000011000001011010;
assign LUT_4[17736] = 32'b00000000000000000110100110110111;
assign LUT_4[17737] = 32'b11111111111111111111110010101111;
assign LUT_4[17738] = 32'b00000000000000000110000001011011;
assign LUT_4[17739] = 32'b11111111111111111111001101010011;
assign LUT_4[17740] = 32'b00000000000000000011100111010011;
assign LUT_4[17741] = 32'b11111111111111111100110011001011;
assign LUT_4[17742] = 32'b00000000000000000011000001110111;
assign LUT_4[17743] = 32'b11111111111111111100001101101111;
assign LUT_4[17744] = 32'b00000000000000001011001100010000;
assign LUT_4[17745] = 32'b00000000000000000100011000001000;
assign LUT_4[17746] = 32'b00000000000000001010100110110100;
assign LUT_4[17747] = 32'b00000000000000000011110010101100;
assign LUT_4[17748] = 32'b00000000000000001000001100101100;
assign LUT_4[17749] = 32'b00000000000000000001011000100100;
assign LUT_4[17750] = 32'b00000000000000000111100111010000;
assign LUT_4[17751] = 32'b00000000000000000000110011001000;
assign LUT_4[17752] = 32'b00000000000000000100011000100101;
assign LUT_4[17753] = 32'b11111111111111111101100100011101;
assign LUT_4[17754] = 32'b00000000000000000011110011001001;
assign LUT_4[17755] = 32'b11111111111111111100111111000001;
assign LUT_4[17756] = 32'b00000000000000000001011001000001;
assign LUT_4[17757] = 32'b11111111111111111010100100111001;
assign LUT_4[17758] = 32'b00000000000000000000110011100101;
assign LUT_4[17759] = 32'b11111111111111111001111111011101;
assign LUT_4[17760] = 32'b00000000000000001011110101101001;
assign LUT_4[17761] = 32'b00000000000000000101000001100001;
assign LUT_4[17762] = 32'b00000000000000001011010000001101;
assign LUT_4[17763] = 32'b00000000000000000100011100000101;
assign LUT_4[17764] = 32'b00000000000000001000110110000101;
assign LUT_4[17765] = 32'b00000000000000000010000001111101;
assign LUT_4[17766] = 32'b00000000000000001000010000101001;
assign LUT_4[17767] = 32'b00000000000000000001011100100001;
assign LUT_4[17768] = 32'b00000000000000000101000001111110;
assign LUT_4[17769] = 32'b11111111111111111110001101110110;
assign LUT_4[17770] = 32'b00000000000000000100011100100010;
assign LUT_4[17771] = 32'b11111111111111111101101000011010;
assign LUT_4[17772] = 32'b00000000000000000010000010011010;
assign LUT_4[17773] = 32'b11111111111111111011001110010010;
assign LUT_4[17774] = 32'b00000000000000000001011100111110;
assign LUT_4[17775] = 32'b11111111111111111010101000110110;
assign LUT_4[17776] = 32'b00000000000000001001100111010111;
assign LUT_4[17777] = 32'b00000000000000000010110011001111;
assign LUT_4[17778] = 32'b00000000000000001001000001111011;
assign LUT_4[17779] = 32'b00000000000000000010001101110011;
assign LUT_4[17780] = 32'b00000000000000000110100111110011;
assign LUT_4[17781] = 32'b11111111111111111111110011101011;
assign LUT_4[17782] = 32'b00000000000000000110000010010111;
assign LUT_4[17783] = 32'b11111111111111111111001110001111;
assign LUT_4[17784] = 32'b00000000000000000010110011101100;
assign LUT_4[17785] = 32'b11111111111111111011111111100100;
assign LUT_4[17786] = 32'b00000000000000000010001110010000;
assign LUT_4[17787] = 32'b11111111111111111011011010001000;
assign LUT_4[17788] = 32'b11111111111111111111110100001000;
assign LUT_4[17789] = 32'b11111111111111111001000000000000;
assign LUT_4[17790] = 32'b11111111111111111111001110101100;
assign LUT_4[17791] = 32'b11111111111111111000011010100100;
assign LUT_4[17792] = 32'b00000000000000001110101001010110;
assign LUT_4[17793] = 32'b00000000000000000111110101001110;
assign LUT_4[17794] = 32'b00000000000000001110000011111010;
assign LUT_4[17795] = 32'b00000000000000000111001111110010;
assign LUT_4[17796] = 32'b00000000000000001011101001110010;
assign LUT_4[17797] = 32'b00000000000000000100110101101010;
assign LUT_4[17798] = 32'b00000000000000001011000100010110;
assign LUT_4[17799] = 32'b00000000000000000100010000001110;
assign LUT_4[17800] = 32'b00000000000000000111110101101011;
assign LUT_4[17801] = 32'b00000000000000000001000001100011;
assign LUT_4[17802] = 32'b00000000000000000111010000001111;
assign LUT_4[17803] = 32'b00000000000000000000011100000111;
assign LUT_4[17804] = 32'b00000000000000000100110110000111;
assign LUT_4[17805] = 32'b11111111111111111110000001111111;
assign LUT_4[17806] = 32'b00000000000000000100010000101011;
assign LUT_4[17807] = 32'b11111111111111111101011100100011;
assign LUT_4[17808] = 32'b00000000000000001100011011000100;
assign LUT_4[17809] = 32'b00000000000000000101100110111100;
assign LUT_4[17810] = 32'b00000000000000001011110101101000;
assign LUT_4[17811] = 32'b00000000000000000101000001100000;
assign LUT_4[17812] = 32'b00000000000000001001011011100000;
assign LUT_4[17813] = 32'b00000000000000000010100111011000;
assign LUT_4[17814] = 32'b00000000000000001000110110000100;
assign LUT_4[17815] = 32'b00000000000000000010000001111100;
assign LUT_4[17816] = 32'b00000000000000000101100111011001;
assign LUT_4[17817] = 32'b11111111111111111110110011010001;
assign LUT_4[17818] = 32'b00000000000000000101000001111101;
assign LUT_4[17819] = 32'b11111111111111111110001101110101;
assign LUT_4[17820] = 32'b00000000000000000010100111110101;
assign LUT_4[17821] = 32'b11111111111111111011110011101101;
assign LUT_4[17822] = 32'b00000000000000000010000010011001;
assign LUT_4[17823] = 32'b11111111111111111011001110010001;
assign LUT_4[17824] = 32'b00000000000000001101000100011101;
assign LUT_4[17825] = 32'b00000000000000000110010000010101;
assign LUT_4[17826] = 32'b00000000000000001100011111000001;
assign LUT_4[17827] = 32'b00000000000000000101101010111001;
assign LUT_4[17828] = 32'b00000000000000001010000100111001;
assign LUT_4[17829] = 32'b00000000000000000011010000110001;
assign LUT_4[17830] = 32'b00000000000000001001011111011101;
assign LUT_4[17831] = 32'b00000000000000000010101011010101;
assign LUT_4[17832] = 32'b00000000000000000110010000110010;
assign LUT_4[17833] = 32'b11111111111111111111011100101010;
assign LUT_4[17834] = 32'b00000000000000000101101011010110;
assign LUT_4[17835] = 32'b11111111111111111110110111001110;
assign LUT_4[17836] = 32'b00000000000000000011010001001110;
assign LUT_4[17837] = 32'b11111111111111111100011101000110;
assign LUT_4[17838] = 32'b00000000000000000010101011110010;
assign LUT_4[17839] = 32'b11111111111111111011110111101010;
assign LUT_4[17840] = 32'b00000000000000001010110110001011;
assign LUT_4[17841] = 32'b00000000000000000100000010000011;
assign LUT_4[17842] = 32'b00000000000000001010010000101111;
assign LUT_4[17843] = 32'b00000000000000000011011100100111;
assign LUT_4[17844] = 32'b00000000000000000111110110100111;
assign LUT_4[17845] = 32'b00000000000000000001000010011111;
assign LUT_4[17846] = 32'b00000000000000000111010001001011;
assign LUT_4[17847] = 32'b00000000000000000000011101000011;
assign LUT_4[17848] = 32'b00000000000000000100000010100000;
assign LUT_4[17849] = 32'b11111111111111111101001110011000;
assign LUT_4[17850] = 32'b00000000000000000011011101000100;
assign LUT_4[17851] = 32'b11111111111111111100101000111100;
assign LUT_4[17852] = 32'b00000000000000000001000010111100;
assign LUT_4[17853] = 32'b11111111111111111010001110110100;
assign LUT_4[17854] = 32'b00000000000000000000011101100000;
assign LUT_4[17855] = 32'b11111111111111111001101001011000;
assign LUT_4[17856] = 32'b00000000000000010000000000101010;
assign LUT_4[17857] = 32'b00000000000000001001001100100010;
assign LUT_4[17858] = 32'b00000000000000001111011011001110;
assign LUT_4[17859] = 32'b00000000000000001000100111000110;
assign LUT_4[17860] = 32'b00000000000000001101000001000110;
assign LUT_4[17861] = 32'b00000000000000000110001100111110;
assign LUT_4[17862] = 32'b00000000000000001100011011101010;
assign LUT_4[17863] = 32'b00000000000000000101100111100010;
assign LUT_4[17864] = 32'b00000000000000001001001100111111;
assign LUT_4[17865] = 32'b00000000000000000010011000110111;
assign LUT_4[17866] = 32'b00000000000000001000100111100011;
assign LUT_4[17867] = 32'b00000000000000000001110011011011;
assign LUT_4[17868] = 32'b00000000000000000110001101011011;
assign LUT_4[17869] = 32'b11111111111111111111011001010011;
assign LUT_4[17870] = 32'b00000000000000000101100111111111;
assign LUT_4[17871] = 32'b11111111111111111110110011110111;
assign LUT_4[17872] = 32'b00000000000000001101110010011000;
assign LUT_4[17873] = 32'b00000000000000000110111110010000;
assign LUT_4[17874] = 32'b00000000000000001101001100111100;
assign LUT_4[17875] = 32'b00000000000000000110011000110100;
assign LUT_4[17876] = 32'b00000000000000001010110010110100;
assign LUT_4[17877] = 32'b00000000000000000011111110101100;
assign LUT_4[17878] = 32'b00000000000000001010001101011000;
assign LUT_4[17879] = 32'b00000000000000000011011001010000;
assign LUT_4[17880] = 32'b00000000000000000110111110101101;
assign LUT_4[17881] = 32'b00000000000000000000001010100101;
assign LUT_4[17882] = 32'b00000000000000000110011001010001;
assign LUT_4[17883] = 32'b11111111111111111111100101001001;
assign LUT_4[17884] = 32'b00000000000000000011111111001001;
assign LUT_4[17885] = 32'b11111111111111111101001011000001;
assign LUT_4[17886] = 32'b00000000000000000011011001101101;
assign LUT_4[17887] = 32'b11111111111111111100100101100101;
assign LUT_4[17888] = 32'b00000000000000001110011011110001;
assign LUT_4[17889] = 32'b00000000000000000111100111101001;
assign LUT_4[17890] = 32'b00000000000000001101110110010101;
assign LUT_4[17891] = 32'b00000000000000000111000010001101;
assign LUT_4[17892] = 32'b00000000000000001011011100001101;
assign LUT_4[17893] = 32'b00000000000000000100101000000101;
assign LUT_4[17894] = 32'b00000000000000001010110110110001;
assign LUT_4[17895] = 32'b00000000000000000100000010101001;
assign LUT_4[17896] = 32'b00000000000000000111101000000110;
assign LUT_4[17897] = 32'b00000000000000000000110011111110;
assign LUT_4[17898] = 32'b00000000000000000111000010101010;
assign LUT_4[17899] = 32'b00000000000000000000001110100010;
assign LUT_4[17900] = 32'b00000000000000000100101000100010;
assign LUT_4[17901] = 32'b11111111111111111101110100011010;
assign LUT_4[17902] = 32'b00000000000000000100000011000110;
assign LUT_4[17903] = 32'b11111111111111111101001110111110;
assign LUT_4[17904] = 32'b00000000000000001100001101011111;
assign LUT_4[17905] = 32'b00000000000000000101011001010111;
assign LUT_4[17906] = 32'b00000000000000001011101000000011;
assign LUT_4[17907] = 32'b00000000000000000100110011111011;
assign LUT_4[17908] = 32'b00000000000000001001001101111011;
assign LUT_4[17909] = 32'b00000000000000000010011001110011;
assign LUT_4[17910] = 32'b00000000000000001000101000011111;
assign LUT_4[17911] = 32'b00000000000000000001110100010111;
assign LUT_4[17912] = 32'b00000000000000000101011001110100;
assign LUT_4[17913] = 32'b11111111111111111110100101101100;
assign LUT_4[17914] = 32'b00000000000000000100110100011000;
assign LUT_4[17915] = 32'b11111111111111111110000000010000;
assign LUT_4[17916] = 32'b00000000000000000010011010010000;
assign LUT_4[17917] = 32'b11111111111111111011100110001000;
assign LUT_4[17918] = 32'b00000000000000000001110100110100;
assign LUT_4[17919] = 32'b11111111111111111011000000101100;
assign LUT_4[17920] = 32'b00000000000000000110001011110011;
assign LUT_4[17921] = 32'b11111111111111111111010111101011;
assign LUT_4[17922] = 32'b00000000000000000101100110010111;
assign LUT_4[17923] = 32'b11111111111111111110110010001111;
assign LUT_4[17924] = 32'b00000000000000000011001100001111;
assign LUT_4[17925] = 32'b11111111111111111100011000000111;
assign LUT_4[17926] = 32'b00000000000000000010100110110011;
assign LUT_4[17927] = 32'b11111111111111111011110010101011;
assign LUT_4[17928] = 32'b11111111111111111111011000001000;
assign LUT_4[17929] = 32'b11111111111111111000100100000000;
assign LUT_4[17930] = 32'b11111111111111111110110010101100;
assign LUT_4[17931] = 32'b11111111111111110111111110100100;
assign LUT_4[17932] = 32'b11111111111111111100011000100100;
assign LUT_4[17933] = 32'b11111111111111110101100100011100;
assign LUT_4[17934] = 32'b11111111111111111011110011001000;
assign LUT_4[17935] = 32'b11111111111111110100111111000000;
assign LUT_4[17936] = 32'b00000000000000000011111101100001;
assign LUT_4[17937] = 32'b11111111111111111101001001011001;
assign LUT_4[17938] = 32'b00000000000000000011011000000101;
assign LUT_4[17939] = 32'b11111111111111111100100011111101;
assign LUT_4[17940] = 32'b00000000000000000000111101111101;
assign LUT_4[17941] = 32'b11111111111111111010001001110101;
assign LUT_4[17942] = 32'b00000000000000000000011000100001;
assign LUT_4[17943] = 32'b11111111111111111001100100011001;
assign LUT_4[17944] = 32'b11111111111111111101001001110110;
assign LUT_4[17945] = 32'b11111111111111110110010101101110;
assign LUT_4[17946] = 32'b11111111111111111100100100011010;
assign LUT_4[17947] = 32'b11111111111111110101110000010010;
assign LUT_4[17948] = 32'b11111111111111111010001010010010;
assign LUT_4[17949] = 32'b11111111111111110011010110001010;
assign LUT_4[17950] = 32'b11111111111111111001100100110110;
assign LUT_4[17951] = 32'b11111111111111110010110000101110;
assign LUT_4[17952] = 32'b00000000000000000100100110111010;
assign LUT_4[17953] = 32'b11111111111111111101110010110010;
assign LUT_4[17954] = 32'b00000000000000000100000001011110;
assign LUT_4[17955] = 32'b11111111111111111101001101010110;
assign LUT_4[17956] = 32'b00000000000000000001100111010110;
assign LUT_4[17957] = 32'b11111111111111111010110011001110;
assign LUT_4[17958] = 32'b00000000000000000001000001111010;
assign LUT_4[17959] = 32'b11111111111111111010001101110010;
assign LUT_4[17960] = 32'b11111111111111111101110011001111;
assign LUT_4[17961] = 32'b11111111111111110110111111000111;
assign LUT_4[17962] = 32'b11111111111111111101001101110011;
assign LUT_4[17963] = 32'b11111111111111110110011001101011;
assign LUT_4[17964] = 32'b11111111111111111010110011101011;
assign LUT_4[17965] = 32'b11111111111111110011111111100011;
assign LUT_4[17966] = 32'b11111111111111111010001110001111;
assign LUT_4[17967] = 32'b11111111111111110011011010000111;
assign LUT_4[17968] = 32'b00000000000000000010011000101000;
assign LUT_4[17969] = 32'b11111111111111111011100100100000;
assign LUT_4[17970] = 32'b00000000000000000001110011001100;
assign LUT_4[17971] = 32'b11111111111111111010111111000100;
assign LUT_4[17972] = 32'b11111111111111111111011001000100;
assign LUT_4[17973] = 32'b11111111111111111000100100111100;
assign LUT_4[17974] = 32'b11111111111111111110110011101000;
assign LUT_4[17975] = 32'b11111111111111110111111111100000;
assign LUT_4[17976] = 32'b11111111111111111011100100111101;
assign LUT_4[17977] = 32'b11111111111111110100110000110101;
assign LUT_4[17978] = 32'b11111111111111111010111111100001;
assign LUT_4[17979] = 32'b11111111111111110100001011011001;
assign LUT_4[17980] = 32'b11111111111111111000100101011001;
assign LUT_4[17981] = 32'b11111111111111110001110001010001;
assign LUT_4[17982] = 32'b11111111111111110111111111111101;
assign LUT_4[17983] = 32'b11111111111111110001001011110101;
assign LUT_4[17984] = 32'b00000000000000000111100011000111;
assign LUT_4[17985] = 32'b00000000000000000000101110111111;
assign LUT_4[17986] = 32'b00000000000000000110111101101011;
assign LUT_4[17987] = 32'b00000000000000000000001001100011;
assign LUT_4[17988] = 32'b00000000000000000100100011100011;
assign LUT_4[17989] = 32'b11111111111111111101101111011011;
assign LUT_4[17990] = 32'b00000000000000000011111110000111;
assign LUT_4[17991] = 32'b11111111111111111101001001111111;
assign LUT_4[17992] = 32'b00000000000000000000101111011100;
assign LUT_4[17993] = 32'b11111111111111111001111011010100;
assign LUT_4[17994] = 32'b00000000000000000000001010000000;
assign LUT_4[17995] = 32'b11111111111111111001010101111000;
assign LUT_4[17996] = 32'b11111111111111111101101111111000;
assign LUT_4[17997] = 32'b11111111111111110110111011110000;
assign LUT_4[17998] = 32'b11111111111111111101001010011100;
assign LUT_4[17999] = 32'b11111111111111110110010110010100;
assign LUT_4[18000] = 32'b00000000000000000101010100110101;
assign LUT_4[18001] = 32'b11111111111111111110100000101101;
assign LUT_4[18002] = 32'b00000000000000000100101111011001;
assign LUT_4[18003] = 32'b11111111111111111101111011010001;
assign LUT_4[18004] = 32'b00000000000000000010010101010001;
assign LUT_4[18005] = 32'b11111111111111111011100001001001;
assign LUT_4[18006] = 32'b00000000000000000001101111110101;
assign LUT_4[18007] = 32'b11111111111111111010111011101101;
assign LUT_4[18008] = 32'b11111111111111111110100001001010;
assign LUT_4[18009] = 32'b11111111111111110111101101000010;
assign LUT_4[18010] = 32'b11111111111111111101111011101110;
assign LUT_4[18011] = 32'b11111111111111110111000111100110;
assign LUT_4[18012] = 32'b11111111111111111011100001100110;
assign LUT_4[18013] = 32'b11111111111111110100101101011110;
assign LUT_4[18014] = 32'b11111111111111111010111100001010;
assign LUT_4[18015] = 32'b11111111111111110100001000000010;
assign LUT_4[18016] = 32'b00000000000000000101111110001110;
assign LUT_4[18017] = 32'b11111111111111111111001010000110;
assign LUT_4[18018] = 32'b00000000000000000101011000110010;
assign LUT_4[18019] = 32'b11111111111111111110100100101010;
assign LUT_4[18020] = 32'b00000000000000000010111110101010;
assign LUT_4[18021] = 32'b11111111111111111100001010100010;
assign LUT_4[18022] = 32'b00000000000000000010011001001110;
assign LUT_4[18023] = 32'b11111111111111111011100101000110;
assign LUT_4[18024] = 32'b11111111111111111111001010100011;
assign LUT_4[18025] = 32'b11111111111111111000010110011011;
assign LUT_4[18026] = 32'b11111111111111111110100101000111;
assign LUT_4[18027] = 32'b11111111111111110111110000111111;
assign LUT_4[18028] = 32'b11111111111111111100001010111111;
assign LUT_4[18029] = 32'b11111111111111110101010110110111;
assign LUT_4[18030] = 32'b11111111111111111011100101100011;
assign LUT_4[18031] = 32'b11111111111111110100110001011011;
assign LUT_4[18032] = 32'b00000000000000000011101111111100;
assign LUT_4[18033] = 32'b11111111111111111100111011110100;
assign LUT_4[18034] = 32'b00000000000000000011001010100000;
assign LUT_4[18035] = 32'b11111111111111111100010110011000;
assign LUT_4[18036] = 32'b00000000000000000000110000011000;
assign LUT_4[18037] = 32'b11111111111111111001111100010000;
assign LUT_4[18038] = 32'b00000000000000000000001010111100;
assign LUT_4[18039] = 32'b11111111111111111001010110110100;
assign LUT_4[18040] = 32'b11111111111111111100111100010001;
assign LUT_4[18041] = 32'b11111111111111110110001000001001;
assign LUT_4[18042] = 32'b11111111111111111100010110110101;
assign LUT_4[18043] = 32'b11111111111111110101100010101101;
assign LUT_4[18044] = 32'b11111111111111111001111100101101;
assign LUT_4[18045] = 32'b11111111111111110011001000100101;
assign LUT_4[18046] = 32'b11111111111111111001010111010001;
assign LUT_4[18047] = 32'b11111111111111110010100011001001;
assign LUT_4[18048] = 32'b00000000000000001000110001111011;
assign LUT_4[18049] = 32'b00000000000000000001111101110011;
assign LUT_4[18050] = 32'b00000000000000001000001100011111;
assign LUT_4[18051] = 32'b00000000000000000001011000010111;
assign LUT_4[18052] = 32'b00000000000000000101110010010111;
assign LUT_4[18053] = 32'b11111111111111111110111110001111;
assign LUT_4[18054] = 32'b00000000000000000101001100111011;
assign LUT_4[18055] = 32'b11111111111111111110011000110011;
assign LUT_4[18056] = 32'b00000000000000000001111110010000;
assign LUT_4[18057] = 32'b11111111111111111011001010001000;
assign LUT_4[18058] = 32'b00000000000000000001011000110100;
assign LUT_4[18059] = 32'b11111111111111111010100100101100;
assign LUT_4[18060] = 32'b11111111111111111110111110101100;
assign LUT_4[18061] = 32'b11111111111111111000001010100100;
assign LUT_4[18062] = 32'b11111111111111111110011001010000;
assign LUT_4[18063] = 32'b11111111111111110111100101001000;
assign LUT_4[18064] = 32'b00000000000000000110100011101001;
assign LUT_4[18065] = 32'b11111111111111111111101111100001;
assign LUT_4[18066] = 32'b00000000000000000101111110001101;
assign LUT_4[18067] = 32'b11111111111111111111001010000101;
assign LUT_4[18068] = 32'b00000000000000000011100100000101;
assign LUT_4[18069] = 32'b11111111111111111100101111111101;
assign LUT_4[18070] = 32'b00000000000000000010111110101001;
assign LUT_4[18071] = 32'b11111111111111111100001010100001;
assign LUT_4[18072] = 32'b11111111111111111111101111111110;
assign LUT_4[18073] = 32'b11111111111111111000111011110110;
assign LUT_4[18074] = 32'b11111111111111111111001010100010;
assign LUT_4[18075] = 32'b11111111111111111000010110011010;
assign LUT_4[18076] = 32'b11111111111111111100110000011010;
assign LUT_4[18077] = 32'b11111111111111110101111100010010;
assign LUT_4[18078] = 32'b11111111111111111100001010111110;
assign LUT_4[18079] = 32'b11111111111111110101010110110110;
assign LUT_4[18080] = 32'b00000000000000000111001101000010;
assign LUT_4[18081] = 32'b00000000000000000000011000111010;
assign LUT_4[18082] = 32'b00000000000000000110100111100110;
assign LUT_4[18083] = 32'b11111111111111111111110011011110;
assign LUT_4[18084] = 32'b00000000000000000100001101011110;
assign LUT_4[18085] = 32'b11111111111111111101011001010110;
assign LUT_4[18086] = 32'b00000000000000000011101000000010;
assign LUT_4[18087] = 32'b11111111111111111100110011111010;
assign LUT_4[18088] = 32'b00000000000000000000011001010111;
assign LUT_4[18089] = 32'b11111111111111111001100101001111;
assign LUT_4[18090] = 32'b11111111111111111111110011111011;
assign LUT_4[18091] = 32'b11111111111111111000111111110011;
assign LUT_4[18092] = 32'b11111111111111111101011001110011;
assign LUT_4[18093] = 32'b11111111111111110110100101101011;
assign LUT_4[18094] = 32'b11111111111111111100110100010111;
assign LUT_4[18095] = 32'b11111111111111110110000000001111;
assign LUT_4[18096] = 32'b00000000000000000100111110110000;
assign LUT_4[18097] = 32'b11111111111111111110001010101000;
assign LUT_4[18098] = 32'b00000000000000000100011001010100;
assign LUT_4[18099] = 32'b11111111111111111101100101001100;
assign LUT_4[18100] = 32'b00000000000000000001111111001100;
assign LUT_4[18101] = 32'b11111111111111111011001011000100;
assign LUT_4[18102] = 32'b00000000000000000001011001110000;
assign LUT_4[18103] = 32'b11111111111111111010100101101000;
assign LUT_4[18104] = 32'b11111111111111111110001011000101;
assign LUT_4[18105] = 32'b11111111111111110111010110111101;
assign LUT_4[18106] = 32'b11111111111111111101100101101001;
assign LUT_4[18107] = 32'b11111111111111110110110001100001;
assign LUT_4[18108] = 32'b11111111111111111011001011100001;
assign LUT_4[18109] = 32'b11111111111111110100010111011001;
assign LUT_4[18110] = 32'b11111111111111111010100110000101;
assign LUT_4[18111] = 32'b11111111111111110011110001111101;
assign LUT_4[18112] = 32'b00000000000000001010001001001111;
assign LUT_4[18113] = 32'b00000000000000000011010101000111;
assign LUT_4[18114] = 32'b00000000000000001001100011110011;
assign LUT_4[18115] = 32'b00000000000000000010101111101011;
assign LUT_4[18116] = 32'b00000000000000000111001001101011;
assign LUT_4[18117] = 32'b00000000000000000000010101100011;
assign LUT_4[18118] = 32'b00000000000000000110100100001111;
assign LUT_4[18119] = 32'b11111111111111111111110000000111;
assign LUT_4[18120] = 32'b00000000000000000011010101100100;
assign LUT_4[18121] = 32'b11111111111111111100100001011100;
assign LUT_4[18122] = 32'b00000000000000000010110000001000;
assign LUT_4[18123] = 32'b11111111111111111011111100000000;
assign LUT_4[18124] = 32'b00000000000000000000010110000000;
assign LUT_4[18125] = 32'b11111111111111111001100001111000;
assign LUT_4[18126] = 32'b11111111111111111111110000100100;
assign LUT_4[18127] = 32'b11111111111111111000111100011100;
assign LUT_4[18128] = 32'b00000000000000000111111010111101;
assign LUT_4[18129] = 32'b00000000000000000001000110110101;
assign LUT_4[18130] = 32'b00000000000000000111010101100001;
assign LUT_4[18131] = 32'b00000000000000000000100001011001;
assign LUT_4[18132] = 32'b00000000000000000100111011011001;
assign LUT_4[18133] = 32'b11111111111111111110000111010001;
assign LUT_4[18134] = 32'b00000000000000000100010101111101;
assign LUT_4[18135] = 32'b11111111111111111101100001110101;
assign LUT_4[18136] = 32'b00000000000000000001000111010010;
assign LUT_4[18137] = 32'b11111111111111111010010011001010;
assign LUT_4[18138] = 32'b00000000000000000000100001110110;
assign LUT_4[18139] = 32'b11111111111111111001101101101110;
assign LUT_4[18140] = 32'b11111111111111111110000111101110;
assign LUT_4[18141] = 32'b11111111111111110111010011100110;
assign LUT_4[18142] = 32'b11111111111111111101100010010010;
assign LUT_4[18143] = 32'b11111111111111110110101110001010;
assign LUT_4[18144] = 32'b00000000000000001000100100010110;
assign LUT_4[18145] = 32'b00000000000000000001110000001110;
assign LUT_4[18146] = 32'b00000000000000000111111110111010;
assign LUT_4[18147] = 32'b00000000000000000001001010110010;
assign LUT_4[18148] = 32'b00000000000000000101100100110010;
assign LUT_4[18149] = 32'b11111111111111111110110000101010;
assign LUT_4[18150] = 32'b00000000000000000100111111010110;
assign LUT_4[18151] = 32'b11111111111111111110001011001110;
assign LUT_4[18152] = 32'b00000000000000000001110000101011;
assign LUT_4[18153] = 32'b11111111111111111010111100100011;
assign LUT_4[18154] = 32'b00000000000000000001001011001111;
assign LUT_4[18155] = 32'b11111111111111111010010111000111;
assign LUT_4[18156] = 32'b11111111111111111110110001000111;
assign LUT_4[18157] = 32'b11111111111111110111111100111111;
assign LUT_4[18158] = 32'b11111111111111111110001011101011;
assign LUT_4[18159] = 32'b11111111111111110111010111100011;
assign LUT_4[18160] = 32'b00000000000000000110010110000100;
assign LUT_4[18161] = 32'b11111111111111111111100001111100;
assign LUT_4[18162] = 32'b00000000000000000101110000101000;
assign LUT_4[18163] = 32'b11111111111111111110111100100000;
assign LUT_4[18164] = 32'b00000000000000000011010110100000;
assign LUT_4[18165] = 32'b11111111111111111100100010011000;
assign LUT_4[18166] = 32'b00000000000000000010110001000100;
assign LUT_4[18167] = 32'b11111111111111111011111100111100;
assign LUT_4[18168] = 32'b11111111111111111111100010011001;
assign LUT_4[18169] = 32'b11111111111111111000101110010001;
assign LUT_4[18170] = 32'b11111111111111111110111100111101;
assign LUT_4[18171] = 32'b11111111111111111000001000110101;
assign LUT_4[18172] = 32'b11111111111111111100100010110101;
assign LUT_4[18173] = 32'b11111111111111110101101110101101;
assign LUT_4[18174] = 32'b11111111111111111011111101011001;
assign LUT_4[18175] = 32'b11111111111111110101001001010001;
assign LUT_4[18176] = 32'b00000000000000001011000111010110;
assign LUT_4[18177] = 32'b00000000000000000100010011001110;
assign LUT_4[18178] = 32'b00000000000000001010100001111010;
assign LUT_4[18179] = 32'b00000000000000000011101101110010;
assign LUT_4[18180] = 32'b00000000000000001000000111110010;
assign LUT_4[18181] = 32'b00000000000000000001010011101010;
assign LUT_4[18182] = 32'b00000000000000000111100010010110;
assign LUT_4[18183] = 32'b00000000000000000000101110001110;
assign LUT_4[18184] = 32'b00000000000000000100010011101011;
assign LUT_4[18185] = 32'b11111111111111111101011111100011;
assign LUT_4[18186] = 32'b00000000000000000011101110001111;
assign LUT_4[18187] = 32'b11111111111111111100111010000111;
assign LUT_4[18188] = 32'b00000000000000000001010100000111;
assign LUT_4[18189] = 32'b11111111111111111010011111111111;
assign LUT_4[18190] = 32'b00000000000000000000101110101011;
assign LUT_4[18191] = 32'b11111111111111111001111010100011;
assign LUT_4[18192] = 32'b00000000000000001000111001000100;
assign LUT_4[18193] = 32'b00000000000000000010000100111100;
assign LUT_4[18194] = 32'b00000000000000001000010011101000;
assign LUT_4[18195] = 32'b00000000000000000001011111100000;
assign LUT_4[18196] = 32'b00000000000000000101111001100000;
assign LUT_4[18197] = 32'b11111111111111111111000101011000;
assign LUT_4[18198] = 32'b00000000000000000101010100000100;
assign LUT_4[18199] = 32'b11111111111111111110011111111100;
assign LUT_4[18200] = 32'b00000000000000000010000101011001;
assign LUT_4[18201] = 32'b11111111111111111011010001010001;
assign LUT_4[18202] = 32'b00000000000000000001011111111101;
assign LUT_4[18203] = 32'b11111111111111111010101011110101;
assign LUT_4[18204] = 32'b11111111111111111111000101110101;
assign LUT_4[18205] = 32'b11111111111111111000010001101101;
assign LUT_4[18206] = 32'b11111111111111111110100000011001;
assign LUT_4[18207] = 32'b11111111111111110111101100010001;
assign LUT_4[18208] = 32'b00000000000000001001100010011101;
assign LUT_4[18209] = 32'b00000000000000000010101110010101;
assign LUT_4[18210] = 32'b00000000000000001000111101000001;
assign LUT_4[18211] = 32'b00000000000000000010001000111001;
assign LUT_4[18212] = 32'b00000000000000000110100010111001;
assign LUT_4[18213] = 32'b11111111111111111111101110110001;
assign LUT_4[18214] = 32'b00000000000000000101111101011101;
assign LUT_4[18215] = 32'b11111111111111111111001001010101;
assign LUT_4[18216] = 32'b00000000000000000010101110110010;
assign LUT_4[18217] = 32'b11111111111111111011111010101010;
assign LUT_4[18218] = 32'b00000000000000000010001001010110;
assign LUT_4[18219] = 32'b11111111111111111011010101001110;
assign LUT_4[18220] = 32'b11111111111111111111101111001110;
assign LUT_4[18221] = 32'b11111111111111111000111011000110;
assign LUT_4[18222] = 32'b11111111111111111111001001110010;
assign LUT_4[18223] = 32'b11111111111111111000010101101010;
assign LUT_4[18224] = 32'b00000000000000000111010100001011;
assign LUT_4[18225] = 32'b00000000000000000000100000000011;
assign LUT_4[18226] = 32'b00000000000000000110101110101111;
assign LUT_4[18227] = 32'b11111111111111111111111010100111;
assign LUT_4[18228] = 32'b00000000000000000100010100100111;
assign LUT_4[18229] = 32'b11111111111111111101100000011111;
assign LUT_4[18230] = 32'b00000000000000000011101111001011;
assign LUT_4[18231] = 32'b11111111111111111100111011000011;
assign LUT_4[18232] = 32'b00000000000000000000100000100000;
assign LUT_4[18233] = 32'b11111111111111111001101100011000;
assign LUT_4[18234] = 32'b11111111111111111111111011000100;
assign LUT_4[18235] = 32'b11111111111111111001000110111100;
assign LUT_4[18236] = 32'b11111111111111111101100000111100;
assign LUT_4[18237] = 32'b11111111111111110110101100110100;
assign LUT_4[18238] = 32'b11111111111111111100111011100000;
assign LUT_4[18239] = 32'b11111111111111110110000111011000;
assign LUT_4[18240] = 32'b00000000000000001100011110101010;
assign LUT_4[18241] = 32'b00000000000000000101101010100010;
assign LUT_4[18242] = 32'b00000000000000001011111001001110;
assign LUT_4[18243] = 32'b00000000000000000101000101000110;
assign LUT_4[18244] = 32'b00000000000000001001011111000110;
assign LUT_4[18245] = 32'b00000000000000000010101010111110;
assign LUT_4[18246] = 32'b00000000000000001000111001101010;
assign LUT_4[18247] = 32'b00000000000000000010000101100010;
assign LUT_4[18248] = 32'b00000000000000000101101010111111;
assign LUT_4[18249] = 32'b11111111111111111110110110110111;
assign LUT_4[18250] = 32'b00000000000000000101000101100011;
assign LUT_4[18251] = 32'b11111111111111111110010001011011;
assign LUT_4[18252] = 32'b00000000000000000010101011011011;
assign LUT_4[18253] = 32'b11111111111111111011110111010011;
assign LUT_4[18254] = 32'b00000000000000000010000101111111;
assign LUT_4[18255] = 32'b11111111111111111011010001110111;
assign LUT_4[18256] = 32'b00000000000000001010010000011000;
assign LUT_4[18257] = 32'b00000000000000000011011100010000;
assign LUT_4[18258] = 32'b00000000000000001001101010111100;
assign LUT_4[18259] = 32'b00000000000000000010110110110100;
assign LUT_4[18260] = 32'b00000000000000000111010000110100;
assign LUT_4[18261] = 32'b00000000000000000000011100101100;
assign LUT_4[18262] = 32'b00000000000000000110101011011000;
assign LUT_4[18263] = 32'b11111111111111111111110111010000;
assign LUT_4[18264] = 32'b00000000000000000011011100101101;
assign LUT_4[18265] = 32'b11111111111111111100101000100101;
assign LUT_4[18266] = 32'b00000000000000000010110111010001;
assign LUT_4[18267] = 32'b11111111111111111100000011001001;
assign LUT_4[18268] = 32'b00000000000000000000011101001001;
assign LUT_4[18269] = 32'b11111111111111111001101001000001;
assign LUT_4[18270] = 32'b11111111111111111111110111101101;
assign LUT_4[18271] = 32'b11111111111111111001000011100101;
assign LUT_4[18272] = 32'b00000000000000001010111001110001;
assign LUT_4[18273] = 32'b00000000000000000100000101101001;
assign LUT_4[18274] = 32'b00000000000000001010010100010101;
assign LUT_4[18275] = 32'b00000000000000000011100000001101;
assign LUT_4[18276] = 32'b00000000000000000111111010001101;
assign LUT_4[18277] = 32'b00000000000000000001000110000101;
assign LUT_4[18278] = 32'b00000000000000000111010100110001;
assign LUT_4[18279] = 32'b00000000000000000000100000101001;
assign LUT_4[18280] = 32'b00000000000000000100000110000110;
assign LUT_4[18281] = 32'b11111111111111111101010001111110;
assign LUT_4[18282] = 32'b00000000000000000011100000101010;
assign LUT_4[18283] = 32'b11111111111111111100101100100010;
assign LUT_4[18284] = 32'b00000000000000000001000110100010;
assign LUT_4[18285] = 32'b11111111111111111010010010011010;
assign LUT_4[18286] = 32'b00000000000000000000100001000110;
assign LUT_4[18287] = 32'b11111111111111111001101100111110;
assign LUT_4[18288] = 32'b00000000000000001000101011011111;
assign LUT_4[18289] = 32'b00000000000000000001110111010111;
assign LUT_4[18290] = 32'b00000000000000001000000110000011;
assign LUT_4[18291] = 32'b00000000000000000001010001111011;
assign LUT_4[18292] = 32'b00000000000000000101101011111011;
assign LUT_4[18293] = 32'b11111111111111111110110111110011;
assign LUT_4[18294] = 32'b00000000000000000101000110011111;
assign LUT_4[18295] = 32'b11111111111111111110010010010111;
assign LUT_4[18296] = 32'b00000000000000000001110111110100;
assign LUT_4[18297] = 32'b11111111111111111011000011101100;
assign LUT_4[18298] = 32'b00000000000000000001010010011000;
assign LUT_4[18299] = 32'b11111111111111111010011110010000;
assign LUT_4[18300] = 32'b11111111111111111110111000010000;
assign LUT_4[18301] = 32'b11111111111111111000000100001000;
assign LUT_4[18302] = 32'b11111111111111111110010010110100;
assign LUT_4[18303] = 32'b11111111111111110111011110101100;
assign LUT_4[18304] = 32'b00000000000000001101101101011110;
assign LUT_4[18305] = 32'b00000000000000000110111001010110;
assign LUT_4[18306] = 32'b00000000000000001101001000000010;
assign LUT_4[18307] = 32'b00000000000000000110010011111010;
assign LUT_4[18308] = 32'b00000000000000001010101101111010;
assign LUT_4[18309] = 32'b00000000000000000011111001110010;
assign LUT_4[18310] = 32'b00000000000000001010001000011110;
assign LUT_4[18311] = 32'b00000000000000000011010100010110;
assign LUT_4[18312] = 32'b00000000000000000110111001110011;
assign LUT_4[18313] = 32'b00000000000000000000000101101011;
assign LUT_4[18314] = 32'b00000000000000000110010100010111;
assign LUT_4[18315] = 32'b11111111111111111111100000001111;
assign LUT_4[18316] = 32'b00000000000000000011111010001111;
assign LUT_4[18317] = 32'b11111111111111111101000110000111;
assign LUT_4[18318] = 32'b00000000000000000011010100110011;
assign LUT_4[18319] = 32'b11111111111111111100100000101011;
assign LUT_4[18320] = 32'b00000000000000001011011111001100;
assign LUT_4[18321] = 32'b00000000000000000100101011000100;
assign LUT_4[18322] = 32'b00000000000000001010111001110000;
assign LUT_4[18323] = 32'b00000000000000000100000101101000;
assign LUT_4[18324] = 32'b00000000000000001000011111101000;
assign LUT_4[18325] = 32'b00000000000000000001101011100000;
assign LUT_4[18326] = 32'b00000000000000000111111010001100;
assign LUT_4[18327] = 32'b00000000000000000001000110000100;
assign LUT_4[18328] = 32'b00000000000000000100101011100001;
assign LUT_4[18329] = 32'b11111111111111111101110111011001;
assign LUT_4[18330] = 32'b00000000000000000100000110000101;
assign LUT_4[18331] = 32'b11111111111111111101010001111101;
assign LUT_4[18332] = 32'b00000000000000000001101011111101;
assign LUT_4[18333] = 32'b11111111111111111010110111110101;
assign LUT_4[18334] = 32'b00000000000000000001000110100001;
assign LUT_4[18335] = 32'b11111111111111111010010010011001;
assign LUT_4[18336] = 32'b00000000000000001100001000100101;
assign LUT_4[18337] = 32'b00000000000000000101010100011101;
assign LUT_4[18338] = 32'b00000000000000001011100011001001;
assign LUT_4[18339] = 32'b00000000000000000100101111000001;
assign LUT_4[18340] = 32'b00000000000000001001001001000001;
assign LUT_4[18341] = 32'b00000000000000000010010100111001;
assign LUT_4[18342] = 32'b00000000000000001000100011100101;
assign LUT_4[18343] = 32'b00000000000000000001101111011101;
assign LUT_4[18344] = 32'b00000000000000000101010100111010;
assign LUT_4[18345] = 32'b11111111111111111110100000110010;
assign LUT_4[18346] = 32'b00000000000000000100101111011110;
assign LUT_4[18347] = 32'b11111111111111111101111011010110;
assign LUT_4[18348] = 32'b00000000000000000010010101010110;
assign LUT_4[18349] = 32'b11111111111111111011100001001110;
assign LUT_4[18350] = 32'b00000000000000000001101111111010;
assign LUT_4[18351] = 32'b11111111111111111010111011110010;
assign LUT_4[18352] = 32'b00000000000000001001111010010011;
assign LUT_4[18353] = 32'b00000000000000000011000110001011;
assign LUT_4[18354] = 32'b00000000000000001001010100110111;
assign LUT_4[18355] = 32'b00000000000000000010100000101111;
assign LUT_4[18356] = 32'b00000000000000000110111010101111;
assign LUT_4[18357] = 32'b00000000000000000000000110100111;
assign LUT_4[18358] = 32'b00000000000000000110010101010011;
assign LUT_4[18359] = 32'b11111111111111111111100001001011;
assign LUT_4[18360] = 32'b00000000000000000011000110101000;
assign LUT_4[18361] = 32'b11111111111111111100010010100000;
assign LUT_4[18362] = 32'b00000000000000000010100001001100;
assign LUT_4[18363] = 32'b11111111111111111011101101000100;
assign LUT_4[18364] = 32'b00000000000000000000000111000100;
assign LUT_4[18365] = 32'b11111111111111111001010010111100;
assign LUT_4[18366] = 32'b11111111111111111111100001101000;
assign LUT_4[18367] = 32'b11111111111111111000101101100000;
assign LUT_4[18368] = 32'b00000000000000001111000100110010;
assign LUT_4[18369] = 32'b00000000000000001000010000101010;
assign LUT_4[18370] = 32'b00000000000000001110011111010110;
assign LUT_4[18371] = 32'b00000000000000000111101011001110;
assign LUT_4[18372] = 32'b00000000000000001100000101001110;
assign LUT_4[18373] = 32'b00000000000000000101010001000110;
assign LUT_4[18374] = 32'b00000000000000001011011111110010;
assign LUT_4[18375] = 32'b00000000000000000100101011101010;
assign LUT_4[18376] = 32'b00000000000000001000010001000111;
assign LUT_4[18377] = 32'b00000000000000000001011100111111;
assign LUT_4[18378] = 32'b00000000000000000111101011101011;
assign LUT_4[18379] = 32'b00000000000000000000110111100011;
assign LUT_4[18380] = 32'b00000000000000000101010001100011;
assign LUT_4[18381] = 32'b11111111111111111110011101011011;
assign LUT_4[18382] = 32'b00000000000000000100101100000111;
assign LUT_4[18383] = 32'b11111111111111111101110111111111;
assign LUT_4[18384] = 32'b00000000000000001100110110100000;
assign LUT_4[18385] = 32'b00000000000000000110000010011000;
assign LUT_4[18386] = 32'b00000000000000001100010001000100;
assign LUT_4[18387] = 32'b00000000000000000101011100111100;
assign LUT_4[18388] = 32'b00000000000000001001110110111100;
assign LUT_4[18389] = 32'b00000000000000000011000010110100;
assign LUT_4[18390] = 32'b00000000000000001001010001100000;
assign LUT_4[18391] = 32'b00000000000000000010011101011000;
assign LUT_4[18392] = 32'b00000000000000000110000010110101;
assign LUT_4[18393] = 32'b11111111111111111111001110101101;
assign LUT_4[18394] = 32'b00000000000000000101011101011001;
assign LUT_4[18395] = 32'b11111111111111111110101001010001;
assign LUT_4[18396] = 32'b00000000000000000011000011010001;
assign LUT_4[18397] = 32'b11111111111111111100001111001001;
assign LUT_4[18398] = 32'b00000000000000000010011101110101;
assign LUT_4[18399] = 32'b11111111111111111011101001101101;
assign LUT_4[18400] = 32'b00000000000000001101011111111001;
assign LUT_4[18401] = 32'b00000000000000000110101011110001;
assign LUT_4[18402] = 32'b00000000000000001100111010011101;
assign LUT_4[18403] = 32'b00000000000000000110000110010101;
assign LUT_4[18404] = 32'b00000000000000001010100000010101;
assign LUT_4[18405] = 32'b00000000000000000011101100001101;
assign LUT_4[18406] = 32'b00000000000000001001111010111001;
assign LUT_4[18407] = 32'b00000000000000000011000110110001;
assign LUT_4[18408] = 32'b00000000000000000110101100001110;
assign LUT_4[18409] = 32'b11111111111111111111111000000110;
assign LUT_4[18410] = 32'b00000000000000000110000110110010;
assign LUT_4[18411] = 32'b11111111111111111111010010101010;
assign LUT_4[18412] = 32'b00000000000000000011101100101010;
assign LUT_4[18413] = 32'b11111111111111111100111000100010;
assign LUT_4[18414] = 32'b00000000000000000011000111001110;
assign LUT_4[18415] = 32'b11111111111111111100010011000110;
assign LUT_4[18416] = 32'b00000000000000001011010001100111;
assign LUT_4[18417] = 32'b00000000000000000100011101011111;
assign LUT_4[18418] = 32'b00000000000000001010101100001011;
assign LUT_4[18419] = 32'b00000000000000000011111000000011;
assign LUT_4[18420] = 32'b00000000000000001000010010000011;
assign LUT_4[18421] = 32'b00000000000000000001011101111011;
assign LUT_4[18422] = 32'b00000000000000000111101100100111;
assign LUT_4[18423] = 32'b00000000000000000000111000011111;
assign LUT_4[18424] = 32'b00000000000000000100011101111100;
assign LUT_4[18425] = 32'b11111111111111111101101001110100;
assign LUT_4[18426] = 32'b00000000000000000011111000100000;
assign LUT_4[18427] = 32'b11111111111111111101000100011000;
assign LUT_4[18428] = 32'b00000000000000000001011110011000;
assign LUT_4[18429] = 32'b11111111111111111010101010010000;
assign LUT_4[18430] = 32'b00000000000000000000111000111100;
assign LUT_4[18431] = 32'b11111111111111111010000100110100;
assign LUT_4[18432] = 32'b00000000000000000000111100010110;
assign LUT_4[18433] = 32'b11111111111111111010001000001110;
assign LUT_4[18434] = 32'b00000000000000000000010110111010;
assign LUT_4[18435] = 32'b11111111111111111001100010110010;
assign LUT_4[18436] = 32'b11111111111111111101111100110010;
assign LUT_4[18437] = 32'b11111111111111110111001000101010;
assign LUT_4[18438] = 32'b11111111111111111101010111010110;
assign LUT_4[18439] = 32'b11111111111111110110100011001110;
assign LUT_4[18440] = 32'b11111111111111111010001000101011;
assign LUT_4[18441] = 32'b11111111111111110011010100100011;
assign LUT_4[18442] = 32'b11111111111111111001100011001111;
assign LUT_4[18443] = 32'b11111111111111110010101111000111;
assign LUT_4[18444] = 32'b11111111111111110111001001000111;
assign LUT_4[18445] = 32'b11111111111111110000010100111111;
assign LUT_4[18446] = 32'b11111111111111110110100011101011;
assign LUT_4[18447] = 32'b11111111111111101111101111100011;
assign LUT_4[18448] = 32'b11111111111111111110101110000100;
assign LUT_4[18449] = 32'b11111111111111110111111001111100;
assign LUT_4[18450] = 32'b11111111111111111110001000101000;
assign LUT_4[18451] = 32'b11111111111111110111010100100000;
assign LUT_4[18452] = 32'b11111111111111111011101110100000;
assign LUT_4[18453] = 32'b11111111111111110100111010011000;
assign LUT_4[18454] = 32'b11111111111111111011001001000100;
assign LUT_4[18455] = 32'b11111111111111110100010100111100;
assign LUT_4[18456] = 32'b11111111111111110111111010011001;
assign LUT_4[18457] = 32'b11111111111111110001000110010001;
assign LUT_4[18458] = 32'b11111111111111110111010100111101;
assign LUT_4[18459] = 32'b11111111111111110000100000110101;
assign LUT_4[18460] = 32'b11111111111111110100111010110101;
assign LUT_4[18461] = 32'b11111111111111101110000110101101;
assign LUT_4[18462] = 32'b11111111111111110100010101011001;
assign LUT_4[18463] = 32'b11111111111111101101100001010001;
assign LUT_4[18464] = 32'b11111111111111111111010111011101;
assign LUT_4[18465] = 32'b11111111111111111000100011010101;
assign LUT_4[18466] = 32'b11111111111111111110110010000001;
assign LUT_4[18467] = 32'b11111111111111110111111101111001;
assign LUT_4[18468] = 32'b11111111111111111100010111111001;
assign LUT_4[18469] = 32'b11111111111111110101100011110001;
assign LUT_4[18470] = 32'b11111111111111111011110010011101;
assign LUT_4[18471] = 32'b11111111111111110100111110010101;
assign LUT_4[18472] = 32'b11111111111111111000100011110010;
assign LUT_4[18473] = 32'b11111111111111110001101111101010;
assign LUT_4[18474] = 32'b11111111111111110111111110010110;
assign LUT_4[18475] = 32'b11111111111111110001001010001110;
assign LUT_4[18476] = 32'b11111111111111110101100100001110;
assign LUT_4[18477] = 32'b11111111111111101110110000000110;
assign LUT_4[18478] = 32'b11111111111111110100111110110010;
assign LUT_4[18479] = 32'b11111111111111101110001010101010;
assign LUT_4[18480] = 32'b11111111111111111101001001001011;
assign LUT_4[18481] = 32'b11111111111111110110010101000011;
assign LUT_4[18482] = 32'b11111111111111111100100011101111;
assign LUT_4[18483] = 32'b11111111111111110101101111100111;
assign LUT_4[18484] = 32'b11111111111111111010001001100111;
assign LUT_4[18485] = 32'b11111111111111110011010101011111;
assign LUT_4[18486] = 32'b11111111111111111001100100001011;
assign LUT_4[18487] = 32'b11111111111111110010110000000011;
assign LUT_4[18488] = 32'b11111111111111110110010101100000;
assign LUT_4[18489] = 32'b11111111111111101111100001011000;
assign LUT_4[18490] = 32'b11111111111111110101110000000100;
assign LUT_4[18491] = 32'b11111111111111101110111011111100;
assign LUT_4[18492] = 32'b11111111111111110011010101111100;
assign LUT_4[18493] = 32'b11111111111111101100100001110100;
assign LUT_4[18494] = 32'b11111111111111110010110000100000;
assign LUT_4[18495] = 32'b11111111111111101011111100011000;
assign LUT_4[18496] = 32'b00000000000000000010010011101010;
assign LUT_4[18497] = 32'b11111111111111111011011111100010;
assign LUT_4[18498] = 32'b00000000000000000001101110001110;
assign LUT_4[18499] = 32'b11111111111111111010111010000110;
assign LUT_4[18500] = 32'b11111111111111111111010100000110;
assign LUT_4[18501] = 32'b11111111111111111000011111111110;
assign LUT_4[18502] = 32'b11111111111111111110101110101010;
assign LUT_4[18503] = 32'b11111111111111110111111010100010;
assign LUT_4[18504] = 32'b11111111111111111011011111111111;
assign LUT_4[18505] = 32'b11111111111111110100101011110111;
assign LUT_4[18506] = 32'b11111111111111111010111010100011;
assign LUT_4[18507] = 32'b11111111111111110100000110011011;
assign LUT_4[18508] = 32'b11111111111111111000100000011011;
assign LUT_4[18509] = 32'b11111111111111110001101100010011;
assign LUT_4[18510] = 32'b11111111111111110111111010111111;
assign LUT_4[18511] = 32'b11111111111111110001000110110111;
assign LUT_4[18512] = 32'b00000000000000000000000101011000;
assign LUT_4[18513] = 32'b11111111111111111001010001010000;
assign LUT_4[18514] = 32'b11111111111111111111011111111100;
assign LUT_4[18515] = 32'b11111111111111111000101011110100;
assign LUT_4[18516] = 32'b11111111111111111101000101110100;
assign LUT_4[18517] = 32'b11111111111111110110010001101100;
assign LUT_4[18518] = 32'b11111111111111111100100000011000;
assign LUT_4[18519] = 32'b11111111111111110101101100010000;
assign LUT_4[18520] = 32'b11111111111111111001010001101101;
assign LUT_4[18521] = 32'b11111111111111110010011101100101;
assign LUT_4[18522] = 32'b11111111111111111000101100010001;
assign LUT_4[18523] = 32'b11111111111111110001111000001001;
assign LUT_4[18524] = 32'b11111111111111110110010010001001;
assign LUT_4[18525] = 32'b11111111111111101111011110000001;
assign LUT_4[18526] = 32'b11111111111111110101101100101101;
assign LUT_4[18527] = 32'b11111111111111101110111000100101;
assign LUT_4[18528] = 32'b00000000000000000000101110110001;
assign LUT_4[18529] = 32'b11111111111111111001111010101001;
assign LUT_4[18530] = 32'b00000000000000000000001001010101;
assign LUT_4[18531] = 32'b11111111111111111001010101001101;
assign LUT_4[18532] = 32'b11111111111111111101101111001101;
assign LUT_4[18533] = 32'b11111111111111110110111011000101;
assign LUT_4[18534] = 32'b11111111111111111101001001110001;
assign LUT_4[18535] = 32'b11111111111111110110010101101001;
assign LUT_4[18536] = 32'b11111111111111111001111011000110;
assign LUT_4[18537] = 32'b11111111111111110011000110111110;
assign LUT_4[18538] = 32'b11111111111111111001010101101010;
assign LUT_4[18539] = 32'b11111111111111110010100001100010;
assign LUT_4[18540] = 32'b11111111111111110110111011100010;
assign LUT_4[18541] = 32'b11111111111111110000000111011010;
assign LUT_4[18542] = 32'b11111111111111110110010110000110;
assign LUT_4[18543] = 32'b11111111111111101111100001111110;
assign LUT_4[18544] = 32'b11111111111111111110100000011111;
assign LUT_4[18545] = 32'b11111111111111110111101100010111;
assign LUT_4[18546] = 32'b11111111111111111101111011000011;
assign LUT_4[18547] = 32'b11111111111111110111000110111011;
assign LUT_4[18548] = 32'b11111111111111111011100000111011;
assign LUT_4[18549] = 32'b11111111111111110100101100110011;
assign LUT_4[18550] = 32'b11111111111111111010111011011111;
assign LUT_4[18551] = 32'b11111111111111110100000111010111;
assign LUT_4[18552] = 32'b11111111111111110111101100110100;
assign LUT_4[18553] = 32'b11111111111111110000111000101100;
assign LUT_4[18554] = 32'b11111111111111110111000111011000;
assign LUT_4[18555] = 32'b11111111111111110000010011010000;
assign LUT_4[18556] = 32'b11111111111111110100101101010000;
assign LUT_4[18557] = 32'b11111111111111101101111001001000;
assign LUT_4[18558] = 32'b11111111111111110100000111110100;
assign LUT_4[18559] = 32'b11111111111111101101010011101100;
assign LUT_4[18560] = 32'b00000000000000000011100010011110;
assign LUT_4[18561] = 32'b11111111111111111100101110010110;
assign LUT_4[18562] = 32'b00000000000000000010111101000010;
assign LUT_4[18563] = 32'b11111111111111111100001000111010;
assign LUT_4[18564] = 32'b00000000000000000000100010111010;
assign LUT_4[18565] = 32'b11111111111111111001101110110010;
assign LUT_4[18566] = 32'b11111111111111111111111101011110;
assign LUT_4[18567] = 32'b11111111111111111001001001010110;
assign LUT_4[18568] = 32'b11111111111111111100101110110011;
assign LUT_4[18569] = 32'b11111111111111110101111010101011;
assign LUT_4[18570] = 32'b11111111111111111100001001010111;
assign LUT_4[18571] = 32'b11111111111111110101010101001111;
assign LUT_4[18572] = 32'b11111111111111111001101111001111;
assign LUT_4[18573] = 32'b11111111111111110010111011000111;
assign LUT_4[18574] = 32'b11111111111111111001001001110011;
assign LUT_4[18575] = 32'b11111111111111110010010101101011;
assign LUT_4[18576] = 32'b00000000000000000001010100001100;
assign LUT_4[18577] = 32'b11111111111111111010100000000100;
assign LUT_4[18578] = 32'b00000000000000000000101110110000;
assign LUT_4[18579] = 32'b11111111111111111001111010101000;
assign LUT_4[18580] = 32'b11111111111111111110010100101000;
assign LUT_4[18581] = 32'b11111111111111110111100000100000;
assign LUT_4[18582] = 32'b11111111111111111101101111001100;
assign LUT_4[18583] = 32'b11111111111111110110111011000100;
assign LUT_4[18584] = 32'b11111111111111111010100000100001;
assign LUT_4[18585] = 32'b11111111111111110011101100011001;
assign LUT_4[18586] = 32'b11111111111111111001111011000101;
assign LUT_4[18587] = 32'b11111111111111110011000110111101;
assign LUT_4[18588] = 32'b11111111111111110111100000111101;
assign LUT_4[18589] = 32'b11111111111111110000101100110101;
assign LUT_4[18590] = 32'b11111111111111110110111011100001;
assign LUT_4[18591] = 32'b11111111111111110000000111011001;
assign LUT_4[18592] = 32'b00000000000000000001111101100101;
assign LUT_4[18593] = 32'b11111111111111111011001001011101;
assign LUT_4[18594] = 32'b00000000000000000001011000001001;
assign LUT_4[18595] = 32'b11111111111111111010100100000001;
assign LUT_4[18596] = 32'b11111111111111111110111110000001;
assign LUT_4[18597] = 32'b11111111111111111000001001111001;
assign LUT_4[18598] = 32'b11111111111111111110011000100101;
assign LUT_4[18599] = 32'b11111111111111110111100100011101;
assign LUT_4[18600] = 32'b11111111111111111011001001111010;
assign LUT_4[18601] = 32'b11111111111111110100010101110010;
assign LUT_4[18602] = 32'b11111111111111111010100100011110;
assign LUT_4[18603] = 32'b11111111111111110011110000010110;
assign LUT_4[18604] = 32'b11111111111111111000001010010110;
assign LUT_4[18605] = 32'b11111111111111110001010110001110;
assign LUT_4[18606] = 32'b11111111111111110111100100111010;
assign LUT_4[18607] = 32'b11111111111111110000110000110010;
assign LUT_4[18608] = 32'b11111111111111111111101111010011;
assign LUT_4[18609] = 32'b11111111111111111000111011001011;
assign LUT_4[18610] = 32'b11111111111111111111001001110111;
assign LUT_4[18611] = 32'b11111111111111111000010101101111;
assign LUT_4[18612] = 32'b11111111111111111100101111101111;
assign LUT_4[18613] = 32'b11111111111111110101111011100111;
assign LUT_4[18614] = 32'b11111111111111111100001010010011;
assign LUT_4[18615] = 32'b11111111111111110101010110001011;
assign LUT_4[18616] = 32'b11111111111111111000111011101000;
assign LUT_4[18617] = 32'b11111111111111110010000111100000;
assign LUT_4[18618] = 32'b11111111111111111000010110001100;
assign LUT_4[18619] = 32'b11111111111111110001100010000100;
assign LUT_4[18620] = 32'b11111111111111110101111100000100;
assign LUT_4[18621] = 32'b11111111111111101111000111111100;
assign LUT_4[18622] = 32'b11111111111111110101010110101000;
assign LUT_4[18623] = 32'b11111111111111101110100010100000;
assign LUT_4[18624] = 32'b00000000000000000100111001110010;
assign LUT_4[18625] = 32'b11111111111111111110000101101010;
assign LUT_4[18626] = 32'b00000000000000000100010100010110;
assign LUT_4[18627] = 32'b11111111111111111101100000001110;
assign LUT_4[18628] = 32'b00000000000000000001111010001110;
assign LUT_4[18629] = 32'b11111111111111111011000110000110;
assign LUT_4[18630] = 32'b00000000000000000001010100110010;
assign LUT_4[18631] = 32'b11111111111111111010100000101010;
assign LUT_4[18632] = 32'b11111111111111111110000110000111;
assign LUT_4[18633] = 32'b11111111111111110111010001111111;
assign LUT_4[18634] = 32'b11111111111111111101100000101011;
assign LUT_4[18635] = 32'b11111111111111110110101100100011;
assign LUT_4[18636] = 32'b11111111111111111011000110100011;
assign LUT_4[18637] = 32'b11111111111111110100010010011011;
assign LUT_4[18638] = 32'b11111111111111111010100001000111;
assign LUT_4[18639] = 32'b11111111111111110011101100111111;
assign LUT_4[18640] = 32'b00000000000000000010101011100000;
assign LUT_4[18641] = 32'b11111111111111111011110111011000;
assign LUT_4[18642] = 32'b00000000000000000010000110000100;
assign LUT_4[18643] = 32'b11111111111111111011010001111100;
assign LUT_4[18644] = 32'b11111111111111111111101011111100;
assign LUT_4[18645] = 32'b11111111111111111000110111110100;
assign LUT_4[18646] = 32'b11111111111111111111000110100000;
assign LUT_4[18647] = 32'b11111111111111111000010010011000;
assign LUT_4[18648] = 32'b11111111111111111011110111110101;
assign LUT_4[18649] = 32'b11111111111111110101000011101101;
assign LUT_4[18650] = 32'b11111111111111111011010010011001;
assign LUT_4[18651] = 32'b11111111111111110100011110010001;
assign LUT_4[18652] = 32'b11111111111111111000111000010001;
assign LUT_4[18653] = 32'b11111111111111110010000100001001;
assign LUT_4[18654] = 32'b11111111111111111000010010110101;
assign LUT_4[18655] = 32'b11111111111111110001011110101101;
assign LUT_4[18656] = 32'b00000000000000000011010100111001;
assign LUT_4[18657] = 32'b11111111111111111100100000110001;
assign LUT_4[18658] = 32'b00000000000000000010101111011101;
assign LUT_4[18659] = 32'b11111111111111111011111011010101;
assign LUT_4[18660] = 32'b00000000000000000000010101010101;
assign LUT_4[18661] = 32'b11111111111111111001100001001101;
assign LUT_4[18662] = 32'b11111111111111111111101111111001;
assign LUT_4[18663] = 32'b11111111111111111000111011110001;
assign LUT_4[18664] = 32'b11111111111111111100100001001110;
assign LUT_4[18665] = 32'b11111111111111110101101101000110;
assign LUT_4[18666] = 32'b11111111111111111011111011110010;
assign LUT_4[18667] = 32'b11111111111111110101000111101010;
assign LUT_4[18668] = 32'b11111111111111111001100001101010;
assign LUT_4[18669] = 32'b11111111111111110010101101100010;
assign LUT_4[18670] = 32'b11111111111111111000111100001110;
assign LUT_4[18671] = 32'b11111111111111110010001000000110;
assign LUT_4[18672] = 32'b00000000000000000001000110100111;
assign LUT_4[18673] = 32'b11111111111111111010010010011111;
assign LUT_4[18674] = 32'b00000000000000000000100001001011;
assign LUT_4[18675] = 32'b11111111111111111001101101000011;
assign LUT_4[18676] = 32'b11111111111111111110000111000011;
assign LUT_4[18677] = 32'b11111111111111110111010010111011;
assign LUT_4[18678] = 32'b11111111111111111101100001100111;
assign LUT_4[18679] = 32'b11111111111111110110101101011111;
assign LUT_4[18680] = 32'b11111111111111111010010010111100;
assign LUT_4[18681] = 32'b11111111111111110011011110110100;
assign LUT_4[18682] = 32'b11111111111111111001101101100000;
assign LUT_4[18683] = 32'b11111111111111110010111001011000;
assign LUT_4[18684] = 32'b11111111111111110111010011011000;
assign LUT_4[18685] = 32'b11111111111111110000011111010000;
assign LUT_4[18686] = 32'b11111111111111110110101101111100;
assign LUT_4[18687] = 32'b11111111111111101111111001110100;
assign LUT_4[18688] = 32'b00000000000000000101110111111001;
assign LUT_4[18689] = 32'b11111111111111111111000011110001;
assign LUT_4[18690] = 32'b00000000000000000101010010011101;
assign LUT_4[18691] = 32'b11111111111111111110011110010101;
assign LUT_4[18692] = 32'b00000000000000000010111000010101;
assign LUT_4[18693] = 32'b11111111111111111100000100001101;
assign LUT_4[18694] = 32'b00000000000000000010010010111001;
assign LUT_4[18695] = 32'b11111111111111111011011110110001;
assign LUT_4[18696] = 32'b11111111111111111111000100001110;
assign LUT_4[18697] = 32'b11111111111111111000010000000110;
assign LUT_4[18698] = 32'b11111111111111111110011110110010;
assign LUT_4[18699] = 32'b11111111111111110111101010101010;
assign LUT_4[18700] = 32'b11111111111111111100000100101010;
assign LUT_4[18701] = 32'b11111111111111110101010000100010;
assign LUT_4[18702] = 32'b11111111111111111011011111001110;
assign LUT_4[18703] = 32'b11111111111111110100101011000110;
assign LUT_4[18704] = 32'b00000000000000000011101001100111;
assign LUT_4[18705] = 32'b11111111111111111100110101011111;
assign LUT_4[18706] = 32'b00000000000000000011000100001011;
assign LUT_4[18707] = 32'b11111111111111111100010000000011;
assign LUT_4[18708] = 32'b00000000000000000000101010000011;
assign LUT_4[18709] = 32'b11111111111111111001110101111011;
assign LUT_4[18710] = 32'b00000000000000000000000100100111;
assign LUT_4[18711] = 32'b11111111111111111001010000011111;
assign LUT_4[18712] = 32'b11111111111111111100110101111100;
assign LUT_4[18713] = 32'b11111111111111110110000001110100;
assign LUT_4[18714] = 32'b11111111111111111100010000100000;
assign LUT_4[18715] = 32'b11111111111111110101011100011000;
assign LUT_4[18716] = 32'b11111111111111111001110110011000;
assign LUT_4[18717] = 32'b11111111111111110011000010010000;
assign LUT_4[18718] = 32'b11111111111111111001010000111100;
assign LUT_4[18719] = 32'b11111111111111110010011100110100;
assign LUT_4[18720] = 32'b00000000000000000100010011000000;
assign LUT_4[18721] = 32'b11111111111111111101011110111000;
assign LUT_4[18722] = 32'b00000000000000000011101101100100;
assign LUT_4[18723] = 32'b11111111111111111100111001011100;
assign LUT_4[18724] = 32'b00000000000000000001010011011100;
assign LUT_4[18725] = 32'b11111111111111111010011111010100;
assign LUT_4[18726] = 32'b00000000000000000000101110000000;
assign LUT_4[18727] = 32'b11111111111111111001111001111000;
assign LUT_4[18728] = 32'b11111111111111111101011111010101;
assign LUT_4[18729] = 32'b11111111111111110110101011001101;
assign LUT_4[18730] = 32'b11111111111111111100111001111001;
assign LUT_4[18731] = 32'b11111111111111110110000101110001;
assign LUT_4[18732] = 32'b11111111111111111010011111110001;
assign LUT_4[18733] = 32'b11111111111111110011101011101001;
assign LUT_4[18734] = 32'b11111111111111111001111010010101;
assign LUT_4[18735] = 32'b11111111111111110011000110001101;
assign LUT_4[18736] = 32'b00000000000000000010000100101110;
assign LUT_4[18737] = 32'b11111111111111111011010000100110;
assign LUT_4[18738] = 32'b00000000000000000001011111010010;
assign LUT_4[18739] = 32'b11111111111111111010101011001010;
assign LUT_4[18740] = 32'b11111111111111111111000101001010;
assign LUT_4[18741] = 32'b11111111111111111000010001000010;
assign LUT_4[18742] = 32'b11111111111111111110011111101110;
assign LUT_4[18743] = 32'b11111111111111110111101011100110;
assign LUT_4[18744] = 32'b11111111111111111011010001000011;
assign LUT_4[18745] = 32'b11111111111111110100011100111011;
assign LUT_4[18746] = 32'b11111111111111111010101011100111;
assign LUT_4[18747] = 32'b11111111111111110011110111011111;
assign LUT_4[18748] = 32'b11111111111111111000010001011111;
assign LUT_4[18749] = 32'b11111111111111110001011101010111;
assign LUT_4[18750] = 32'b11111111111111110111101100000011;
assign LUT_4[18751] = 32'b11111111111111110000110111111011;
assign LUT_4[18752] = 32'b00000000000000000111001111001101;
assign LUT_4[18753] = 32'b00000000000000000000011011000101;
assign LUT_4[18754] = 32'b00000000000000000110101001110001;
assign LUT_4[18755] = 32'b11111111111111111111110101101001;
assign LUT_4[18756] = 32'b00000000000000000100001111101001;
assign LUT_4[18757] = 32'b11111111111111111101011011100001;
assign LUT_4[18758] = 32'b00000000000000000011101010001101;
assign LUT_4[18759] = 32'b11111111111111111100110110000101;
assign LUT_4[18760] = 32'b00000000000000000000011011100010;
assign LUT_4[18761] = 32'b11111111111111111001100111011010;
assign LUT_4[18762] = 32'b11111111111111111111110110000110;
assign LUT_4[18763] = 32'b11111111111111111001000001111110;
assign LUT_4[18764] = 32'b11111111111111111101011011111110;
assign LUT_4[18765] = 32'b11111111111111110110100111110110;
assign LUT_4[18766] = 32'b11111111111111111100110110100010;
assign LUT_4[18767] = 32'b11111111111111110110000010011010;
assign LUT_4[18768] = 32'b00000000000000000101000000111011;
assign LUT_4[18769] = 32'b11111111111111111110001100110011;
assign LUT_4[18770] = 32'b00000000000000000100011011011111;
assign LUT_4[18771] = 32'b11111111111111111101100111010111;
assign LUT_4[18772] = 32'b00000000000000000010000001010111;
assign LUT_4[18773] = 32'b11111111111111111011001101001111;
assign LUT_4[18774] = 32'b00000000000000000001011011111011;
assign LUT_4[18775] = 32'b11111111111111111010100111110011;
assign LUT_4[18776] = 32'b11111111111111111110001101010000;
assign LUT_4[18777] = 32'b11111111111111110111011001001000;
assign LUT_4[18778] = 32'b11111111111111111101100111110100;
assign LUT_4[18779] = 32'b11111111111111110110110011101100;
assign LUT_4[18780] = 32'b11111111111111111011001101101100;
assign LUT_4[18781] = 32'b11111111111111110100011001100100;
assign LUT_4[18782] = 32'b11111111111111111010101000010000;
assign LUT_4[18783] = 32'b11111111111111110011110100001000;
assign LUT_4[18784] = 32'b00000000000000000101101010010100;
assign LUT_4[18785] = 32'b11111111111111111110110110001100;
assign LUT_4[18786] = 32'b00000000000000000101000100111000;
assign LUT_4[18787] = 32'b11111111111111111110010000110000;
assign LUT_4[18788] = 32'b00000000000000000010101010110000;
assign LUT_4[18789] = 32'b11111111111111111011110110101000;
assign LUT_4[18790] = 32'b00000000000000000010000101010100;
assign LUT_4[18791] = 32'b11111111111111111011010001001100;
assign LUT_4[18792] = 32'b11111111111111111110110110101001;
assign LUT_4[18793] = 32'b11111111111111111000000010100001;
assign LUT_4[18794] = 32'b11111111111111111110010001001101;
assign LUT_4[18795] = 32'b11111111111111110111011101000101;
assign LUT_4[18796] = 32'b11111111111111111011110111000101;
assign LUT_4[18797] = 32'b11111111111111110101000010111101;
assign LUT_4[18798] = 32'b11111111111111111011010001101001;
assign LUT_4[18799] = 32'b11111111111111110100011101100001;
assign LUT_4[18800] = 32'b00000000000000000011011100000010;
assign LUT_4[18801] = 32'b11111111111111111100100111111010;
assign LUT_4[18802] = 32'b00000000000000000010110110100110;
assign LUT_4[18803] = 32'b11111111111111111100000010011110;
assign LUT_4[18804] = 32'b00000000000000000000011100011110;
assign LUT_4[18805] = 32'b11111111111111111001101000010110;
assign LUT_4[18806] = 32'b11111111111111111111110111000010;
assign LUT_4[18807] = 32'b11111111111111111001000010111010;
assign LUT_4[18808] = 32'b11111111111111111100101000010111;
assign LUT_4[18809] = 32'b11111111111111110101110100001111;
assign LUT_4[18810] = 32'b11111111111111111100000010111011;
assign LUT_4[18811] = 32'b11111111111111110101001110110011;
assign LUT_4[18812] = 32'b11111111111111111001101000110011;
assign LUT_4[18813] = 32'b11111111111111110010110100101011;
assign LUT_4[18814] = 32'b11111111111111111001000011010111;
assign LUT_4[18815] = 32'b11111111111111110010001111001111;
assign LUT_4[18816] = 32'b00000000000000001000011110000001;
assign LUT_4[18817] = 32'b00000000000000000001101001111001;
assign LUT_4[18818] = 32'b00000000000000000111111000100101;
assign LUT_4[18819] = 32'b00000000000000000001000100011101;
assign LUT_4[18820] = 32'b00000000000000000101011110011101;
assign LUT_4[18821] = 32'b11111111111111111110101010010101;
assign LUT_4[18822] = 32'b00000000000000000100111001000001;
assign LUT_4[18823] = 32'b11111111111111111110000100111001;
assign LUT_4[18824] = 32'b00000000000000000001101010010110;
assign LUT_4[18825] = 32'b11111111111111111010110110001110;
assign LUT_4[18826] = 32'b00000000000000000001000100111010;
assign LUT_4[18827] = 32'b11111111111111111010010000110010;
assign LUT_4[18828] = 32'b11111111111111111110101010110010;
assign LUT_4[18829] = 32'b11111111111111110111110110101010;
assign LUT_4[18830] = 32'b11111111111111111110000101010110;
assign LUT_4[18831] = 32'b11111111111111110111010001001110;
assign LUT_4[18832] = 32'b00000000000000000110001111101111;
assign LUT_4[18833] = 32'b11111111111111111111011011100111;
assign LUT_4[18834] = 32'b00000000000000000101101010010011;
assign LUT_4[18835] = 32'b11111111111111111110110110001011;
assign LUT_4[18836] = 32'b00000000000000000011010000001011;
assign LUT_4[18837] = 32'b11111111111111111100011100000011;
assign LUT_4[18838] = 32'b00000000000000000010101010101111;
assign LUT_4[18839] = 32'b11111111111111111011110110100111;
assign LUT_4[18840] = 32'b11111111111111111111011100000100;
assign LUT_4[18841] = 32'b11111111111111111000100111111100;
assign LUT_4[18842] = 32'b11111111111111111110110110101000;
assign LUT_4[18843] = 32'b11111111111111111000000010100000;
assign LUT_4[18844] = 32'b11111111111111111100011100100000;
assign LUT_4[18845] = 32'b11111111111111110101101000011000;
assign LUT_4[18846] = 32'b11111111111111111011110111000100;
assign LUT_4[18847] = 32'b11111111111111110101000010111100;
assign LUT_4[18848] = 32'b00000000000000000110111001001000;
assign LUT_4[18849] = 32'b00000000000000000000000101000000;
assign LUT_4[18850] = 32'b00000000000000000110010011101100;
assign LUT_4[18851] = 32'b11111111111111111111011111100100;
assign LUT_4[18852] = 32'b00000000000000000011111001100100;
assign LUT_4[18853] = 32'b11111111111111111101000101011100;
assign LUT_4[18854] = 32'b00000000000000000011010100001000;
assign LUT_4[18855] = 32'b11111111111111111100100000000000;
assign LUT_4[18856] = 32'b00000000000000000000000101011101;
assign LUT_4[18857] = 32'b11111111111111111001010001010101;
assign LUT_4[18858] = 32'b11111111111111111111100000000001;
assign LUT_4[18859] = 32'b11111111111111111000101011111001;
assign LUT_4[18860] = 32'b11111111111111111101000101111001;
assign LUT_4[18861] = 32'b11111111111111110110010001110001;
assign LUT_4[18862] = 32'b11111111111111111100100000011101;
assign LUT_4[18863] = 32'b11111111111111110101101100010101;
assign LUT_4[18864] = 32'b00000000000000000100101010110110;
assign LUT_4[18865] = 32'b11111111111111111101110110101110;
assign LUT_4[18866] = 32'b00000000000000000100000101011010;
assign LUT_4[18867] = 32'b11111111111111111101010001010010;
assign LUT_4[18868] = 32'b00000000000000000001101011010010;
assign LUT_4[18869] = 32'b11111111111111111010110111001010;
assign LUT_4[18870] = 32'b00000000000000000001000101110110;
assign LUT_4[18871] = 32'b11111111111111111010010001101110;
assign LUT_4[18872] = 32'b11111111111111111101110111001011;
assign LUT_4[18873] = 32'b11111111111111110111000011000011;
assign LUT_4[18874] = 32'b11111111111111111101010001101111;
assign LUT_4[18875] = 32'b11111111111111110110011101100111;
assign LUT_4[18876] = 32'b11111111111111111010110111100111;
assign LUT_4[18877] = 32'b11111111111111110100000011011111;
assign LUT_4[18878] = 32'b11111111111111111010010010001011;
assign LUT_4[18879] = 32'b11111111111111110011011110000011;
assign LUT_4[18880] = 32'b00000000000000001001110101010101;
assign LUT_4[18881] = 32'b00000000000000000011000001001101;
assign LUT_4[18882] = 32'b00000000000000001001001111111001;
assign LUT_4[18883] = 32'b00000000000000000010011011110001;
assign LUT_4[18884] = 32'b00000000000000000110110101110001;
assign LUT_4[18885] = 32'b00000000000000000000000001101001;
assign LUT_4[18886] = 32'b00000000000000000110010000010101;
assign LUT_4[18887] = 32'b11111111111111111111011100001101;
assign LUT_4[18888] = 32'b00000000000000000011000001101010;
assign LUT_4[18889] = 32'b11111111111111111100001101100010;
assign LUT_4[18890] = 32'b00000000000000000010011100001110;
assign LUT_4[18891] = 32'b11111111111111111011101000000110;
assign LUT_4[18892] = 32'b00000000000000000000000010000110;
assign LUT_4[18893] = 32'b11111111111111111001001101111110;
assign LUT_4[18894] = 32'b11111111111111111111011100101010;
assign LUT_4[18895] = 32'b11111111111111111000101000100010;
assign LUT_4[18896] = 32'b00000000000000000111100111000011;
assign LUT_4[18897] = 32'b00000000000000000000110010111011;
assign LUT_4[18898] = 32'b00000000000000000111000001100111;
assign LUT_4[18899] = 32'b00000000000000000000001101011111;
assign LUT_4[18900] = 32'b00000000000000000100100111011111;
assign LUT_4[18901] = 32'b11111111111111111101110011010111;
assign LUT_4[18902] = 32'b00000000000000000100000010000011;
assign LUT_4[18903] = 32'b11111111111111111101001101111011;
assign LUT_4[18904] = 32'b00000000000000000000110011011000;
assign LUT_4[18905] = 32'b11111111111111111001111111010000;
assign LUT_4[18906] = 32'b00000000000000000000001101111100;
assign LUT_4[18907] = 32'b11111111111111111001011001110100;
assign LUT_4[18908] = 32'b11111111111111111101110011110100;
assign LUT_4[18909] = 32'b11111111111111110110111111101100;
assign LUT_4[18910] = 32'b11111111111111111101001110011000;
assign LUT_4[18911] = 32'b11111111111111110110011010010000;
assign LUT_4[18912] = 32'b00000000000000001000010000011100;
assign LUT_4[18913] = 32'b00000000000000000001011100010100;
assign LUT_4[18914] = 32'b00000000000000000111101011000000;
assign LUT_4[18915] = 32'b00000000000000000000110110111000;
assign LUT_4[18916] = 32'b00000000000000000101010000111000;
assign LUT_4[18917] = 32'b11111111111111111110011100110000;
assign LUT_4[18918] = 32'b00000000000000000100101011011100;
assign LUT_4[18919] = 32'b11111111111111111101110111010100;
assign LUT_4[18920] = 32'b00000000000000000001011100110001;
assign LUT_4[18921] = 32'b11111111111111111010101000101001;
assign LUT_4[18922] = 32'b00000000000000000000110111010101;
assign LUT_4[18923] = 32'b11111111111111111010000011001101;
assign LUT_4[18924] = 32'b11111111111111111110011101001101;
assign LUT_4[18925] = 32'b11111111111111110111101001000101;
assign LUT_4[18926] = 32'b11111111111111111101110111110001;
assign LUT_4[18927] = 32'b11111111111111110111000011101001;
assign LUT_4[18928] = 32'b00000000000000000110000010001010;
assign LUT_4[18929] = 32'b11111111111111111111001110000010;
assign LUT_4[18930] = 32'b00000000000000000101011100101110;
assign LUT_4[18931] = 32'b11111111111111111110101000100110;
assign LUT_4[18932] = 32'b00000000000000000011000010100110;
assign LUT_4[18933] = 32'b11111111111111111100001110011110;
assign LUT_4[18934] = 32'b00000000000000000010011101001010;
assign LUT_4[18935] = 32'b11111111111111111011101001000010;
assign LUT_4[18936] = 32'b11111111111111111111001110011111;
assign LUT_4[18937] = 32'b11111111111111111000011010010111;
assign LUT_4[18938] = 32'b11111111111111111110101001000011;
assign LUT_4[18939] = 32'b11111111111111110111110100111011;
assign LUT_4[18940] = 32'b11111111111111111100001110111011;
assign LUT_4[18941] = 32'b11111111111111110101011010110011;
assign LUT_4[18942] = 32'b11111111111111111011101001011111;
assign LUT_4[18943] = 32'b11111111111111110100110101010111;
assign LUT_4[18944] = 32'b00000000000000000000000000011110;
assign LUT_4[18945] = 32'b11111111111111111001001100010110;
assign LUT_4[18946] = 32'b11111111111111111111011011000010;
assign LUT_4[18947] = 32'b11111111111111111000100110111010;
assign LUT_4[18948] = 32'b11111111111111111101000000111010;
assign LUT_4[18949] = 32'b11111111111111110110001100110010;
assign LUT_4[18950] = 32'b11111111111111111100011011011110;
assign LUT_4[18951] = 32'b11111111111111110101100111010110;
assign LUT_4[18952] = 32'b11111111111111111001001100110011;
assign LUT_4[18953] = 32'b11111111111111110010011000101011;
assign LUT_4[18954] = 32'b11111111111111111000100111010111;
assign LUT_4[18955] = 32'b11111111111111110001110011001111;
assign LUT_4[18956] = 32'b11111111111111110110001101001111;
assign LUT_4[18957] = 32'b11111111111111101111011001000111;
assign LUT_4[18958] = 32'b11111111111111110101100111110011;
assign LUT_4[18959] = 32'b11111111111111101110110011101011;
assign LUT_4[18960] = 32'b11111111111111111101110010001100;
assign LUT_4[18961] = 32'b11111111111111110110111110000100;
assign LUT_4[18962] = 32'b11111111111111111101001100110000;
assign LUT_4[18963] = 32'b11111111111111110110011000101000;
assign LUT_4[18964] = 32'b11111111111111111010110010101000;
assign LUT_4[18965] = 32'b11111111111111110011111110100000;
assign LUT_4[18966] = 32'b11111111111111111010001101001100;
assign LUT_4[18967] = 32'b11111111111111110011011001000100;
assign LUT_4[18968] = 32'b11111111111111110110111110100001;
assign LUT_4[18969] = 32'b11111111111111110000001010011001;
assign LUT_4[18970] = 32'b11111111111111110110011001000101;
assign LUT_4[18971] = 32'b11111111111111101111100100111101;
assign LUT_4[18972] = 32'b11111111111111110011111110111101;
assign LUT_4[18973] = 32'b11111111111111101101001010110101;
assign LUT_4[18974] = 32'b11111111111111110011011001100001;
assign LUT_4[18975] = 32'b11111111111111101100100101011001;
assign LUT_4[18976] = 32'b11111111111111111110011011100101;
assign LUT_4[18977] = 32'b11111111111111110111100111011101;
assign LUT_4[18978] = 32'b11111111111111111101110110001001;
assign LUT_4[18979] = 32'b11111111111111110111000010000001;
assign LUT_4[18980] = 32'b11111111111111111011011100000001;
assign LUT_4[18981] = 32'b11111111111111110100100111111001;
assign LUT_4[18982] = 32'b11111111111111111010110110100101;
assign LUT_4[18983] = 32'b11111111111111110100000010011101;
assign LUT_4[18984] = 32'b11111111111111110111100111111010;
assign LUT_4[18985] = 32'b11111111111111110000110011110010;
assign LUT_4[18986] = 32'b11111111111111110111000010011110;
assign LUT_4[18987] = 32'b11111111111111110000001110010110;
assign LUT_4[18988] = 32'b11111111111111110100101000010110;
assign LUT_4[18989] = 32'b11111111111111101101110100001110;
assign LUT_4[18990] = 32'b11111111111111110100000010111010;
assign LUT_4[18991] = 32'b11111111111111101101001110110010;
assign LUT_4[18992] = 32'b11111111111111111100001101010011;
assign LUT_4[18993] = 32'b11111111111111110101011001001011;
assign LUT_4[18994] = 32'b11111111111111111011100111110111;
assign LUT_4[18995] = 32'b11111111111111110100110011101111;
assign LUT_4[18996] = 32'b11111111111111111001001101101111;
assign LUT_4[18997] = 32'b11111111111111110010011001100111;
assign LUT_4[18998] = 32'b11111111111111111000101000010011;
assign LUT_4[18999] = 32'b11111111111111110001110100001011;
assign LUT_4[19000] = 32'b11111111111111110101011001101000;
assign LUT_4[19001] = 32'b11111111111111101110100101100000;
assign LUT_4[19002] = 32'b11111111111111110100110100001100;
assign LUT_4[19003] = 32'b11111111111111101110000000000100;
assign LUT_4[19004] = 32'b11111111111111110010011010000100;
assign LUT_4[19005] = 32'b11111111111111101011100101111100;
assign LUT_4[19006] = 32'b11111111111111110001110100101000;
assign LUT_4[19007] = 32'b11111111111111101011000000100000;
assign LUT_4[19008] = 32'b00000000000000000001010111110010;
assign LUT_4[19009] = 32'b11111111111111111010100011101010;
assign LUT_4[19010] = 32'b00000000000000000000110010010110;
assign LUT_4[19011] = 32'b11111111111111111001111110001110;
assign LUT_4[19012] = 32'b11111111111111111110011000001110;
assign LUT_4[19013] = 32'b11111111111111110111100100000110;
assign LUT_4[19014] = 32'b11111111111111111101110010110010;
assign LUT_4[19015] = 32'b11111111111111110110111110101010;
assign LUT_4[19016] = 32'b11111111111111111010100100000111;
assign LUT_4[19017] = 32'b11111111111111110011101111111111;
assign LUT_4[19018] = 32'b11111111111111111001111110101011;
assign LUT_4[19019] = 32'b11111111111111110011001010100011;
assign LUT_4[19020] = 32'b11111111111111110111100100100011;
assign LUT_4[19021] = 32'b11111111111111110000110000011011;
assign LUT_4[19022] = 32'b11111111111111110110111111000111;
assign LUT_4[19023] = 32'b11111111111111110000001010111111;
assign LUT_4[19024] = 32'b11111111111111111111001001100000;
assign LUT_4[19025] = 32'b11111111111111111000010101011000;
assign LUT_4[19026] = 32'b11111111111111111110100100000100;
assign LUT_4[19027] = 32'b11111111111111110111101111111100;
assign LUT_4[19028] = 32'b11111111111111111100001001111100;
assign LUT_4[19029] = 32'b11111111111111110101010101110100;
assign LUT_4[19030] = 32'b11111111111111111011100100100000;
assign LUT_4[19031] = 32'b11111111111111110100110000011000;
assign LUT_4[19032] = 32'b11111111111111111000010101110101;
assign LUT_4[19033] = 32'b11111111111111110001100001101101;
assign LUT_4[19034] = 32'b11111111111111110111110000011001;
assign LUT_4[19035] = 32'b11111111111111110000111100010001;
assign LUT_4[19036] = 32'b11111111111111110101010110010001;
assign LUT_4[19037] = 32'b11111111111111101110100010001001;
assign LUT_4[19038] = 32'b11111111111111110100110000110101;
assign LUT_4[19039] = 32'b11111111111111101101111100101101;
assign LUT_4[19040] = 32'b11111111111111111111110010111001;
assign LUT_4[19041] = 32'b11111111111111111000111110110001;
assign LUT_4[19042] = 32'b11111111111111111111001101011101;
assign LUT_4[19043] = 32'b11111111111111111000011001010101;
assign LUT_4[19044] = 32'b11111111111111111100110011010101;
assign LUT_4[19045] = 32'b11111111111111110101111111001101;
assign LUT_4[19046] = 32'b11111111111111111100001101111001;
assign LUT_4[19047] = 32'b11111111111111110101011001110001;
assign LUT_4[19048] = 32'b11111111111111111000111111001110;
assign LUT_4[19049] = 32'b11111111111111110010001011000110;
assign LUT_4[19050] = 32'b11111111111111111000011001110010;
assign LUT_4[19051] = 32'b11111111111111110001100101101010;
assign LUT_4[19052] = 32'b11111111111111110101111111101010;
assign LUT_4[19053] = 32'b11111111111111101111001011100010;
assign LUT_4[19054] = 32'b11111111111111110101011010001110;
assign LUT_4[19055] = 32'b11111111111111101110100110000110;
assign LUT_4[19056] = 32'b11111111111111111101100100100111;
assign LUT_4[19057] = 32'b11111111111111110110110000011111;
assign LUT_4[19058] = 32'b11111111111111111100111111001011;
assign LUT_4[19059] = 32'b11111111111111110110001011000011;
assign LUT_4[19060] = 32'b11111111111111111010100101000011;
assign LUT_4[19061] = 32'b11111111111111110011110000111011;
assign LUT_4[19062] = 32'b11111111111111111001111111100111;
assign LUT_4[19063] = 32'b11111111111111110011001011011111;
assign LUT_4[19064] = 32'b11111111111111110110110000111100;
assign LUT_4[19065] = 32'b11111111111111101111111100110100;
assign LUT_4[19066] = 32'b11111111111111110110001011100000;
assign LUT_4[19067] = 32'b11111111111111101111010111011000;
assign LUT_4[19068] = 32'b11111111111111110011110001011000;
assign LUT_4[19069] = 32'b11111111111111101100111101010000;
assign LUT_4[19070] = 32'b11111111111111110011001011111100;
assign LUT_4[19071] = 32'b11111111111111101100010111110100;
assign LUT_4[19072] = 32'b00000000000000000010100110100110;
assign LUT_4[19073] = 32'b11111111111111111011110010011110;
assign LUT_4[19074] = 32'b00000000000000000010000001001010;
assign LUT_4[19075] = 32'b11111111111111111011001101000010;
assign LUT_4[19076] = 32'b11111111111111111111100111000010;
assign LUT_4[19077] = 32'b11111111111111111000110010111010;
assign LUT_4[19078] = 32'b11111111111111111111000001100110;
assign LUT_4[19079] = 32'b11111111111111111000001101011110;
assign LUT_4[19080] = 32'b11111111111111111011110010111011;
assign LUT_4[19081] = 32'b11111111111111110100111110110011;
assign LUT_4[19082] = 32'b11111111111111111011001101011111;
assign LUT_4[19083] = 32'b11111111111111110100011001010111;
assign LUT_4[19084] = 32'b11111111111111111000110011010111;
assign LUT_4[19085] = 32'b11111111111111110001111111001111;
assign LUT_4[19086] = 32'b11111111111111111000001101111011;
assign LUT_4[19087] = 32'b11111111111111110001011001110011;
assign LUT_4[19088] = 32'b00000000000000000000011000010100;
assign LUT_4[19089] = 32'b11111111111111111001100100001100;
assign LUT_4[19090] = 32'b11111111111111111111110010111000;
assign LUT_4[19091] = 32'b11111111111111111000111110110000;
assign LUT_4[19092] = 32'b11111111111111111101011000110000;
assign LUT_4[19093] = 32'b11111111111111110110100100101000;
assign LUT_4[19094] = 32'b11111111111111111100110011010100;
assign LUT_4[19095] = 32'b11111111111111110101111111001100;
assign LUT_4[19096] = 32'b11111111111111111001100100101001;
assign LUT_4[19097] = 32'b11111111111111110010110000100001;
assign LUT_4[19098] = 32'b11111111111111111000111111001101;
assign LUT_4[19099] = 32'b11111111111111110010001011000101;
assign LUT_4[19100] = 32'b11111111111111110110100101000101;
assign LUT_4[19101] = 32'b11111111111111101111110000111101;
assign LUT_4[19102] = 32'b11111111111111110101111111101001;
assign LUT_4[19103] = 32'b11111111111111101111001011100001;
assign LUT_4[19104] = 32'b00000000000000000001000001101101;
assign LUT_4[19105] = 32'b11111111111111111010001101100101;
assign LUT_4[19106] = 32'b00000000000000000000011100010001;
assign LUT_4[19107] = 32'b11111111111111111001101000001001;
assign LUT_4[19108] = 32'b11111111111111111110000010001001;
assign LUT_4[19109] = 32'b11111111111111110111001110000001;
assign LUT_4[19110] = 32'b11111111111111111101011100101101;
assign LUT_4[19111] = 32'b11111111111111110110101000100101;
assign LUT_4[19112] = 32'b11111111111111111010001110000010;
assign LUT_4[19113] = 32'b11111111111111110011011001111010;
assign LUT_4[19114] = 32'b11111111111111111001101000100110;
assign LUT_4[19115] = 32'b11111111111111110010110100011110;
assign LUT_4[19116] = 32'b11111111111111110111001110011110;
assign LUT_4[19117] = 32'b11111111111111110000011010010110;
assign LUT_4[19118] = 32'b11111111111111110110101001000010;
assign LUT_4[19119] = 32'b11111111111111101111110100111010;
assign LUT_4[19120] = 32'b11111111111111111110110011011011;
assign LUT_4[19121] = 32'b11111111111111110111111111010011;
assign LUT_4[19122] = 32'b11111111111111111110001101111111;
assign LUT_4[19123] = 32'b11111111111111110111011001110111;
assign LUT_4[19124] = 32'b11111111111111111011110011110111;
assign LUT_4[19125] = 32'b11111111111111110100111111101111;
assign LUT_4[19126] = 32'b11111111111111111011001110011011;
assign LUT_4[19127] = 32'b11111111111111110100011010010011;
assign LUT_4[19128] = 32'b11111111111111110111111111110000;
assign LUT_4[19129] = 32'b11111111111111110001001011101000;
assign LUT_4[19130] = 32'b11111111111111110111011010010100;
assign LUT_4[19131] = 32'b11111111111111110000100110001100;
assign LUT_4[19132] = 32'b11111111111111110101000000001100;
assign LUT_4[19133] = 32'b11111111111111101110001100000100;
assign LUT_4[19134] = 32'b11111111111111110100011010110000;
assign LUT_4[19135] = 32'b11111111111111101101100110101000;
assign LUT_4[19136] = 32'b00000000000000000011111101111010;
assign LUT_4[19137] = 32'b11111111111111111101001001110010;
assign LUT_4[19138] = 32'b00000000000000000011011000011110;
assign LUT_4[19139] = 32'b11111111111111111100100100010110;
assign LUT_4[19140] = 32'b00000000000000000000111110010110;
assign LUT_4[19141] = 32'b11111111111111111010001010001110;
assign LUT_4[19142] = 32'b00000000000000000000011000111010;
assign LUT_4[19143] = 32'b11111111111111111001100100110010;
assign LUT_4[19144] = 32'b11111111111111111101001010001111;
assign LUT_4[19145] = 32'b11111111111111110110010110000111;
assign LUT_4[19146] = 32'b11111111111111111100100100110011;
assign LUT_4[19147] = 32'b11111111111111110101110000101011;
assign LUT_4[19148] = 32'b11111111111111111010001010101011;
assign LUT_4[19149] = 32'b11111111111111110011010110100011;
assign LUT_4[19150] = 32'b11111111111111111001100101001111;
assign LUT_4[19151] = 32'b11111111111111110010110001000111;
assign LUT_4[19152] = 32'b00000000000000000001101111101000;
assign LUT_4[19153] = 32'b11111111111111111010111011100000;
assign LUT_4[19154] = 32'b00000000000000000001001010001100;
assign LUT_4[19155] = 32'b11111111111111111010010110000100;
assign LUT_4[19156] = 32'b11111111111111111110110000000100;
assign LUT_4[19157] = 32'b11111111111111110111111011111100;
assign LUT_4[19158] = 32'b11111111111111111110001010101000;
assign LUT_4[19159] = 32'b11111111111111110111010110100000;
assign LUT_4[19160] = 32'b11111111111111111010111011111101;
assign LUT_4[19161] = 32'b11111111111111110100000111110101;
assign LUT_4[19162] = 32'b11111111111111111010010110100001;
assign LUT_4[19163] = 32'b11111111111111110011100010011001;
assign LUT_4[19164] = 32'b11111111111111110111111100011001;
assign LUT_4[19165] = 32'b11111111111111110001001000010001;
assign LUT_4[19166] = 32'b11111111111111110111010110111101;
assign LUT_4[19167] = 32'b11111111111111110000100010110101;
assign LUT_4[19168] = 32'b00000000000000000010011001000001;
assign LUT_4[19169] = 32'b11111111111111111011100100111001;
assign LUT_4[19170] = 32'b00000000000000000001110011100101;
assign LUT_4[19171] = 32'b11111111111111111010111111011101;
assign LUT_4[19172] = 32'b11111111111111111111011001011101;
assign LUT_4[19173] = 32'b11111111111111111000100101010101;
assign LUT_4[19174] = 32'b11111111111111111110110100000001;
assign LUT_4[19175] = 32'b11111111111111110111111111111001;
assign LUT_4[19176] = 32'b11111111111111111011100101010110;
assign LUT_4[19177] = 32'b11111111111111110100110001001110;
assign LUT_4[19178] = 32'b11111111111111111010111111111010;
assign LUT_4[19179] = 32'b11111111111111110100001011110010;
assign LUT_4[19180] = 32'b11111111111111111000100101110010;
assign LUT_4[19181] = 32'b11111111111111110001110001101010;
assign LUT_4[19182] = 32'b11111111111111111000000000010110;
assign LUT_4[19183] = 32'b11111111111111110001001100001110;
assign LUT_4[19184] = 32'b00000000000000000000001010101111;
assign LUT_4[19185] = 32'b11111111111111111001010110100111;
assign LUT_4[19186] = 32'b11111111111111111111100101010011;
assign LUT_4[19187] = 32'b11111111111111111000110001001011;
assign LUT_4[19188] = 32'b11111111111111111101001011001011;
assign LUT_4[19189] = 32'b11111111111111110110010111000011;
assign LUT_4[19190] = 32'b11111111111111111100100101101111;
assign LUT_4[19191] = 32'b11111111111111110101110001100111;
assign LUT_4[19192] = 32'b11111111111111111001010111000100;
assign LUT_4[19193] = 32'b11111111111111110010100010111100;
assign LUT_4[19194] = 32'b11111111111111111000110001101000;
assign LUT_4[19195] = 32'b11111111111111110001111101100000;
assign LUT_4[19196] = 32'b11111111111111110110010111100000;
assign LUT_4[19197] = 32'b11111111111111101111100011011000;
assign LUT_4[19198] = 32'b11111111111111110101110010000100;
assign LUT_4[19199] = 32'b11111111111111101110111101111100;
assign LUT_4[19200] = 32'b00000000000000000100111100000001;
assign LUT_4[19201] = 32'b11111111111111111110000111111001;
assign LUT_4[19202] = 32'b00000000000000000100010110100101;
assign LUT_4[19203] = 32'b11111111111111111101100010011101;
assign LUT_4[19204] = 32'b00000000000000000001111100011101;
assign LUT_4[19205] = 32'b11111111111111111011001000010101;
assign LUT_4[19206] = 32'b00000000000000000001010111000001;
assign LUT_4[19207] = 32'b11111111111111111010100010111001;
assign LUT_4[19208] = 32'b11111111111111111110001000010110;
assign LUT_4[19209] = 32'b11111111111111110111010100001110;
assign LUT_4[19210] = 32'b11111111111111111101100010111010;
assign LUT_4[19211] = 32'b11111111111111110110101110110010;
assign LUT_4[19212] = 32'b11111111111111111011001000110010;
assign LUT_4[19213] = 32'b11111111111111110100010100101010;
assign LUT_4[19214] = 32'b11111111111111111010100011010110;
assign LUT_4[19215] = 32'b11111111111111110011101111001110;
assign LUT_4[19216] = 32'b00000000000000000010101101101111;
assign LUT_4[19217] = 32'b11111111111111111011111001100111;
assign LUT_4[19218] = 32'b00000000000000000010001000010011;
assign LUT_4[19219] = 32'b11111111111111111011010100001011;
assign LUT_4[19220] = 32'b11111111111111111111101110001011;
assign LUT_4[19221] = 32'b11111111111111111000111010000011;
assign LUT_4[19222] = 32'b11111111111111111111001000101111;
assign LUT_4[19223] = 32'b11111111111111111000010100100111;
assign LUT_4[19224] = 32'b11111111111111111011111010000100;
assign LUT_4[19225] = 32'b11111111111111110101000101111100;
assign LUT_4[19226] = 32'b11111111111111111011010100101000;
assign LUT_4[19227] = 32'b11111111111111110100100000100000;
assign LUT_4[19228] = 32'b11111111111111111000111010100000;
assign LUT_4[19229] = 32'b11111111111111110010000110011000;
assign LUT_4[19230] = 32'b11111111111111111000010101000100;
assign LUT_4[19231] = 32'b11111111111111110001100000111100;
assign LUT_4[19232] = 32'b00000000000000000011010111001000;
assign LUT_4[19233] = 32'b11111111111111111100100011000000;
assign LUT_4[19234] = 32'b00000000000000000010110001101100;
assign LUT_4[19235] = 32'b11111111111111111011111101100100;
assign LUT_4[19236] = 32'b00000000000000000000010111100100;
assign LUT_4[19237] = 32'b11111111111111111001100011011100;
assign LUT_4[19238] = 32'b11111111111111111111110010001000;
assign LUT_4[19239] = 32'b11111111111111111000111110000000;
assign LUT_4[19240] = 32'b11111111111111111100100011011101;
assign LUT_4[19241] = 32'b11111111111111110101101111010101;
assign LUT_4[19242] = 32'b11111111111111111011111110000001;
assign LUT_4[19243] = 32'b11111111111111110101001001111001;
assign LUT_4[19244] = 32'b11111111111111111001100011111001;
assign LUT_4[19245] = 32'b11111111111111110010101111110001;
assign LUT_4[19246] = 32'b11111111111111111000111110011101;
assign LUT_4[19247] = 32'b11111111111111110010001010010101;
assign LUT_4[19248] = 32'b00000000000000000001001000110110;
assign LUT_4[19249] = 32'b11111111111111111010010100101110;
assign LUT_4[19250] = 32'b00000000000000000000100011011010;
assign LUT_4[19251] = 32'b11111111111111111001101111010010;
assign LUT_4[19252] = 32'b11111111111111111110001001010010;
assign LUT_4[19253] = 32'b11111111111111110111010101001010;
assign LUT_4[19254] = 32'b11111111111111111101100011110110;
assign LUT_4[19255] = 32'b11111111111111110110101111101110;
assign LUT_4[19256] = 32'b11111111111111111010010101001011;
assign LUT_4[19257] = 32'b11111111111111110011100001000011;
assign LUT_4[19258] = 32'b11111111111111111001101111101111;
assign LUT_4[19259] = 32'b11111111111111110010111011100111;
assign LUT_4[19260] = 32'b11111111111111110111010101100111;
assign LUT_4[19261] = 32'b11111111111111110000100001011111;
assign LUT_4[19262] = 32'b11111111111111110110110000001011;
assign LUT_4[19263] = 32'b11111111111111101111111100000011;
assign LUT_4[19264] = 32'b00000000000000000110010011010101;
assign LUT_4[19265] = 32'b11111111111111111111011111001101;
assign LUT_4[19266] = 32'b00000000000000000101101101111001;
assign LUT_4[19267] = 32'b11111111111111111110111001110001;
assign LUT_4[19268] = 32'b00000000000000000011010011110001;
assign LUT_4[19269] = 32'b11111111111111111100011111101001;
assign LUT_4[19270] = 32'b00000000000000000010101110010101;
assign LUT_4[19271] = 32'b11111111111111111011111010001101;
assign LUT_4[19272] = 32'b11111111111111111111011111101010;
assign LUT_4[19273] = 32'b11111111111111111000101011100010;
assign LUT_4[19274] = 32'b11111111111111111110111010001110;
assign LUT_4[19275] = 32'b11111111111111111000000110000110;
assign LUT_4[19276] = 32'b11111111111111111100100000000110;
assign LUT_4[19277] = 32'b11111111111111110101101011111110;
assign LUT_4[19278] = 32'b11111111111111111011111010101010;
assign LUT_4[19279] = 32'b11111111111111110101000110100010;
assign LUT_4[19280] = 32'b00000000000000000100000101000011;
assign LUT_4[19281] = 32'b11111111111111111101010000111011;
assign LUT_4[19282] = 32'b00000000000000000011011111100111;
assign LUT_4[19283] = 32'b11111111111111111100101011011111;
assign LUT_4[19284] = 32'b00000000000000000001000101011111;
assign LUT_4[19285] = 32'b11111111111111111010010001010111;
assign LUT_4[19286] = 32'b00000000000000000000100000000011;
assign LUT_4[19287] = 32'b11111111111111111001101011111011;
assign LUT_4[19288] = 32'b11111111111111111101010001011000;
assign LUT_4[19289] = 32'b11111111111111110110011101010000;
assign LUT_4[19290] = 32'b11111111111111111100101011111100;
assign LUT_4[19291] = 32'b11111111111111110101110111110100;
assign LUT_4[19292] = 32'b11111111111111111010010001110100;
assign LUT_4[19293] = 32'b11111111111111110011011101101100;
assign LUT_4[19294] = 32'b11111111111111111001101100011000;
assign LUT_4[19295] = 32'b11111111111111110010111000010000;
assign LUT_4[19296] = 32'b00000000000000000100101110011100;
assign LUT_4[19297] = 32'b11111111111111111101111010010100;
assign LUT_4[19298] = 32'b00000000000000000100001001000000;
assign LUT_4[19299] = 32'b11111111111111111101010100111000;
assign LUT_4[19300] = 32'b00000000000000000001101110111000;
assign LUT_4[19301] = 32'b11111111111111111010111010110000;
assign LUT_4[19302] = 32'b00000000000000000001001001011100;
assign LUT_4[19303] = 32'b11111111111111111010010101010100;
assign LUT_4[19304] = 32'b11111111111111111101111010110001;
assign LUT_4[19305] = 32'b11111111111111110111000110101001;
assign LUT_4[19306] = 32'b11111111111111111101010101010101;
assign LUT_4[19307] = 32'b11111111111111110110100001001101;
assign LUT_4[19308] = 32'b11111111111111111010111011001101;
assign LUT_4[19309] = 32'b11111111111111110100000111000101;
assign LUT_4[19310] = 32'b11111111111111111010010101110001;
assign LUT_4[19311] = 32'b11111111111111110011100001101001;
assign LUT_4[19312] = 32'b00000000000000000010100000001010;
assign LUT_4[19313] = 32'b11111111111111111011101100000010;
assign LUT_4[19314] = 32'b00000000000000000001111010101110;
assign LUT_4[19315] = 32'b11111111111111111011000110100110;
assign LUT_4[19316] = 32'b11111111111111111111100000100110;
assign LUT_4[19317] = 32'b11111111111111111000101100011110;
assign LUT_4[19318] = 32'b11111111111111111110111011001010;
assign LUT_4[19319] = 32'b11111111111111111000000111000010;
assign LUT_4[19320] = 32'b11111111111111111011101100011111;
assign LUT_4[19321] = 32'b11111111111111110100111000010111;
assign LUT_4[19322] = 32'b11111111111111111011000111000011;
assign LUT_4[19323] = 32'b11111111111111110100010010111011;
assign LUT_4[19324] = 32'b11111111111111111000101100111011;
assign LUT_4[19325] = 32'b11111111111111110001111000110011;
assign LUT_4[19326] = 32'b11111111111111111000000111011111;
assign LUT_4[19327] = 32'b11111111111111110001010011010111;
assign LUT_4[19328] = 32'b00000000000000000111100010001001;
assign LUT_4[19329] = 32'b00000000000000000000101110000001;
assign LUT_4[19330] = 32'b00000000000000000110111100101101;
assign LUT_4[19331] = 32'b00000000000000000000001000100101;
assign LUT_4[19332] = 32'b00000000000000000100100010100101;
assign LUT_4[19333] = 32'b11111111111111111101101110011101;
assign LUT_4[19334] = 32'b00000000000000000011111101001001;
assign LUT_4[19335] = 32'b11111111111111111101001001000001;
assign LUT_4[19336] = 32'b00000000000000000000101110011110;
assign LUT_4[19337] = 32'b11111111111111111001111010010110;
assign LUT_4[19338] = 32'b00000000000000000000001001000010;
assign LUT_4[19339] = 32'b11111111111111111001010100111010;
assign LUT_4[19340] = 32'b11111111111111111101101110111010;
assign LUT_4[19341] = 32'b11111111111111110110111010110010;
assign LUT_4[19342] = 32'b11111111111111111101001001011110;
assign LUT_4[19343] = 32'b11111111111111110110010101010110;
assign LUT_4[19344] = 32'b00000000000000000101010011110111;
assign LUT_4[19345] = 32'b11111111111111111110011111101111;
assign LUT_4[19346] = 32'b00000000000000000100101110011011;
assign LUT_4[19347] = 32'b11111111111111111101111010010011;
assign LUT_4[19348] = 32'b00000000000000000010010100010011;
assign LUT_4[19349] = 32'b11111111111111111011100000001011;
assign LUT_4[19350] = 32'b00000000000000000001101110110111;
assign LUT_4[19351] = 32'b11111111111111111010111010101111;
assign LUT_4[19352] = 32'b11111111111111111110100000001100;
assign LUT_4[19353] = 32'b11111111111111110111101100000100;
assign LUT_4[19354] = 32'b11111111111111111101111010110000;
assign LUT_4[19355] = 32'b11111111111111110111000110101000;
assign LUT_4[19356] = 32'b11111111111111111011100000101000;
assign LUT_4[19357] = 32'b11111111111111110100101100100000;
assign LUT_4[19358] = 32'b11111111111111111010111011001100;
assign LUT_4[19359] = 32'b11111111111111110100000111000100;
assign LUT_4[19360] = 32'b00000000000000000101111101010000;
assign LUT_4[19361] = 32'b11111111111111111111001001001000;
assign LUT_4[19362] = 32'b00000000000000000101010111110100;
assign LUT_4[19363] = 32'b11111111111111111110100011101100;
assign LUT_4[19364] = 32'b00000000000000000010111101101100;
assign LUT_4[19365] = 32'b11111111111111111100001001100100;
assign LUT_4[19366] = 32'b00000000000000000010011000010000;
assign LUT_4[19367] = 32'b11111111111111111011100100001000;
assign LUT_4[19368] = 32'b11111111111111111111001001100101;
assign LUT_4[19369] = 32'b11111111111111111000010101011101;
assign LUT_4[19370] = 32'b11111111111111111110100100001001;
assign LUT_4[19371] = 32'b11111111111111110111110000000001;
assign LUT_4[19372] = 32'b11111111111111111100001010000001;
assign LUT_4[19373] = 32'b11111111111111110101010101111001;
assign LUT_4[19374] = 32'b11111111111111111011100100100101;
assign LUT_4[19375] = 32'b11111111111111110100110000011101;
assign LUT_4[19376] = 32'b00000000000000000011101110111110;
assign LUT_4[19377] = 32'b11111111111111111100111010110110;
assign LUT_4[19378] = 32'b00000000000000000011001001100010;
assign LUT_4[19379] = 32'b11111111111111111100010101011010;
assign LUT_4[19380] = 32'b00000000000000000000101111011010;
assign LUT_4[19381] = 32'b11111111111111111001111011010010;
assign LUT_4[19382] = 32'b00000000000000000000001001111110;
assign LUT_4[19383] = 32'b11111111111111111001010101110110;
assign LUT_4[19384] = 32'b11111111111111111100111011010011;
assign LUT_4[19385] = 32'b11111111111111110110000111001011;
assign LUT_4[19386] = 32'b11111111111111111100010101110111;
assign LUT_4[19387] = 32'b11111111111111110101100001101111;
assign LUT_4[19388] = 32'b11111111111111111001111011101111;
assign LUT_4[19389] = 32'b11111111111111110011000111100111;
assign LUT_4[19390] = 32'b11111111111111111001010110010011;
assign LUT_4[19391] = 32'b11111111111111110010100010001011;
assign LUT_4[19392] = 32'b00000000000000001000111001011101;
assign LUT_4[19393] = 32'b00000000000000000010000101010101;
assign LUT_4[19394] = 32'b00000000000000001000010100000001;
assign LUT_4[19395] = 32'b00000000000000000001011111111001;
assign LUT_4[19396] = 32'b00000000000000000101111001111001;
assign LUT_4[19397] = 32'b11111111111111111111000101110001;
assign LUT_4[19398] = 32'b00000000000000000101010100011101;
assign LUT_4[19399] = 32'b11111111111111111110100000010101;
assign LUT_4[19400] = 32'b00000000000000000010000101110010;
assign LUT_4[19401] = 32'b11111111111111111011010001101010;
assign LUT_4[19402] = 32'b00000000000000000001100000010110;
assign LUT_4[19403] = 32'b11111111111111111010101100001110;
assign LUT_4[19404] = 32'b11111111111111111111000110001110;
assign LUT_4[19405] = 32'b11111111111111111000010010000110;
assign LUT_4[19406] = 32'b11111111111111111110100000110010;
assign LUT_4[19407] = 32'b11111111111111110111101100101010;
assign LUT_4[19408] = 32'b00000000000000000110101011001011;
assign LUT_4[19409] = 32'b11111111111111111111110111000011;
assign LUT_4[19410] = 32'b00000000000000000110000101101111;
assign LUT_4[19411] = 32'b11111111111111111111010001100111;
assign LUT_4[19412] = 32'b00000000000000000011101011100111;
assign LUT_4[19413] = 32'b11111111111111111100110111011111;
assign LUT_4[19414] = 32'b00000000000000000011000110001011;
assign LUT_4[19415] = 32'b11111111111111111100010010000011;
assign LUT_4[19416] = 32'b11111111111111111111110111100000;
assign LUT_4[19417] = 32'b11111111111111111001000011011000;
assign LUT_4[19418] = 32'b11111111111111111111010010000100;
assign LUT_4[19419] = 32'b11111111111111111000011101111100;
assign LUT_4[19420] = 32'b11111111111111111100110111111100;
assign LUT_4[19421] = 32'b11111111111111110110000011110100;
assign LUT_4[19422] = 32'b11111111111111111100010010100000;
assign LUT_4[19423] = 32'b11111111111111110101011110011000;
assign LUT_4[19424] = 32'b00000000000000000111010100100100;
assign LUT_4[19425] = 32'b00000000000000000000100000011100;
assign LUT_4[19426] = 32'b00000000000000000110101111001000;
assign LUT_4[19427] = 32'b11111111111111111111111011000000;
assign LUT_4[19428] = 32'b00000000000000000100010101000000;
assign LUT_4[19429] = 32'b11111111111111111101100000111000;
assign LUT_4[19430] = 32'b00000000000000000011101111100100;
assign LUT_4[19431] = 32'b11111111111111111100111011011100;
assign LUT_4[19432] = 32'b00000000000000000000100000111001;
assign LUT_4[19433] = 32'b11111111111111111001101100110001;
assign LUT_4[19434] = 32'b11111111111111111111111011011101;
assign LUT_4[19435] = 32'b11111111111111111001000111010101;
assign LUT_4[19436] = 32'b11111111111111111101100001010101;
assign LUT_4[19437] = 32'b11111111111111110110101101001101;
assign LUT_4[19438] = 32'b11111111111111111100111011111001;
assign LUT_4[19439] = 32'b11111111111111110110000111110001;
assign LUT_4[19440] = 32'b00000000000000000101000110010010;
assign LUT_4[19441] = 32'b11111111111111111110010010001010;
assign LUT_4[19442] = 32'b00000000000000000100100000110110;
assign LUT_4[19443] = 32'b11111111111111111101101100101110;
assign LUT_4[19444] = 32'b00000000000000000010000110101110;
assign LUT_4[19445] = 32'b11111111111111111011010010100110;
assign LUT_4[19446] = 32'b00000000000000000001100001010010;
assign LUT_4[19447] = 32'b11111111111111111010101101001010;
assign LUT_4[19448] = 32'b11111111111111111110010010100111;
assign LUT_4[19449] = 32'b11111111111111110111011110011111;
assign LUT_4[19450] = 32'b11111111111111111101101101001011;
assign LUT_4[19451] = 32'b11111111111111110110111001000011;
assign LUT_4[19452] = 32'b11111111111111111011010011000011;
assign LUT_4[19453] = 32'b11111111111111110100011110111011;
assign LUT_4[19454] = 32'b11111111111111111010101101100111;
assign LUT_4[19455] = 32'b11111111111111110011111001011111;
assign LUT_4[19456] = 32'b00000000000000000010100110110101;
assign LUT_4[19457] = 32'b11111111111111111011110010101101;
assign LUT_4[19458] = 32'b00000000000000000010000001011001;
assign LUT_4[19459] = 32'b11111111111111111011001101010001;
assign LUT_4[19460] = 32'b11111111111111111111100111010001;
assign LUT_4[19461] = 32'b11111111111111111000110011001001;
assign LUT_4[19462] = 32'b11111111111111111111000001110101;
assign LUT_4[19463] = 32'b11111111111111111000001101101101;
assign LUT_4[19464] = 32'b11111111111111111011110011001010;
assign LUT_4[19465] = 32'b11111111111111110100111111000010;
assign LUT_4[19466] = 32'b11111111111111111011001101101110;
assign LUT_4[19467] = 32'b11111111111111110100011001100110;
assign LUT_4[19468] = 32'b11111111111111111000110011100110;
assign LUT_4[19469] = 32'b11111111111111110001111111011110;
assign LUT_4[19470] = 32'b11111111111111111000001110001010;
assign LUT_4[19471] = 32'b11111111111111110001011010000010;
assign LUT_4[19472] = 32'b00000000000000000000011000100011;
assign LUT_4[19473] = 32'b11111111111111111001100100011011;
assign LUT_4[19474] = 32'b11111111111111111111110011000111;
assign LUT_4[19475] = 32'b11111111111111111000111110111111;
assign LUT_4[19476] = 32'b11111111111111111101011000111111;
assign LUT_4[19477] = 32'b11111111111111110110100100110111;
assign LUT_4[19478] = 32'b11111111111111111100110011100011;
assign LUT_4[19479] = 32'b11111111111111110101111111011011;
assign LUT_4[19480] = 32'b11111111111111111001100100111000;
assign LUT_4[19481] = 32'b11111111111111110010110000110000;
assign LUT_4[19482] = 32'b11111111111111111000111111011100;
assign LUT_4[19483] = 32'b11111111111111110010001011010100;
assign LUT_4[19484] = 32'b11111111111111110110100101010100;
assign LUT_4[19485] = 32'b11111111111111101111110001001100;
assign LUT_4[19486] = 32'b11111111111111110101111111111000;
assign LUT_4[19487] = 32'b11111111111111101111001011110000;
assign LUT_4[19488] = 32'b00000000000000000001000001111100;
assign LUT_4[19489] = 32'b11111111111111111010001101110100;
assign LUT_4[19490] = 32'b00000000000000000000011100100000;
assign LUT_4[19491] = 32'b11111111111111111001101000011000;
assign LUT_4[19492] = 32'b11111111111111111110000010011000;
assign LUT_4[19493] = 32'b11111111111111110111001110010000;
assign LUT_4[19494] = 32'b11111111111111111101011100111100;
assign LUT_4[19495] = 32'b11111111111111110110101000110100;
assign LUT_4[19496] = 32'b11111111111111111010001110010001;
assign LUT_4[19497] = 32'b11111111111111110011011010001001;
assign LUT_4[19498] = 32'b11111111111111111001101000110101;
assign LUT_4[19499] = 32'b11111111111111110010110100101101;
assign LUT_4[19500] = 32'b11111111111111110111001110101101;
assign LUT_4[19501] = 32'b11111111111111110000011010100101;
assign LUT_4[19502] = 32'b11111111111111110110101001010001;
assign LUT_4[19503] = 32'b11111111111111101111110101001001;
assign LUT_4[19504] = 32'b11111111111111111110110011101010;
assign LUT_4[19505] = 32'b11111111111111110111111111100010;
assign LUT_4[19506] = 32'b11111111111111111110001110001110;
assign LUT_4[19507] = 32'b11111111111111110111011010000110;
assign LUT_4[19508] = 32'b11111111111111111011110100000110;
assign LUT_4[19509] = 32'b11111111111111110100111111111110;
assign LUT_4[19510] = 32'b11111111111111111011001110101010;
assign LUT_4[19511] = 32'b11111111111111110100011010100010;
assign LUT_4[19512] = 32'b11111111111111110111111111111111;
assign LUT_4[19513] = 32'b11111111111111110001001011110111;
assign LUT_4[19514] = 32'b11111111111111110111011010100011;
assign LUT_4[19515] = 32'b11111111111111110000100110011011;
assign LUT_4[19516] = 32'b11111111111111110101000000011011;
assign LUT_4[19517] = 32'b11111111111111101110001100010011;
assign LUT_4[19518] = 32'b11111111111111110100011010111111;
assign LUT_4[19519] = 32'b11111111111111101101100110110111;
assign LUT_4[19520] = 32'b00000000000000000011111110001001;
assign LUT_4[19521] = 32'b11111111111111111101001010000001;
assign LUT_4[19522] = 32'b00000000000000000011011000101101;
assign LUT_4[19523] = 32'b11111111111111111100100100100101;
assign LUT_4[19524] = 32'b00000000000000000000111110100101;
assign LUT_4[19525] = 32'b11111111111111111010001010011101;
assign LUT_4[19526] = 32'b00000000000000000000011001001001;
assign LUT_4[19527] = 32'b11111111111111111001100101000001;
assign LUT_4[19528] = 32'b11111111111111111101001010011110;
assign LUT_4[19529] = 32'b11111111111111110110010110010110;
assign LUT_4[19530] = 32'b11111111111111111100100101000010;
assign LUT_4[19531] = 32'b11111111111111110101110000111010;
assign LUT_4[19532] = 32'b11111111111111111010001010111010;
assign LUT_4[19533] = 32'b11111111111111110011010110110010;
assign LUT_4[19534] = 32'b11111111111111111001100101011110;
assign LUT_4[19535] = 32'b11111111111111110010110001010110;
assign LUT_4[19536] = 32'b00000000000000000001101111110111;
assign LUT_4[19537] = 32'b11111111111111111010111011101111;
assign LUT_4[19538] = 32'b00000000000000000001001010011011;
assign LUT_4[19539] = 32'b11111111111111111010010110010011;
assign LUT_4[19540] = 32'b11111111111111111110110000010011;
assign LUT_4[19541] = 32'b11111111111111110111111100001011;
assign LUT_4[19542] = 32'b11111111111111111110001010110111;
assign LUT_4[19543] = 32'b11111111111111110111010110101111;
assign LUT_4[19544] = 32'b11111111111111111010111100001100;
assign LUT_4[19545] = 32'b11111111111111110100001000000100;
assign LUT_4[19546] = 32'b11111111111111111010010110110000;
assign LUT_4[19547] = 32'b11111111111111110011100010101000;
assign LUT_4[19548] = 32'b11111111111111110111111100101000;
assign LUT_4[19549] = 32'b11111111111111110001001000100000;
assign LUT_4[19550] = 32'b11111111111111110111010111001100;
assign LUT_4[19551] = 32'b11111111111111110000100011000100;
assign LUT_4[19552] = 32'b00000000000000000010011001010000;
assign LUT_4[19553] = 32'b11111111111111111011100101001000;
assign LUT_4[19554] = 32'b00000000000000000001110011110100;
assign LUT_4[19555] = 32'b11111111111111111010111111101100;
assign LUT_4[19556] = 32'b11111111111111111111011001101100;
assign LUT_4[19557] = 32'b11111111111111111000100101100100;
assign LUT_4[19558] = 32'b11111111111111111110110100010000;
assign LUT_4[19559] = 32'b11111111111111111000000000001000;
assign LUT_4[19560] = 32'b11111111111111111011100101100101;
assign LUT_4[19561] = 32'b11111111111111110100110001011101;
assign LUT_4[19562] = 32'b11111111111111111011000000001001;
assign LUT_4[19563] = 32'b11111111111111110100001100000001;
assign LUT_4[19564] = 32'b11111111111111111000100110000001;
assign LUT_4[19565] = 32'b11111111111111110001110001111001;
assign LUT_4[19566] = 32'b11111111111111111000000000100101;
assign LUT_4[19567] = 32'b11111111111111110001001100011101;
assign LUT_4[19568] = 32'b00000000000000000000001010111110;
assign LUT_4[19569] = 32'b11111111111111111001010110110110;
assign LUT_4[19570] = 32'b11111111111111111111100101100010;
assign LUT_4[19571] = 32'b11111111111111111000110001011010;
assign LUT_4[19572] = 32'b11111111111111111101001011011010;
assign LUT_4[19573] = 32'b11111111111111110110010111010010;
assign LUT_4[19574] = 32'b11111111111111111100100101111110;
assign LUT_4[19575] = 32'b11111111111111110101110001110110;
assign LUT_4[19576] = 32'b11111111111111111001010111010011;
assign LUT_4[19577] = 32'b11111111111111110010100011001011;
assign LUT_4[19578] = 32'b11111111111111111000110001110111;
assign LUT_4[19579] = 32'b11111111111111110001111101101111;
assign LUT_4[19580] = 32'b11111111111111110110010111101111;
assign LUT_4[19581] = 32'b11111111111111101111100011100111;
assign LUT_4[19582] = 32'b11111111111111110101110010010011;
assign LUT_4[19583] = 32'b11111111111111101110111110001011;
assign LUT_4[19584] = 32'b00000000000000000101001100111101;
assign LUT_4[19585] = 32'b11111111111111111110011000110101;
assign LUT_4[19586] = 32'b00000000000000000100100111100001;
assign LUT_4[19587] = 32'b11111111111111111101110011011001;
assign LUT_4[19588] = 32'b00000000000000000010001101011001;
assign LUT_4[19589] = 32'b11111111111111111011011001010001;
assign LUT_4[19590] = 32'b00000000000000000001100111111101;
assign LUT_4[19591] = 32'b11111111111111111010110011110101;
assign LUT_4[19592] = 32'b11111111111111111110011001010010;
assign LUT_4[19593] = 32'b11111111111111110111100101001010;
assign LUT_4[19594] = 32'b11111111111111111101110011110110;
assign LUT_4[19595] = 32'b11111111111111110110111111101110;
assign LUT_4[19596] = 32'b11111111111111111011011001101110;
assign LUT_4[19597] = 32'b11111111111111110100100101100110;
assign LUT_4[19598] = 32'b11111111111111111010110100010010;
assign LUT_4[19599] = 32'b11111111111111110100000000001010;
assign LUT_4[19600] = 32'b00000000000000000010111110101011;
assign LUT_4[19601] = 32'b11111111111111111100001010100011;
assign LUT_4[19602] = 32'b00000000000000000010011001001111;
assign LUT_4[19603] = 32'b11111111111111111011100101000111;
assign LUT_4[19604] = 32'b11111111111111111111111111000111;
assign LUT_4[19605] = 32'b11111111111111111001001010111111;
assign LUT_4[19606] = 32'b11111111111111111111011001101011;
assign LUT_4[19607] = 32'b11111111111111111000100101100011;
assign LUT_4[19608] = 32'b11111111111111111100001011000000;
assign LUT_4[19609] = 32'b11111111111111110101010110111000;
assign LUT_4[19610] = 32'b11111111111111111011100101100100;
assign LUT_4[19611] = 32'b11111111111111110100110001011100;
assign LUT_4[19612] = 32'b11111111111111111001001011011100;
assign LUT_4[19613] = 32'b11111111111111110010010111010100;
assign LUT_4[19614] = 32'b11111111111111111000100110000000;
assign LUT_4[19615] = 32'b11111111111111110001110001111000;
assign LUT_4[19616] = 32'b00000000000000000011101000000100;
assign LUT_4[19617] = 32'b11111111111111111100110011111100;
assign LUT_4[19618] = 32'b00000000000000000011000010101000;
assign LUT_4[19619] = 32'b11111111111111111100001110100000;
assign LUT_4[19620] = 32'b00000000000000000000101000100000;
assign LUT_4[19621] = 32'b11111111111111111001110100011000;
assign LUT_4[19622] = 32'b00000000000000000000000011000100;
assign LUT_4[19623] = 32'b11111111111111111001001110111100;
assign LUT_4[19624] = 32'b11111111111111111100110100011001;
assign LUT_4[19625] = 32'b11111111111111110110000000010001;
assign LUT_4[19626] = 32'b11111111111111111100001110111101;
assign LUT_4[19627] = 32'b11111111111111110101011010110101;
assign LUT_4[19628] = 32'b11111111111111111001110100110101;
assign LUT_4[19629] = 32'b11111111111111110011000000101101;
assign LUT_4[19630] = 32'b11111111111111111001001111011001;
assign LUT_4[19631] = 32'b11111111111111110010011011010001;
assign LUT_4[19632] = 32'b00000000000000000001011001110010;
assign LUT_4[19633] = 32'b11111111111111111010100101101010;
assign LUT_4[19634] = 32'b00000000000000000000110100010110;
assign LUT_4[19635] = 32'b11111111111111111010000000001110;
assign LUT_4[19636] = 32'b11111111111111111110011010001110;
assign LUT_4[19637] = 32'b11111111111111110111100110000110;
assign LUT_4[19638] = 32'b11111111111111111101110100110010;
assign LUT_4[19639] = 32'b11111111111111110111000000101010;
assign LUT_4[19640] = 32'b11111111111111111010100110000111;
assign LUT_4[19641] = 32'b11111111111111110011110001111111;
assign LUT_4[19642] = 32'b11111111111111111010000000101011;
assign LUT_4[19643] = 32'b11111111111111110011001100100011;
assign LUT_4[19644] = 32'b11111111111111110111100110100011;
assign LUT_4[19645] = 32'b11111111111111110000110010011011;
assign LUT_4[19646] = 32'b11111111111111110111000001000111;
assign LUT_4[19647] = 32'b11111111111111110000001100111111;
assign LUT_4[19648] = 32'b00000000000000000110100100010001;
assign LUT_4[19649] = 32'b11111111111111111111110000001001;
assign LUT_4[19650] = 32'b00000000000000000101111110110101;
assign LUT_4[19651] = 32'b11111111111111111111001010101101;
assign LUT_4[19652] = 32'b00000000000000000011100100101101;
assign LUT_4[19653] = 32'b11111111111111111100110000100101;
assign LUT_4[19654] = 32'b00000000000000000010111111010001;
assign LUT_4[19655] = 32'b11111111111111111100001011001001;
assign LUT_4[19656] = 32'b11111111111111111111110000100110;
assign LUT_4[19657] = 32'b11111111111111111000111100011110;
assign LUT_4[19658] = 32'b11111111111111111111001011001010;
assign LUT_4[19659] = 32'b11111111111111111000010111000010;
assign LUT_4[19660] = 32'b11111111111111111100110001000010;
assign LUT_4[19661] = 32'b11111111111111110101111100111010;
assign LUT_4[19662] = 32'b11111111111111111100001011100110;
assign LUT_4[19663] = 32'b11111111111111110101010111011110;
assign LUT_4[19664] = 32'b00000000000000000100010101111111;
assign LUT_4[19665] = 32'b11111111111111111101100001110111;
assign LUT_4[19666] = 32'b00000000000000000011110000100011;
assign LUT_4[19667] = 32'b11111111111111111100111100011011;
assign LUT_4[19668] = 32'b00000000000000000001010110011011;
assign LUT_4[19669] = 32'b11111111111111111010100010010011;
assign LUT_4[19670] = 32'b00000000000000000000110000111111;
assign LUT_4[19671] = 32'b11111111111111111001111100110111;
assign LUT_4[19672] = 32'b11111111111111111101100010010100;
assign LUT_4[19673] = 32'b11111111111111110110101110001100;
assign LUT_4[19674] = 32'b11111111111111111100111100111000;
assign LUT_4[19675] = 32'b11111111111111110110001000110000;
assign LUT_4[19676] = 32'b11111111111111111010100010110000;
assign LUT_4[19677] = 32'b11111111111111110011101110101000;
assign LUT_4[19678] = 32'b11111111111111111001111101010100;
assign LUT_4[19679] = 32'b11111111111111110011001001001100;
assign LUT_4[19680] = 32'b00000000000000000100111111011000;
assign LUT_4[19681] = 32'b11111111111111111110001011010000;
assign LUT_4[19682] = 32'b00000000000000000100011001111100;
assign LUT_4[19683] = 32'b11111111111111111101100101110100;
assign LUT_4[19684] = 32'b00000000000000000001111111110100;
assign LUT_4[19685] = 32'b11111111111111111011001011101100;
assign LUT_4[19686] = 32'b00000000000000000001011010011000;
assign LUT_4[19687] = 32'b11111111111111111010100110010000;
assign LUT_4[19688] = 32'b11111111111111111110001011101101;
assign LUT_4[19689] = 32'b11111111111111110111010111100101;
assign LUT_4[19690] = 32'b11111111111111111101100110010001;
assign LUT_4[19691] = 32'b11111111111111110110110010001001;
assign LUT_4[19692] = 32'b11111111111111111011001100001001;
assign LUT_4[19693] = 32'b11111111111111110100011000000001;
assign LUT_4[19694] = 32'b11111111111111111010100110101101;
assign LUT_4[19695] = 32'b11111111111111110011110010100101;
assign LUT_4[19696] = 32'b00000000000000000010110001000110;
assign LUT_4[19697] = 32'b11111111111111111011111100111110;
assign LUT_4[19698] = 32'b00000000000000000010001011101010;
assign LUT_4[19699] = 32'b11111111111111111011010111100010;
assign LUT_4[19700] = 32'b11111111111111111111110001100010;
assign LUT_4[19701] = 32'b11111111111111111000111101011010;
assign LUT_4[19702] = 32'b11111111111111111111001100000110;
assign LUT_4[19703] = 32'b11111111111111111000010111111110;
assign LUT_4[19704] = 32'b11111111111111111011111101011011;
assign LUT_4[19705] = 32'b11111111111111110101001001010011;
assign LUT_4[19706] = 32'b11111111111111111011010111111111;
assign LUT_4[19707] = 32'b11111111111111110100100011110111;
assign LUT_4[19708] = 32'b11111111111111111000111101110111;
assign LUT_4[19709] = 32'b11111111111111110010001001101111;
assign LUT_4[19710] = 32'b11111111111111111000011000011011;
assign LUT_4[19711] = 32'b11111111111111110001100100010011;
assign LUT_4[19712] = 32'b00000000000000000111100010011000;
assign LUT_4[19713] = 32'b00000000000000000000101110010000;
assign LUT_4[19714] = 32'b00000000000000000110111100111100;
assign LUT_4[19715] = 32'b00000000000000000000001000110100;
assign LUT_4[19716] = 32'b00000000000000000100100010110100;
assign LUT_4[19717] = 32'b11111111111111111101101110101100;
assign LUT_4[19718] = 32'b00000000000000000011111101011000;
assign LUT_4[19719] = 32'b11111111111111111101001001010000;
assign LUT_4[19720] = 32'b00000000000000000000101110101101;
assign LUT_4[19721] = 32'b11111111111111111001111010100101;
assign LUT_4[19722] = 32'b00000000000000000000001001010001;
assign LUT_4[19723] = 32'b11111111111111111001010101001001;
assign LUT_4[19724] = 32'b11111111111111111101101111001001;
assign LUT_4[19725] = 32'b11111111111111110110111011000001;
assign LUT_4[19726] = 32'b11111111111111111101001001101101;
assign LUT_4[19727] = 32'b11111111111111110110010101100101;
assign LUT_4[19728] = 32'b00000000000000000101010100000110;
assign LUT_4[19729] = 32'b11111111111111111110011111111110;
assign LUT_4[19730] = 32'b00000000000000000100101110101010;
assign LUT_4[19731] = 32'b11111111111111111101111010100010;
assign LUT_4[19732] = 32'b00000000000000000010010100100010;
assign LUT_4[19733] = 32'b11111111111111111011100000011010;
assign LUT_4[19734] = 32'b00000000000000000001101111000110;
assign LUT_4[19735] = 32'b11111111111111111010111010111110;
assign LUT_4[19736] = 32'b11111111111111111110100000011011;
assign LUT_4[19737] = 32'b11111111111111110111101100010011;
assign LUT_4[19738] = 32'b11111111111111111101111010111111;
assign LUT_4[19739] = 32'b11111111111111110111000110110111;
assign LUT_4[19740] = 32'b11111111111111111011100000110111;
assign LUT_4[19741] = 32'b11111111111111110100101100101111;
assign LUT_4[19742] = 32'b11111111111111111010111011011011;
assign LUT_4[19743] = 32'b11111111111111110100000111010011;
assign LUT_4[19744] = 32'b00000000000000000101111101011111;
assign LUT_4[19745] = 32'b11111111111111111111001001010111;
assign LUT_4[19746] = 32'b00000000000000000101011000000011;
assign LUT_4[19747] = 32'b11111111111111111110100011111011;
assign LUT_4[19748] = 32'b00000000000000000010111101111011;
assign LUT_4[19749] = 32'b11111111111111111100001001110011;
assign LUT_4[19750] = 32'b00000000000000000010011000011111;
assign LUT_4[19751] = 32'b11111111111111111011100100010111;
assign LUT_4[19752] = 32'b11111111111111111111001001110100;
assign LUT_4[19753] = 32'b11111111111111111000010101101100;
assign LUT_4[19754] = 32'b11111111111111111110100100011000;
assign LUT_4[19755] = 32'b11111111111111110111110000010000;
assign LUT_4[19756] = 32'b11111111111111111100001010010000;
assign LUT_4[19757] = 32'b11111111111111110101010110001000;
assign LUT_4[19758] = 32'b11111111111111111011100100110100;
assign LUT_4[19759] = 32'b11111111111111110100110000101100;
assign LUT_4[19760] = 32'b00000000000000000011101111001101;
assign LUT_4[19761] = 32'b11111111111111111100111011000101;
assign LUT_4[19762] = 32'b00000000000000000011001001110001;
assign LUT_4[19763] = 32'b11111111111111111100010101101001;
assign LUT_4[19764] = 32'b00000000000000000000101111101001;
assign LUT_4[19765] = 32'b11111111111111111001111011100001;
assign LUT_4[19766] = 32'b00000000000000000000001010001101;
assign LUT_4[19767] = 32'b11111111111111111001010110000101;
assign LUT_4[19768] = 32'b11111111111111111100111011100010;
assign LUT_4[19769] = 32'b11111111111111110110000111011010;
assign LUT_4[19770] = 32'b11111111111111111100010110000110;
assign LUT_4[19771] = 32'b11111111111111110101100001111110;
assign LUT_4[19772] = 32'b11111111111111111001111011111110;
assign LUT_4[19773] = 32'b11111111111111110011000111110110;
assign LUT_4[19774] = 32'b11111111111111111001010110100010;
assign LUT_4[19775] = 32'b11111111111111110010100010011010;
assign LUT_4[19776] = 32'b00000000000000001000111001101100;
assign LUT_4[19777] = 32'b00000000000000000010000101100100;
assign LUT_4[19778] = 32'b00000000000000001000010100010000;
assign LUT_4[19779] = 32'b00000000000000000001100000001000;
assign LUT_4[19780] = 32'b00000000000000000101111010001000;
assign LUT_4[19781] = 32'b11111111111111111111000110000000;
assign LUT_4[19782] = 32'b00000000000000000101010100101100;
assign LUT_4[19783] = 32'b11111111111111111110100000100100;
assign LUT_4[19784] = 32'b00000000000000000010000110000001;
assign LUT_4[19785] = 32'b11111111111111111011010001111001;
assign LUT_4[19786] = 32'b00000000000000000001100000100101;
assign LUT_4[19787] = 32'b11111111111111111010101100011101;
assign LUT_4[19788] = 32'b11111111111111111111000110011101;
assign LUT_4[19789] = 32'b11111111111111111000010010010101;
assign LUT_4[19790] = 32'b11111111111111111110100001000001;
assign LUT_4[19791] = 32'b11111111111111110111101100111001;
assign LUT_4[19792] = 32'b00000000000000000110101011011010;
assign LUT_4[19793] = 32'b11111111111111111111110111010010;
assign LUT_4[19794] = 32'b00000000000000000110000101111110;
assign LUT_4[19795] = 32'b11111111111111111111010001110110;
assign LUT_4[19796] = 32'b00000000000000000011101011110110;
assign LUT_4[19797] = 32'b11111111111111111100110111101110;
assign LUT_4[19798] = 32'b00000000000000000011000110011010;
assign LUT_4[19799] = 32'b11111111111111111100010010010010;
assign LUT_4[19800] = 32'b11111111111111111111110111101111;
assign LUT_4[19801] = 32'b11111111111111111001000011100111;
assign LUT_4[19802] = 32'b11111111111111111111010010010011;
assign LUT_4[19803] = 32'b11111111111111111000011110001011;
assign LUT_4[19804] = 32'b11111111111111111100111000001011;
assign LUT_4[19805] = 32'b11111111111111110110000100000011;
assign LUT_4[19806] = 32'b11111111111111111100010010101111;
assign LUT_4[19807] = 32'b11111111111111110101011110100111;
assign LUT_4[19808] = 32'b00000000000000000111010100110011;
assign LUT_4[19809] = 32'b00000000000000000000100000101011;
assign LUT_4[19810] = 32'b00000000000000000110101111010111;
assign LUT_4[19811] = 32'b11111111111111111111111011001111;
assign LUT_4[19812] = 32'b00000000000000000100010101001111;
assign LUT_4[19813] = 32'b11111111111111111101100001000111;
assign LUT_4[19814] = 32'b00000000000000000011101111110011;
assign LUT_4[19815] = 32'b11111111111111111100111011101011;
assign LUT_4[19816] = 32'b00000000000000000000100001001000;
assign LUT_4[19817] = 32'b11111111111111111001101101000000;
assign LUT_4[19818] = 32'b11111111111111111111111011101100;
assign LUT_4[19819] = 32'b11111111111111111001000111100100;
assign LUT_4[19820] = 32'b11111111111111111101100001100100;
assign LUT_4[19821] = 32'b11111111111111110110101101011100;
assign LUT_4[19822] = 32'b11111111111111111100111100001000;
assign LUT_4[19823] = 32'b11111111111111110110001000000000;
assign LUT_4[19824] = 32'b00000000000000000101000110100001;
assign LUT_4[19825] = 32'b11111111111111111110010010011001;
assign LUT_4[19826] = 32'b00000000000000000100100001000101;
assign LUT_4[19827] = 32'b11111111111111111101101100111101;
assign LUT_4[19828] = 32'b00000000000000000010000110111101;
assign LUT_4[19829] = 32'b11111111111111111011010010110101;
assign LUT_4[19830] = 32'b00000000000000000001100001100001;
assign LUT_4[19831] = 32'b11111111111111111010101101011001;
assign LUT_4[19832] = 32'b11111111111111111110010010110110;
assign LUT_4[19833] = 32'b11111111111111110111011110101110;
assign LUT_4[19834] = 32'b11111111111111111101101101011010;
assign LUT_4[19835] = 32'b11111111111111110110111001010010;
assign LUT_4[19836] = 32'b11111111111111111011010011010010;
assign LUT_4[19837] = 32'b11111111111111110100011111001010;
assign LUT_4[19838] = 32'b11111111111111111010101101110110;
assign LUT_4[19839] = 32'b11111111111111110011111001101110;
assign LUT_4[19840] = 32'b00000000000000001010001000100000;
assign LUT_4[19841] = 32'b00000000000000000011010100011000;
assign LUT_4[19842] = 32'b00000000000000001001100011000100;
assign LUT_4[19843] = 32'b00000000000000000010101110111100;
assign LUT_4[19844] = 32'b00000000000000000111001000111100;
assign LUT_4[19845] = 32'b00000000000000000000010100110100;
assign LUT_4[19846] = 32'b00000000000000000110100011100000;
assign LUT_4[19847] = 32'b11111111111111111111101111011000;
assign LUT_4[19848] = 32'b00000000000000000011010100110101;
assign LUT_4[19849] = 32'b11111111111111111100100000101101;
assign LUT_4[19850] = 32'b00000000000000000010101111011001;
assign LUT_4[19851] = 32'b11111111111111111011111011010001;
assign LUT_4[19852] = 32'b00000000000000000000010101010001;
assign LUT_4[19853] = 32'b11111111111111111001100001001001;
assign LUT_4[19854] = 32'b11111111111111111111101111110101;
assign LUT_4[19855] = 32'b11111111111111111000111011101101;
assign LUT_4[19856] = 32'b00000000000000000111111010001110;
assign LUT_4[19857] = 32'b00000000000000000001000110000110;
assign LUT_4[19858] = 32'b00000000000000000111010100110010;
assign LUT_4[19859] = 32'b00000000000000000000100000101010;
assign LUT_4[19860] = 32'b00000000000000000100111010101010;
assign LUT_4[19861] = 32'b11111111111111111110000110100010;
assign LUT_4[19862] = 32'b00000000000000000100010101001110;
assign LUT_4[19863] = 32'b11111111111111111101100001000110;
assign LUT_4[19864] = 32'b00000000000000000001000110100011;
assign LUT_4[19865] = 32'b11111111111111111010010010011011;
assign LUT_4[19866] = 32'b00000000000000000000100001000111;
assign LUT_4[19867] = 32'b11111111111111111001101100111111;
assign LUT_4[19868] = 32'b11111111111111111110000110111111;
assign LUT_4[19869] = 32'b11111111111111110111010010110111;
assign LUT_4[19870] = 32'b11111111111111111101100001100011;
assign LUT_4[19871] = 32'b11111111111111110110101101011011;
assign LUT_4[19872] = 32'b00000000000000001000100011100111;
assign LUT_4[19873] = 32'b00000000000000000001101111011111;
assign LUT_4[19874] = 32'b00000000000000000111111110001011;
assign LUT_4[19875] = 32'b00000000000000000001001010000011;
assign LUT_4[19876] = 32'b00000000000000000101100100000011;
assign LUT_4[19877] = 32'b11111111111111111110101111111011;
assign LUT_4[19878] = 32'b00000000000000000100111110100111;
assign LUT_4[19879] = 32'b11111111111111111110001010011111;
assign LUT_4[19880] = 32'b00000000000000000001101111111100;
assign LUT_4[19881] = 32'b11111111111111111010111011110100;
assign LUT_4[19882] = 32'b00000000000000000001001010100000;
assign LUT_4[19883] = 32'b11111111111111111010010110011000;
assign LUT_4[19884] = 32'b11111111111111111110110000011000;
assign LUT_4[19885] = 32'b11111111111111110111111100010000;
assign LUT_4[19886] = 32'b11111111111111111110001010111100;
assign LUT_4[19887] = 32'b11111111111111110111010110110100;
assign LUT_4[19888] = 32'b00000000000000000110010101010101;
assign LUT_4[19889] = 32'b11111111111111111111100001001101;
assign LUT_4[19890] = 32'b00000000000000000101101111111001;
assign LUT_4[19891] = 32'b11111111111111111110111011110001;
assign LUT_4[19892] = 32'b00000000000000000011010101110001;
assign LUT_4[19893] = 32'b11111111111111111100100001101001;
assign LUT_4[19894] = 32'b00000000000000000010110000010101;
assign LUT_4[19895] = 32'b11111111111111111011111100001101;
assign LUT_4[19896] = 32'b11111111111111111111100001101010;
assign LUT_4[19897] = 32'b11111111111111111000101101100010;
assign LUT_4[19898] = 32'b11111111111111111110111100001110;
assign LUT_4[19899] = 32'b11111111111111111000001000000110;
assign LUT_4[19900] = 32'b11111111111111111100100010000110;
assign LUT_4[19901] = 32'b11111111111111110101101101111110;
assign LUT_4[19902] = 32'b11111111111111111011111100101010;
assign LUT_4[19903] = 32'b11111111111111110101001000100010;
assign LUT_4[19904] = 32'b00000000000000001011011111110100;
assign LUT_4[19905] = 32'b00000000000000000100101011101100;
assign LUT_4[19906] = 32'b00000000000000001010111010011000;
assign LUT_4[19907] = 32'b00000000000000000100000110010000;
assign LUT_4[19908] = 32'b00000000000000001000100000010000;
assign LUT_4[19909] = 32'b00000000000000000001101100001000;
assign LUT_4[19910] = 32'b00000000000000000111111010110100;
assign LUT_4[19911] = 32'b00000000000000000001000110101100;
assign LUT_4[19912] = 32'b00000000000000000100101100001001;
assign LUT_4[19913] = 32'b11111111111111111101111000000001;
assign LUT_4[19914] = 32'b00000000000000000100000110101101;
assign LUT_4[19915] = 32'b11111111111111111101010010100101;
assign LUT_4[19916] = 32'b00000000000000000001101100100101;
assign LUT_4[19917] = 32'b11111111111111111010111000011101;
assign LUT_4[19918] = 32'b00000000000000000001000111001001;
assign LUT_4[19919] = 32'b11111111111111111010010011000001;
assign LUT_4[19920] = 32'b00000000000000001001010001100010;
assign LUT_4[19921] = 32'b00000000000000000010011101011010;
assign LUT_4[19922] = 32'b00000000000000001000101100000110;
assign LUT_4[19923] = 32'b00000000000000000001110111111110;
assign LUT_4[19924] = 32'b00000000000000000110010001111110;
assign LUT_4[19925] = 32'b11111111111111111111011101110110;
assign LUT_4[19926] = 32'b00000000000000000101101100100010;
assign LUT_4[19927] = 32'b11111111111111111110111000011010;
assign LUT_4[19928] = 32'b00000000000000000010011101110111;
assign LUT_4[19929] = 32'b11111111111111111011101001101111;
assign LUT_4[19930] = 32'b00000000000000000001111000011011;
assign LUT_4[19931] = 32'b11111111111111111011000100010011;
assign LUT_4[19932] = 32'b11111111111111111111011110010011;
assign LUT_4[19933] = 32'b11111111111111111000101010001011;
assign LUT_4[19934] = 32'b11111111111111111110111000110111;
assign LUT_4[19935] = 32'b11111111111111111000000100101111;
assign LUT_4[19936] = 32'b00000000000000001001111010111011;
assign LUT_4[19937] = 32'b00000000000000000011000110110011;
assign LUT_4[19938] = 32'b00000000000000001001010101011111;
assign LUT_4[19939] = 32'b00000000000000000010100001010111;
assign LUT_4[19940] = 32'b00000000000000000110111011010111;
assign LUT_4[19941] = 32'b00000000000000000000000111001111;
assign LUT_4[19942] = 32'b00000000000000000110010101111011;
assign LUT_4[19943] = 32'b11111111111111111111100001110011;
assign LUT_4[19944] = 32'b00000000000000000011000111010000;
assign LUT_4[19945] = 32'b11111111111111111100010011001000;
assign LUT_4[19946] = 32'b00000000000000000010100001110100;
assign LUT_4[19947] = 32'b11111111111111111011101101101100;
assign LUT_4[19948] = 32'b00000000000000000000000111101100;
assign LUT_4[19949] = 32'b11111111111111111001010011100100;
assign LUT_4[19950] = 32'b11111111111111111111100010010000;
assign LUT_4[19951] = 32'b11111111111111111000101110001000;
assign LUT_4[19952] = 32'b00000000000000000111101100101001;
assign LUT_4[19953] = 32'b00000000000000000000111000100001;
assign LUT_4[19954] = 32'b00000000000000000111000111001101;
assign LUT_4[19955] = 32'b00000000000000000000010011000101;
assign LUT_4[19956] = 32'b00000000000000000100101101000101;
assign LUT_4[19957] = 32'b11111111111111111101111000111101;
assign LUT_4[19958] = 32'b00000000000000000100000111101001;
assign LUT_4[19959] = 32'b11111111111111111101010011100001;
assign LUT_4[19960] = 32'b00000000000000000000111000111110;
assign LUT_4[19961] = 32'b11111111111111111010000100110110;
assign LUT_4[19962] = 32'b00000000000000000000010011100010;
assign LUT_4[19963] = 32'b11111111111111111001011111011010;
assign LUT_4[19964] = 32'b11111111111111111101111001011010;
assign LUT_4[19965] = 32'b11111111111111110111000101010010;
assign LUT_4[19966] = 32'b11111111111111111101010011111110;
assign LUT_4[19967] = 32'b11111111111111110110011111110110;
assign LUT_4[19968] = 32'b00000000000000000001101010111101;
assign LUT_4[19969] = 32'b11111111111111111010110110110101;
assign LUT_4[19970] = 32'b00000000000000000001000101100001;
assign LUT_4[19971] = 32'b11111111111111111010010001011001;
assign LUT_4[19972] = 32'b11111111111111111110101011011001;
assign LUT_4[19973] = 32'b11111111111111110111110111010001;
assign LUT_4[19974] = 32'b11111111111111111110000101111101;
assign LUT_4[19975] = 32'b11111111111111110111010001110101;
assign LUT_4[19976] = 32'b11111111111111111010110111010010;
assign LUT_4[19977] = 32'b11111111111111110100000011001010;
assign LUT_4[19978] = 32'b11111111111111111010010001110110;
assign LUT_4[19979] = 32'b11111111111111110011011101101110;
assign LUT_4[19980] = 32'b11111111111111110111110111101110;
assign LUT_4[19981] = 32'b11111111111111110001000011100110;
assign LUT_4[19982] = 32'b11111111111111110111010010010010;
assign LUT_4[19983] = 32'b11111111111111110000011110001010;
assign LUT_4[19984] = 32'b11111111111111111111011100101011;
assign LUT_4[19985] = 32'b11111111111111111000101000100011;
assign LUT_4[19986] = 32'b11111111111111111110110111001111;
assign LUT_4[19987] = 32'b11111111111111111000000011000111;
assign LUT_4[19988] = 32'b11111111111111111100011101000111;
assign LUT_4[19989] = 32'b11111111111111110101101000111111;
assign LUT_4[19990] = 32'b11111111111111111011110111101011;
assign LUT_4[19991] = 32'b11111111111111110101000011100011;
assign LUT_4[19992] = 32'b11111111111111111000101001000000;
assign LUT_4[19993] = 32'b11111111111111110001110100111000;
assign LUT_4[19994] = 32'b11111111111111111000000011100100;
assign LUT_4[19995] = 32'b11111111111111110001001111011100;
assign LUT_4[19996] = 32'b11111111111111110101101001011100;
assign LUT_4[19997] = 32'b11111111111111101110110101010100;
assign LUT_4[19998] = 32'b11111111111111110101000100000000;
assign LUT_4[19999] = 32'b11111111111111101110001111111000;
assign LUT_4[20000] = 32'b00000000000000000000000110000100;
assign LUT_4[20001] = 32'b11111111111111111001010001111100;
assign LUT_4[20002] = 32'b11111111111111111111100000101000;
assign LUT_4[20003] = 32'b11111111111111111000101100100000;
assign LUT_4[20004] = 32'b11111111111111111101000110100000;
assign LUT_4[20005] = 32'b11111111111111110110010010011000;
assign LUT_4[20006] = 32'b11111111111111111100100001000100;
assign LUT_4[20007] = 32'b11111111111111110101101100111100;
assign LUT_4[20008] = 32'b11111111111111111001010010011001;
assign LUT_4[20009] = 32'b11111111111111110010011110010001;
assign LUT_4[20010] = 32'b11111111111111111000101100111101;
assign LUT_4[20011] = 32'b11111111111111110001111000110101;
assign LUT_4[20012] = 32'b11111111111111110110010010110101;
assign LUT_4[20013] = 32'b11111111111111101111011110101101;
assign LUT_4[20014] = 32'b11111111111111110101101101011001;
assign LUT_4[20015] = 32'b11111111111111101110111001010001;
assign LUT_4[20016] = 32'b11111111111111111101110111110010;
assign LUT_4[20017] = 32'b11111111111111110111000011101010;
assign LUT_4[20018] = 32'b11111111111111111101010010010110;
assign LUT_4[20019] = 32'b11111111111111110110011110001110;
assign LUT_4[20020] = 32'b11111111111111111010111000001110;
assign LUT_4[20021] = 32'b11111111111111110100000100000110;
assign LUT_4[20022] = 32'b11111111111111111010010010110010;
assign LUT_4[20023] = 32'b11111111111111110011011110101010;
assign LUT_4[20024] = 32'b11111111111111110111000100000111;
assign LUT_4[20025] = 32'b11111111111111110000001111111111;
assign LUT_4[20026] = 32'b11111111111111110110011110101011;
assign LUT_4[20027] = 32'b11111111111111101111101010100011;
assign LUT_4[20028] = 32'b11111111111111110100000100100011;
assign LUT_4[20029] = 32'b11111111111111101101010000011011;
assign LUT_4[20030] = 32'b11111111111111110011011111000111;
assign LUT_4[20031] = 32'b11111111111111101100101010111111;
assign LUT_4[20032] = 32'b00000000000000000011000010010001;
assign LUT_4[20033] = 32'b11111111111111111100001110001001;
assign LUT_4[20034] = 32'b00000000000000000010011100110101;
assign LUT_4[20035] = 32'b11111111111111111011101000101101;
assign LUT_4[20036] = 32'b00000000000000000000000010101101;
assign LUT_4[20037] = 32'b11111111111111111001001110100101;
assign LUT_4[20038] = 32'b11111111111111111111011101010001;
assign LUT_4[20039] = 32'b11111111111111111000101001001001;
assign LUT_4[20040] = 32'b11111111111111111100001110100110;
assign LUT_4[20041] = 32'b11111111111111110101011010011110;
assign LUT_4[20042] = 32'b11111111111111111011101001001010;
assign LUT_4[20043] = 32'b11111111111111110100110101000010;
assign LUT_4[20044] = 32'b11111111111111111001001111000010;
assign LUT_4[20045] = 32'b11111111111111110010011010111010;
assign LUT_4[20046] = 32'b11111111111111111000101001100110;
assign LUT_4[20047] = 32'b11111111111111110001110101011110;
assign LUT_4[20048] = 32'b00000000000000000000110011111111;
assign LUT_4[20049] = 32'b11111111111111111001111111110111;
assign LUT_4[20050] = 32'b00000000000000000000001110100011;
assign LUT_4[20051] = 32'b11111111111111111001011010011011;
assign LUT_4[20052] = 32'b11111111111111111101110100011011;
assign LUT_4[20053] = 32'b11111111111111110111000000010011;
assign LUT_4[20054] = 32'b11111111111111111101001110111111;
assign LUT_4[20055] = 32'b11111111111111110110011010110111;
assign LUT_4[20056] = 32'b11111111111111111010000000010100;
assign LUT_4[20057] = 32'b11111111111111110011001100001100;
assign LUT_4[20058] = 32'b11111111111111111001011010111000;
assign LUT_4[20059] = 32'b11111111111111110010100110110000;
assign LUT_4[20060] = 32'b11111111111111110111000000110000;
assign LUT_4[20061] = 32'b11111111111111110000001100101000;
assign LUT_4[20062] = 32'b11111111111111110110011011010100;
assign LUT_4[20063] = 32'b11111111111111101111100111001100;
assign LUT_4[20064] = 32'b00000000000000000001011101011000;
assign LUT_4[20065] = 32'b11111111111111111010101001010000;
assign LUT_4[20066] = 32'b00000000000000000000110111111100;
assign LUT_4[20067] = 32'b11111111111111111010000011110100;
assign LUT_4[20068] = 32'b11111111111111111110011101110100;
assign LUT_4[20069] = 32'b11111111111111110111101001101100;
assign LUT_4[20070] = 32'b11111111111111111101111000011000;
assign LUT_4[20071] = 32'b11111111111111110111000100010000;
assign LUT_4[20072] = 32'b11111111111111111010101001101101;
assign LUT_4[20073] = 32'b11111111111111110011110101100101;
assign LUT_4[20074] = 32'b11111111111111111010000100010001;
assign LUT_4[20075] = 32'b11111111111111110011010000001001;
assign LUT_4[20076] = 32'b11111111111111110111101010001001;
assign LUT_4[20077] = 32'b11111111111111110000110110000001;
assign LUT_4[20078] = 32'b11111111111111110111000100101101;
assign LUT_4[20079] = 32'b11111111111111110000010000100101;
assign LUT_4[20080] = 32'b11111111111111111111001111000110;
assign LUT_4[20081] = 32'b11111111111111111000011010111110;
assign LUT_4[20082] = 32'b11111111111111111110101001101010;
assign LUT_4[20083] = 32'b11111111111111110111110101100010;
assign LUT_4[20084] = 32'b11111111111111111100001111100010;
assign LUT_4[20085] = 32'b11111111111111110101011011011010;
assign LUT_4[20086] = 32'b11111111111111111011101010000110;
assign LUT_4[20087] = 32'b11111111111111110100110101111110;
assign LUT_4[20088] = 32'b11111111111111111000011011011011;
assign LUT_4[20089] = 32'b11111111111111110001100111010011;
assign LUT_4[20090] = 32'b11111111111111110111110101111111;
assign LUT_4[20091] = 32'b11111111111111110001000001110111;
assign LUT_4[20092] = 32'b11111111111111110101011011110111;
assign LUT_4[20093] = 32'b11111111111111101110100111101111;
assign LUT_4[20094] = 32'b11111111111111110100110110011011;
assign LUT_4[20095] = 32'b11111111111111101110000010010011;
assign LUT_4[20096] = 32'b00000000000000000100010001000101;
assign LUT_4[20097] = 32'b11111111111111111101011100111101;
assign LUT_4[20098] = 32'b00000000000000000011101011101001;
assign LUT_4[20099] = 32'b11111111111111111100110111100001;
assign LUT_4[20100] = 32'b00000000000000000001010001100001;
assign LUT_4[20101] = 32'b11111111111111111010011101011001;
assign LUT_4[20102] = 32'b00000000000000000000101100000101;
assign LUT_4[20103] = 32'b11111111111111111001110111111101;
assign LUT_4[20104] = 32'b11111111111111111101011101011010;
assign LUT_4[20105] = 32'b11111111111111110110101001010010;
assign LUT_4[20106] = 32'b11111111111111111100110111111110;
assign LUT_4[20107] = 32'b11111111111111110110000011110110;
assign LUT_4[20108] = 32'b11111111111111111010011101110110;
assign LUT_4[20109] = 32'b11111111111111110011101001101110;
assign LUT_4[20110] = 32'b11111111111111111001111000011010;
assign LUT_4[20111] = 32'b11111111111111110011000100010010;
assign LUT_4[20112] = 32'b00000000000000000010000010110011;
assign LUT_4[20113] = 32'b11111111111111111011001110101011;
assign LUT_4[20114] = 32'b00000000000000000001011101010111;
assign LUT_4[20115] = 32'b11111111111111111010101001001111;
assign LUT_4[20116] = 32'b11111111111111111111000011001111;
assign LUT_4[20117] = 32'b11111111111111111000001111000111;
assign LUT_4[20118] = 32'b11111111111111111110011101110011;
assign LUT_4[20119] = 32'b11111111111111110111101001101011;
assign LUT_4[20120] = 32'b11111111111111111011001111001000;
assign LUT_4[20121] = 32'b11111111111111110100011011000000;
assign LUT_4[20122] = 32'b11111111111111111010101001101100;
assign LUT_4[20123] = 32'b11111111111111110011110101100100;
assign LUT_4[20124] = 32'b11111111111111111000001111100100;
assign LUT_4[20125] = 32'b11111111111111110001011011011100;
assign LUT_4[20126] = 32'b11111111111111110111101010001000;
assign LUT_4[20127] = 32'b11111111111111110000110110000000;
assign LUT_4[20128] = 32'b00000000000000000010101100001100;
assign LUT_4[20129] = 32'b11111111111111111011111000000100;
assign LUT_4[20130] = 32'b00000000000000000010000110110000;
assign LUT_4[20131] = 32'b11111111111111111011010010101000;
assign LUT_4[20132] = 32'b11111111111111111111101100101000;
assign LUT_4[20133] = 32'b11111111111111111000111000100000;
assign LUT_4[20134] = 32'b11111111111111111111000111001100;
assign LUT_4[20135] = 32'b11111111111111111000010011000100;
assign LUT_4[20136] = 32'b11111111111111111011111000100001;
assign LUT_4[20137] = 32'b11111111111111110101000100011001;
assign LUT_4[20138] = 32'b11111111111111111011010011000101;
assign LUT_4[20139] = 32'b11111111111111110100011110111101;
assign LUT_4[20140] = 32'b11111111111111111000111000111101;
assign LUT_4[20141] = 32'b11111111111111110010000100110101;
assign LUT_4[20142] = 32'b11111111111111111000010011100001;
assign LUT_4[20143] = 32'b11111111111111110001011111011001;
assign LUT_4[20144] = 32'b00000000000000000000011101111010;
assign LUT_4[20145] = 32'b11111111111111111001101001110010;
assign LUT_4[20146] = 32'b11111111111111111111111000011110;
assign LUT_4[20147] = 32'b11111111111111111001000100010110;
assign LUT_4[20148] = 32'b11111111111111111101011110010110;
assign LUT_4[20149] = 32'b11111111111111110110101010001110;
assign LUT_4[20150] = 32'b11111111111111111100111000111010;
assign LUT_4[20151] = 32'b11111111111111110110000100110010;
assign LUT_4[20152] = 32'b11111111111111111001101010001111;
assign LUT_4[20153] = 32'b11111111111111110010110110000111;
assign LUT_4[20154] = 32'b11111111111111111001000100110011;
assign LUT_4[20155] = 32'b11111111111111110010010000101011;
assign LUT_4[20156] = 32'b11111111111111110110101010101011;
assign LUT_4[20157] = 32'b11111111111111101111110110100011;
assign LUT_4[20158] = 32'b11111111111111110110000101001111;
assign LUT_4[20159] = 32'b11111111111111101111010001000111;
assign LUT_4[20160] = 32'b00000000000000000101101000011001;
assign LUT_4[20161] = 32'b11111111111111111110110100010001;
assign LUT_4[20162] = 32'b00000000000000000101000010111101;
assign LUT_4[20163] = 32'b11111111111111111110001110110101;
assign LUT_4[20164] = 32'b00000000000000000010101000110101;
assign LUT_4[20165] = 32'b11111111111111111011110100101101;
assign LUT_4[20166] = 32'b00000000000000000010000011011001;
assign LUT_4[20167] = 32'b11111111111111111011001111010001;
assign LUT_4[20168] = 32'b11111111111111111110110100101110;
assign LUT_4[20169] = 32'b11111111111111111000000000100110;
assign LUT_4[20170] = 32'b11111111111111111110001111010010;
assign LUT_4[20171] = 32'b11111111111111110111011011001010;
assign LUT_4[20172] = 32'b11111111111111111011110101001010;
assign LUT_4[20173] = 32'b11111111111111110101000001000010;
assign LUT_4[20174] = 32'b11111111111111111011001111101110;
assign LUT_4[20175] = 32'b11111111111111110100011011100110;
assign LUT_4[20176] = 32'b00000000000000000011011010000111;
assign LUT_4[20177] = 32'b11111111111111111100100101111111;
assign LUT_4[20178] = 32'b00000000000000000010110100101011;
assign LUT_4[20179] = 32'b11111111111111111100000000100011;
assign LUT_4[20180] = 32'b00000000000000000000011010100011;
assign LUT_4[20181] = 32'b11111111111111111001100110011011;
assign LUT_4[20182] = 32'b11111111111111111111110101000111;
assign LUT_4[20183] = 32'b11111111111111111001000000111111;
assign LUT_4[20184] = 32'b11111111111111111100100110011100;
assign LUT_4[20185] = 32'b11111111111111110101110010010100;
assign LUT_4[20186] = 32'b11111111111111111100000001000000;
assign LUT_4[20187] = 32'b11111111111111110101001100111000;
assign LUT_4[20188] = 32'b11111111111111111001100110111000;
assign LUT_4[20189] = 32'b11111111111111110010110010110000;
assign LUT_4[20190] = 32'b11111111111111111001000001011100;
assign LUT_4[20191] = 32'b11111111111111110010001101010100;
assign LUT_4[20192] = 32'b00000000000000000100000011100000;
assign LUT_4[20193] = 32'b11111111111111111101001111011000;
assign LUT_4[20194] = 32'b00000000000000000011011110000100;
assign LUT_4[20195] = 32'b11111111111111111100101001111100;
assign LUT_4[20196] = 32'b00000000000000000001000011111100;
assign LUT_4[20197] = 32'b11111111111111111010001111110100;
assign LUT_4[20198] = 32'b00000000000000000000011110100000;
assign LUT_4[20199] = 32'b11111111111111111001101010011000;
assign LUT_4[20200] = 32'b11111111111111111101001111110101;
assign LUT_4[20201] = 32'b11111111111111110110011011101101;
assign LUT_4[20202] = 32'b11111111111111111100101010011001;
assign LUT_4[20203] = 32'b11111111111111110101110110010001;
assign LUT_4[20204] = 32'b11111111111111111010010000010001;
assign LUT_4[20205] = 32'b11111111111111110011011100001001;
assign LUT_4[20206] = 32'b11111111111111111001101010110101;
assign LUT_4[20207] = 32'b11111111111111110010110110101101;
assign LUT_4[20208] = 32'b00000000000000000001110101001110;
assign LUT_4[20209] = 32'b11111111111111111011000001000110;
assign LUT_4[20210] = 32'b00000000000000000001001111110010;
assign LUT_4[20211] = 32'b11111111111111111010011011101010;
assign LUT_4[20212] = 32'b11111111111111111110110101101010;
assign LUT_4[20213] = 32'b11111111111111111000000001100010;
assign LUT_4[20214] = 32'b11111111111111111110010000001110;
assign LUT_4[20215] = 32'b11111111111111110111011100000110;
assign LUT_4[20216] = 32'b11111111111111111011000001100011;
assign LUT_4[20217] = 32'b11111111111111110100001101011011;
assign LUT_4[20218] = 32'b11111111111111111010011100000111;
assign LUT_4[20219] = 32'b11111111111111110011100111111111;
assign LUT_4[20220] = 32'b11111111111111111000000001111111;
assign LUT_4[20221] = 32'b11111111111111110001001101110111;
assign LUT_4[20222] = 32'b11111111111111110111011100100011;
assign LUT_4[20223] = 32'b11111111111111110000101000011011;
assign LUT_4[20224] = 32'b00000000000000000110100110100000;
assign LUT_4[20225] = 32'b11111111111111111111110010011000;
assign LUT_4[20226] = 32'b00000000000000000110000001000100;
assign LUT_4[20227] = 32'b11111111111111111111001100111100;
assign LUT_4[20228] = 32'b00000000000000000011100110111100;
assign LUT_4[20229] = 32'b11111111111111111100110010110100;
assign LUT_4[20230] = 32'b00000000000000000011000001100000;
assign LUT_4[20231] = 32'b11111111111111111100001101011000;
assign LUT_4[20232] = 32'b11111111111111111111110010110101;
assign LUT_4[20233] = 32'b11111111111111111000111110101101;
assign LUT_4[20234] = 32'b11111111111111111111001101011001;
assign LUT_4[20235] = 32'b11111111111111111000011001010001;
assign LUT_4[20236] = 32'b11111111111111111100110011010001;
assign LUT_4[20237] = 32'b11111111111111110101111111001001;
assign LUT_4[20238] = 32'b11111111111111111100001101110101;
assign LUT_4[20239] = 32'b11111111111111110101011001101101;
assign LUT_4[20240] = 32'b00000000000000000100011000001110;
assign LUT_4[20241] = 32'b11111111111111111101100100000110;
assign LUT_4[20242] = 32'b00000000000000000011110010110010;
assign LUT_4[20243] = 32'b11111111111111111100111110101010;
assign LUT_4[20244] = 32'b00000000000000000001011000101010;
assign LUT_4[20245] = 32'b11111111111111111010100100100010;
assign LUT_4[20246] = 32'b00000000000000000000110011001110;
assign LUT_4[20247] = 32'b11111111111111111001111111000110;
assign LUT_4[20248] = 32'b11111111111111111101100100100011;
assign LUT_4[20249] = 32'b11111111111111110110110000011011;
assign LUT_4[20250] = 32'b11111111111111111100111111000111;
assign LUT_4[20251] = 32'b11111111111111110110001010111111;
assign LUT_4[20252] = 32'b11111111111111111010100100111111;
assign LUT_4[20253] = 32'b11111111111111110011110000110111;
assign LUT_4[20254] = 32'b11111111111111111001111111100011;
assign LUT_4[20255] = 32'b11111111111111110011001011011011;
assign LUT_4[20256] = 32'b00000000000000000101000001100111;
assign LUT_4[20257] = 32'b11111111111111111110001101011111;
assign LUT_4[20258] = 32'b00000000000000000100011100001011;
assign LUT_4[20259] = 32'b11111111111111111101101000000011;
assign LUT_4[20260] = 32'b00000000000000000010000010000011;
assign LUT_4[20261] = 32'b11111111111111111011001101111011;
assign LUT_4[20262] = 32'b00000000000000000001011100100111;
assign LUT_4[20263] = 32'b11111111111111111010101000011111;
assign LUT_4[20264] = 32'b11111111111111111110001101111100;
assign LUT_4[20265] = 32'b11111111111111110111011001110100;
assign LUT_4[20266] = 32'b11111111111111111101101000100000;
assign LUT_4[20267] = 32'b11111111111111110110110100011000;
assign LUT_4[20268] = 32'b11111111111111111011001110011000;
assign LUT_4[20269] = 32'b11111111111111110100011010010000;
assign LUT_4[20270] = 32'b11111111111111111010101000111100;
assign LUT_4[20271] = 32'b11111111111111110011110100110100;
assign LUT_4[20272] = 32'b00000000000000000010110011010101;
assign LUT_4[20273] = 32'b11111111111111111011111111001101;
assign LUT_4[20274] = 32'b00000000000000000010001101111001;
assign LUT_4[20275] = 32'b11111111111111111011011001110001;
assign LUT_4[20276] = 32'b11111111111111111111110011110001;
assign LUT_4[20277] = 32'b11111111111111111000111111101001;
assign LUT_4[20278] = 32'b11111111111111111111001110010101;
assign LUT_4[20279] = 32'b11111111111111111000011010001101;
assign LUT_4[20280] = 32'b11111111111111111011111111101010;
assign LUT_4[20281] = 32'b11111111111111110101001011100010;
assign LUT_4[20282] = 32'b11111111111111111011011010001110;
assign LUT_4[20283] = 32'b11111111111111110100100110000110;
assign LUT_4[20284] = 32'b11111111111111111001000000000110;
assign LUT_4[20285] = 32'b11111111111111110010001011111110;
assign LUT_4[20286] = 32'b11111111111111111000011010101010;
assign LUT_4[20287] = 32'b11111111111111110001100110100010;
assign LUT_4[20288] = 32'b00000000000000000111111101110100;
assign LUT_4[20289] = 32'b00000000000000000001001001101100;
assign LUT_4[20290] = 32'b00000000000000000111011000011000;
assign LUT_4[20291] = 32'b00000000000000000000100100010000;
assign LUT_4[20292] = 32'b00000000000000000100111110010000;
assign LUT_4[20293] = 32'b11111111111111111110001010001000;
assign LUT_4[20294] = 32'b00000000000000000100011000110100;
assign LUT_4[20295] = 32'b11111111111111111101100100101100;
assign LUT_4[20296] = 32'b00000000000000000001001010001001;
assign LUT_4[20297] = 32'b11111111111111111010010110000001;
assign LUT_4[20298] = 32'b00000000000000000000100100101101;
assign LUT_4[20299] = 32'b11111111111111111001110000100101;
assign LUT_4[20300] = 32'b11111111111111111110001010100101;
assign LUT_4[20301] = 32'b11111111111111110111010110011101;
assign LUT_4[20302] = 32'b11111111111111111101100101001001;
assign LUT_4[20303] = 32'b11111111111111110110110001000001;
assign LUT_4[20304] = 32'b00000000000000000101101111100010;
assign LUT_4[20305] = 32'b11111111111111111110111011011010;
assign LUT_4[20306] = 32'b00000000000000000101001010000110;
assign LUT_4[20307] = 32'b11111111111111111110010101111110;
assign LUT_4[20308] = 32'b00000000000000000010101111111110;
assign LUT_4[20309] = 32'b11111111111111111011111011110110;
assign LUT_4[20310] = 32'b00000000000000000010001010100010;
assign LUT_4[20311] = 32'b11111111111111111011010110011010;
assign LUT_4[20312] = 32'b11111111111111111110111011110111;
assign LUT_4[20313] = 32'b11111111111111111000000111101111;
assign LUT_4[20314] = 32'b11111111111111111110010110011011;
assign LUT_4[20315] = 32'b11111111111111110111100010010011;
assign LUT_4[20316] = 32'b11111111111111111011111100010011;
assign LUT_4[20317] = 32'b11111111111111110101001000001011;
assign LUT_4[20318] = 32'b11111111111111111011010110110111;
assign LUT_4[20319] = 32'b11111111111111110100100010101111;
assign LUT_4[20320] = 32'b00000000000000000110011000111011;
assign LUT_4[20321] = 32'b11111111111111111111100100110011;
assign LUT_4[20322] = 32'b00000000000000000101110011011111;
assign LUT_4[20323] = 32'b11111111111111111110111111010111;
assign LUT_4[20324] = 32'b00000000000000000011011001010111;
assign LUT_4[20325] = 32'b11111111111111111100100101001111;
assign LUT_4[20326] = 32'b00000000000000000010110011111011;
assign LUT_4[20327] = 32'b11111111111111111011111111110011;
assign LUT_4[20328] = 32'b11111111111111111111100101010000;
assign LUT_4[20329] = 32'b11111111111111111000110001001000;
assign LUT_4[20330] = 32'b11111111111111111110111111110100;
assign LUT_4[20331] = 32'b11111111111111111000001011101100;
assign LUT_4[20332] = 32'b11111111111111111100100101101100;
assign LUT_4[20333] = 32'b11111111111111110101110001100100;
assign LUT_4[20334] = 32'b11111111111111111100000000010000;
assign LUT_4[20335] = 32'b11111111111111110101001100001000;
assign LUT_4[20336] = 32'b00000000000000000100001010101001;
assign LUT_4[20337] = 32'b11111111111111111101010110100001;
assign LUT_4[20338] = 32'b00000000000000000011100101001101;
assign LUT_4[20339] = 32'b11111111111111111100110001000101;
assign LUT_4[20340] = 32'b00000000000000000001001011000101;
assign LUT_4[20341] = 32'b11111111111111111010010110111101;
assign LUT_4[20342] = 32'b00000000000000000000100101101001;
assign LUT_4[20343] = 32'b11111111111111111001110001100001;
assign LUT_4[20344] = 32'b11111111111111111101010110111110;
assign LUT_4[20345] = 32'b11111111111111110110100010110110;
assign LUT_4[20346] = 32'b11111111111111111100110001100010;
assign LUT_4[20347] = 32'b11111111111111110101111101011010;
assign LUT_4[20348] = 32'b11111111111111111010010111011010;
assign LUT_4[20349] = 32'b11111111111111110011100011010010;
assign LUT_4[20350] = 32'b11111111111111111001110001111110;
assign LUT_4[20351] = 32'b11111111111111110010111101110110;
assign LUT_4[20352] = 32'b00000000000000001001001100101000;
assign LUT_4[20353] = 32'b00000000000000000010011000100000;
assign LUT_4[20354] = 32'b00000000000000001000100111001100;
assign LUT_4[20355] = 32'b00000000000000000001110011000100;
assign LUT_4[20356] = 32'b00000000000000000110001101000100;
assign LUT_4[20357] = 32'b11111111111111111111011000111100;
assign LUT_4[20358] = 32'b00000000000000000101100111101000;
assign LUT_4[20359] = 32'b11111111111111111110110011100000;
assign LUT_4[20360] = 32'b00000000000000000010011000111101;
assign LUT_4[20361] = 32'b11111111111111111011100100110101;
assign LUT_4[20362] = 32'b00000000000000000001110011100001;
assign LUT_4[20363] = 32'b11111111111111111010111111011001;
assign LUT_4[20364] = 32'b11111111111111111111011001011001;
assign LUT_4[20365] = 32'b11111111111111111000100101010001;
assign LUT_4[20366] = 32'b11111111111111111110110011111101;
assign LUT_4[20367] = 32'b11111111111111110111111111110101;
assign LUT_4[20368] = 32'b00000000000000000110111110010110;
assign LUT_4[20369] = 32'b00000000000000000000001010001110;
assign LUT_4[20370] = 32'b00000000000000000110011000111010;
assign LUT_4[20371] = 32'b11111111111111111111100100110010;
assign LUT_4[20372] = 32'b00000000000000000011111110110010;
assign LUT_4[20373] = 32'b11111111111111111101001010101010;
assign LUT_4[20374] = 32'b00000000000000000011011001010110;
assign LUT_4[20375] = 32'b11111111111111111100100101001110;
assign LUT_4[20376] = 32'b00000000000000000000001010101011;
assign LUT_4[20377] = 32'b11111111111111111001010110100011;
assign LUT_4[20378] = 32'b11111111111111111111100101001111;
assign LUT_4[20379] = 32'b11111111111111111000110001000111;
assign LUT_4[20380] = 32'b11111111111111111101001011000111;
assign LUT_4[20381] = 32'b11111111111111110110010110111111;
assign LUT_4[20382] = 32'b11111111111111111100100101101011;
assign LUT_4[20383] = 32'b11111111111111110101110001100011;
assign LUT_4[20384] = 32'b00000000000000000111100111101111;
assign LUT_4[20385] = 32'b00000000000000000000110011100111;
assign LUT_4[20386] = 32'b00000000000000000111000010010011;
assign LUT_4[20387] = 32'b00000000000000000000001110001011;
assign LUT_4[20388] = 32'b00000000000000000100101000001011;
assign LUT_4[20389] = 32'b11111111111111111101110100000011;
assign LUT_4[20390] = 32'b00000000000000000100000010101111;
assign LUT_4[20391] = 32'b11111111111111111101001110100111;
assign LUT_4[20392] = 32'b00000000000000000000110100000100;
assign LUT_4[20393] = 32'b11111111111111111001111111111100;
assign LUT_4[20394] = 32'b00000000000000000000001110101000;
assign LUT_4[20395] = 32'b11111111111111111001011010100000;
assign LUT_4[20396] = 32'b11111111111111111101110100100000;
assign LUT_4[20397] = 32'b11111111111111110111000000011000;
assign LUT_4[20398] = 32'b11111111111111111101001111000100;
assign LUT_4[20399] = 32'b11111111111111110110011010111100;
assign LUT_4[20400] = 32'b00000000000000000101011001011101;
assign LUT_4[20401] = 32'b11111111111111111110100101010101;
assign LUT_4[20402] = 32'b00000000000000000100110100000001;
assign LUT_4[20403] = 32'b11111111111111111101111111111001;
assign LUT_4[20404] = 32'b00000000000000000010011001111001;
assign LUT_4[20405] = 32'b11111111111111111011100101110001;
assign LUT_4[20406] = 32'b00000000000000000001110100011101;
assign LUT_4[20407] = 32'b11111111111111111011000000010101;
assign LUT_4[20408] = 32'b11111111111111111110100101110010;
assign LUT_4[20409] = 32'b11111111111111110111110001101010;
assign LUT_4[20410] = 32'b11111111111111111110000000010110;
assign LUT_4[20411] = 32'b11111111111111110111001100001110;
assign LUT_4[20412] = 32'b11111111111111111011100110001110;
assign LUT_4[20413] = 32'b11111111111111110100110010000110;
assign LUT_4[20414] = 32'b11111111111111111011000000110010;
assign LUT_4[20415] = 32'b11111111111111110100001100101010;
assign LUT_4[20416] = 32'b00000000000000001010100011111100;
assign LUT_4[20417] = 32'b00000000000000000011101111110100;
assign LUT_4[20418] = 32'b00000000000000001001111110100000;
assign LUT_4[20419] = 32'b00000000000000000011001010011000;
assign LUT_4[20420] = 32'b00000000000000000111100100011000;
assign LUT_4[20421] = 32'b00000000000000000000110000010000;
assign LUT_4[20422] = 32'b00000000000000000110111110111100;
assign LUT_4[20423] = 32'b00000000000000000000001010110100;
assign LUT_4[20424] = 32'b00000000000000000011110000010001;
assign LUT_4[20425] = 32'b11111111111111111100111100001001;
assign LUT_4[20426] = 32'b00000000000000000011001010110101;
assign LUT_4[20427] = 32'b11111111111111111100010110101101;
assign LUT_4[20428] = 32'b00000000000000000000110000101101;
assign LUT_4[20429] = 32'b11111111111111111001111100100101;
assign LUT_4[20430] = 32'b00000000000000000000001011010001;
assign LUT_4[20431] = 32'b11111111111111111001010111001001;
assign LUT_4[20432] = 32'b00000000000000001000010101101010;
assign LUT_4[20433] = 32'b00000000000000000001100001100010;
assign LUT_4[20434] = 32'b00000000000000000111110000001110;
assign LUT_4[20435] = 32'b00000000000000000000111100000110;
assign LUT_4[20436] = 32'b00000000000000000101010110000110;
assign LUT_4[20437] = 32'b11111111111111111110100001111110;
assign LUT_4[20438] = 32'b00000000000000000100110000101010;
assign LUT_4[20439] = 32'b11111111111111111101111100100010;
assign LUT_4[20440] = 32'b00000000000000000001100001111111;
assign LUT_4[20441] = 32'b11111111111111111010101101110111;
assign LUT_4[20442] = 32'b00000000000000000000111100100011;
assign LUT_4[20443] = 32'b11111111111111111010001000011011;
assign LUT_4[20444] = 32'b11111111111111111110100010011011;
assign LUT_4[20445] = 32'b11111111111111110111101110010011;
assign LUT_4[20446] = 32'b11111111111111111101111100111111;
assign LUT_4[20447] = 32'b11111111111111110111001000110111;
assign LUT_4[20448] = 32'b00000000000000001000111111000011;
assign LUT_4[20449] = 32'b00000000000000000010001010111011;
assign LUT_4[20450] = 32'b00000000000000001000011001100111;
assign LUT_4[20451] = 32'b00000000000000000001100101011111;
assign LUT_4[20452] = 32'b00000000000000000101111111011111;
assign LUT_4[20453] = 32'b11111111111111111111001011010111;
assign LUT_4[20454] = 32'b00000000000000000101011010000011;
assign LUT_4[20455] = 32'b11111111111111111110100101111011;
assign LUT_4[20456] = 32'b00000000000000000010001011011000;
assign LUT_4[20457] = 32'b11111111111111111011010111010000;
assign LUT_4[20458] = 32'b00000000000000000001100101111100;
assign LUT_4[20459] = 32'b11111111111111111010110001110100;
assign LUT_4[20460] = 32'b11111111111111111111001011110100;
assign LUT_4[20461] = 32'b11111111111111111000010111101100;
assign LUT_4[20462] = 32'b11111111111111111110100110011000;
assign LUT_4[20463] = 32'b11111111111111110111110010010000;
assign LUT_4[20464] = 32'b00000000000000000110110000110001;
assign LUT_4[20465] = 32'b11111111111111111111111100101001;
assign LUT_4[20466] = 32'b00000000000000000110001011010101;
assign LUT_4[20467] = 32'b11111111111111111111010111001101;
assign LUT_4[20468] = 32'b00000000000000000011110001001101;
assign LUT_4[20469] = 32'b11111111111111111100111101000101;
assign LUT_4[20470] = 32'b00000000000000000011001011110001;
assign LUT_4[20471] = 32'b11111111111111111100010111101001;
assign LUT_4[20472] = 32'b11111111111111111111111101000110;
assign LUT_4[20473] = 32'b11111111111111111001001000111110;
assign LUT_4[20474] = 32'b11111111111111111111010111101010;
assign LUT_4[20475] = 32'b11111111111111111000100011100010;
assign LUT_4[20476] = 32'b11111111111111111100111101100010;
assign LUT_4[20477] = 32'b11111111111111110110001001011010;
assign LUT_4[20478] = 32'b11111111111111111100011000000110;
assign LUT_4[20479] = 32'b11111111111111110101100011111110;
assign LUT_4[20480] = 32'b00000000000000000001101100111101;
assign LUT_4[20481] = 32'b11111111111111111010111000110101;
assign LUT_4[20482] = 32'b00000000000000000001000111100001;
assign LUT_4[20483] = 32'b11111111111111111010010011011001;
assign LUT_4[20484] = 32'b11111111111111111110101101011001;
assign LUT_4[20485] = 32'b11111111111111110111111001010001;
assign LUT_4[20486] = 32'b11111111111111111110000111111101;
assign LUT_4[20487] = 32'b11111111111111110111010011110101;
assign LUT_4[20488] = 32'b11111111111111111010111001010010;
assign LUT_4[20489] = 32'b11111111111111110100000101001010;
assign LUT_4[20490] = 32'b11111111111111111010010011110110;
assign LUT_4[20491] = 32'b11111111111111110011011111101110;
assign LUT_4[20492] = 32'b11111111111111110111111001101110;
assign LUT_4[20493] = 32'b11111111111111110001000101100110;
assign LUT_4[20494] = 32'b11111111111111110111010100010010;
assign LUT_4[20495] = 32'b11111111111111110000100000001010;
assign LUT_4[20496] = 32'b11111111111111111111011110101011;
assign LUT_4[20497] = 32'b11111111111111111000101010100011;
assign LUT_4[20498] = 32'b11111111111111111110111001001111;
assign LUT_4[20499] = 32'b11111111111111111000000101000111;
assign LUT_4[20500] = 32'b11111111111111111100011111000111;
assign LUT_4[20501] = 32'b11111111111111110101101010111111;
assign LUT_4[20502] = 32'b11111111111111111011111001101011;
assign LUT_4[20503] = 32'b11111111111111110101000101100011;
assign LUT_4[20504] = 32'b11111111111111111000101011000000;
assign LUT_4[20505] = 32'b11111111111111110001110110111000;
assign LUT_4[20506] = 32'b11111111111111111000000101100100;
assign LUT_4[20507] = 32'b11111111111111110001010001011100;
assign LUT_4[20508] = 32'b11111111111111110101101011011100;
assign LUT_4[20509] = 32'b11111111111111101110110111010100;
assign LUT_4[20510] = 32'b11111111111111110101000110000000;
assign LUT_4[20511] = 32'b11111111111111101110010001111000;
assign LUT_4[20512] = 32'b00000000000000000000001000000100;
assign LUT_4[20513] = 32'b11111111111111111001010011111100;
assign LUT_4[20514] = 32'b11111111111111111111100010101000;
assign LUT_4[20515] = 32'b11111111111111111000101110100000;
assign LUT_4[20516] = 32'b11111111111111111101001000100000;
assign LUT_4[20517] = 32'b11111111111111110110010100011000;
assign LUT_4[20518] = 32'b11111111111111111100100011000100;
assign LUT_4[20519] = 32'b11111111111111110101101110111100;
assign LUT_4[20520] = 32'b11111111111111111001010100011001;
assign LUT_4[20521] = 32'b11111111111111110010100000010001;
assign LUT_4[20522] = 32'b11111111111111111000101110111101;
assign LUT_4[20523] = 32'b11111111111111110001111010110101;
assign LUT_4[20524] = 32'b11111111111111110110010100110101;
assign LUT_4[20525] = 32'b11111111111111101111100000101101;
assign LUT_4[20526] = 32'b11111111111111110101101111011001;
assign LUT_4[20527] = 32'b11111111111111101110111011010001;
assign LUT_4[20528] = 32'b11111111111111111101111001110010;
assign LUT_4[20529] = 32'b11111111111111110111000101101010;
assign LUT_4[20530] = 32'b11111111111111111101010100010110;
assign LUT_4[20531] = 32'b11111111111111110110100000001110;
assign LUT_4[20532] = 32'b11111111111111111010111010001110;
assign LUT_4[20533] = 32'b11111111111111110100000110000110;
assign LUT_4[20534] = 32'b11111111111111111010010100110010;
assign LUT_4[20535] = 32'b11111111111111110011100000101010;
assign LUT_4[20536] = 32'b11111111111111110111000110000111;
assign LUT_4[20537] = 32'b11111111111111110000010001111111;
assign LUT_4[20538] = 32'b11111111111111110110100000101011;
assign LUT_4[20539] = 32'b11111111111111101111101100100011;
assign LUT_4[20540] = 32'b11111111111111110100000110100011;
assign LUT_4[20541] = 32'b11111111111111101101010010011011;
assign LUT_4[20542] = 32'b11111111111111110011100001000111;
assign LUT_4[20543] = 32'b11111111111111101100101100111111;
assign LUT_4[20544] = 32'b00000000000000000011000100010001;
assign LUT_4[20545] = 32'b11111111111111111100010000001001;
assign LUT_4[20546] = 32'b00000000000000000010011110110101;
assign LUT_4[20547] = 32'b11111111111111111011101010101101;
assign LUT_4[20548] = 32'b00000000000000000000000100101101;
assign LUT_4[20549] = 32'b11111111111111111001010000100101;
assign LUT_4[20550] = 32'b11111111111111111111011111010001;
assign LUT_4[20551] = 32'b11111111111111111000101011001001;
assign LUT_4[20552] = 32'b11111111111111111100010000100110;
assign LUT_4[20553] = 32'b11111111111111110101011100011110;
assign LUT_4[20554] = 32'b11111111111111111011101011001010;
assign LUT_4[20555] = 32'b11111111111111110100110111000010;
assign LUT_4[20556] = 32'b11111111111111111001010001000010;
assign LUT_4[20557] = 32'b11111111111111110010011100111010;
assign LUT_4[20558] = 32'b11111111111111111000101011100110;
assign LUT_4[20559] = 32'b11111111111111110001110111011110;
assign LUT_4[20560] = 32'b00000000000000000000110101111111;
assign LUT_4[20561] = 32'b11111111111111111010000001110111;
assign LUT_4[20562] = 32'b00000000000000000000010000100011;
assign LUT_4[20563] = 32'b11111111111111111001011100011011;
assign LUT_4[20564] = 32'b11111111111111111101110110011011;
assign LUT_4[20565] = 32'b11111111111111110111000010010011;
assign LUT_4[20566] = 32'b11111111111111111101010000111111;
assign LUT_4[20567] = 32'b11111111111111110110011100110111;
assign LUT_4[20568] = 32'b11111111111111111010000010010100;
assign LUT_4[20569] = 32'b11111111111111110011001110001100;
assign LUT_4[20570] = 32'b11111111111111111001011100111000;
assign LUT_4[20571] = 32'b11111111111111110010101000110000;
assign LUT_4[20572] = 32'b11111111111111110111000010110000;
assign LUT_4[20573] = 32'b11111111111111110000001110101000;
assign LUT_4[20574] = 32'b11111111111111110110011101010100;
assign LUT_4[20575] = 32'b11111111111111101111101001001100;
assign LUT_4[20576] = 32'b00000000000000000001011111011000;
assign LUT_4[20577] = 32'b11111111111111111010101011010000;
assign LUT_4[20578] = 32'b00000000000000000000111001111100;
assign LUT_4[20579] = 32'b11111111111111111010000101110100;
assign LUT_4[20580] = 32'b11111111111111111110011111110100;
assign LUT_4[20581] = 32'b11111111111111110111101011101100;
assign LUT_4[20582] = 32'b11111111111111111101111010011000;
assign LUT_4[20583] = 32'b11111111111111110111000110010000;
assign LUT_4[20584] = 32'b11111111111111111010101011101101;
assign LUT_4[20585] = 32'b11111111111111110011110111100101;
assign LUT_4[20586] = 32'b11111111111111111010000110010001;
assign LUT_4[20587] = 32'b11111111111111110011010010001001;
assign LUT_4[20588] = 32'b11111111111111110111101100001001;
assign LUT_4[20589] = 32'b11111111111111110000111000000001;
assign LUT_4[20590] = 32'b11111111111111110111000110101101;
assign LUT_4[20591] = 32'b11111111111111110000010010100101;
assign LUT_4[20592] = 32'b11111111111111111111010001000110;
assign LUT_4[20593] = 32'b11111111111111111000011100111110;
assign LUT_4[20594] = 32'b11111111111111111110101011101010;
assign LUT_4[20595] = 32'b11111111111111110111110111100010;
assign LUT_4[20596] = 32'b11111111111111111100010001100010;
assign LUT_4[20597] = 32'b11111111111111110101011101011010;
assign LUT_4[20598] = 32'b11111111111111111011101100000110;
assign LUT_4[20599] = 32'b11111111111111110100110111111110;
assign LUT_4[20600] = 32'b11111111111111111000011101011011;
assign LUT_4[20601] = 32'b11111111111111110001101001010011;
assign LUT_4[20602] = 32'b11111111111111110111110111111111;
assign LUT_4[20603] = 32'b11111111111111110001000011110111;
assign LUT_4[20604] = 32'b11111111111111110101011101110111;
assign LUT_4[20605] = 32'b11111111111111101110101001101111;
assign LUT_4[20606] = 32'b11111111111111110100111000011011;
assign LUT_4[20607] = 32'b11111111111111101110000100010011;
assign LUT_4[20608] = 32'b00000000000000000100010011000101;
assign LUT_4[20609] = 32'b11111111111111111101011110111101;
assign LUT_4[20610] = 32'b00000000000000000011101101101001;
assign LUT_4[20611] = 32'b11111111111111111100111001100001;
assign LUT_4[20612] = 32'b00000000000000000001010011100001;
assign LUT_4[20613] = 32'b11111111111111111010011111011001;
assign LUT_4[20614] = 32'b00000000000000000000101110000101;
assign LUT_4[20615] = 32'b11111111111111111001111001111101;
assign LUT_4[20616] = 32'b11111111111111111101011111011010;
assign LUT_4[20617] = 32'b11111111111111110110101011010010;
assign LUT_4[20618] = 32'b11111111111111111100111001111110;
assign LUT_4[20619] = 32'b11111111111111110110000101110110;
assign LUT_4[20620] = 32'b11111111111111111010011111110110;
assign LUT_4[20621] = 32'b11111111111111110011101011101110;
assign LUT_4[20622] = 32'b11111111111111111001111010011010;
assign LUT_4[20623] = 32'b11111111111111110011000110010010;
assign LUT_4[20624] = 32'b00000000000000000010000100110011;
assign LUT_4[20625] = 32'b11111111111111111011010000101011;
assign LUT_4[20626] = 32'b00000000000000000001011111010111;
assign LUT_4[20627] = 32'b11111111111111111010101011001111;
assign LUT_4[20628] = 32'b11111111111111111111000101001111;
assign LUT_4[20629] = 32'b11111111111111111000010001000111;
assign LUT_4[20630] = 32'b11111111111111111110011111110011;
assign LUT_4[20631] = 32'b11111111111111110111101011101011;
assign LUT_4[20632] = 32'b11111111111111111011010001001000;
assign LUT_4[20633] = 32'b11111111111111110100011101000000;
assign LUT_4[20634] = 32'b11111111111111111010101011101100;
assign LUT_4[20635] = 32'b11111111111111110011110111100100;
assign LUT_4[20636] = 32'b11111111111111111000010001100100;
assign LUT_4[20637] = 32'b11111111111111110001011101011100;
assign LUT_4[20638] = 32'b11111111111111110111101100001000;
assign LUT_4[20639] = 32'b11111111111111110000111000000000;
assign LUT_4[20640] = 32'b00000000000000000010101110001100;
assign LUT_4[20641] = 32'b11111111111111111011111010000100;
assign LUT_4[20642] = 32'b00000000000000000010001000110000;
assign LUT_4[20643] = 32'b11111111111111111011010100101000;
assign LUT_4[20644] = 32'b11111111111111111111101110101000;
assign LUT_4[20645] = 32'b11111111111111111000111010100000;
assign LUT_4[20646] = 32'b11111111111111111111001001001100;
assign LUT_4[20647] = 32'b11111111111111111000010101000100;
assign LUT_4[20648] = 32'b11111111111111111011111010100001;
assign LUT_4[20649] = 32'b11111111111111110101000110011001;
assign LUT_4[20650] = 32'b11111111111111111011010101000101;
assign LUT_4[20651] = 32'b11111111111111110100100000111101;
assign LUT_4[20652] = 32'b11111111111111111000111010111101;
assign LUT_4[20653] = 32'b11111111111111110010000110110101;
assign LUT_4[20654] = 32'b11111111111111111000010101100001;
assign LUT_4[20655] = 32'b11111111111111110001100001011001;
assign LUT_4[20656] = 32'b00000000000000000000011111111010;
assign LUT_4[20657] = 32'b11111111111111111001101011110010;
assign LUT_4[20658] = 32'b11111111111111111111111010011110;
assign LUT_4[20659] = 32'b11111111111111111001000110010110;
assign LUT_4[20660] = 32'b11111111111111111101100000010110;
assign LUT_4[20661] = 32'b11111111111111110110101100001110;
assign LUT_4[20662] = 32'b11111111111111111100111010111010;
assign LUT_4[20663] = 32'b11111111111111110110000110110010;
assign LUT_4[20664] = 32'b11111111111111111001101100001111;
assign LUT_4[20665] = 32'b11111111111111110010111000000111;
assign LUT_4[20666] = 32'b11111111111111111001000110110011;
assign LUT_4[20667] = 32'b11111111111111110010010010101011;
assign LUT_4[20668] = 32'b11111111111111110110101100101011;
assign LUT_4[20669] = 32'b11111111111111101111111000100011;
assign LUT_4[20670] = 32'b11111111111111110110000111001111;
assign LUT_4[20671] = 32'b11111111111111101111010011000111;
assign LUT_4[20672] = 32'b00000000000000000101101010011001;
assign LUT_4[20673] = 32'b11111111111111111110110110010001;
assign LUT_4[20674] = 32'b00000000000000000101000100111101;
assign LUT_4[20675] = 32'b11111111111111111110010000110101;
assign LUT_4[20676] = 32'b00000000000000000010101010110101;
assign LUT_4[20677] = 32'b11111111111111111011110110101101;
assign LUT_4[20678] = 32'b00000000000000000010000101011001;
assign LUT_4[20679] = 32'b11111111111111111011010001010001;
assign LUT_4[20680] = 32'b11111111111111111110110110101110;
assign LUT_4[20681] = 32'b11111111111111111000000010100110;
assign LUT_4[20682] = 32'b11111111111111111110010001010010;
assign LUT_4[20683] = 32'b11111111111111110111011101001010;
assign LUT_4[20684] = 32'b11111111111111111011110111001010;
assign LUT_4[20685] = 32'b11111111111111110101000011000010;
assign LUT_4[20686] = 32'b11111111111111111011010001101110;
assign LUT_4[20687] = 32'b11111111111111110100011101100110;
assign LUT_4[20688] = 32'b00000000000000000011011100000111;
assign LUT_4[20689] = 32'b11111111111111111100100111111111;
assign LUT_4[20690] = 32'b00000000000000000010110110101011;
assign LUT_4[20691] = 32'b11111111111111111100000010100011;
assign LUT_4[20692] = 32'b00000000000000000000011100100011;
assign LUT_4[20693] = 32'b11111111111111111001101000011011;
assign LUT_4[20694] = 32'b11111111111111111111110111000111;
assign LUT_4[20695] = 32'b11111111111111111001000010111111;
assign LUT_4[20696] = 32'b11111111111111111100101000011100;
assign LUT_4[20697] = 32'b11111111111111110101110100010100;
assign LUT_4[20698] = 32'b11111111111111111100000011000000;
assign LUT_4[20699] = 32'b11111111111111110101001110111000;
assign LUT_4[20700] = 32'b11111111111111111001101000111000;
assign LUT_4[20701] = 32'b11111111111111110010110100110000;
assign LUT_4[20702] = 32'b11111111111111111001000011011100;
assign LUT_4[20703] = 32'b11111111111111110010001111010100;
assign LUT_4[20704] = 32'b00000000000000000100000101100000;
assign LUT_4[20705] = 32'b11111111111111111101010001011000;
assign LUT_4[20706] = 32'b00000000000000000011100000000100;
assign LUT_4[20707] = 32'b11111111111111111100101011111100;
assign LUT_4[20708] = 32'b00000000000000000001000101111100;
assign LUT_4[20709] = 32'b11111111111111111010010001110100;
assign LUT_4[20710] = 32'b00000000000000000000100000100000;
assign LUT_4[20711] = 32'b11111111111111111001101100011000;
assign LUT_4[20712] = 32'b11111111111111111101010001110101;
assign LUT_4[20713] = 32'b11111111111111110110011101101101;
assign LUT_4[20714] = 32'b11111111111111111100101100011001;
assign LUT_4[20715] = 32'b11111111111111110101111000010001;
assign LUT_4[20716] = 32'b11111111111111111010010010010001;
assign LUT_4[20717] = 32'b11111111111111110011011110001001;
assign LUT_4[20718] = 32'b11111111111111111001101100110101;
assign LUT_4[20719] = 32'b11111111111111110010111000101101;
assign LUT_4[20720] = 32'b00000000000000000001110111001110;
assign LUT_4[20721] = 32'b11111111111111111011000011000110;
assign LUT_4[20722] = 32'b00000000000000000001010001110010;
assign LUT_4[20723] = 32'b11111111111111111010011101101010;
assign LUT_4[20724] = 32'b11111111111111111110110111101010;
assign LUT_4[20725] = 32'b11111111111111111000000011100010;
assign LUT_4[20726] = 32'b11111111111111111110010010001110;
assign LUT_4[20727] = 32'b11111111111111110111011110000110;
assign LUT_4[20728] = 32'b11111111111111111011000011100011;
assign LUT_4[20729] = 32'b11111111111111110100001111011011;
assign LUT_4[20730] = 32'b11111111111111111010011110000111;
assign LUT_4[20731] = 32'b11111111111111110011101001111111;
assign LUT_4[20732] = 32'b11111111111111111000000011111111;
assign LUT_4[20733] = 32'b11111111111111110001001111110111;
assign LUT_4[20734] = 32'b11111111111111110111011110100011;
assign LUT_4[20735] = 32'b11111111111111110000101010011011;
assign LUT_4[20736] = 32'b00000000000000000110101000100000;
assign LUT_4[20737] = 32'b11111111111111111111110100011000;
assign LUT_4[20738] = 32'b00000000000000000110000011000100;
assign LUT_4[20739] = 32'b11111111111111111111001110111100;
assign LUT_4[20740] = 32'b00000000000000000011101000111100;
assign LUT_4[20741] = 32'b11111111111111111100110100110100;
assign LUT_4[20742] = 32'b00000000000000000011000011100000;
assign LUT_4[20743] = 32'b11111111111111111100001111011000;
assign LUT_4[20744] = 32'b11111111111111111111110100110101;
assign LUT_4[20745] = 32'b11111111111111111001000000101101;
assign LUT_4[20746] = 32'b11111111111111111111001111011001;
assign LUT_4[20747] = 32'b11111111111111111000011011010001;
assign LUT_4[20748] = 32'b11111111111111111100110101010001;
assign LUT_4[20749] = 32'b11111111111111110110000001001001;
assign LUT_4[20750] = 32'b11111111111111111100001111110101;
assign LUT_4[20751] = 32'b11111111111111110101011011101101;
assign LUT_4[20752] = 32'b00000000000000000100011010001110;
assign LUT_4[20753] = 32'b11111111111111111101100110000110;
assign LUT_4[20754] = 32'b00000000000000000011110100110010;
assign LUT_4[20755] = 32'b11111111111111111101000000101010;
assign LUT_4[20756] = 32'b00000000000000000001011010101010;
assign LUT_4[20757] = 32'b11111111111111111010100110100010;
assign LUT_4[20758] = 32'b00000000000000000000110101001110;
assign LUT_4[20759] = 32'b11111111111111111010000001000110;
assign LUT_4[20760] = 32'b11111111111111111101100110100011;
assign LUT_4[20761] = 32'b11111111111111110110110010011011;
assign LUT_4[20762] = 32'b11111111111111111101000001000111;
assign LUT_4[20763] = 32'b11111111111111110110001100111111;
assign LUT_4[20764] = 32'b11111111111111111010100110111111;
assign LUT_4[20765] = 32'b11111111111111110011110010110111;
assign LUT_4[20766] = 32'b11111111111111111010000001100011;
assign LUT_4[20767] = 32'b11111111111111110011001101011011;
assign LUT_4[20768] = 32'b00000000000000000101000011100111;
assign LUT_4[20769] = 32'b11111111111111111110001111011111;
assign LUT_4[20770] = 32'b00000000000000000100011110001011;
assign LUT_4[20771] = 32'b11111111111111111101101010000011;
assign LUT_4[20772] = 32'b00000000000000000010000100000011;
assign LUT_4[20773] = 32'b11111111111111111011001111111011;
assign LUT_4[20774] = 32'b00000000000000000001011110100111;
assign LUT_4[20775] = 32'b11111111111111111010101010011111;
assign LUT_4[20776] = 32'b11111111111111111110001111111100;
assign LUT_4[20777] = 32'b11111111111111110111011011110100;
assign LUT_4[20778] = 32'b11111111111111111101101010100000;
assign LUT_4[20779] = 32'b11111111111111110110110110011000;
assign LUT_4[20780] = 32'b11111111111111111011010000011000;
assign LUT_4[20781] = 32'b11111111111111110100011100010000;
assign LUT_4[20782] = 32'b11111111111111111010101010111100;
assign LUT_4[20783] = 32'b11111111111111110011110110110100;
assign LUT_4[20784] = 32'b00000000000000000010110101010101;
assign LUT_4[20785] = 32'b11111111111111111100000001001101;
assign LUT_4[20786] = 32'b00000000000000000010001111111001;
assign LUT_4[20787] = 32'b11111111111111111011011011110001;
assign LUT_4[20788] = 32'b11111111111111111111110101110001;
assign LUT_4[20789] = 32'b11111111111111111001000001101001;
assign LUT_4[20790] = 32'b11111111111111111111010000010101;
assign LUT_4[20791] = 32'b11111111111111111000011100001101;
assign LUT_4[20792] = 32'b11111111111111111100000001101010;
assign LUT_4[20793] = 32'b11111111111111110101001101100010;
assign LUT_4[20794] = 32'b11111111111111111011011100001110;
assign LUT_4[20795] = 32'b11111111111111110100101000000110;
assign LUT_4[20796] = 32'b11111111111111111001000010000110;
assign LUT_4[20797] = 32'b11111111111111110010001101111110;
assign LUT_4[20798] = 32'b11111111111111111000011100101010;
assign LUT_4[20799] = 32'b11111111111111110001101000100010;
assign LUT_4[20800] = 32'b00000000000000000111111111110100;
assign LUT_4[20801] = 32'b00000000000000000001001011101100;
assign LUT_4[20802] = 32'b00000000000000000111011010011000;
assign LUT_4[20803] = 32'b00000000000000000000100110010000;
assign LUT_4[20804] = 32'b00000000000000000101000000010000;
assign LUT_4[20805] = 32'b11111111111111111110001100001000;
assign LUT_4[20806] = 32'b00000000000000000100011010110100;
assign LUT_4[20807] = 32'b11111111111111111101100110101100;
assign LUT_4[20808] = 32'b00000000000000000001001100001001;
assign LUT_4[20809] = 32'b11111111111111111010011000000001;
assign LUT_4[20810] = 32'b00000000000000000000100110101101;
assign LUT_4[20811] = 32'b11111111111111111001110010100101;
assign LUT_4[20812] = 32'b11111111111111111110001100100101;
assign LUT_4[20813] = 32'b11111111111111110111011000011101;
assign LUT_4[20814] = 32'b11111111111111111101100111001001;
assign LUT_4[20815] = 32'b11111111111111110110110011000001;
assign LUT_4[20816] = 32'b00000000000000000101110001100010;
assign LUT_4[20817] = 32'b11111111111111111110111101011010;
assign LUT_4[20818] = 32'b00000000000000000101001100000110;
assign LUT_4[20819] = 32'b11111111111111111110010111111110;
assign LUT_4[20820] = 32'b00000000000000000010110001111110;
assign LUT_4[20821] = 32'b11111111111111111011111101110110;
assign LUT_4[20822] = 32'b00000000000000000010001100100010;
assign LUT_4[20823] = 32'b11111111111111111011011000011010;
assign LUT_4[20824] = 32'b11111111111111111110111101110111;
assign LUT_4[20825] = 32'b11111111111111111000001001101111;
assign LUT_4[20826] = 32'b11111111111111111110011000011011;
assign LUT_4[20827] = 32'b11111111111111110111100100010011;
assign LUT_4[20828] = 32'b11111111111111111011111110010011;
assign LUT_4[20829] = 32'b11111111111111110101001010001011;
assign LUT_4[20830] = 32'b11111111111111111011011000110111;
assign LUT_4[20831] = 32'b11111111111111110100100100101111;
assign LUT_4[20832] = 32'b00000000000000000110011010111011;
assign LUT_4[20833] = 32'b11111111111111111111100110110011;
assign LUT_4[20834] = 32'b00000000000000000101110101011111;
assign LUT_4[20835] = 32'b11111111111111111111000001010111;
assign LUT_4[20836] = 32'b00000000000000000011011011010111;
assign LUT_4[20837] = 32'b11111111111111111100100111001111;
assign LUT_4[20838] = 32'b00000000000000000010110101111011;
assign LUT_4[20839] = 32'b11111111111111111100000001110011;
assign LUT_4[20840] = 32'b11111111111111111111100111010000;
assign LUT_4[20841] = 32'b11111111111111111000110011001000;
assign LUT_4[20842] = 32'b11111111111111111111000001110100;
assign LUT_4[20843] = 32'b11111111111111111000001101101100;
assign LUT_4[20844] = 32'b11111111111111111100100111101100;
assign LUT_4[20845] = 32'b11111111111111110101110011100100;
assign LUT_4[20846] = 32'b11111111111111111100000010010000;
assign LUT_4[20847] = 32'b11111111111111110101001110001000;
assign LUT_4[20848] = 32'b00000000000000000100001100101001;
assign LUT_4[20849] = 32'b11111111111111111101011000100001;
assign LUT_4[20850] = 32'b00000000000000000011100111001101;
assign LUT_4[20851] = 32'b11111111111111111100110011000101;
assign LUT_4[20852] = 32'b00000000000000000001001101000101;
assign LUT_4[20853] = 32'b11111111111111111010011000111101;
assign LUT_4[20854] = 32'b00000000000000000000100111101001;
assign LUT_4[20855] = 32'b11111111111111111001110011100001;
assign LUT_4[20856] = 32'b11111111111111111101011000111110;
assign LUT_4[20857] = 32'b11111111111111110110100100110110;
assign LUT_4[20858] = 32'b11111111111111111100110011100010;
assign LUT_4[20859] = 32'b11111111111111110101111111011010;
assign LUT_4[20860] = 32'b11111111111111111010011001011010;
assign LUT_4[20861] = 32'b11111111111111110011100101010010;
assign LUT_4[20862] = 32'b11111111111111111001110011111110;
assign LUT_4[20863] = 32'b11111111111111110010111111110110;
assign LUT_4[20864] = 32'b00000000000000001001001110101000;
assign LUT_4[20865] = 32'b00000000000000000010011010100000;
assign LUT_4[20866] = 32'b00000000000000001000101001001100;
assign LUT_4[20867] = 32'b00000000000000000001110101000100;
assign LUT_4[20868] = 32'b00000000000000000110001111000100;
assign LUT_4[20869] = 32'b11111111111111111111011010111100;
assign LUT_4[20870] = 32'b00000000000000000101101001101000;
assign LUT_4[20871] = 32'b11111111111111111110110101100000;
assign LUT_4[20872] = 32'b00000000000000000010011010111101;
assign LUT_4[20873] = 32'b11111111111111111011100110110101;
assign LUT_4[20874] = 32'b00000000000000000001110101100001;
assign LUT_4[20875] = 32'b11111111111111111011000001011001;
assign LUT_4[20876] = 32'b11111111111111111111011011011001;
assign LUT_4[20877] = 32'b11111111111111111000100111010001;
assign LUT_4[20878] = 32'b11111111111111111110110101111101;
assign LUT_4[20879] = 32'b11111111111111111000000001110101;
assign LUT_4[20880] = 32'b00000000000000000111000000010110;
assign LUT_4[20881] = 32'b00000000000000000000001100001110;
assign LUT_4[20882] = 32'b00000000000000000110011010111010;
assign LUT_4[20883] = 32'b11111111111111111111100110110010;
assign LUT_4[20884] = 32'b00000000000000000100000000110010;
assign LUT_4[20885] = 32'b11111111111111111101001100101010;
assign LUT_4[20886] = 32'b00000000000000000011011011010110;
assign LUT_4[20887] = 32'b11111111111111111100100111001110;
assign LUT_4[20888] = 32'b00000000000000000000001100101011;
assign LUT_4[20889] = 32'b11111111111111111001011000100011;
assign LUT_4[20890] = 32'b11111111111111111111100111001111;
assign LUT_4[20891] = 32'b11111111111111111000110011000111;
assign LUT_4[20892] = 32'b11111111111111111101001101000111;
assign LUT_4[20893] = 32'b11111111111111110110011000111111;
assign LUT_4[20894] = 32'b11111111111111111100100111101011;
assign LUT_4[20895] = 32'b11111111111111110101110011100011;
assign LUT_4[20896] = 32'b00000000000000000111101001101111;
assign LUT_4[20897] = 32'b00000000000000000000110101100111;
assign LUT_4[20898] = 32'b00000000000000000111000100010011;
assign LUT_4[20899] = 32'b00000000000000000000010000001011;
assign LUT_4[20900] = 32'b00000000000000000100101010001011;
assign LUT_4[20901] = 32'b11111111111111111101110110000011;
assign LUT_4[20902] = 32'b00000000000000000100000100101111;
assign LUT_4[20903] = 32'b11111111111111111101010000100111;
assign LUT_4[20904] = 32'b00000000000000000000110110000100;
assign LUT_4[20905] = 32'b11111111111111111010000001111100;
assign LUT_4[20906] = 32'b00000000000000000000010000101000;
assign LUT_4[20907] = 32'b11111111111111111001011100100000;
assign LUT_4[20908] = 32'b11111111111111111101110110100000;
assign LUT_4[20909] = 32'b11111111111111110111000010011000;
assign LUT_4[20910] = 32'b11111111111111111101010001000100;
assign LUT_4[20911] = 32'b11111111111111110110011100111100;
assign LUT_4[20912] = 32'b00000000000000000101011011011101;
assign LUT_4[20913] = 32'b11111111111111111110100111010101;
assign LUT_4[20914] = 32'b00000000000000000100110110000001;
assign LUT_4[20915] = 32'b11111111111111111110000001111001;
assign LUT_4[20916] = 32'b00000000000000000010011011111001;
assign LUT_4[20917] = 32'b11111111111111111011100111110001;
assign LUT_4[20918] = 32'b00000000000000000001110110011101;
assign LUT_4[20919] = 32'b11111111111111111011000010010101;
assign LUT_4[20920] = 32'b11111111111111111110100111110010;
assign LUT_4[20921] = 32'b11111111111111110111110011101010;
assign LUT_4[20922] = 32'b11111111111111111110000010010110;
assign LUT_4[20923] = 32'b11111111111111110111001110001110;
assign LUT_4[20924] = 32'b11111111111111111011101000001110;
assign LUT_4[20925] = 32'b11111111111111110100110100000110;
assign LUT_4[20926] = 32'b11111111111111111011000010110010;
assign LUT_4[20927] = 32'b11111111111111110100001110101010;
assign LUT_4[20928] = 32'b00000000000000001010100101111100;
assign LUT_4[20929] = 32'b00000000000000000011110001110100;
assign LUT_4[20930] = 32'b00000000000000001010000000100000;
assign LUT_4[20931] = 32'b00000000000000000011001100011000;
assign LUT_4[20932] = 32'b00000000000000000111100110011000;
assign LUT_4[20933] = 32'b00000000000000000000110010010000;
assign LUT_4[20934] = 32'b00000000000000000111000000111100;
assign LUT_4[20935] = 32'b00000000000000000000001100110100;
assign LUT_4[20936] = 32'b00000000000000000011110010010001;
assign LUT_4[20937] = 32'b11111111111111111100111110001001;
assign LUT_4[20938] = 32'b00000000000000000011001100110101;
assign LUT_4[20939] = 32'b11111111111111111100011000101101;
assign LUT_4[20940] = 32'b00000000000000000000110010101101;
assign LUT_4[20941] = 32'b11111111111111111001111110100101;
assign LUT_4[20942] = 32'b00000000000000000000001101010001;
assign LUT_4[20943] = 32'b11111111111111111001011001001001;
assign LUT_4[20944] = 32'b00000000000000001000010111101010;
assign LUT_4[20945] = 32'b00000000000000000001100011100010;
assign LUT_4[20946] = 32'b00000000000000000111110010001110;
assign LUT_4[20947] = 32'b00000000000000000000111110000110;
assign LUT_4[20948] = 32'b00000000000000000101011000000110;
assign LUT_4[20949] = 32'b11111111111111111110100011111110;
assign LUT_4[20950] = 32'b00000000000000000100110010101010;
assign LUT_4[20951] = 32'b11111111111111111101111110100010;
assign LUT_4[20952] = 32'b00000000000000000001100011111111;
assign LUT_4[20953] = 32'b11111111111111111010101111110111;
assign LUT_4[20954] = 32'b00000000000000000000111110100011;
assign LUT_4[20955] = 32'b11111111111111111010001010011011;
assign LUT_4[20956] = 32'b11111111111111111110100100011011;
assign LUT_4[20957] = 32'b11111111111111110111110000010011;
assign LUT_4[20958] = 32'b11111111111111111101111110111111;
assign LUT_4[20959] = 32'b11111111111111110111001010110111;
assign LUT_4[20960] = 32'b00000000000000001001000001000011;
assign LUT_4[20961] = 32'b00000000000000000010001100111011;
assign LUT_4[20962] = 32'b00000000000000001000011011100111;
assign LUT_4[20963] = 32'b00000000000000000001100111011111;
assign LUT_4[20964] = 32'b00000000000000000110000001011111;
assign LUT_4[20965] = 32'b11111111111111111111001101010111;
assign LUT_4[20966] = 32'b00000000000000000101011100000011;
assign LUT_4[20967] = 32'b11111111111111111110100111111011;
assign LUT_4[20968] = 32'b00000000000000000010001101011000;
assign LUT_4[20969] = 32'b11111111111111111011011001010000;
assign LUT_4[20970] = 32'b00000000000000000001100111111100;
assign LUT_4[20971] = 32'b11111111111111111010110011110100;
assign LUT_4[20972] = 32'b11111111111111111111001101110100;
assign LUT_4[20973] = 32'b11111111111111111000011001101100;
assign LUT_4[20974] = 32'b11111111111111111110101000011000;
assign LUT_4[20975] = 32'b11111111111111110111110100010000;
assign LUT_4[20976] = 32'b00000000000000000110110010110001;
assign LUT_4[20977] = 32'b11111111111111111111111110101001;
assign LUT_4[20978] = 32'b00000000000000000110001101010101;
assign LUT_4[20979] = 32'b11111111111111111111011001001101;
assign LUT_4[20980] = 32'b00000000000000000011110011001101;
assign LUT_4[20981] = 32'b11111111111111111100111111000101;
assign LUT_4[20982] = 32'b00000000000000000011001101110001;
assign LUT_4[20983] = 32'b11111111111111111100011001101001;
assign LUT_4[20984] = 32'b11111111111111111111111111000110;
assign LUT_4[20985] = 32'b11111111111111111001001010111110;
assign LUT_4[20986] = 32'b11111111111111111111011001101010;
assign LUT_4[20987] = 32'b11111111111111111000100101100010;
assign LUT_4[20988] = 32'b11111111111111111100111111100010;
assign LUT_4[20989] = 32'b11111111111111110110001011011010;
assign LUT_4[20990] = 32'b11111111111111111100011010000110;
assign LUT_4[20991] = 32'b11111111111111110101100101111110;
assign LUT_4[20992] = 32'b00000000000000000000110001000101;
assign LUT_4[20993] = 32'b11111111111111111001111100111101;
assign LUT_4[20994] = 32'b00000000000000000000001011101001;
assign LUT_4[20995] = 32'b11111111111111111001010111100001;
assign LUT_4[20996] = 32'b11111111111111111101110001100001;
assign LUT_4[20997] = 32'b11111111111111110110111101011001;
assign LUT_4[20998] = 32'b11111111111111111101001100000101;
assign LUT_4[20999] = 32'b11111111111111110110010111111101;
assign LUT_4[21000] = 32'b11111111111111111001111101011010;
assign LUT_4[21001] = 32'b11111111111111110011001001010010;
assign LUT_4[21002] = 32'b11111111111111111001010111111110;
assign LUT_4[21003] = 32'b11111111111111110010100011110110;
assign LUT_4[21004] = 32'b11111111111111110110111101110110;
assign LUT_4[21005] = 32'b11111111111111110000001001101110;
assign LUT_4[21006] = 32'b11111111111111110110011000011010;
assign LUT_4[21007] = 32'b11111111111111101111100100010010;
assign LUT_4[21008] = 32'b11111111111111111110100010110011;
assign LUT_4[21009] = 32'b11111111111111110111101110101011;
assign LUT_4[21010] = 32'b11111111111111111101111101010111;
assign LUT_4[21011] = 32'b11111111111111110111001001001111;
assign LUT_4[21012] = 32'b11111111111111111011100011001111;
assign LUT_4[21013] = 32'b11111111111111110100101111000111;
assign LUT_4[21014] = 32'b11111111111111111010111101110011;
assign LUT_4[21015] = 32'b11111111111111110100001001101011;
assign LUT_4[21016] = 32'b11111111111111110111101111001000;
assign LUT_4[21017] = 32'b11111111111111110000111011000000;
assign LUT_4[21018] = 32'b11111111111111110111001001101100;
assign LUT_4[21019] = 32'b11111111111111110000010101100100;
assign LUT_4[21020] = 32'b11111111111111110100101111100100;
assign LUT_4[21021] = 32'b11111111111111101101111011011100;
assign LUT_4[21022] = 32'b11111111111111110100001010001000;
assign LUT_4[21023] = 32'b11111111111111101101010110000000;
assign LUT_4[21024] = 32'b11111111111111111111001100001100;
assign LUT_4[21025] = 32'b11111111111111111000011000000100;
assign LUT_4[21026] = 32'b11111111111111111110100110110000;
assign LUT_4[21027] = 32'b11111111111111110111110010101000;
assign LUT_4[21028] = 32'b11111111111111111100001100101000;
assign LUT_4[21029] = 32'b11111111111111110101011000100000;
assign LUT_4[21030] = 32'b11111111111111111011100111001100;
assign LUT_4[21031] = 32'b11111111111111110100110011000100;
assign LUT_4[21032] = 32'b11111111111111111000011000100001;
assign LUT_4[21033] = 32'b11111111111111110001100100011001;
assign LUT_4[21034] = 32'b11111111111111110111110011000101;
assign LUT_4[21035] = 32'b11111111111111110000111110111101;
assign LUT_4[21036] = 32'b11111111111111110101011000111101;
assign LUT_4[21037] = 32'b11111111111111101110100100110101;
assign LUT_4[21038] = 32'b11111111111111110100110011100001;
assign LUT_4[21039] = 32'b11111111111111101101111111011001;
assign LUT_4[21040] = 32'b11111111111111111100111101111010;
assign LUT_4[21041] = 32'b11111111111111110110001001110010;
assign LUT_4[21042] = 32'b11111111111111111100011000011110;
assign LUT_4[21043] = 32'b11111111111111110101100100010110;
assign LUT_4[21044] = 32'b11111111111111111001111110010110;
assign LUT_4[21045] = 32'b11111111111111110011001010001110;
assign LUT_4[21046] = 32'b11111111111111111001011000111010;
assign LUT_4[21047] = 32'b11111111111111110010100100110010;
assign LUT_4[21048] = 32'b11111111111111110110001010001111;
assign LUT_4[21049] = 32'b11111111111111101111010110000111;
assign LUT_4[21050] = 32'b11111111111111110101100100110011;
assign LUT_4[21051] = 32'b11111111111111101110110000101011;
assign LUT_4[21052] = 32'b11111111111111110011001010101011;
assign LUT_4[21053] = 32'b11111111111111101100010110100011;
assign LUT_4[21054] = 32'b11111111111111110010100101001111;
assign LUT_4[21055] = 32'b11111111111111101011110001000111;
assign LUT_4[21056] = 32'b00000000000000000010001000011001;
assign LUT_4[21057] = 32'b11111111111111111011010100010001;
assign LUT_4[21058] = 32'b00000000000000000001100010111101;
assign LUT_4[21059] = 32'b11111111111111111010101110110101;
assign LUT_4[21060] = 32'b11111111111111111111001000110101;
assign LUT_4[21061] = 32'b11111111111111111000010100101101;
assign LUT_4[21062] = 32'b11111111111111111110100011011001;
assign LUT_4[21063] = 32'b11111111111111110111101111010001;
assign LUT_4[21064] = 32'b11111111111111111011010100101110;
assign LUT_4[21065] = 32'b11111111111111110100100000100110;
assign LUT_4[21066] = 32'b11111111111111111010101111010010;
assign LUT_4[21067] = 32'b11111111111111110011111011001010;
assign LUT_4[21068] = 32'b11111111111111111000010101001010;
assign LUT_4[21069] = 32'b11111111111111110001100001000010;
assign LUT_4[21070] = 32'b11111111111111110111101111101110;
assign LUT_4[21071] = 32'b11111111111111110000111011100110;
assign LUT_4[21072] = 32'b11111111111111111111111010000111;
assign LUT_4[21073] = 32'b11111111111111111001000101111111;
assign LUT_4[21074] = 32'b11111111111111111111010100101011;
assign LUT_4[21075] = 32'b11111111111111111000100000100011;
assign LUT_4[21076] = 32'b11111111111111111100111010100011;
assign LUT_4[21077] = 32'b11111111111111110110000110011011;
assign LUT_4[21078] = 32'b11111111111111111100010101000111;
assign LUT_4[21079] = 32'b11111111111111110101100000111111;
assign LUT_4[21080] = 32'b11111111111111111001000110011100;
assign LUT_4[21081] = 32'b11111111111111110010010010010100;
assign LUT_4[21082] = 32'b11111111111111111000100001000000;
assign LUT_4[21083] = 32'b11111111111111110001101100111000;
assign LUT_4[21084] = 32'b11111111111111110110000110111000;
assign LUT_4[21085] = 32'b11111111111111101111010010110000;
assign LUT_4[21086] = 32'b11111111111111110101100001011100;
assign LUT_4[21087] = 32'b11111111111111101110101101010100;
assign LUT_4[21088] = 32'b00000000000000000000100011100000;
assign LUT_4[21089] = 32'b11111111111111111001101111011000;
assign LUT_4[21090] = 32'b11111111111111111111111110000100;
assign LUT_4[21091] = 32'b11111111111111111001001001111100;
assign LUT_4[21092] = 32'b11111111111111111101100011111100;
assign LUT_4[21093] = 32'b11111111111111110110101111110100;
assign LUT_4[21094] = 32'b11111111111111111100111110100000;
assign LUT_4[21095] = 32'b11111111111111110110001010011000;
assign LUT_4[21096] = 32'b11111111111111111001101111110101;
assign LUT_4[21097] = 32'b11111111111111110010111011101101;
assign LUT_4[21098] = 32'b11111111111111111001001010011001;
assign LUT_4[21099] = 32'b11111111111111110010010110010001;
assign LUT_4[21100] = 32'b11111111111111110110110000010001;
assign LUT_4[21101] = 32'b11111111111111101111111100001001;
assign LUT_4[21102] = 32'b11111111111111110110001010110101;
assign LUT_4[21103] = 32'b11111111111111101111010110101101;
assign LUT_4[21104] = 32'b11111111111111111110010101001110;
assign LUT_4[21105] = 32'b11111111111111110111100001000110;
assign LUT_4[21106] = 32'b11111111111111111101101111110010;
assign LUT_4[21107] = 32'b11111111111111110110111011101010;
assign LUT_4[21108] = 32'b11111111111111111011010101101010;
assign LUT_4[21109] = 32'b11111111111111110100100001100010;
assign LUT_4[21110] = 32'b11111111111111111010110000001110;
assign LUT_4[21111] = 32'b11111111111111110011111100000110;
assign LUT_4[21112] = 32'b11111111111111110111100001100011;
assign LUT_4[21113] = 32'b11111111111111110000101101011011;
assign LUT_4[21114] = 32'b11111111111111110110111100000111;
assign LUT_4[21115] = 32'b11111111111111110000000111111111;
assign LUT_4[21116] = 32'b11111111111111110100100001111111;
assign LUT_4[21117] = 32'b11111111111111101101101101110111;
assign LUT_4[21118] = 32'b11111111111111110011111100100011;
assign LUT_4[21119] = 32'b11111111111111101101001000011011;
assign LUT_4[21120] = 32'b00000000000000000011010111001101;
assign LUT_4[21121] = 32'b11111111111111111100100011000101;
assign LUT_4[21122] = 32'b00000000000000000010110001110001;
assign LUT_4[21123] = 32'b11111111111111111011111101101001;
assign LUT_4[21124] = 32'b00000000000000000000010111101001;
assign LUT_4[21125] = 32'b11111111111111111001100011100001;
assign LUT_4[21126] = 32'b11111111111111111111110010001101;
assign LUT_4[21127] = 32'b11111111111111111000111110000101;
assign LUT_4[21128] = 32'b11111111111111111100100011100010;
assign LUT_4[21129] = 32'b11111111111111110101101111011010;
assign LUT_4[21130] = 32'b11111111111111111011111110000110;
assign LUT_4[21131] = 32'b11111111111111110101001001111110;
assign LUT_4[21132] = 32'b11111111111111111001100011111110;
assign LUT_4[21133] = 32'b11111111111111110010101111110110;
assign LUT_4[21134] = 32'b11111111111111111000111110100010;
assign LUT_4[21135] = 32'b11111111111111110010001010011010;
assign LUT_4[21136] = 32'b00000000000000000001001000111011;
assign LUT_4[21137] = 32'b11111111111111111010010100110011;
assign LUT_4[21138] = 32'b00000000000000000000100011011111;
assign LUT_4[21139] = 32'b11111111111111111001101111010111;
assign LUT_4[21140] = 32'b11111111111111111110001001010111;
assign LUT_4[21141] = 32'b11111111111111110111010101001111;
assign LUT_4[21142] = 32'b11111111111111111101100011111011;
assign LUT_4[21143] = 32'b11111111111111110110101111110011;
assign LUT_4[21144] = 32'b11111111111111111010010101010000;
assign LUT_4[21145] = 32'b11111111111111110011100001001000;
assign LUT_4[21146] = 32'b11111111111111111001101111110100;
assign LUT_4[21147] = 32'b11111111111111110010111011101100;
assign LUT_4[21148] = 32'b11111111111111110111010101101100;
assign LUT_4[21149] = 32'b11111111111111110000100001100100;
assign LUT_4[21150] = 32'b11111111111111110110110000010000;
assign LUT_4[21151] = 32'b11111111111111101111111100001000;
assign LUT_4[21152] = 32'b00000000000000000001110010010100;
assign LUT_4[21153] = 32'b11111111111111111010111110001100;
assign LUT_4[21154] = 32'b00000000000000000001001100111000;
assign LUT_4[21155] = 32'b11111111111111111010011000110000;
assign LUT_4[21156] = 32'b11111111111111111110110010110000;
assign LUT_4[21157] = 32'b11111111111111110111111110101000;
assign LUT_4[21158] = 32'b11111111111111111110001101010100;
assign LUT_4[21159] = 32'b11111111111111110111011001001100;
assign LUT_4[21160] = 32'b11111111111111111010111110101001;
assign LUT_4[21161] = 32'b11111111111111110100001010100001;
assign LUT_4[21162] = 32'b11111111111111111010011001001101;
assign LUT_4[21163] = 32'b11111111111111110011100101000101;
assign LUT_4[21164] = 32'b11111111111111110111111111000101;
assign LUT_4[21165] = 32'b11111111111111110001001010111101;
assign LUT_4[21166] = 32'b11111111111111110111011001101001;
assign LUT_4[21167] = 32'b11111111111111110000100101100001;
assign LUT_4[21168] = 32'b11111111111111111111100100000010;
assign LUT_4[21169] = 32'b11111111111111111000101111111010;
assign LUT_4[21170] = 32'b11111111111111111110111110100110;
assign LUT_4[21171] = 32'b11111111111111111000001010011110;
assign LUT_4[21172] = 32'b11111111111111111100100100011110;
assign LUT_4[21173] = 32'b11111111111111110101110000010110;
assign LUT_4[21174] = 32'b11111111111111111011111111000010;
assign LUT_4[21175] = 32'b11111111111111110101001010111010;
assign LUT_4[21176] = 32'b11111111111111111000110000010111;
assign LUT_4[21177] = 32'b11111111111111110001111100001111;
assign LUT_4[21178] = 32'b11111111111111111000001010111011;
assign LUT_4[21179] = 32'b11111111111111110001010110110011;
assign LUT_4[21180] = 32'b11111111111111110101110000110011;
assign LUT_4[21181] = 32'b11111111111111101110111100101011;
assign LUT_4[21182] = 32'b11111111111111110101001011010111;
assign LUT_4[21183] = 32'b11111111111111101110010111001111;
assign LUT_4[21184] = 32'b00000000000000000100101110100001;
assign LUT_4[21185] = 32'b11111111111111111101111010011001;
assign LUT_4[21186] = 32'b00000000000000000100001001000101;
assign LUT_4[21187] = 32'b11111111111111111101010100111101;
assign LUT_4[21188] = 32'b00000000000000000001101110111101;
assign LUT_4[21189] = 32'b11111111111111111010111010110101;
assign LUT_4[21190] = 32'b00000000000000000001001001100001;
assign LUT_4[21191] = 32'b11111111111111111010010101011001;
assign LUT_4[21192] = 32'b11111111111111111101111010110110;
assign LUT_4[21193] = 32'b11111111111111110111000110101110;
assign LUT_4[21194] = 32'b11111111111111111101010101011010;
assign LUT_4[21195] = 32'b11111111111111110110100001010010;
assign LUT_4[21196] = 32'b11111111111111111010111011010010;
assign LUT_4[21197] = 32'b11111111111111110100000111001010;
assign LUT_4[21198] = 32'b11111111111111111010010101110110;
assign LUT_4[21199] = 32'b11111111111111110011100001101110;
assign LUT_4[21200] = 32'b00000000000000000010100000001111;
assign LUT_4[21201] = 32'b11111111111111111011101100000111;
assign LUT_4[21202] = 32'b00000000000000000001111010110011;
assign LUT_4[21203] = 32'b11111111111111111011000110101011;
assign LUT_4[21204] = 32'b11111111111111111111100000101011;
assign LUT_4[21205] = 32'b11111111111111111000101100100011;
assign LUT_4[21206] = 32'b11111111111111111110111011001111;
assign LUT_4[21207] = 32'b11111111111111111000000111000111;
assign LUT_4[21208] = 32'b11111111111111111011101100100100;
assign LUT_4[21209] = 32'b11111111111111110100111000011100;
assign LUT_4[21210] = 32'b11111111111111111011000111001000;
assign LUT_4[21211] = 32'b11111111111111110100010011000000;
assign LUT_4[21212] = 32'b11111111111111111000101101000000;
assign LUT_4[21213] = 32'b11111111111111110001111000111000;
assign LUT_4[21214] = 32'b11111111111111111000000111100100;
assign LUT_4[21215] = 32'b11111111111111110001010011011100;
assign LUT_4[21216] = 32'b00000000000000000011001001101000;
assign LUT_4[21217] = 32'b11111111111111111100010101100000;
assign LUT_4[21218] = 32'b00000000000000000010100100001100;
assign LUT_4[21219] = 32'b11111111111111111011110000000100;
assign LUT_4[21220] = 32'b00000000000000000000001010000100;
assign LUT_4[21221] = 32'b11111111111111111001010101111100;
assign LUT_4[21222] = 32'b11111111111111111111100100101000;
assign LUT_4[21223] = 32'b11111111111111111000110000100000;
assign LUT_4[21224] = 32'b11111111111111111100010101111101;
assign LUT_4[21225] = 32'b11111111111111110101100001110101;
assign LUT_4[21226] = 32'b11111111111111111011110000100001;
assign LUT_4[21227] = 32'b11111111111111110100111100011001;
assign LUT_4[21228] = 32'b11111111111111111001010110011001;
assign LUT_4[21229] = 32'b11111111111111110010100010010001;
assign LUT_4[21230] = 32'b11111111111111111000110000111101;
assign LUT_4[21231] = 32'b11111111111111110001111100110101;
assign LUT_4[21232] = 32'b00000000000000000000111011010110;
assign LUT_4[21233] = 32'b11111111111111111010000111001110;
assign LUT_4[21234] = 32'b00000000000000000000010101111010;
assign LUT_4[21235] = 32'b11111111111111111001100001110010;
assign LUT_4[21236] = 32'b11111111111111111101111011110010;
assign LUT_4[21237] = 32'b11111111111111110111000111101010;
assign LUT_4[21238] = 32'b11111111111111111101010110010110;
assign LUT_4[21239] = 32'b11111111111111110110100010001110;
assign LUT_4[21240] = 32'b11111111111111111010000111101011;
assign LUT_4[21241] = 32'b11111111111111110011010011100011;
assign LUT_4[21242] = 32'b11111111111111111001100010001111;
assign LUT_4[21243] = 32'b11111111111111110010101110000111;
assign LUT_4[21244] = 32'b11111111111111110111001000000111;
assign LUT_4[21245] = 32'b11111111111111110000010011111111;
assign LUT_4[21246] = 32'b11111111111111110110100010101011;
assign LUT_4[21247] = 32'b11111111111111101111101110100011;
assign LUT_4[21248] = 32'b00000000000000000101101100101000;
assign LUT_4[21249] = 32'b11111111111111111110111000100000;
assign LUT_4[21250] = 32'b00000000000000000101000111001100;
assign LUT_4[21251] = 32'b11111111111111111110010011000100;
assign LUT_4[21252] = 32'b00000000000000000010101101000100;
assign LUT_4[21253] = 32'b11111111111111111011111000111100;
assign LUT_4[21254] = 32'b00000000000000000010000111101000;
assign LUT_4[21255] = 32'b11111111111111111011010011100000;
assign LUT_4[21256] = 32'b11111111111111111110111000111101;
assign LUT_4[21257] = 32'b11111111111111111000000100110101;
assign LUT_4[21258] = 32'b11111111111111111110010011100001;
assign LUT_4[21259] = 32'b11111111111111110111011111011001;
assign LUT_4[21260] = 32'b11111111111111111011111001011001;
assign LUT_4[21261] = 32'b11111111111111110101000101010001;
assign LUT_4[21262] = 32'b11111111111111111011010011111101;
assign LUT_4[21263] = 32'b11111111111111110100011111110101;
assign LUT_4[21264] = 32'b00000000000000000011011110010110;
assign LUT_4[21265] = 32'b11111111111111111100101010001110;
assign LUT_4[21266] = 32'b00000000000000000010111000111010;
assign LUT_4[21267] = 32'b11111111111111111100000100110010;
assign LUT_4[21268] = 32'b00000000000000000000011110110010;
assign LUT_4[21269] = 32'b11111111111111111001101010101010;
assign LUT_4[21270] = 32'b11111111111111111111111001010110;
assign LUT_4[21271] = 32'b11111111111111111001000101001110;
assign LUT_4[21272] = 32'b11111111111111111100101010101011;
assign LUT_4[21273] = 32'b11111111111111110101110110100011;
assign LUT_4[21274] = 32'b11111111111111111100000101001111;
assign LUT_4[21275] = 32'b11111111111111110101010001000111;
assign LUT_4[21276] = 32'b11111111111111111001101011000111;
assign LUT_4[21277] = 32'b11111111111111110010110110111111;
assign LUT_4[21278] = 32'b11111111111111111001000101101011;
assign LUT_4[21279] = 32'b11111111111111110010010001100011;
assign LUT_4[21280] = 32'b00000000000000000100000111101111;
assign LUT_4[21281] = 32'b11111111111111111101010011100111;
assign LUT_4[21282] = 32'b00000000000000000011100010010011;
assign LUT_4[21283] = 32'b11111111111111111100101110001011;
assign LUT_4[21284] = 32'b00000000000000000001001000001011;
assign LUT_4[21285] = 32'b11111111111111111010010100000011;
assign LUT_4[21286] = 32'b00000000000000000000100010101111;
assign LUT_4[21287] = 32'b11111111111111111001101110100111;
assign LUT_4[21288] = 32'b11111111111111111101010100000100;
assign LUT_4[21289] = 32'b11111111111111110110011111111100;
assign LUT_4[21290] = 32'b11111111111111111100101110101000;
assign LUT_4[21291] = 32'b11111111111111110101111010100000;
assign LUT_4[21292] = 32'b11111111111111111010010100100000;
assign LUT_4[21293] = 32'b11111111111111110011100000011000;
assign LUT_4[21294] = 32'b11111111111111111001101111000100;
assign LUT_4[21295] = 32'b11111111111111110010111010111100;
assign LUT_4[21296] = 32'b00000000000000000001111001011101;
assign LUT_4[21297] = 32'b11111111111111111011000101010101;
assign LUT_4[21298] = 32'b00000000000000000001010100000001;
assign LUT_4[21299] = 32'b11111111111111111010011111111001;
assign LUT_4[21300] = 32'b11111111111111111110111001111001;
assign LUT_4[21301] = 32'b11111111111111111000000101110001;
assign LUT_4[21302] = 32'b11111111111111111110010100011101;
assign LUT_4[21303] = 32'b11111111111111110111100000010101;
assign LUT_4[21304] = 32'b11111111111111111011000101110010;
assign LUT_4[21305] = 32'b11111111111111110100010001101010;
assign LUT_4[21306] = 32'b11111111111111111010100000010110;
assign LUT_4[21307] = 32'b11111111111111110011101100001110;
assign LUT_4[21308] = 32'b11111111111111111000000110001110;
assign LUT_4[21309] = 32'b11111111111111110001010010000110;
assign LUT_4[21310] = 32'b11111111111111110111100000110010;
assign LUT_4[21311] = 32'b11111111111111110000101100101010;
assign LUT_4[21312] = 32'b00000000000000000111000011111100;
assign LUT_4[21313] = 32'b00000000000000000000001111110100;
assign LUT_4[21314] = 32'b00000000000000000110011110100000;
assign LUT_4[21315] = 32'b11111111111111111111101010011000;
assign LUT_4[21316] = 32'b00000000000000000100000100011000;
assign LUT_4[21317] = 32'b11111111111111111101010000010000;
assign LUT_4[21318] = 32'b00000000000000000011011110111100;
assign LUT_4[21319] = 32'b11111111111111111100101010110100;
assign LUT_4[21320] = 32'b00000000000000000000010000010001;
assign LUT_4[21321] = 32'b11111111111111111001011100001001;
assign LUT_4[21322] = 32'b11111111111111111111101010110101;
assign LUT_4[21323] = 32'b11111111111111111000110110101101;
assign LUT_4[21324] = 32'b11111111111111111101010000101101;
assign LUT_4[21325] = 32'b11111111111111110110011100100101;
assign LUT_4[21326] = 32'b11111111111111111100101011010001;
assign LUT_4[21327] = 32'b11111111111111110101110111001001;
assign LUT_4[21328] = 32'b00000000000000000100110101101010;
assign LUT_4[21329] = 32'b11111111111111111110000001100010;
assign LUT_4[21330] = 32'b00000000000000000100010000001110;
assign LUT_4[21331] = 32'b11111111111111111101011100000110;
assign LUT_4[21332] = 32'b00000000000000000001110110000110;
assign LUT_4[21333] = 32'b11111111111111111011000001111110;
assign LUT_4[21334] = 32'b00000000000000000001010000101010;
assign LUT_4[21335] = 32'b11111111111111111010011100100010;
assign LUT_4[21336] = 32'b11111111111111111110000001111111;
assign LUT_4[21337] = 32'b11111111111111110111001101110111;
assign LUT_4[21338] = 32'b11111111111111111101011100100011;
assign LUT_4[21339] = 32'b11111111111111110110101000011011;
assign LUT_4[21340] = 32'b11111111111111111011000010011011;
assign LUT_4[21341] = 32'b11111111111111110100001110010011;
assign LUT_4[21342] = 32'b11111111111111111010011100111111;
assign LUT_4[21343] = 32'b11111111111111110011101000110111;
assign LUT_4[21344] = 32'b00000000000000000101011111000011;
assign LUT_4[21345] = 32'b11111111111111111110101010111011;
assign LUT_4[21346] = 32'b00000000000000000100111001100111;
assign LUT_4[21347] = 32'b11111111111111111110000101011111;
assign LUT_4[21348] = 32'b00000000000000000010011111011111;
assign LUT_4[21349] = 32'b11111111111111111011101011010111;
assign LUT_4[21350] = 32'b00000000000000000001111010000011;
assign LUT_4[21351] = 32'b11111111111111111011000101111011;
assign LUT_4[21352] = 32'b11111111111111111110101011011000;
assign LUT_4[21353] = 32'b11111111111111110111110111010000;
assign LUT_4[21354] = 32'b11111111111111111110000101111100;
assign LUT_4[21355] = 32'b11111111111111110111010001110100;
assign LUT_4[21356] = 32'b11111111111111111011101011110100;
assign LUT_4[21357] = 32'b11111111111111110100110111101100;
assign LUT_4[21358] = 32'b11111111111111111011000110011000;
assign LUT_4[21359] = 32'b11111111111111110100010010010000;
assign LUT_4[21360] = 32'b00000000000000000011010000110001;
assign LUT_4[21361] = 32'b11111111111111111100011100101001;
assign LUT_4[21362] = 32'b00000000000000000010101011010101;
assign LUT_4[21363] = 32'b11111111111111111011110111001101;
assign LUT_4[21364] = 32'b00000000000000000000010001001101;
assign LUT_4[21365] = 32'b11111111111111111001011101000101;
assign LUT_4[21366] = 32'b11111111111111111111101011110001;
assign LUT_4[21367] = 32'b11111111111111111000110111101001;
assign LUT_4[21368] = 32'b11111111111111111100011101000110;
assign LUT_4[21369] = 32'b11111111111111110101101000111110;
assign LUT_4[21370] = 32'b11111111111111111011110111101010;
assign LUT_4[21371] = 32'b11111111111111110101000011100010;
assign LUT_4[21372] = 32'b11111111111111111001011101100010;
assign LUT_4[21373] = 32'b11111111111111110010101001011010;
assign LUT_4[21374] = 32'b11111111111111111000111000000110;
assign LUT_4[21375] = 32'b11111111111111110010000011111110;
assign LUT_4[21376] = 32'b00000000000000001000010010110000;
assign LUT_4[21377] = 32'b00000000000000000001011110101000;
assign LUT_4[21378] = 32'b00000000000000000111101101010100;
assign LUT_4[21379] = 32'b00000000000000000000111001001100;
assign LUT_4[21380] = 32'b00000000000000000101010011001100;
assign LUT_4[21381] = 32'b11111111111111111110011111000100;
assign LUT_4[21382] = 32'b00000000000000000100101101110000;
assign LUT_4[21383] = 32'b11111111111111111101111001101000;
assign LUT_4[21384] = 32'b00000000000000000001011111000101;
assign LUT_4[21385] = 32'b11111111111111111010101010111101;
assign LUT_4[21386] = 32'b00000000000000000000111001101001;
assign LUT_4[21387] = 32'b11111111111111111010000101100001;
assign LUT_4[21388] = 32'b11111111111111111110011111100001;
assign LUT_4[21389] = 32'b11111111111111110111101011011001;
assign LUT_4[21390] = 32'b11111111111111111101111010000101;
assign LUT_4[21391] = 32'b11111111111111110111000101111101;
assign LUT_4[21392] = 32'b00000000000000000110000100011110;
assign LUT_4[21393] = 32'b11111111111111111111010000010110;
assign LUT_4[21394] = 32'b00000000000000000101011111000010;
assign LUT_4[21395] = 32'b11111111111111111110101010111010;
assign LUT_4[21396] = 32'b00000000000000000011000100111010;
assign LUT_4[21397] = 32'b11111111111111111100010000110010;
assign LUT_4[21398] = 32'b00000000000000000010011111011110;
assign LUT_4[21399] = 32'b11111111111111111011101011010110;
assign LUT_4[21400] = 32'b11111111111111111111010000110011;
assign LUT_4[21401] = 32'b11111111111111111000011100101011;
assign LUT_4[21402] = 32'b11111111111111111110101011010111;
assign LUT_4[21403] = 32'b11111111111111110111110111001111;
assign LUT_4[21404] = 32'b11111111111111111100010001001111;
assign LUT_4[21405] = 32'b11111111111111110101011101000111;
assign LUT_4[21406] = 32'b11111111111111111011101011110011;
assign LUT_4[21407] = 32'b11111111111111110100110111101011;
assign LUT_4[21408] = 32'b00000000000000000110101101110111;
assign LUT_4[21409] = 32'b11111111111111111111111001101111;
assign LUT_4[21410] = 32'b00000000000000000110001000011011;
assign LUT_4[21411] = 32'b11111111111111111111010100010011;
assign LUT_4[21412] = 32'b00000000000000000011101110010011;
assign LUT_4[21413] = 32'b11111111111111111100111010001011;
assign LUT_4[21414] = 32'b00000000000000000011001000110111;
assign LUT_4[21415] = 32'b11111111111111111100010100101111;
assign LUT_4[21416] = 32'b11111111111111111111111010001100;
assign LUT_4[21417] = 32'b11111111111111111001000110000100;
assign LUT_4[21418] = 32'b11111111111111111111010100110000;
assign LUT_4[21419] = 32'b11111111111111111000100000101000;
assign LUT_4[21420] = 32'b11111111111111111100111010101000;
assign LUT_4[21421] = 32'b11111111111111110110000110100000;
assign LUT_4[21422] = 32'b11111111111111111100010101001100;
assign LUT_4[21423] = 32'b11111111111111110101100001000100;
assign LUT_4[21424] = 32'b00000000000000000100011111100101;
assign LUT_4[21425] = 32'b11111111111111111101101011011101;
assign LUT_4[21426] = 32'b00000000000000000011111010001001;
assign LUT_4[21427] = 32'b11111111111111111101000110000001;
assign LUT_4[21428] = 32'b00000000000000000001100000000001;
assign LUT_4[21429] = 32'b11111111111111111010101011111001;
assign LUT_4[21430] = 32'b00000000000000000000111010100101;
assign LUT_4[21431] = 32'b11111111111111111010000110011101;
assign LUT_4[21432] = 32'b11111111111111111101101011111010;
assign LUT_4[21433] = 32'b11111111111111110110110111110010;
assign LUT_4[21434] = 32'b11111111111111111101000110011110;
assign LUT_4[21435] = 32'b11111111111111110110010010010110;
assign LUT_4[21436] = 32'b11111111111111111010101100010110;
assign LUT_4[21437] = 32'b11111111111111110011111000001110;
assign LUT_4[21438] = 32'b11111111111111111010000110111010;
assign LUT_4[21439] = 32'b11111111111111110011010010110010;
assign LUT_4[21440] = 32'b00000000000000001001101010000100;
assign LUT_4[21441] = 32'b00000000000000000010110101111100;
assign LUT_4[21442] = 32'b00000000000000001001000100101000;
assign LUT_4[21443] = 32'b00000000000000000010010000100000;
assign LUT_4[21444] = 32'b00000000000000000110101010100000;
assign LUT_4[21445] = 32'b11111111111111111111110110011000;
assign LUT_4[21446] = 32'b00000000000000000110000101000100;
assign LUT_4[21447] = 32'b11111111111111111111010000111100;
assign LUT_4[21448] = 32'b00000000000000000010110110011001;
assign LUT_4[21449] = 32'b11111111111111111100000010010001;
assign LUT_4[21450] = 32'b00000000000000000010010000111101;
assign LUT_4[21451] = 32'b11111111111111111011011100110101;
assign LUT_4[21452] = 32'b11111111111111111111110110110101;
assign LUT_4[21453] = 32'b11111111111111111001000010101101;
assign LUT_4[21454] = 32'b11111111111111111111010001011001;
assign LUT_4[21455] = 32'b11111111111111111000011101010001;
assign LUT_4[21456] = 32'b00000000000000000111011011110010;
assign LUT_4[21457] = 32'b00000000000000000000100111101010;
assign LUT_4[21458] = 32'b00000000000000000110110110010110;
assign LUT_4[21459] = 32'b00000000000000000000000010001110;
assign LUT_4[21460] = 32'b00000000000000000100011100001110;
assign LUT_4[21461] = 32'b11111111111111111101101000000110;
assign LUT_4[21462] = 32'b00000000000000000011110110110010;
assign LUT_4[21463] = 32'b11111111111111111101000010101010;
assign LUT_4[21464] = 32'b00000000000000000000101000000111;
assign LUT_4[21465] = 32'b11111111111111111001110011111111;
assign LUT_4[21466] = 32'b00000000000000000000000010101011;
assign LUT_4[21467] = 32'b11111111111111111001001110100011;
assign LUT_4[21468] = 32'b11111111111111111101101000100011;
assign LUT_4[21469] = 32'b11111111111111110110110100011011;
assign LUT_4[21470] = 32'b11111111111111111101000011000111;
assign LUT_4[21471] = 32'b11111111111111110110001110111111;
assign LUT_4[21472] = 32'b00000000000000001000000101001011;
assign LUT_4[21473] = 32'b00000000000000000001010001000011;
assign LUT_4[21474] = 32'b00000000000000000111011111101111;
assign LUT_4[21475] = 32'b00000000000000000000101011100111;
assign LUT_4[21476] = 32'b00000000000000000101000101100111;
assign LUT_4[21477] = 32'b11111111111111111110010001011111;
assign LUT_4[21478] = 32'b00000000000000000100100000001011;
assign LUT_4[21479] = 32'b11111111111111111101101100000011;
assign LUT_4[21480] = 32'b00000000000000000001010001100000;
assign LUT_4[21481] = 32'b11111111111111111010011101011000;
assign LUT_4[21482] = 32'b00000000000000000000101100000100;
assign LUT_4[21483] = 32'b11111111111111111001110111111100;
assign LUT_4[21484] = 32'b11111111111111111110010001111100;
assign LUT_4[21485] = 32'b11111111111111110111011101110100;
assign LUT_4[21486] = 32'b11111111111111111101101100100000;
assign LUT_4[21487] = 32'b11111111111111110110111000011000;
assign LUT_4[21488] = 32'b00000000000000000101110110111001;
assign LUT_4[21489] = 32'b11111111111111111111000010110001;
assign LUT_4[21490] = 32'b00000000000000000101010001011101;
assign LUT_4[21491] = 32'b11111111111111111110011101010101;
assign LUT_4[21492] = 32'b00000000000000000010110111010101;
assign LUT_4[21493] = 32'b11111111111111111100000011001101;
assign LUT_4[21494] = 32'b00000000000000000010010001111001;
assign LUT_4[21495] = 32'b11111111111111111011011101110001;
assign LUT_4[21496] = 32'b11111111111111111111000011001110;
assign LUT_4[21497] = 32'b11111111111111111000001111000110;
assign LUT_4[21498] = 32'b11111111111111111110011101110010;
assign LUT_4[21499] = 32'b11111111111111110111101001101010;
assign LUT_4[21500] = 32'b11111111111111111100000011101010;
assign LUT_4[21501] = 32'b11111111111111110101001111100010;
assign LUT_4[21502] = 32'b11111111111111111011011110001110;
assign LUT_4[21503] = 32'b11111111111111110100101010000110;
assign LUT_4[21504] = 32'b00000000000000000011010111011100;
assign LUT_4[21505] = 32'b11111111111111111100100011010100;
assign LUT_4[21506] = 32'b00000000000000000010110010000000;
assign LUT_4[21507] = 32'b11111111111111111011111101111000;
assign LUT_4[21508] = 32'b00000000000000000000010111111000;
assign LUT_4[21509] = 32'b11111111111111111001100011110000;
assign LUT_4[21510] = 32'b11111111111111111111110010011100;
assign LUT_4[21511] = 32'b11111111111111111000111110010100;
assign LUT_4[21512] = 32'b11111111111111111100100011110001;
assign LUT_4[21513] = 32'b11111111111111110101101111101001;
assign LUT_4[21514] = 32'b11111111111111111011111110010101;
assign LUT_4[21515] = 32'b11111111111111110101001010001101;
assign LUT_4[21516] = 32'b11111111111111111001100100001101;
assign LUT_4[21517] = 32'b11111111111111110010110000000101;
assign LUT_4[21518] = 32'b11111111111111111000111110110001;
assign LUT_4[21519] = 32'b11111111111111110010001010101001;
assign LUT_4[21520] = 32'b00000000000000000001001001001010;
assign LUT_4[21521] = 32'b11111111111111111010010101000010;
assign LUT_4[21522] = 32'b00000000000000000000100011101110;
assign LUT_4[21523] = 32'b11111111111111111001101111100110;
assign LUT_4[21524] = 32'b11111111111111111110001001100110;
assign LUT_4[21525] = 32'b11111111111111110111010101011110;
assign LUT_4[21526] = 32'b11111111111111111101100100001010;
assign LUT_4[21527] = 32'b11111111111111110110110000000010;
assign LUT_4[21528] = 32'b11111111111111111010010101011111;
assign LUT_4[21529] = 32'b11111111111111110011100001010111;
assign LUT_4[21530] = 32'b11111111111111111001110000000011;
assign LUT_4[21531] = 32'b11111111111111110010111011111011;
assign LUT_4[21532] = 32'b11111111111111110111010101111011;
assign LUT_4[21533] = 32'b11111111111111110000100001110011;
assign LUT_4[21534] = 32'b11111111111111110110110000011111;
assign LUT_4[21535] = 32'b11111111111111101111111100010111;
assign LUT_4[21536] = 32'b00000000000000000001110010100011;
assign LUT_4[21537] = 32'b11111111111111111010111110011011;
assign LUT_4[21538] = 32'b00000000000000000001001101000111;
assign LUT_4[21539] = 32'b11111111111111111010011000111111;
assign LUT_4[21540] = 32'b11111111111111111110110010111111;
assign LUT_4[21541] = 32'b11111111111111110111111110110111;
assign LUT_4[21542] = 32'b11111111111111111110001101100011;
assign LUT_4[21543] = 32'b11111111111111110111011001011011;
assign LUT_4[21544] = 32'b11111111111111111010111110111000;
assign LUT_4[21545] = 32'b11111111111111110100001010110000;
assign LUT_4[21546] = 32'b11111111111111111010011001011100;
assign LUT_4[21547] = 32'b11111111111111110011100101010100;
assign LUT_4[21548] = 32'b11111111111111110111111111010100;
assign LUT_4[21549] = 32'b11111111111111110001001011001100;
assign LUT_4[21550] = 32'b11111111111111110111011001111000;
assign LUT_4[21551] = 32'b11111111111111110000100101110000;
assign LUT_4[21552] = 32'b11111111111111111111100100010001;
assign LUT_4[21553] = 32'b11111111111111111000110000001001;
assign LUT_4[21554] = 32'b11111111111111111110111110110101;
assign LUT_4[21555] = 32'b11111111111111111000001010101101;
assign LUT_4[21556] = 32'b11111111111111111100100100101101;
assign LUT_4[21557] = 32'b11111111111111110101110000100101;
assign LUT_4[21558] = 32'b11111111111111111011111111010001;
assign LUT_4[21559] = 32'b11111111111111110101001011001001;
assign LUT_4[21560] = 32'b11111111111111111000110000100110;
assign LUT_4[21561] = 32'b11111111111111110001111100011110;
assign LUT_4[21562] = 32'b11111111111111111000001011001010;
assign LUT_4[21563] = 32'b11111111111111110001010111000010;
assign LUT_4[21564] = 32'b11111111111111110101110001000010;
assign LUT_4[21565] = 32'b11111111111111101110111100111010;
assign LUT_4[21566] = 32'b11111111111111110101001011100110;
assign LUT_4[21567] = 32'b11111111111111101110010111011110;
assign LUT_4[21568] = 32'b00000000000000000100101110110000;
assign LUT_4[21569] = 32'b11111111111111111101111010101000;
assign LUT_4[21570] = 32'b00000000000000000100001001010100;
assign LUT_4[21571] = 32'b11111111111111111101010101001100;
assign LUT_4[21572] = 32'b00000000000000000001101111001100;
assign LUT_4[21573] = 32'b11111111111111111010111011000100;
assign LUT_4[21574] = 32'b00000000000000000001001001110000;
assign LUT_4[21575] = 32'b11111111111111111010010101101000;
assign LUT_4[21576] = 32'b11111111111111111101111011000101;
assign LUT_4[21577] = 32'b11111111111111110111000110111101;
assign LUT_4[21578] = 32'b11111111111111111101010101101001;
assign LUT_4[21579] = 32'b11111111111111110110100001100001;
assign LUT_4[21580] = 32'b11111111111111111010111011100001;
assign LUT_4[21581] = 32'b11111111111111110100000111011001;
assign LUT_4[21582] = 32'b11111111111111111010010110000101;
assign LUT_4[21583] = 32'b11111111111111110011100001111101;
assign LUT_4[21584] = 32'b00000000000000000010100000011110;
assign LUT_4[21585] = 32'b11111111111111111011101100010110;
assign LUT_4[21586] = 32'b00000000000000000001111011000010;
assign LUT_4[21587] = 32'b11111111111111111011000110111010;
assign LUT_4[21588] = 32'b11111111111111111111100000111010;
assign LUT_4[21589] = 32'b11111111111111111000101100110010;
assign LUT_4[21590] = 32'b11111111111111111110111011011110;
assign LUT_4[21591] = 32'b11111111111111111000000111010110;
assign LUT_4[21592] = 32'b11111111111111111011101100110011;
assign LUT_4[21593] = 32'b11111111111111110100111000101011;
assign LUT_4[21594] = 32'b11111111111111111011000111010111;
assign LUT_4[21595] = 32'b11111111111111110100010011001111;
assign LUT_4[21596] = 32'b11111111111111111000101101001111;
assign LUT_4[21597] = 32'b11111111111111110001111001000111;
assign LUT_4[21598] = 32'b11111111111111111000000111110011;
assign LUT_4[21599] = 32'b11111111111111110001010011101011;
assign LUT_4[21600] = 32'b00000000000000000011001001110111;
assign LUT_4[21601] = 32'b11111111111111111100010101101111;
assign LUT_4[21602] = 32'b00000000000000000010100100011011;
assign LUT_4[21603] = 32'b11111111111111111011110000010011;
assign LUT_4[21604] = 32'b00000000000000000000001010010011;
assign LUT_4[21605] = 32'b11111111111111111001010110001011;
assign LUT_4[21606] = 32'b11111111111111111111100100110111;
assign LUT_4[21607] = 32'b11111111111111111000110000101111;
assign LUT_4[21608] = 32'b11111111111111111100010110001100;
assign LUT_4[21609] = 32'b11111111111111110101100010000100;
assign LUT_4[21610] = 32'b11111111111111111011110000110000;
assign LUT_4[21611] = 32'b11111111111111110100111100101000;
assign LUT_4[21612] = 32'b11111111111111111001010110101000;
assign LUT_4[21613] = 32'b11111111111111110010100010100000;
assign LUT_4[21614] = 32'b11111111111111111000110001001100;
assign LUT_4[21615] = 32'b11111111111111110001111101000100;
assign LUT_4[21616] = 32'b00000000000000000000111011100101;
assign LUT_4[21617] = 32'b11111111111111111010000111011101;
assign LUT_4[21618] = 32'b00000000000000000000010110001001;
assign LUT_4[21619] = 32'b11111111111111111001100010000001;
assign LUT_4[21620] = 32'b11111111111111111101111100000001;
assign LUT_4[21621] = 32'b11111111111111110111000111111001;
assign LUT_4[21622] = 32'b11111111111111111101010110100101;
assign LUT_4[21623] = 32'b11111111111111110110100010011101;
assign LUT_4[21624] = 32'b11111111111111111010000111111010;
assign LUT_4[21625] = 32'b11111111111111110011010011110010;
assign LUT_4[21626] = 32'b11111111111111111001100010011110;
assign LUT_4[21627] = 32'b11111111111111110010101110010110;
assign LUT_4[21628] = 32'b11111111111111110111001000010110;
assign LUT_4[21629] = 32'b11111111111111110000010100001110;
assign LUT_4[21630] = 32'b11111111111111110110100010111010;
assign LUT_4[21631] = 32'b11111111111111101111101110110010;
assign LUT_4[21632] = 32'b00000000000000000101111101100100;
assign LUT_4[21633] = 32'b11111111111111111111001001011100;
assign LUT_4[21634] = 32'b00000000000000000101011000001000;
assign LUT_4[21635] = 32'b11111111111111111110100100000000;
assign LUT_4[21636] = 32'b00000000000000000010111110000000;
assign LUT_4[21637] = 32'b11111111111111111100001001111000;
assign LUT_4[21638] = 32'b00000000000000000010011000100100;
assign LUT_4[21639] = 32'b11111111111111111011100100011100;
assign LUT_4[21640] = 32'b11111111111111111111001001111001;
assign LUT_4[21641] = 32'b11111111111111111000010101110001;
assign LUT_4[21642] = 32'b11111111111111111110100100011101;
assign LUT_4[21643] = 32'b11111111111111110111110000010101;
assign LUT_4[21644] = 32'b11111111111111111100001010010101;
assign LUT_4[21645] = 32'b11111111111111110101010110001101;
assign LUT_4[21646] = 32'b11111111111111111011100100111001;
assign LUT_4[21647] = 32'b11111111111111110100110000110001;
assign LUT_4[21648] = 32'b00000000000000000011101111010010;
assign LUT_4[21649] = 32'b11111111111111111100111011001010;
assign LUT_4[21650] = 32'b00000000000000000011001001110110;
assign LUT_4[21651] = 32'b11111111111111111100010101101110;
assign LUT_4[21652] = 32'b00000000000000000000101111101110;
assign LUT_4[21653] = 32'b11111111111111111001111011100110;
assign LUT_4[21654] = 32'b00000000000000000000001010010010;
assign LUT_4[21655] = 32'b11111111111111111001010110001010;
assign LUT_4[21656] = 32'b11111111111111111100111011100111;
assign LUT_4[21657] = 32'b11111111111111110110000111011111;
assign LUT_4[21658] = 32'b11111111111111111100010110001011;
assign LUT_4[21659] = 32'b11111111111111110101100010000011;
assign LUT_4[21660] = 32'b11111111111111111001111100000011;
assign LUT_4[21661] = 32'b11111111111111110011000111111011;
assign LUT_4[21662] = 32'b11111111111111111001010110100111;
assign LUT_4[21663] = 32'b11111111111111110010100010011111;
assign LUT_4[21664] = 32'b00000000000000000100011000101011;
assign LUT_4[21665] = 32'b11111111111111111101100100100011;
assign LUT_4[21666] = 32'b00000000000000000011110011001111;
assign LUT_4[21667] = 32'b11111111111111111100111111000111;
assign LUT_4[21668] = 32'b00000000000000000001011001000111;
assign LUT_4[21669] = 32'b11111111111111111010100100111111;
assign LUT_4[21670] = 32'b00000000000000000000110011101011;
assign LUT_4[21671] = 32'b11111111111111111001111111100011;
assign LUT_4[21672] = 32'b11111111111111111101100101000000;
assign LUT_4[21673] = 32'b11111111111111110110110000111000;
assign LUT_4[21674] = 32'b11111111111111111100111111100100;
assign LUT_4[21675] = 32'b11111111111111110110001011011100;
assign LUT_4[21676] = 32'b11111111111111111010100101011100;
assign LUT_4[21677] = 32'b11111111111111110011110001010100;
assign LUT_4[21678] = 32'b11111111111111111010000000000000;
assign LUT_4[21679] = 32'b11111111111111110011001011111000;
assign LUT_4[21680] = 32'b00000000000000000010001010011001;
assign LUT_4[21681] = 32'b11111111111111111011010110010001;
assign LUT_4[21682] = 32'b00000000000000000001100100111101;
assign LUT_4[21683] = 32'b11111111111111111010110000110101;
assign LUT_4[21684] = 32'b11111111111111111111001010110101;
assign LUT_4[21685] = 32'b11111111111111111000010110101101;
assign LUT_4[21686] = 32'b11111111111111111110100101011001;
assign LUT_4[21687] = 32'b11111111111111110111110001010001;
assign LUT_4[21688] = 32'b11111111111111111011010110101110;
assign LUT_4[21689] = 32'b11111111111111110100100010100110;
assign LUT_4[21690] = 32'b11111111111111111010110001010010;
assign LUT_4[21691] = 32'b11111111111111110011111101001010;
assign LUT_4[21692] = 32'b11111111111111111000010111001010;
assign LUT_4[21693] = 32'b11111111111111110001100011000010;
assign LUT_4[21694] = 32'b11111111111111110111110001101110;
assign LUT_4[21695] = 32'b11111111111111110000111101100110;
assign LUT_4[21696] = 32'b00000000000000000111010100111000;
assign LUT_4[21697] = 32'b00000000000000000000100000110000;
assign LUT_4[21698] = 32'b00000000000000000110101111011100;
assign LUT_4[21699] = 32'b11111111111111111111111011010100;
assign LUT_4[21700] = 32'b00000000000000000100010101010100;
assign LUT_4[21701] = 32'b11111111111111111101100001001100;
assign LUT_4[21702] = 32'b00000000000000000011101111111000;
assign LUT_4[21703] = 32'b11111111111111111100111011110000;
assign LUT_4[21704] = 32'b00000000000000000000100001001101;
assign LUT_4[21705] = 32'b11111111111111111001101101000101;
assign LUT_4[21706] = 32'b11111111111111111111111011110001;
assign LUT_4[21707] = 32'b11111111111111111001000111101001;
assign LUT_4[21708] = 32'b11111111111111111101100001101001;
assign LUT_4[21709] = 32'b11111111111111110110101101100001;
assign LUT_4[21710] = 32'b11111111111111111100111100001101;
assign LUT_4[21711] = 32'b11111111111111110110001000000101;
assign LUT_4[21712] = 32'b00000000000000000101000110100110;
assign LUT_4[21713] = 32'b11111111111111111110010010011110;
assign LUT_4[21714] = 32'b00000000000000000100100001001010;
assign LUT_4[21715] = 32'b11111111111111111101101101000010;
assign LUT_4[21716] = 32'b00000000000000000010000111000010;
assign LUT_4[21717] = 32'b11111111111111111011010010111010;
assign LUT_4[21718] = 32'b00000000000000000001100001100110;
assign LUT_4[21719] = 32'b11111111111111111010101101011110;
assign LUT_4[21720] = 32'b11111111111111111110010010111011;
assign LUT_4[21721] = 32'b11111111111111110111011110110011;
assign LUT_4[21722] = 32'b11111111111111111101101101011111;
assign LUT_4[21723] = 32'b11111111111111110110111001010111;
assign LUT_4[21724] = 32'b11111111111111111011010011010111;
assign LUT_4[21725] = 32'b11111111111111110100011111001111;
assign LUT_4[21726] = 32'b11111111111111111010101101111011;
assign LUT_4[21727] = 32'b11111111111111110011111001110011;
assign LUT_4[21728] = 32'b00000000000000000101101111111111;
assign LUT_4[21729] = 32'b11111111111111111110111011110111;
assign LUT_4[21730] = 32'b00000000000000000101001010100011;
assign LUT_4[21731] = 32'b11111111111111111110010110011011;
assign LUT_4[21732] = 32'b00000000000000000010110000011011;
assign LUT_4[21733] = 32'b11111111111111111011111100010011;
assign LUT_4[21734] = 32'b00000000000000000010001010111111;
assign LUT_4[21735] = 32'b11111111111111111011010110110111;
assign LUT_4[21736] = 32'b11111111111111111110111100010100;
assign LUT_4[21737] = 32'b11111111111111111000001000001100;
assign LUT_4[21738] = 32'b11111111111111111110010110111000;
assign LUT_4[21739] = 32'b11111111111111110111100010110000;
assign LUT_4[21740] = 32'b11111111111111111011111100110000;
assign LUT_4[21741] = 32'b11111111111111110101001000101000;
assign LUT_4[21742] = 32'b11111111111111111011010111010100;
assign LUT_4[21743] = 32'b11111111111111110100100011001100;
assign LUT_4[21744] = 32'b00000000000000000011100001101101;
assign LUT_4[21745] = 32'b11111111111111111100101101100101;
assign LUT_4[21746] = 32'b00000000000000000010111100010001;
assign LUT_4[21747] = 32'b11111111111111111100001000001001;
assign LUT_4[21748] = 32'b00000000000000000000100010001001;
assign LUT_4[21749] = 32'b11111111111111111001101110000001;
assign LUT_4[21750] = 32'b11111111111111111111111100101101;
assign LUT_4[21751] = 32'b11111111111111111001001000100101;
assign LUT_4[21752] = 32'b11111111111111111100101110000010;
assign LUT_4[21753] = 32'b11111111111111110101111001111010;
assign LUT_4[21754] = 32'b11111111111111111100001000100110;
assign LUT_4[21755] = 32'b11111111111111110101010100011110;
assign LUT_4[21756] = 32'b11111111111111111001101110011110;
assign LUT_4[21757] = 32'b11111111111111110010111010010110;
assign LUT_4[21758] = 32'b11111111111111111001001001000010;
assign LUT_4[21759] = 32'b11111111111111110010010100111010;
assign LUT_4[21760] = 32'b00000000000000001000010010111111;
assign LUT_4[21761] = 32'b00000000000000000001011110110111;
assign LUT_4[21762] = 32'b00000000000000000111101101100011;
assign LUT_4[21763] = 32'b00000000000000000000111001011011;
assign LUT_4[21764] = 32'b00000000000000000101010011011011;
assign LUT_4[21765] = 32'b11111111111111111110011111010011;
assign LUT_4[21766] = 32'b00000000000000000100101101111111;
assign LUT_4[21767] = 32'b11111111111111111101111001110111;
assign LUT_4[21768] = 32'b00000000000000000001011111010100;
assign LUT_4[21769] = 32'b11111111111111111010101011001100;
assign LUT_4[21770] = 32'b00000000000000000000111001111000;
assign LUT_4[21771] = 32'b11111111111111111010000101110000;
assign LUT_4[21772] = 32'b11111111111111111110011111110000;
assign LUT_4[21773] = 32'b11111111111111110111101011101000;
assign LUT_4[21774] = 32'b11111111111111111101111010010100;
assign LUT_4[21775] = 32'b11111111111111110111000110001100;
assign LUT_4[21776] = 32'b00000000000000000110000100101101;
assign LUT_4[21777] = 32'b11111111111111111111010000100101;
assign LUT_4[21778] = 32'b00000000000000000101011111010001;
assign LUT_4[21779] = 32'b11111111111111111110101011001001;
assign LUT_4[21780] = 32'b00000000000000000011000101001001;
assign LUT_4[21781] = 32'b11111111111111111100010001000001;
assign LUT_4[21782] = 32'b00000000000000000010011111101101;
assign LUT_4[21783] = 32'b11111111111111111011101011100101;
assign LUT_4[21784] = 32'b11111111111111111111010001000010;
assign LUT_4[21785] = 32'b11111111111111111000011100111010;
assign LUT_4[21786] = 32'b11111111111111111110101011100110;
assign LUT_4[21787] = 32'b11111111111111110111110111011110;
assign LUT_4[21788] = 32'b11111111111111111100010001011110;
assign LUT_4[21789] = 32'b11111111111111110101011101010110;
assign LUT_4[21790] = 32'b11111111111111111011101100000010;
assign LUT_4[21791] = 32'b11111111111111110100110111111010;
assign LUT_4[21792] = 32'b00000000000000000110101110000110;
assign LUT_4[21793] = 32'b11111111111111111111111001111110;
assign LUT_4[21794] = 32'b00000000000000000110001000101010;
assign LUT_4[21795] = 32'b11111111111111111111010100100010;
assign LUT_4[21796] = 32'b00000000000000000011101110100010;
assign LUT_4[21797] = 32'b11111111111111111100111010011010;
assign LUT_4[21798] = 32'b00000000000000000011001001000110;
assign LUT_4[21799] = 32'b11111111111111111100010100111110;
assign LUT_4[21800] = 32'b11111111111111111111111010011011;
assign LUT_4[21801] = 32'b11111111111111111001000110010011;
assign LUT_4[21802] = 32'b11111111111111111111010100111111;
assign LUT_4[21803] = 32'b11111111111111111000100000110111;
assign LUT_4[21804] = 32'b11111111111111111100111010110111;
assign LUT_4[21805] = 32'b11111111111111110110000110101111;
assign LUT_4[21806] = 32'b11111111111111111100010101011011;
assign LUT_4[21807] = 32'b11111111111111110101100001010011;
assign LUT_4[21808] = 32'b00000000000000000100011111110100;
assign LUT_4[21809] = 32'b11111111111111111101101011101100;
assign LUT_4[21810] = 32'b00000000000000000011111010011000;
assign LUT_4[21811] = 32'b11111111111111111101000110010000;
assign LUT_4[21812] = 32'b00000000000000000001100000010000;
assign LUT_4[21813] = 32'b11111111111111111010101100001000;
assign LUT_4[21814] = 32'b00000000000000000000111010110100;
assign LUT_4[21815] = 32'b11111111111111111010000110101100;
assign LUT_4[21816] = 32'b11111111111111111101101100001001;
assign LUT_4[21817] = 32'b11111111111111110110111000000001;
assign LUT_4[21818] = 32'b11111111111111111101000110101101;
assign LUT_4[21819] = 32'b11111111111111110110010010100101;
assign LUT_4[21820] = 32'b11111111111111111010101100100101;
assign LUT_4[21821] = 32'b11111111111111110011111000011101;
assign LUT_4[21822] = 32'b11111111111111111010000111001001;
assign LUT_4[21823] = 32'b11111111111111110011010011000001;
assign LUT_4[21824] = 32'b00000000000000001001101010010011;
assign LUT_4[21825] = 32'b00000000000000000010110110001011;
assign LUT_4[21826] = 32'b00000000000000001001000100110111;
assign LUT_4[21827] = 32'b00000000000000000010010000101111;
assign LUT_4[21828] = 32'b00000000000000000110101010101111;
assign LUT_4[21829] = 32'b11111111111111111111110110100111;
assign LUT_4[21830] = 32'b00000000000000000110000101010011;
assign LUT_4[21831] = 32'b11111111111111111111010001001011;
assign LUT_4[21832] = 32'b00000000000000000010110110101000;
assign LUT_4[21833] = 32'b11111111111111111100000010100000;
assign LUT_4[21834] = 32'b00000000000000000010010001001100;
assign LUT_4[21835] = 32'b11111111111111111011011101000100;
assign LUT_4[21836] = 32'b11111111111111111111110111000100;
assign LUT_4[21837] = 32'b11111111111111111001000010111100;
assign LUT_4[21838] = 32'b11111111111111111111010001101000;
assign LUT_4[21839] = 32'b11111111111111111000011101100000;
assign LUT_4[21840] = 32'b00000000000000000111011100000001;
assign LUT_4[21841] = 32'b00000000000000000000100111111001;
assign LUT_4[21842] = 32'b00000000000000000110110110100101;
assign LUT_4[21843] = 32'b00000000000000000000000010011101;
assign LUT_4[21844] = 32'b00000000000000000100011100011101;
assign LUT_4[21845] = 32'b11111111111111111101101000010101;
assign LUT_4[21846] = 32'b00000000000000000011110111000001;
assign LUT_4[21847] = 32'b11111111111111111101000010111001;
assign LUT_4[21848] = 32'b00000000000000000000101000010110;
assign LUT_4[21849] = 32'b11111111111111111001110100001110;
assign LUT_4[21850] = 32'b00000000000000000000000010111010;
assign LUT_4[21851] = 32'b11111111111111111001001110110010;
assign LUT_4[21852] = 32'b11111111111111111101101000110010;
assign LUT_4[21853] = 32'b11111111111111110110110100101010;
assign LUT_4[21854] = 32'b11111111111111111101000011010110;
assign LUT_4[21855] = 32'b11111111111111110110001111001110;
assign LUT_4[21856] = 32'b00000000000000001000000101011010;
assign LUT_4[21857] = 32'b00000000000000000001010001010010;
assign LUT_4[21858] = 32'b00000000000000000111011111111110;
assign LUT_4[21859] = 32'b00000000000000000000101011110110;
assign LUT_4[21860] = 32'b00000000000000000101000101110110;
assign LUT_4[21861] = 32'b11111111111111111110010001101110;
assign LUT_4[21862] = 32'b00000000000000000100100000011010;
assign LUT_4[21863] = 32'b11111111111111111101101100010010;
assign LUT_4[21864] = 32'b00000000000000000001010001101111;
assign LUT_4[21865] = 32'b11111111111111111010011101100111;
assign LUT_4[21866] = 32'b00000000000000000000101100010011;
assign LUT_4[21867] = 32'b11111111111111111001111000001011;
assign LUT_4[21868] = 32'b11111111111111111110010010001011;
assign LUT_4[21869] = 32'b11111111111111110111011110000011;
assign LUT_4[21870] = 32'b11111111111111111101101100101111;
assign LUT_4[21871] = 32'b11111111111111110110111000100111;
assign LUT_4[21872] = 32'b00000000000000000101110111001000;
assign LUT_4[21873] = 32'b11111111111111111111000011000000;
assign LUT_4[21874] = 32'b00000000000000000101010001101100;
assign LUT_4[21875] = 32'b11111111111111111110011101100100;
assign LUT_4[21876] = 32'b00000000000000000010110111100100;
assign LUT_4[21877] = 32'b11111111111111111100000011011100;
assign LUT_4[21878] = 32'b00000000000000000010010010001000;
assign LUT_4[21879] = 32'b11111111111111111011011110000000;
assign LUT_4[21880] = 32'b11111111111111111111000011011101;
assign LUT_4[21881] = 32'b11111111111111111000001111010101;
assign LUT_4[21882] = 32'b11111111111111111110011110000001;
assign LUT_4[21883] = 32'b11111111111111110111101001111001;
assign LUT_4[21884] = 32'b11111111111111111100000011111001;
assign LUT_4[21885] = 32'b11111111111111110101001111110001;
assign LUT_4[21886] = 32'b11111111111111111011011110011101;
assign LUT_4[21887] = 32'b11111111111111110100101010010101;
assign LUT_4[21888] = 32'b00000000000000001010111001000111;
assign LUT_4[21889] = 32'b00000000000000000100000100111111;
assign LUT_4[21890] = 32'b00000000000000001010010011101011;
assign LUT_4[21891] = 32'b00000000000000000011011111100011;
assign LUT_4[21892] = 32'b00000000000000000111111001100011;
assign LUT_4[21893] = 32'b00000000000000000001000101011011;
assign LUT_4[21894] = 32'b00000000000000000111010100000111;
assign LUT_4[21895] = 32'b00000000000000000000011111111111;
assign LUT_4[21896] = 32'b00000000000000000100000101011100;
assign LUT_4[21897] = 32'b11111111111111111101010001010100;
assign LUT_4[21898] = 32'b00000000000000000011100000000000;
assign LUT_4[21899] = 32'b11111111111111111100101011111000;
assign LUT_4[21900] = 32'b00000000000000000001000101111000;
assign LUT_4[21901] = 32'b11111111111111111010010001110000;
assign LUT_4[21902] = 32'b00000000000000000000100000011100;
assign LUT_4[21903] = 32'b11111111111111111001101100010100;
assign LUT_4[21904] = 32'b00000000000000001000101010110101;
assign LUT_4[21905] = 32'b00000000000000000001110110101101;
assign LUT_4[21906] = 32'b00000000000000001000000101011001;
assign LUT_4[21907] = 32'b00000000000000000001010001010001;
assign LUT_4[21908] = 32'b00000000000000000101101011010001;
assign LUT_4[21909] = 32'b11111111111111111110110111001001;
assign LUT_4[21910] = 32'b00000000000000000101000101110101;
assign LUT_4[21911] = 32'b11111111111111111110010001101101;
assign LUT_4[21912] = 32'b00000000000000000001110111001010;
assign LUT_4[21913] = 32'b11111111111111111011000011000010;
assign LUT_4[21914] = 32'b00000000000000000001010001101110;
assign LUT_4[21915] = 32'b11111111111111111010011101100110;
assign LUT_4[21916] = 32'b11111111111111111110110111100110;
assign LUT_4[21917] = 32'b11111111111111111000000011011110;
assign LUT_4[21918] = 32'b11111111111111111110010010001010;
assign LUT_4[21919] = 32'b11111111111111110111011110000010;
assign LUT_4[21920] = 32'b00000000000000001001010100001110;
assign LUT_4[21921] = 32'b00000000000000000010100000000110;
assign LUT_4[21922] = 32'b00000000000000001000101110110010;
assign LUT_4[21923] = 32'b00000000000000000001111010101010;
assign LUT_4[21924] = 32'b00000000000000000110010100101010;
assign LUT_4[21925] = 32'b11111111111111111111100000100010;
assign LUT_4[21926] = 32'b00000000000000000101101111001110;
assign LUT_4[21927] = 32'b11111111111111111110111011000110;
assign LUT_4[21928] = 32'b00000000000000000010100000100011;
assign LUT_4[21929] = 32'b11111111111111111011101100011011;
assign LUT_4[21930] = 32'b00000000000000000001111011000111;
assign LUT_4[21931] = 32'b11111111111111111011000110111111;
assign LUT_4[21932] = 32'b11111111111111111111100000111111;
assign LUT_4[21933] = 32'b11111111111111111000101100110111;
assign LUT_4[21934] = 32'b11111111111111111110111011100011;
assign LUT_4[21935] = 32'b11111111111111111000000111011011;
assign LUT_4[21936] = 32'b00000000000000000111000101111100;
assign LUT_4[21937] = 32'b00000000000000000000010001110100;
assign LUT_4[21938] = 32'b00000000000000000110100000100000;
assign LUT_4[21939] = 32'b11111111111111111111101100011000;
assign LUT_4[21940] = 32'b00000000000000000100000110011000;
assign LUT_4[21941] = 32'b11111111111111111101010010010000;
assign LUT_4[21942] = 32'b00000000000000000011100000111100;
assign LUT_4[21943] = 32'b11111111111111111100101100110100;
assign LUT_4[21944] = 32'b00000000000000000000010010010001;
assign LUT_4[21945] = 32'b11111111111111111001011110001001;
assign LUT_4[21946] = 32'b11111111111111111111101100110101;
assign LUT_4[21947] = 32'b11111111111111111000111000101101;
assign LUT_4[21948] = 32'b11111111111111111101010010101101;
assign LUT_4[21949] = 32'b11111111111111110110011110100101;
assign LUT_4[21950] = 32'b11111111111111111100101101010001;
assign LUT_4[21951] = 32'b11111111111111110101111001001001;
assign LUT_4[21952] = 32'b00000000000000001100010000011011;
assign LUT_4[21953] = 32'b00000000000000000101011100010011;
assign LUT_4[21954] = 32'b00000000000000001011101010111111;
assign LUT_4[21955] = 32'b00000000000000000100110110110111;
assign LUT_4[21956] = 32'b00000000000000001001010000110111;
assign LUT_4[21957] = 32'b00000000000000000010011100101111;
assign LUT_4[21958] = 32'b00000000000000001000101011011011;
assign LUT_4[21959] = 32'b00000000000000000001110111010011;
assign LUT_4[21960] = 32'b00000000000000000101011100110000;
assign LUT_4[21961] = 32'b11111111111111111110101000101000;
assign LUT_4[21962] = 32'b00000000000000000100110111010100;
assign LUT_4[21963] = 32'b11111111111111111110000011001100;
assign LUT_4[21964] = 32'b00000000000000000010011101001100;
assign LUT_4[21965] = 32'b11111111111111111011101001000100;
assign LUT_4[21966] = 32'b00000000000000000001110111110000;
assign LUT_4[21967] = 32'b11111111111111111011000011101000;
assign LUT_4[21968] = 32'b00000000000000001010000010001001;
assign LUT_4[21969] = 32'b00000000000000000011001110000001;
assign LUT_4[21970] = 32'b00000000000000001001011100101101;
assign LUT_4[21971] = 32'b00000000000000000010101000100101;
assign LUT_4[21972] = 32'b00000000000000000111000010100101;
assign LUT_4[21973] = 32'b00000000000000000000001110011101;
assign LUT_4[21974] = 32'b00000000000000000110011101001001;
assign LUT_4[21975] = 32'b11111111111111111111101001000001;
assign LUT_4[21976] = 32'b00000000000000000011001110011110;
assign LUT_4[21977] = 32'b11111111111111111100011010010110;
assign LUT_4[21978] = 32'b00000000000000000010101001000010;
assign LUT_4[21979] = 32'b11111111111111111011110100111010;
assign LUT_4[21980] = 32'b00000000000000000000001110111010;
assign LUT_4[21981] = 32'b11111111111111111001011010110010;
assign LUT_4[21982] = 32'b11111111111111111111101001011110;
assign LUT_4[21983] = 32'b11111111111111111000110101010110;
assign LUT_4[21984] = 32'b00000000000000001010101011100010;
assign LUT_4[21985] = 32'b00000000000000000011110111011010;
assign LUT_4[21986] = 32'b00000000000000001010000110000110;
assign LUT_4[21987] = 32'b00000000000000000011010001111110;
assign LUT_4[21988] = 32'b00000000000000000111101011111110;
assign LUT_4[21989] = 32'b00000000000000000000110111110110;
assign LUT_4[21990] = 32'b00000000000000000111000110100010;
assign LUT_4[21991] = 32'b00000000000000000000010010011010;
assign LUT_4[21992] = 32'b00000000000000000011110111110111;
assign LUT_4[21993] = 32'b11111111111111111101000011101111;
assign LUT_4[21994] = 32'b00000000000000000011010010011011;
assign LUT_4[21995] = 32'b11111111111111111100011110010011;
assign LUT_4[21996] = 32'b00000000000000000000111000010011;
assign LUT_4[21997] = 32'b11111111111111111010000100001011;
assign LUT_4[21998] = 32'b00000000000000000000010010110111;
assign LUT_4[21999] = 32'b11111111111111111001011110101111;
assign LUT_4[22000] = 32'b00000000000000001000011101010000;
assign LUT_4[22001] = 32'b00000000000000000001101001001000;
assign LUT_4[22002] = 32'b00000000000000000111110111110100;
assign LUT_4[22003] = 32'b00000000000000000001000011101100;
assign LUT_4[22004] = 32'b00000000000000000101011101101100;
assign LUT_4[22005] = 32'b11111111111111111110101001100100;
assign LUT_4[22006] = 32'b00000000000000000100111000010000;
assign LUT_4[22007] = 32'b11111111111111111110000100001000;
assign LUT_4[22008] = 32'b00000000000000000001101001100101;
assign LUT_4[22009] = 32'b11111111111111111010110101011101;
assign LUT_4[22010] = 32'b00000000000000000001000100001001;
assign LUT_4[22011] = 32'b11111111111111111010010000000001;
assign LUT_4[22012] = 32'b11111111111111111110101010000001;
assign LUT_4[22013] = 32'b11111111111111110111110101111001;
assign LUT_4[22014] = 32'b11111111111111111110000100100101;
assign LUT_4[22015] = 32'b11111111111111110111010000011101;
assign LUT_4[22016] = 32'b00000000000000000010011011100100;
assign LUT_4[22017] = 32'b11111111111111111011100111011100;
assign LUT_4[22018] = 32'b00000000000000000001110110001000;
assign LUT_4[22019] = 32'b11111111111111111011000010000000;
assign LUT_4[22020] = 32'b11111111111111111111011100000000;
assign LUT_4[22021] = 32'b11111111111111111000100111111000;
assign LUT_4[22022] = 32'b11111111111111111110110110100100;
assign LUT_4[22023] = 32'b11111111111111111000000010011100;
assign LUT_4[22024] = 32'b11111111111111111011100111111001;
assign LUT_4[22025] = 32'b11111111111111110100110011110001;
assign LUT_4[22026] = 32'b11111111111111111011000010011101;
assign LUT_4[22027] = 32'b11111111111111110100001110010101;
assign LUT_4[22028] = 32'b11111111111111111000101000010101;
assign LUT_4[22029] = 32'b11111111111111110001110100001101;
assign LUT_4[22030] = 32'b11111111111111111000000010111001;
assign LUT_4[22031] = 32'b11111111111111110001001110110001;
assign LUT_4[22032] = 32'b00000000000000000000001101010010;
assign LUT_4[22033] = 32'b11111111111111111001011001001010;
assign LUT_4[22034] = 32'b11111111111111111111100111110110;
assign LUT_4[22035] = 32'b11111111111111111000110011101110;
assign LUT_4[22036] = 32'b11111111111111111101001101101110;
assign LUT_4[22037] = 32'b11111111111111110110011001100110;
assign LUT_4[22038] = 32'b11111111111111111100101000010010;
assign LUT_4[22039] = 32'b11111111111111110101110100001010;
assign LUT_4[22040] = 32'b11111111111111111001011001100111;
assign LUT_4[22041] = 32'b11111111111111110010100101011111;
assign LUT_4[22042] = 32'b11111111111111111000110100001011;
assign LUT_4[22043] = 32'b11111111111111110010000000000011;
assign LUT_4[22044] = 32'b11111111111111110110011010000011;
assign LUT_4[22045] = 32'b11111111111111101111100101111011;
assign LUT_4[22046] = 32'b11111111111111110101110100100111;
assign LUT_4[22047] = 32'b11111111111111101111000000011111;
assign LUT_4[22048] = 32'b00000000000000000000110110101011;
assign LUT_4[22049] = 32'b11111111111111111010000010100011;
assign LUT_4[22050] = 32'b00000000000000000000010001001111;
assign LUT_4[22051] = 32'b11111111111111111001011101000111;
assign LUT_4[22052] = 32'b11111111111111111101110111000111;
assign LUT_4[22053] = 32'b11111111111111110111000010111111;
assign LUT_4[22054] = 32'b11111111111111111101010001101011;
assign LUT_4[22055] = 32'b11111111111111110110011101100011;
assign LUT_4[22056] = 32'b11111111111111111010000011000000;
assign LUT_4[22057] = 32'b11111111111111110011001110111000;
assign LUT_4[22058] = 32'b11111111111111111001011101100100;
assign LUT_4[22059] = 32'b11111111111111110010101001011100;
assign LUT_4[22060] = 32'b11111111111111110111000011011100;
assign LUT_4[22061] = 32'b11111111111111110000001111010100;
assign LUT_4[22062] = 32'b11111111111111110110011110000000;
assign LUT_4[22063] = 32'b11111111111111101111101001111000;
assign LUT_4[22064] = 32'b11111111111111111110101000011001;
assign LUT_4[22065] = 32'b11111111111111110111110100010001;
assign LUT_4[22066] = 32'b11111111111111111110000010111101;
assign LUT_4[22067] = 32'b11111111111111110111001110110101;
assign LUT_4[22068] = 32'b11111111111111111011101000110101;
assign LUT_4[22069] = 32'b11111111111111110100110100101101;
assign LUT_4[22070] = 32'b11111111111111111011000011011001;
assign LUT_4[22071] = 32'b11111111111111110100001111010001;
assign LUT_4[22072] = 32'b11111111111111110111110100101110;
assign LUT_4[22073] = 32'b11111111111111110001000000100110;
assign LUT_4[22074] = 32'b11111111111111110111001111010010;
assign LUT_4[22075] = 32'b11111111111111110000011011001010;
assign LUT_4[22076] = 32'b11111111111111110100110101001010;
assign LUT_4[22077] = 32'b11111111111111101110000001000010;
assign LUT_4[22078] = 32'b11111111111111110100001111101110;
assign LUT_4[22079] = 32'b11111111111111101101011011100110;
assign LUT_4[22080] = 32'b00000000000000000011110010111000;
assign LUT_4[22081] = 32'b11111111111111111100111110110000;
assign LUT_4[22082] = 32'b00000000000000000011001101011100;
assign LUT_4[22083] = 32'b11111111111111111100011001010100;
assign LUT_4[22084] = 32'b00000000000000000000110011010100;
assign LUT_4[22085] = 32'b11111111111111111001111111001100;
assign LUT_4[22086] = 32'b00000000000000000000001101111000;
assign LUT_4[22087] = 32'b11111111111111111001011001110000;
assign LUT_4[22088] = 32'b11111111111111111100111111001101;
assign LUT_4[22089] = 32'b11111111111111110110001011000101;
assign LUT_4[22090] = 32'b11111111111111111100011001110001;
assign LUT_4[22091] = 32'b11111111111111110101100101101001;
assign LUT_4[22092] = 32'b11111111111111111001111111101001;
assign LUT_4[22093] = 32'b11111111111111110011001011100001;
assign LUT_4[22094] = 32'b11111111111111111001011010001101;
assign LUT_4[22095] = 32'b11111111111111110010100110000101;
assign LUT_4[22096] = 32'b00000000000000000001100100100110;
assign LUT_4[22097] = 32'b11111111111111111010110000011110;
assign LUT_4[22098] = 32'b00000000000000000000111111001010;
assign LUT_4[22099] = 32'b11111111111111111010001011000010;
assign LUT_4[22100] = 32'b11111111111111111110100101000010;
assign LUT_4[22101] = 32'b11111111111111110111110000111010;
assign LUT_4[22102] = 32'b11111111111111111101111111100110;
assign LUT_4[22103] = 32'b11111111111111110111001011011110;
assign LUT_4[22104] = 32'b11111111111111111010110000111011;
assign LUT_4[22105] = 32'b11111111111111110011111100110011;
assign LUT_4[22106] = 32'b11111111111111111010001011011111;
assign LUT_4[22107] = 32'b11111111111111110011010111010111;
assign LUT_4[22108] = 32'b11111111111111110111110001010111;
assign LUT_4[22109] = 32'b11111111111111110000111101001111;
assign LUT_4[22110] = 32'b11111111111111110111001011111011;
assign LUT_4[22111] = 32'b11111111111111110000010111110011;
assign LUT_4[22112] = 32'b00000000000000000010001101111111;
assign LUT_4[22113] = 32'b11111111111111111011011001110111;
assign LUT_4[22114] = 32'b00000000000000000001101000100011;
assign LUT_4[22115] = 32'b11111111111111111010110100011011;
assign LUT_4[22116] = 32'b11111111111111111111001110011011;
assign LUT_4[22117] = 32'b11111111111111111000011010010011;
assign LUT_4[22118] = 32'b11111111111111111110101000111111;
assign LUT_4[22119] = 32'b11111111111111110111110100110111;
assign LUT_4[22120] = 32'b11111111111111111011011010010100;
assign LUT_4[22121] = 32'b11111111111111110100100110001100;
assign LUT_4[22122] = 32'b11111111111111111010110100111000;
assign LUT_4[22123] = 32'b11111111111111110100000000110000;
assign LUT_4[22124] = 32'b11111111111111111000011010110000;
assign LUT_4[22125] = 32'b11111111111111110001100110101000;
assign LUT_4[22126] = 32'b11111111111111110111110101010100;
assign LUT_4[22127] = 32'b11111111111111110001000001001100;
assign LUT_4[22128] = 32'b11111111111111111111111111101101;
assign LUT_4[22129] = 32'b11111111111111111001001011100101;
assign LUT_4[22130] = 32'b11111111111111111111011010010001;
assign LUT_4[22131] = 32'b11111111111111111000100110001001;
assign LUT_4[22132] = 32'b11111111111111111101000000001001;
assign LUT_4[22133] = 32'b11111111111111110110001100000001;
assign LUT_4[22134] = 32'b11111111111111111100011010101101;
assign LUT_4[22135] = 32'b11111111111111110101100110100101;
assign LUT_4[22136] = 32'b11111111111111111001001100000010;
assign LUT_4[22137] = 32'b11111111111111110010010111111010;
assign LUT_4[22138] = 32'b11111111111111111000100110100110;
assign LUT_4[22139] = 32'b11111111111111110001110010011110;
assign LUT_4[22140] = 32'b11111111111111110110001100011110;
assign LUT_4[22141] = 32'b11111111111111101111011000010110;
assign LUT_4[22142] = 32'b11111111111111110101100111000010;
assign LUT_4[22143] = 32'b11111111111111101110110010111010;
assign LUT_4[22144] = 32'b00000000000000000101000001101100;
assign LUT_4[22145] = 32'b11111111111111111110001101100100;
assign LUT_4[22146] = 32'b00000000000000000100011100010000;
assign LUT_4[22147] = 32'b11111111111111111101101000001000;
assign LUT_4[22148] = 32'b00000000000000000010000010001000;
assign LUT_4[22149] = 32'b11111111111111111011001110000000;
assign LUT_4[22150] = 32'b00000000000000000001011100101100;
assign LUT_4[22151] = 32'b11111111111111111010101000100100;
assign LUT_4[22152] = 32'b11111111111111111110001110000001;
assign LUT_4[22153] = 32'b11111111111111110111011001111001;
assign LUT_4[22154] = 32'b11111111111111111101101000100101;
assign LUT_4[22155] = 32'b11111111111111110110110100011101;
assign LUT_4[22156] = 32'b11111111111111111011001110011101;
assign LUT_4[22157] = 32'b11111111111111110100011010010101;
assign LUT_4[22158] = 32'b11111111111111111010101001000001;
assign LUT_4[22159] = 32'b11111111111111110011110100111001;
assign LUT_4[22160] = 32'b00000000000000000010110011011010;
assign LUT_4[22161] = 32'b11111111111111111011111111010010;
assign LUT_4[22162] = 32'b00000000000000000010001101111110;
assign LUT_4[22163] = 32'b11111111111111111011011001110110;
assign LUT_4[22164] = 32'b11111111111111111111110011110110;
assign LUT_4[22165] = 32'b11111111111111111000111111101110;
assign LUT_4[22166] = 32'b11111111111111111111001110011010;
assign LUT_4[22167] = 32'b11111111111111111000011010010010;
assign LUT_4[22168] = 32'b11111111111111111011111111101111;
assign LUT_4[22169] = 32'b11111111111111110101001011100111;
assign LUT_4[22170] = 32'b11111111111111111011011010010011;
assign LUT_4[22171] = 32'b11111111111111110100100110001011;
assign LUT_4[22172] = 32'b11111111111111111001000000001011;
assign LUT_4[22173] = 32'b11111111111111110010001100000011;
assign LUT_4[22174] = 32'b11111111111111111000011010101111;
assign LUT_4[22175] = 32'b11111111111111110001100110100111;
assign LUT_4[22176] = 32'b00000000000000000011011100110011;
assign LUT_4[22177] = 32'b11111111111111111100101000101011;
assign LUT_4[22178] = 32'b00000000000000000010110111010111;
assign LUT_4[22179] = 32'b11111111111111111100000011001111;
assign LUT_4[22180] = 32'b00000000000000000000011101001111;
assign LUT_4[22181] = 32'b11111111111111111001101001000111;
assign LUT_4[22182] = 32'b11111111111111111111110111110011;
assign LUT_4[22183] = 32'b11111111111111111001000011101011;
assign LUT_4[22184] = 32'b11111111111111111100101001001000;
assign LUT_4[22185] = 32'b11111111111111110101110101000000;
assign LUT_4[22186] = 32'b11111111111111111100000011101100;
assign LUT_4[22187] = 32'b11111111111111110101001111100100;
assign LUT_4[22188] = 32'b11111111111111111001101001100100;
assign LUT_4[22189] = 32'b11111111111111110010110101011100;
assign LUT_4[22190] = 32'b11111111111111111001000100001000;
assign LUT_4[22191] = 32'b11111111111111110010010000000000;
assign LUT_4[22192] = 32'b00000000000000000001001110100001;
assign LUT_4[22193] = 32'b11111111111111111010011010011001;
assign LUT_4[22194] = 32'b00000000000000000000101001000101;
assign LUT_4[22195] = 32'b11111111111111111001110100111101;
assign LUT_4[22196] = 32'b11111111111111111110001110111101;
assign LUT_4[22197] = 32'b11111111111111110111011010110101;
assign LUT_4[22198] = 32'b11111111111111111101101001100001;
assign LUT_4[22199] = 32'b11111111111111110110110101011001;
assign LUT_4[22200] = 32'b11111111111111111010011010110110;
assign LUT_4[22201] = 32'b11111111111111110011100110101110;
assign LUT_4[22202] = 32'b11111111111111111001110101011010;
assign LUT_4[22203] = 32'b11111111111111110011000001010010;
assign LUT_4[22204] = 32'b11111111111111110111011011010010;
assign LUT_4[22205] = 32'b11111111111111110000100111001010;
assign LUT_4[22206] = 32'b11111111111111110110110101110110;
assign LUT_4[22207] = 32'b11111111111111110000000001101110;
assign LUT_4[22208] = 32'b00000000000000000110011001000000;
assign LUT_4[22209] = 32'b11111111111111111111100100111000;
assign LUT_4[22210] = 32'b00000000000000000101110011100100;
assign LUT_4[22211] = 32'b11111111111111111110111111011100;
assign LUT_4[22212] = 32'b00000000000000000011011001011100;
assign LUT_4[22213] = 32'b11111111111111111100100101010100;
assign LUT_4[22214] = 32'b00000000000000000010110100000000;
assign LUT_4[22215] = 32'b11111111111111111011111111111000;
assign LUT_4[22216] = 32'b11111111111111111111100101010101;
assign LUT_4[22217] = 32'b11111111111111111000110001001101;
assign LUT_4[22218] = 32'b11111111111111111110111111111001;
assign LUT_4[22219] = 32'b11111111111111111000001011110001;
assign LUT_4[22220] = 32'b11111111111111111100100101110001;
assign LUT_4[22221] = 32'b11111111111111110101110001101001;
assign LUT_4[22222] = 32'b11111111111111111100000000010101;
assign LUT_4[22223] = 32'b11111111111111110101001100001101;
assign LUT_4[22224] = 32'b00000000000000000100001010101110;
assign LUT_4[22225] = 32'b11111111111111111101010110100110;
assign LUT_4[22226] = 32'b00000000000000000011100101010010;
assign LUT_4[22227] = 32'b11111111111111111100110001001010;
assign LUT_4[22228] = 32'b00000000000000000001001011001010;
assign LUT_4[22229] = 32'b11111111111111111010010111000010;
assign LUT_4[22230] = 32'b00000000000000000000100101101110;
assign LUT_4[22231] = 32'b11111111111111111001110001100110;
assign LUT_4[22232] = 32'b11111111111111111101010111000011;
assign LUT_4[22233] = 32'b11111111111111110110100010111011;
assign LUT_4[22234] = 32'b11111111111111111100110001100111;
assign LUT_4[22235] = 32'b11111111111111110101111101011111;
assign LUT_4[22236] = 32'b11111111111111111010010111011111;
assign LUT_4[22237] = 32'b11111111111111110011100011010111;
assign LUT_4[22238] = 32'b11111111111111111001110010000011;
assign LUT_4[22239] = 32'b11111111111111110010111101111011;
assign LUT_4[22240] = 32'b00000000000000000100110100000111;
assign LUT_4[22241] = 32'b11111111111111111101111111111111;
assign LUT_4[22242] = 32'b00000000000000000100001110101011;
assign LUT_4[22243] = 32'b11111111111111111101011010100011;
assign LUT_4[22244] = 32'b00000000000000000001110100100011;
assign LUT_4[22245] = 32'b11111111111111111011000000011011;
assign LUT_4[22246] = 32'b00000000000000000001001111000111;
assign LUT_4[22247] = 32'b11111111111111111010011010111111;
assign LUT_4[22248] = 32'b11111111111111111110000000011100;
assign LUT_4[22249] = 32'b11111111111111110111001100010100;
assign LUT_4[22250] = 32'b11111111111111111101011011000000;
assign LUT_4[22251] = 32'b11111111111111110110100110111000;
assign LUT_4[22252] = 32'b11111111111111111011000000111000;
assign LUT_4[22253] = 32'b11111111111111110100001100110000;
assign LUT_4[22254] = 32'b11111111111111111010011011011100;
assign LUT_4[22255] = 32'b11111111111111110011100111010100;
assign LUT_4[22256] = 32'b00000000000000000010100101110101;
assign LUT_4[22257] = 32'b11111111111111111011110001101101;
assign LUT_4[22258] = 32'b00000000000000000010000000011001;
assign LUT_4[22259] = 32'b11111111111111111011001100010001;
assign LUT_4[22260] = 32'b11111111111111111111100110010001;
assign LUT_4[22261] = 32'b11111111111111111000110010001001;
assign LUT_4[22262] = 32'b11111111111111111111000000110101;
assign LUT_4[22263] = 32'b11111111111111111000001100101101;
assign LUT_4[22264] = 32'b11111111111111111011110010001010;
assign LUT_4[22265] = 32'b11111111111111110100111110000010;
assign LUT_4[22266] = 32'b11111111111111111011001100101110;
assign LUT_4[22267] = 32'b11111111111111110100011000100110;
assign LUT_4[22268] = 32'b11111111111111111000110010100110;
assign LUT_4[22269] = 32'b11111111111111110001111110011110;
assign LUT_4[22270] = 32'b11111111111111111000001101001010;
assign LUT_4[22271] = 32'b11111111111111110001011001000010;
assign LUT_4[22272] = 32'b00000000000000000111010111000111;
assign LUT_4[22273] = 32'b00000000000000000000100010111111;
assign LUT_4[22274] = 32'b00000000000000000110110001101011;
assign LUT_4[22275] = 32'b11111111111111111111111101100011;
assign LUT_4[22276] = 32'b00000000000000000100010111100011;
assign LUT_4[22277] = 32'b11111111111111111101100011011011;
assign LUT_4[22278] = 32'b00000000000000000011110010000111;
assign LUT_4[22279] = 32'b11111111111111111100111101111111;
assign LUT_4[22280] = 32'b00000000000000000000100011011100;
assign LUT_4[22281] = 32'b11111111111111111001101111010100;
assign LUT_4[22282] = 32'b11111111111111111111111110000000;
assign LUT_4[22283] = 32'b11111111111111111001001001111000;
assign LUT_4[22284] = 32'b11111111111111111101100011111000;
assign LUT_4[22285] = 32'b11111111111111110110101111110000;
assign LUT_4[22286] = 32'b11111111111111111100111110011100;
assign LUT_4[22287] = 32'b11111111111111110110001010010100;
assign LUT_4[22288] = 32'b00000000000000000101001000110101;
assign LUT_4[22289] = 32'b11111111111111111110010100101101;
assign LUT_4[22290] = 32'b00000000000000000100100011011001;
assign LUT_4[22291] = 32'b11111111111111111101101111010001;
assign LUT_4[22292] = 32'b00000000000000000010001001010001;
assign LUT_4[22293] = 32'b11111111111111111011010101001001;
assign LUT_4[22294] = 32'b00000000000000000001100011110101;
assign LUT_4[22295] = 32'b11111111111111111010101111101101;
assign LUT_4[22296] = 32'b11111111111111111110010101001010;
assign LUT_4[22297] = 32'b11111111111111110111100001000010;
assign LUT_4[22298] = 32'b11111111111111111101101111101110;
assign LUT_4[22299] = 32'b11111111111111110110111011100110;
assign LUT_4[22300] = 32'b11111111111111111011010101100110;
assign LUT_4[22301] = 32'b11111111111111110100100001011110;
assign LUT_4[22302] = 32'b11111111111111111010110000001010;
assign LUT_4[22303] = 32'b11111111111111110011111100000010;
assign LUT_4[22304] = 32'b00000000000000000101110010001110;
assign LUT_4[22305] = 32'b11111111111111111110111110000110;
assign LUT_4[22306] = 32'b00000000000000000101001100110010;
assign LUT_4[22307] = 32'b11111111111111111110011000101010;
assign LUT_4[22308] = 32'b00000000000000000010110010101010;
assign LUT_4[22309] = 32'b11111111111111111011111110100010;
assign LUT_4[22310] = 32'b00000000000000000010001101001110;
assign LUT_4[22311] = 32'b11111111111111111011011001000110;
assign LUT_4[22312] = 32'b11111111111111111110111110100011;
assign LUT_4[22313] = 32'b11111111111111111000001010011011;
assign LUT_4[22314] = 32'b11111111111111111110011001000111;
assign LUT_4[22315] = 32'b11111111111111110111100100111111;
assign LUT_4[22316] = 32'b11111111111111111011111110111111;
assign LUT_4[22317] = 32'b11111111111111110101001010110111;
assign LUT_4[22318] = 32'b11111111111111111011011001100011;
assign LUT_4[22319] = 32'b11111111111111110100100101011011;
assign LUT_4[22320] = 32'b00000000000000000011100011111100;
assign LUT_4[22321] = 32'b11111111111111111100101111110100;
assign LUT_4[22322] = 32'b00000000000000000010111110100000;
assign LUT_4[22323] = 32'b11111111111111111100001010011000;
assign LUT_4[22324] = 32'b00000000000000000000100100011000;
assign LUT_4[22325] = 32'b11111111111111111001110000010000;
assign LUT_4[22326] = 32'b11111111111111111111111110111100;
assign LUT_4[22327] = 32'b11111111111111111001001010110100;
assign LUT_4[22328] = 32'b11111111111111111100110000010001;
assign LUT_4[22329] = 32'b11111111111111110101111100001001;
assign LUT_4[22330] = 32'b11111111111111111100001010110101;
assign LUT_4[22331] = 32'b11111111111111110101010110101101;
assign LUT_4[22332] = 32'b11111111111111111001110000101101;
assign LUT_4[22333] = 32'b11111111111111110010111100100101;
assign LUT_4[22334] = 32'b11111111111111111001001011010001;
assign LUT_4[22335] = 32'b11111111111111110010010111001001;
assign LUT_4[22336] = 32'b00000000000000001000101110011011;
assign LUT_4[22337] = 32'b00000000000000000001111010010011;
assign LUT_4[22338] = 32'b00000000000000001000001000111111;
assign LUT_4[22339] = 32'b00000000000000000001010100110111;
assign LUT_4[22340] = 32'b00000000000000000101101110110111;
assign LUT_4[22341] = 32'b11111111111111111110111010101111;
assign LUT_4[22342] = 32'b00000000000000000101001001011011;
assign LUT_4[22343] = 32'b11111111111111111110010101010011;
assign LUT_4[22344] = 32'b00000000000000000001111010110000;
assign LUT_4[22345] = 32'b11111111111111111011000110101000;
assign LUT_4[22346] = 32'b00000000000000000001010101010100;
assign LUT_4[22347] = 32'b11111111111111111010100001001100;
assign LUT_4[22348] = 32'b11111111111111111110111011001100;
assign LUT_4[22349] = 32'b11111111111111111000000111000100;
assign LUT_4[22350] = 32'b11111111111111111110010101110000;
assign LUT_4[22351] = 32'b11111111111111110111100001101000;
assign LUT_4[22352] = 32'b00000000000000000110100000001001;
assign LUT_4[22353] = 32'b11111111111111111111101100000001;
assign LUT_4[22354] = 32'b00000000000000000101111010101101;
assign LUT_4[22355] = 32'b11111111111111111111000110100101;
assign LUT_4[22356] = 32'b00000000000000000011100000100101;
assign LUT_4[22357] = 32'b11111111111111111100101100011101;
assign LUT_4[22358] = 32'b00000000000000000010111011001001;
assign LUT_4[22359] = 32'b11111111111111111100000111000001;
assign LUT_4[22360] = 32'b11111111111111111111101100011110;
assign LUT_4[22361] = 32'b11111111111111111000111000010110;
assign LUT_4[22362] = 32'b11111111111111111111000111000010;
assign LUT_4[22363] = 32'b11111111111111111000010010111010;
assign LUT_4[22364] = 32'b11111111111111111100101100111010;
assign LUT_4[22365] = 32'b11111111111111110101111000110010;
assign LUT_4[22366] = 32'b11111111111111111100000111011110;
assign LUT_4[22367] = 32'b11111111111111110101010011010110;
assign LUT_4[22368] = 32'b00000000000000000111001001100010;
assign LUT_4[22369] = 32'b00000000000000000000010101011010;
assign LUT_4[22370] = 32'b00000000000000000110100100000110;
assign LUT_4[22371] = 32'b11111111111111111111101111111110;
assign LUT_4[22372] = 32'b00000000000000000100001001111110;
assign LUT_4[22373] = 32'b11111111111111111101010101110110;
assign LUT_4[22374] = 32'b00000000000000000011100100100010;
assign LUT_4[22375] = 32'b11111111111111111100110000011010;
assign LUT_4[22376] = 32'b00000000000000000000010101110111;
assign LUT_4[22377] = 32'b11111111111111111001100001101111;
assign LUT_4[22378] = 32'b11111111111111111111110000011011;
assign LUT_4[22379] = 32'b11111111111111111000111100010011;
assign LUT_4[22380] = 32'b11111111111111111101010110010011;
assign LUT_4[22381] = 32'b11111111111111110110100010001011;
assign LUT_4[22382] = 32'b11111111111111111100110000110111;
assign LUT_4[22383] = 32'b11111111111111110101111100101111;
assign LUT_4[22384] = 32'b00000000000000000100111011010000;
assign LUT_4[22385] = 32'b11111111111111111110000111001000;
assign LUT_4[22386] = 32'b00000000000000000100010101110100;
assign LUT_4[22387] = 32'b11111111111111111101100001101100;
assign LUT_4[22388] = 32'b00000000000000000001111011101100;
assign LUT_4[22389] = 32'b11111111111111111011000111100100;
assign LUT_4[22390] = 32'b00000000000000000001010110010000;
assign LUT_4[22391] = 32'b11111111111111111010100010001000;
assign LUT_4[22392] = 32'b11111111111111111110000111100101;
assign LUT_4[22393] = 32'b11111111111111110111010011011101;
assign LUT_4[22394] = 32'b11111111111111111101100010001001;
assign LUT_4[22395] = 32'b11111111111111110110101110000001;
assign LUT_4[22396] = 32'b11111111111111111011001000000001;
assign LUT_4[22397] = 32'b11111111111111110100010011111001;
assign LUT_4[22398] = 32'b11111111111111111010100010100101;
assign LUT_4[22399] = 32'b11111111111111110011101110011101;
assign LUT_4[22400] = 32'b00000000000000001001111101001111;
assign LUT_4[22401] = 32'b00000000000000000011001001000111;
assign LUT_4[22402] = 32'b00000000000000001001010111110011;
assign LUT_4[22403] = 32'b00000000000000000010100011101011;
assign LUT_4[22404] = 32'b00000000000000000110111101101011;
assign LUT_4[22405] = 32'b00000000000000000000001001100011;
assign LUT_4[22406] = 32'b00000000000000000110011000001111;
assign LUT_4[22407] = 32'b11111111111111111111100100000111;
assign LUT_4[22408] = 32'b00000000000000000011001001100100;
assign LUT_4[22409] = 32'b11111111111111111100010101011100;
assign LUT_4[22410] = 32'b00000000000000000010100100001000;
assign LUT_4[22411] = 32'b11111111111111111011110000000000;
assign LUT_4[22412] = 32'b00000000000000000000001010000000;
assign LUT_4[22413] = 32'b11111111111111111001010101111000;
assign LUT_4[22414] = 32'b11111111111111111111100100100100;
assign LUT_4[22415] = 32'b11111111111111111000110000011100;
assign LUT_4[22416] = 32'b00000000000000000111101110111101;
assign LUT_4[22417] = 32'b00000000000000000000111010110101;
assign LUT_4[22418] = 32'b00000000000000000111001001100001;
assign LUT_4[22419] = 32'b00000000000000000000010101011001;
assign LUT_4[22420] = 32'b00000000000000000100101111011001;
assign LUT_4[22421] = 32'b11111111111111111101111011010001;
assign LUT_4[22422] = 32'b00000000000000000100001001111101;
assign LUT_4[22423] = 32'b11111111111111111101010101110101;
assign LUT_4[22424] = 32'b00000000000000000000111011010010;
assign LUT_4[22425] = 32'b11111111111111111010000111001010;
assign LUT_4[22426] = 32'b00000000000000000000010101110110;
assign LUT_4[22427] = 32'b11111111111111111001100001101110;
assign LUT_4[22428] = 32'b11111111111111111101111011101110;
assign LUT_4[22429] = 32'b11111111111111110111000111100110;
assign LUT_4[22430] = 32'b11111111111111111101010110010010;
assign LUT_4[22431] = 32'b11111111111111110110100010001010;
assign LUT_4[22432] = 32'b00000000000000001000011000010110;
assign LUT_4[22433] = 32'b00000000000000000001100100001110;
assign LUT_4[22434] = 32'b00000000000000000111110010111010;
assign LUT_4[22435] = 32'b00000000000000000000111110110010;
assign LUT_4[22436] = 32'b00000000000000000101011000110010;
assign LUT_4[22437] = 32'b11111111111111111110100100101010;
assign LUT_4[22438] = 32'b00000000000000000100110011010110;
assign LUT_4[22439] = 32'b11111111111111111101111111001110;
assign LUT_4[22440] = 32'b00000000000000000001100100101011;
assign LUT_4[22441] = 32'b11111111111111111010110000100011;
assign LUT_4[22442] = 32'b00000000000000000000111111001111;
assign LUT_4[22443] = 32'b11111111111111111010001011000111;
assign LUT_4[22444] = 32'b11111111111111111110100101000111;
assign LUT_4[22445] = 32'b11111111111111110111110000111111;
assign LUT_4[22446] = 32'b11111111111111111101111111101011;
assign LUT_4[22447] = 32'b11111111111111110111001011100011;
assign LUT_4[22448] = 32'b00000000000000000110001010000100;
assign LUT_4[22449] = 32'b11111111111111111111010101111100;
assign LUT_4[22450] = 32'b00000000000000000101100100101000;
assign LUT_4[22451] = 32'b11111111111111111110110000100000;
assign LUT_4[22452] = 32'b00000000000000000011001010100000;
assign LUT_4[22453] = 32'b11111111111111111100010110011000;
assign LUT_4[22454] = 32'b00000000000000000010100101000100;
assign LUT_4[22455] = 32'b11111111111111111011110000111100;
assign LUT_4[22456] = 32'b11111111111111111111010110011001;
assign LUT_4[22457] = 32'b11111111111111111000100010010001;
assign LUT_4[22458] = 32'b11111111111111111110110000111101;
assign LUT_4[22459] = 32'b11111111111111110111111100110101;
assign LUT_4[22460] = 32'b11111111111111111100010110110101;
assign LUT_4[22461] = 32'b11111111111111110101100010101101;
assign LUT_4[22462] = 32'b11111111111111111011110001011001;
assign LUT_4[22463] = 32'b11111111111111110100111101010001;
assign LUT_4[22464] = 32'b00000000000000001011010100100011;
assign LUT_4[22465] = 32'b00000000000000000100100000011011;
assign LUT_4[22466] = 32'b00000000000000001010101111000111;
assign LUT_4[22467] = 32'b00000000000000000011111010111111;
assign LUT_4[22468] = 32'b00000000000000001000010100111111;
assign LUT_4[22469] = 32'b00000000000000000001100000110111;
assign LUT_4[22470] = 32'b00000000000000000111101111100011;
assign LUT_4[22471] = 32'b00000000000000000000111011011011;
assign LUT_4[22472] = 32'b00000000000000000100100000111000;
assign LUT_4[22473] = 32'b11111111111111111101101100110000;
assign LUT_4[22474] = 32'b00000000000000000011111011011100;
assign LUT_4[22475] = 32'b11111111111111111101000111010100;
assign LUT_4[22476] = 32'b00000000000000000001100001010100;
assign LUT_4[22477] = 32'b11111111111111111010101101001100;
assign LUT_4[22478] = 32'b00000000000000000000111011111000;
assign LUT_4[22479] = 32'b11111111111111111010000111110000;
assign LUT_4[22480] = 32'b00000000000000001001000110010001;
assign LUT_4[22481] = 32'b00000000000000000010010010001001;
assign LUT_4[22482] = 32'b00000000000000001000100000110101;
assign LUT_4[22483] = 32'b00000000000000000001101100101101;
assign LUT_4[22484] = 32'b00000000000000000110000110101101;
assign LUT_4[22485] = 32'b11111111111111111111010010100101;
assign LUT_4[22486] = 32'b00000000000000000101100001010001;
assign LUT_4[22487] = 32'b11111111111111111110101101001001;
assign LUT_4[22488] = 32'b00000000000000000010010010100110;
assign LUT_4[22489] = 32'b11111111111111111011011110011110;
assign LUT_4[22490] = 32'b00000000000000000001101101001010;
assign LUT_4[22491] = 32'b11111111111111111010111001000010;
assign LUT_4[22492] = 32'b11111111111111111111010011000010;
assign LUT_4[22493] = 32'b11111111111111111000011110111010;
assign LUT_4[22494] = 32'b11111111111111111110101101100110;
assign LUT_4[22495] = 32'b11111111111111110111111001011110;
assign LUT_4[22496] = 32'b00000000000000001001101111101010;
assign LUT_4[22497] = 32'b00000000000000000010111011100010;
assign LUT_4[22498] = 32'b00000000000000001001001010001110;
assign LUT_4[22499] = 32'b00000000000000000010010110000110;
assign LUT_4[22500] = 32'b00000000000000000110110000000110;
assign LUT_4[22501] = 32'b11111111111111111111111011111110;
assign LUT_4[22502] = 32'b00000000000000000110001010101010;
assign LUT_4[22503] = 32'b11111111111111111111010110100010;
assign LUT_4[22504] = 32'b00000000000000000010111011111111;
assign LUT_4[22505] = 32'b11111111111111111100000111110111;
assign LUT_4[22506] = 32'b00000000000000000010010110100011;
assign LUT_4[22507] = 32'b11111111111111111011100010011011;
assign LUT_4[22508] = 32'b11111111111111111111111100011011;
assign LUT_4[22509] = 32'b11111111111111111001001000010011;
assign LUT_4[22510] = 32'b11111111111111111111010110111111;
assign LUT_4[22511] = 32'b11111111111111111000100010110111;
assign LUT_4[22512] = 32'b00000000000000000111100001011000;
assign LUT_4[22513] = 32'b00000000000000000000101101010000;
assign LUT_4[22514] = 32'b00000000000000000110111011111100;
assign LUT_4[22515] = 32'b00000000000000000000000111110100;
assign LUT_4[22516] = 32'b00000000000000000100100001110100;
assign LUT_4[22517] = 32'b11111111111111111101101101101100;
assign LUT_4[22518] = 32'b00000000000000000011111100011000;
assign LUT_4[22519] = 32'b11111111111111111101001000010000;
assign LUT_4[22520] = 32'b00000000000000000000101101101101;
assign LUT_4[22521] = 32'b11111111111111111001111001100101;
assign LUT_4[22522] = 32'b00000000000000000000001000010001;
assign LUT_4[22523] = 32'b11111111111111111001010100001001;
assign LUT_4[22524] = 32'b11111111111111111101101110001001;
assign LUT_4[22525] = 32'b11111111111111110110111010000001;
assign LUT_4[22526] = 32'b11111111111111111101001000101101;
assign LUT_4[22527] = 32'b11111111111111110110010100100101;
assign LUT_4[22528] = 32'b11111111111111111101001100000111;
assign LUT_4[22529] = 32'b11111111111111110110010111111111;
assign LUT_4[22530] = 32'b11111111111111111100100110101011;
assign LUT_4[22531] = 32'b11111111111111110101110010100011;
assign LUT_4[22532] = 32'b11111111111111111010001100100011;
assign LUT_4[22533] = 32'b11111111111111110011011000011011;
assign LUT_4[22534] = 32'b11111111111111111001100111000111;
assign LUT_4[22535] = 32'b11111111111111110010110010111111;
assign LUT_4[22536] = 32'b11111111111111110110011000011100;
assign LUT_4[22537] = 32'b11111111111111101111100100010100;
assign LUT_4[22538] = 32'b11111111111111110101110011000000;
assign LUT_4[22539] = 32'b11111111111111101110111110111000;
assign LUT_4[22540] = 32'b11111111111111110011011000111000;
assign LUT_4[22541] = 32'b11111111111111101100100100110000;
assign LUT_4[22542] = 32'b11111111111111110010110011011100;
assign LUT_4[22543] = 32'b11111111111111101011111111010100;
assign LUT_4[22544] = 32'b11111111111111111010111101110101;
assign LUT_4[22545] = 32'b11111111111111110100001001101101;
assign LUT_4[22546] = 32'b11111111111111111010011000011001;
assign LUT_4[22547] = 32'b11111111111111110011100100010001;
assign LUT_4[22548] = 32'b11111111111111110111111110010001;
assign LUT_4[22549] = 32'b11111111111111110001001010001001;
assign LUT_4[22550] = 32'b11111111111111110111011000110101;
assign LUT_4[22551] = 32'b11111111111111110000100100101101;
assign LUT_4[22552] = 32'b11111111111111110100001010001010;
assign LUT_4[22553] = 32'b11111111111111101101010110000010;
assign LUT_4[22554] = 32'b11111111111111110011100100101110;
assign LUT_4[22555] = 32'b11111111111111101100110000100110;
assign LUT_4[22556] = 32'b11111111111111110001001010100110;
assign LUT_4[22557] = 32'b11111111111111101010010110011110;
assign LUT_4[22558] = 32'b11111111111111110000100101001010;
assign LUT_4[22559] = 32'b11111111111111101001110001000010;
assign LUT_4[22560] = 32'b11111111111111111011100111001110;
assign LUT_4[22561] = 32'b11111111111111110100110011000110;
assign LUT_4[22562] = 32'b11111111111111111011000001110010;
assign LUT_4[22563] = 32'b11111111111111110100001101101010;
assign LUT_4[22564] = 32'b11111111111111111000100111101010;
assign LUT_4[22565] = 32'b11111111111111110001110011100010;
assign LUT_4[22566] = 32'b11111111111111111000000010001110;
assign LUT_4[22567] = 32'b11111111111111110001001110000110;
assign LUT_4[22568] = 32'b11111111111111110100110011100011;
assign LUT_4[22569] = 32'b11111111111111101101111111011011;
assign LUT_4[22570] = 32'b11111111111111110100001110000111;
assign LUT_4[22571] = 32'b11111111111111101101011001111111;
assign LUT_4[22572] = 32'b11111111111111110001110011111111;
assign LUT_4[22573] = 32'b11111111111111101010111111110111;
assign LUT_4[22574] = 32'b11111111111111110001001110100011;
assign LUT_4[22575] = 32'b11111111111111101010011010011011;
assign LUT_4[22576] = 32'b11111111111111111001011000111100;
assign LUT_4[22577] = 32'b11111111111111110010100100110100;
assign LUT_4[22578] = 32'b11111111111111111000110011100000;
assign LUT_4[22579] = 32'b11111111111111110001111111011000;
assign LUT_4[22580] = 32'b11111111111111110110011001011000;
assign LUT_4[22581] = 32'b11111111111111101111100101010000;
assign LUT_4[22582] = 32'b11111111111111110101110011111100;
assign LUT_4[22583] = 32'b11111111111111101110111111110100;
assign LUT_4[22584] = 32'b11111111111111110010100101010001;
assign LUT_4[22585] = 32'b11111111111111101011110001001001;
assign LUT_4[22586] = 32'b11111111111111110001111111110101;
assign LUT_4[22587] = 32'b11111111111111101011001011101101;
assign LUT_4[22588] = 32'b11111111111111101111100101101101;
assign LUT_4[22589] = 32'b11111111111111101000110001100101;
assign LUT_4[22590] = 32'b11111111111111101111000000010001;
assign LUT_4[22591] = 32'b11111111111111101000001100001001;
assign LUT_4[22592] = 32'b11111111111111111110100011011011;
assign LUT_4[22593] = 32'b11111111111111110111101111010011;
assign LUT_4[22594] = 32'b11111111111111111101111101111111;
assign LUT_4[22595] = 32'b11111111111111110111001001110111;
assign LUT_4[22596] = 32'b11111111111111111011100011110111;
assign LUT_4[22597] = 32'b11111111111111110100101111101111;
assign LUT_4[22598] = 32'b11111111111111111010111110011011;
assign LUT_4[22599] = 32'b11111111111111110100001010010011;
assign LUT_4[22600] = 32'b11111111111111110111101111110000;
assign LUT_4[22601] = 32'b11111111111111110000111011101000;
assign LUT_4[22602] = 32'b11111111111111110111001010010100;
assign LUT_4[22603] = 32'b11111111111111110000010110001100;
assign LUT_4[22604] = 32'b11111111111111110100110000001100;
assign LUT_4[22605] = 32'b11111111111111101101111100000100;
assign LUT_4[22606] = 32'b11111111111111110100001010110000;
assign LUT_4[22607] = 32'b11111111111111101101010110101000;
assign LUT_4[22608] = 32'b11111111111111111100010101001001;
assign LUT_4[22609] = 32'b11111111111111110101100001000001;
assign LUT_4[22610] = 32'b11111111111111111011101111101101;
assign LUT_4[22611] = 32'b11111111111111110100111011100101;
assign LUT_4[22612] = 32'b11111111111111111001010101100101;
assign LUT_4[22613] = 32'b11111111111111110010100001011101;
assign LUT_4[22614] = 32'b11111111111111111000110000001001;
assign LUT_4[22615] = 32'b11111111111111110001111100000001;
assign LUT_4[22616] = 32'b11111111111111110101100001011110;
assign LUT_4[22617] = 32'b11111111111111101110101101010110;
assign LUT_4[22618] = 32'b11111111111111110100111100000010;
assign LUT_4[22619] = 32'b11111111111111101110000111111010;
assign LUT_4[22620] = 32'b11111111111111110010100001111010;
assign LUT_4[22621] = 32'b11111111111111101011101101110010;
assign LUT_4[22622] = 32'b11111111111111110001111100011110;
assign LUT_4[22623] = 32'b11111111111111101011001000010110;
assign LUT_4[22624] = 32'b11111111111111111100111110100010;
assign LUT_4[22625] = 32'b11111111111111110110001010011010;
assign LUT_4[22626] = 32'b11111111111111111100011001000110;
assign LUT_4[22627] = 32'b11111111111111110101100100111110;
assign LUT_4[22628] = 32'b11111111111111111001111110111110;
assign LUT_4[22629] = 32'b11111111111111110011001010110110;
assign LUT_4[22630] = 32'b11111111111111111001011001100010;
assign LUT_4[22631] = 32'b11111111111111110010100101011010;
assign LUT_4[22632] = 32'b11111111111111110110001010110111;
assign LUT_4[22633] = 32'b11111111111111101111010110101111;
assign LUT_4[22634] = 32'b11111111111111110101100101011011;
assign LUT_4[22635] = 32'b11111111111111101110110001010011;
assign LUT_4[22636] = 32'b11111111111111110011001011010011;
assign LUT_4[22637] = 32'b11111111111111101100010111001011;
assign LUT_4[22638] = 32'b11111111111111110010100101110111;
assign LUT_4[22639] = 32'b11111111111111101011110001101111;
assign LUT_4[22640] = 32'b11111111111111111010110000010000;
assign LUT_4[22641] = 32'b11111111111111110011111100001000;
assign LUT_4[22642] = 32'b11111111111111111010001010110100;
assign LUT_4[22643] = 32'b11111111111111110011010110101100;
assign LUT_4[22644] = 32'b11111111111111110111110000101100;
assign LUT_4[22645] = 32'b11111111111111110000111100100100;
assign LUT_4[22646] = 32'b11111111111111110111001011010000;
assign LUT_4[22647] = 32'b11111111111111110000010111001000;
assign LUT_4[22648] = 32'b11111111111111110011111100100101;
assign LUT_4[22649] = 32'b11111111111111101101001000011101;
assign LUT_4[22650] = 32'b11111111111111110011010111001001;
assign LUT_4[22651] = 32'b11111111111111101100100011000001;
assign LUT_4[22652] = 32'b11111111111111110000111101000001;
assign LUT_4[22653] = 32'b11111111111111101010001000111001;
assign LUT_4[22654] = 32'b11111111111111110000010111100101;
assign LUT_4[22655] = 32'b11111111111111101001100011011101;
assign LUT_4[22656] = 32'b11111111111111111111110010001111;
assign LUT_4[22657] = 32'b11111111111111111000111110000111;
assign LUT_4[22658] = 32'b11111111111111111111001100110011;
assign LUT_4[22659] = 32'b11111111111111111000011000101011;
assign LUT_4[22660] = 32'b11111111111111111100110010101011;
assign LUT_4[22661] = 32'b11111111111111110101111110100011;
assign LUT_4[22662] = 32'b11111111111111111100001101001111;
assign LUT_4[22663] = 32'b11111111111111110101011001000111;
assign LUT_4[22664] = 32'b11111111111111111000111110100100;
assign LUT_4[22665] = 32'b11111111111111110010001010011100;
assign LUT_4[22666] = 32'b11111111111111111000011001001000;
assign LUT_4[22667] = 32'b11111111111111110001100101000000;
assign LUT_4[22668] = 32'b11111111111111110101111111000000;
assign LUT_4[22669] = 32'b11111111111111101111001010111000;
assign LUT_4[22670] = 32'b11111111111111110101011001100100;
assign LUT_4[22671] = 32'b11111111111111101110100101011100;
assign LUT_4[22672] = 32'b11111111111111111101100011111101;
assign LUT_4[22673] = 32'b11111111111111110110101111110101;
assign LUT_4[22674] = 32'b11111111111111111100111110100001;
assign LUT_4[22675] = 32'b11111111111111110110001010011001;
assign LUT_4[22676] = 32'b11111111111111111010100100011001;
assign LUT_4[22677] = 32'b11111111111111110011110000010001;
assign LUT_4[22678] = 32'b11111111111111111001111110111101;
assign LUT_4[22679] = 32'b11111111111111110011001010110101;
assign LUT_4[22680] = 32'b11111111111111110110110000010010;
assign LUT_4[22681] = 32'b11111111111111101111111100001010;
assign LUT_4[22682] = 32'b11111111111111110110001010110110;
assign LUT_4[22683] = 32'b11111111111111101111010110101110;
assign LUT_4[22684] = 32'b11111111111111110011110000101110;
assign LUT_4[22685] = 32'b11111111111111101100111100100110;
assign LUT_4[22686] = 32'b11111111111111110011001011010010;
assign LUT_4[22687] = 32'b11111111111111101100010111001010;
assign LUT_4[22688] = 32'b11111111111111111110001101010110;
assign LUT_4[22689] = 32'b11111111111111110111011001001110;
assign LUT_4[22690] = 32'b11111111111111111101100111111010;
assign LUT_4[22691] = 32'b11111111111111110110110011110010;
assign LUT_4[22692] = 32'b11111111111111111011001101110010;
assign LUT_4[22693] = 32'b11111111111111110100011001101010;
assign LUT_4[22694] = 32'b11111111111111111010101000010110;
assign LUT_4[22695] = 32'b11111111111111110011110100001110;
assign LUT_4[22696] = 32'b11111111111111110111011001101011;
assign LUT_4[22697] = 32'b11111111111111110000100101100011;
assign LUT_4[22698] = 32'b11111111111111110110110100001111;
assign LUT_4[22699] = 32'b11111111111111110000000000000111;
assign LUT_4[22700] = 32'b11111111111111110100011010000111;
assign LUT_4[22701] = 32'b11111111111111101101100101111111;
assign LUT_4[22702] = 32'b11111111111111110011110100101011;
assign LUT_4[22703] = 32'b11111111111111101101000000100011;
assign LUT_4[22704] = 32'b11111111111111111011111111000100;
assign LUT_4[22705] = 32'b11111111111111110101001010111100;
assign LUT_4[22706] = 32'b11111111111111111011011001101000;
assign LUT_4[22707] = 32'b11111111111111110100100101100000;
assign LUT_4[22708] = 32'b11111111111111111000111111100000;
assign LUT_4[22709] = 32'b11111111111111110010001011011000;
assign LUT_4[22710] = 32'b11111111111111111000011010000100;
assign LUT_4[22711] = 32'b11111111111111110001100101111100;
assign LUT_4[22712] = 32'b11111111111111110101001011011001;
assign LUT_4[22713] = 32'b11111111111111101110010111010001;
assign LUT_4[22714] = 32'b11111111111111110100100101111101;
assign LUT_4[22715] = 32'b11111111111111101101110001110101;
assign LUT_4[22716] = 32'b11111111111111110010001011110101;
assign LUT_4[22717] = 32'b11111111111111101011010111101101;
assign LUT_4[22718] = 32'b11111111111111110001100110011001;
assign LUT_4[22719] = 32'b11111111111111101010110010010001;
assign LUT_4[22720] = 32'b00000000000000000001001001100011;
assign LUT_4[22721] = 32'b11111111111111111010010101011011;
assign LUT_4[22722] = 32'b00000000000000000000100100000111;
assign LUT_4[22723] = 32'b11111111111111111001101111111111;
assign LUT_4[22724] = 32'b11111111111111111110001001111111;
assign LUT_4[22725] = 32'b11111111111111110111010101110111;
assign LUT_4[22726] = 32'b11111111111111111101100100100011;
assign LUT_4[22727] = 32'b11111111111111110110110000011011;
assign LUT_4[22728] = 32'b11111111111111111010010101111000;
assign LUT_4[22729] = 32'b11111111111111110011100001110000;
assign LUT_4[22730] = 32'b11111111111111111001110000011100;
assign LUT_4[22731] = 32'b11111111111111110010111100010100;
assign LUT_4[22732] = 32'b11111111111111110111010110010100;
assign LUT_4[22733] = 32'b11111111111111110000100010001100;
assign LUT_4[22734] = 32'b11111111111111110110110000111000;
assign LUT_4[22735] = 32'b11111111111111101111111100110000;
assign LUT_4[22736] = 32'b11111111111111111110111011010001;
assign LUT_4[22737] = 32'b11111111111111111000000111001001;
assign LUT_4[22738] = 32'b11111111111111111110010101110101;
assign LUT_4[22739] = 32'b11111111111111110111100001101101;
assign LUT_4[22740] = 32'b11111111111111111011111011101101;
assign LUT_4[22741] = 32'b11111111111111110101000111100101;
assign LUT_4[22742] = 32'b11111111111111111011010110010001;
assign LUT_4[22743] = 32'b11111111111111110100100010001001;
assign LUT_4[22744] = 32'b11111111111111111000000111100110;
assign LUT_4[22745] = 32'b11111111111111110001010011011110;
assign LUT_4[22746] = 32'b11111111111111110111100010001010;
assign LUT_4[22747] = 32'b11111111111111110000101110000010;
assign LUT_4[22748] = 32'b11111111111111110101001000000010;
assign LUT_4[22749] = 32'b11111111111111101110010011111010;
assign LUT_4[22750] = 32'b11111111111111110100100010100110;
assign LUT_4[22751] = 32'b11111111111111101101101110011110;
assign LUT_4[22752] = 32'b11111111111111111111100100101010;
assign LUT_4[22753] = 32'b11111111111111111000110000100010;
assign LUT_4[22754] = 32'b11111111111111111110111111001110;
assign LUT_4[22755] = 32'b11111111111111111000001011000110;
assign LUT_4[22756] = 32'b11111111111111111100100101000110;
assign LUT_4[22757] = 32'b11111111111111110101110000111110;
assign LUT_4[22758] = 32'b11111111111111111011111111101010;
assign LUT_4[22759] = 32'b11111111111111110101001011100010;
assign LUT_4[22760] = 32'b11111111111111111000110000111111;
assign LUT_4[22761] = 32'b11111111111111110001111100110111;
assign LUT_4[22762] = 32'b11111111111111111000001011100011;
assign LUT_4[22763] = 32'b11111111111111110001010111011011;
assign LUT_4[22764] = 32'b11111111111111110101110001011011;
assign LUT_4[22765] = 32'b11111111111111101110111101010011;
assign LUT_4[22766] = 32'b11111111111111110101001011111111;
assign LUT_4[22767] = 32'b11111111111111101110010111110111;
assign LUT_4[22768] = 32'b11111111111111111101010110011000;
assign LUT_4[22769] = 32'b11111111111111110110100010010000;
assign LUT_4[22770] = 32'b11111111111111111100110000111100;
assign LUT_4[22771] = 32'b11111111111111110101111100110100;
assign LUT_4[22772] = 32'b11111111111111111010010110110100;
assign LUT_4[22773] = 32'b11111111111111110011100010101100;
assign LUT_4[22774] = 32'b11111111111111111001110001011000;
assign LUT_4[22775] = 32'b11111111111111110010111101010000;
assign LUT_4[22776] = 32'b11111111111111110110100010101101;
assign LUT_4[22777] = 32'b11111111111111101111101110100101;
assign LUT_4[22778] = 32'b11111111111111110101111101010001;
assign LUT_4[22779] = 32'b11111111111111101111001001001001;
assign LUT_4[22780] = 32'b11111111111111110011100011001001;
assign LUT_4[22781] = 32'b11111111111111101100101111000001;
assign LUT_4[22782] = 32'b11111111111111110010111101101101;
assign LUT_4[22783] = 32'b11111111111111101100001001100101;
assign LUT_4[22784] = 32'b00000000000000000010000111101010;
assign LUT_4[22785] = 32'b11111111111111111011010011100010;
assign LUT_4[22786] = 32'b00000000000000000001100010001110;
assign LUT_4[22787] = 32'b11111111111111111010101110000110;
assign LUT_4[22788] = 32'b11111111111111111111001000000110;
assign LUT_4[22789] = 32'b11111111111111111000010011111110;
assign LUT_4[22790] = 32'b11111111111111111110100010101010;
assign LUT_4[22791] = 32'b11111111111111110111101110100010;
assign LUT_4[22792] = 32'b11111111111111111011010011111111;
assign LUT_4[22793] = 32'b11111111111111110100011111110111;
assign LUT_4[22794] = 32'b11111111111111111010101110100011;
assign LUT_4[22795] = 32'b11111111111111110011111010011011;
assign LUT_4[22796] = 32'b11111111111111111000010100011011;
assign LUT_4[22797] = 32'b11111111111111110001100000010011;
assign LUT_4[22798] = 32'b11111111111111110111101110111111;
assign LUT_4[22799] = 32'b11111111111111110000111010110111;
assign LUT_4[22800] = 32'b11111111111111111111111001011000;
assign LUT_4[22801] = 32'b11111111111111111001000101010000;
assign LUT_4[22802] = 32'b11111111111111111111010011111100;
assign LUT_4[22803] = 32'b11111111111111111000011111110100;
assign LUT_4[22804] = 32'b11111111111111111100111001110100;
assign LUT_4[22805] = 32'b11111111111111110110000101101100;
assign LUT_4[22806] = 32'b11111111111111111100010100011000;
assign LUT_4[22807] = 32'b11111111111111110101100000010000;
assign LUT_4[22808] = 32'b11111111111111111001000101101101;
assign LUT_4[22809] = 32'b11111111111111110010010001100101;
assign LUT_4[22810] = 32'b11111111111111111000100000010001;
assign LUT_4[22811] = 32'b11111111111111110001101100001001;
assign LUT_4[22812] = 32'b11111111111111110110000110001001;
assign LUT_4[22813] = 32'b11111111111111101111010010000001;
assign LUT_4[22814] = 32'b11111111111111110101100000101101;
assign LUT_4[22815] = 32'b11111111111111101110101100100101;
assign LUT_4[22816] = 32'b00000000000000000000100010110001;
assign LUT_4[22817] = 32'b11111111111111111001101110101001;
assign LUT_4[22818] = 32'b11111111111111111111111101010101;
assign LUT_4[22819] = 32'b11111111111111111001001001001101;
assign LUT_4[22820] = 32'b11111111111111111101100011001101;
assign LUT_4[22821] = 32'b11111111111111110110101111000101;
assign LUT_4[22822] = 32'b11111111111111111100111101110001;
assign LUT_4[22823] = 32'b11111111111111110110001001101001;
assign LUT_4[22824] = 32'b11111111111111111001101111000110;
assign LUT_4[22825] = 32'b11111111111111110010111010111110;
assign LUT_4[22826] = 32'b11111111111111111001001001101010;
assign LUT_4[22827] = 32'b11111111111111110010010101100010;
assign LUT_4[22828] = 32'b11111111111111110110101111100010;
assign LUT_4[22829] = 32'b11111111111111101111111011011010;
assign LUT_4[22830] = 32'b11111111111111110110001010000110;
assign LUT_4[22831] = 32'b11111111111111101111010101111110;
assign LUT_4[22832] = 32'b11111111111111111110010100011111;
assign LUT_4[22833] = 32'b11111111111111110111100000010111;
assign LUT_4[22834] = 32'b11111111111111111101101111000011;
assign LUT_4[22835] = 32'b11111111111111110110111010111011;
assign LUT_4[22836] = 32'b11111111111111111011010100111011;
assign LUT_4[22837] = 32'b11111111111111110100100000110011;
assign LUT_4[22838] = 32'b11111111111111111010101111011111;
assign LUT_4[22839] = 32'b11111111111111110011111011010111;
assign LUT_4[22840] = 32'b11111111111111110111100000110100;
assign LUT_4[22841] = 32'b11111111111111110000101100101100;
assign LUT_4[22842] = 32'b11111111111111110110111011011000;
assign LUT_4[22843] = 32'b11111111111111110000000111010000;
assign LUT_4[22844] = 32'b11111111111111110100100001010000;
assign LUT_4[22845] = 32'b11111111111111101101101101001000;
assign LUT_4[22846] = 32'b11111111111111110011111011110100;
assign LUT_4[22847] = 32'b11111111111111101101000111101100;
assign LUT_4[22848] = 32'b00000000000000000011011110111110;
assign LUT_4[22849] = 32'b11111111111111111100101010110110;
assign LUT_4[22850] = 32'b00000000000000000010111001100010;
assign LUT_4[22851] = 32'b11111111111111111100000101011010;
assign LUT_4[22852] = 32'b00000000000000000000011111011010;
assign LUT_4[22853] = 32'b11111111111111111001101011010010;
assign LUT_4[22854] = 32'b11111111111111111111111001111110;
assign LUT_4[22855] = 32'b11111111111111111001000101110110;
assign LUT_4[22856] = 32'b11111111111111111100101011010011;
assign LUT_4[22857] = 32'b11111111111111110101110111001011;
assign LUT_4[22858] = 32'b11111111111111111100000101110111;
assign LUT_4[22859] = 32'b11111111111111110101010001101111;
assign LUT_4[22860] = 32'b11111111111111111001101011101111;
assign LUT_4[22861] = 32'b11111111111111110010110111100111;
assign LUT_4[22862] = 32'b11111111111111111001000110010011;
assign LUT_4[22863] = 32'b11111111111111110010010010001011;
assign LUT_4[22864] = 32'b00000000000000000001010000101100;
assign LUT_4[22865] = 32'b11111111111111111010011100100100;
assign LUT_4[22866] = 32'b00000000000000000000101011010000;
assign LUT_4[22867] = 32'b11111111111111111001110111001000;
assign LUT_4[22868] = 32'b11111111111111111110010001001000;
assign LUT_4[22869] = 32'b11111111111111110111011101000000;
assign LUT_4[22870] = 32'b11111111111111111101101011101100;
assign LUT_4[22871] = 32'b11111111111111110110110111100100;
assign LUT_4[22872] = 32'b11111111111111111010011101000001;
assign LUT_4[22873] = 32'b11111111111111110011101000111001;
assign LUT_4[22874] = 32'b11111111111111111001110111100101;
assign LUT_4[22875] = 32'b11111111111111110011000011011101;
assign LUT_4[22876] = 32'b11111111111111110111011101011101;
assign LUT_4[22877] = 32'b11111111111111110000101001010101;
assign LUT_4[22878] = 32'b11111111111111110110111000000001;
assign LUT_4[22879] = 32'b11111111111111110000000011111001;
assign LUT_4[22880] = 32'b00000000000000000001111010000101;
assign LUT_4[22881] = 32'b11111111111111111011000101111101;
assign LUT_4[22882] = 32'b00000000000000000001010100101001;
assign LUT_4[22883] = 32'b11111111111111111010100000100001;
assign LUT_4[22884] = 32'b11111111111111111110111010100001;
assign LUT_4[22885] = 32'b11111111111111111000000110011001;
assign LUT_4[22886] = 32'b11111111111111111110010101000101;
assign LUT_4[22887] = 32'b11111111111111110111100000111101;
assign LUT_4[22888] = 32'b11111111111111111011000110011010;
assign LUT_4[22889] = 32'b11111111111111110100010010010010;
assign LUT_4[22890] = 32'b11111111111111111010100000111110;
assign LUT_4[22891] = 32'b11111111111111110011101100110110;
assign LUT_4[22892] = 32'b11111111111111111000000110110110;
assign LUT_4[22893] = 32'b11111111111111110001010010101110;
assign LUT_4[22894] = 32'b11111111111111110111100001011010;
assign LUT_4[22895] = 32'b11111111111111110000101101010010;
assign LUT_4[22896] = 32'b11111111111111111111101011110011;
assign LUT_4[22897] = 32'b11111111111111111000110111101011;
assign LUT_4[22898] = 32'b11111111111111111111000110010111;
assign LUT_4[22899] = 32'b11111111111111111000010010001111;
assign LUT_4[22900] = 32'b11111111111111111100101100001111;
assign LUT_4[22901] = 32'b11111111111111110101111000000111;
assign LUT_4[22902] = 32'b11111111111111111100000110110011;
assign LUT_4[22903] = 32'b11111111111111110101010010101011;
assign LUT_4[22904] = 32'b11111111111111111000111000001000;
assign LUT_4[22905] = 32'b11111111111111110010000100000000;
assign LUT_4[22906] = 32'b11111111111111111000010010101100;
assign LUT_4[22907] = 32'b11111111111111110001011110100100;
assign LUT_4[22908] = 32'b11111111111111110101111000100100;
assign LUT_4[22909] = 32'b11111111111111101111000100011100;
assign LUT_4[22910] = 32'b11111111111111110101010011001000;
assign LUT_4[22911] = 32'b11111111111111101110011111000000;
assign LUT_4[22912] = 32'b00000000000000000100101101110010;
assign LUT_4[22913] = 32'b11111111111111111101111001101010;
assign LUT_4[22914] = 32'b00000000000000000100001000010110;
assign LUT_4[22915] = 32'b11111111111111111101010100001110;
assign LUT_4[22916] = 32'b00000000000000000001101110001110;
assign LUT_4[22917] = 32'b11111111111111111010111010000110;
assign LUT_4[22918] = 32'b00000000000000000001001000110010;
assign LUT_4[22919] = 32'b11111111111111111010010100101010;
assign LUT_4[22920] = 32'b11111111111111111101111010000111;
assign LUT_4[22921] = 32'b11111111111111110111000101111111;
assign LUT_4[22922] = 32'b11111111111111111101010100101011;
assign LUT_4[22923] = 32'b11111111111111110110100000100011;
assign LUT_4[22924] = 32'b11111111111111111010111010100011;
assign LUT_4[22925] = 32'b11111111111111110100000110011011;
assign LUT_4[22926] = 32'b11111111111111111010010101000111;
assign LUT_4[22927] = 32'b11111111111111110011100000111111;
assign LUT_4[22928] = 32'b00000000000000000010011111100000;
assign LUT_4[22929] = 32'b11111111111111111011101011011000;
assign LUT_4[22930] = 32'b00000000000000000001111010000100;
assign LUT_4[22931] = 32'b11111111111111111011000101111100;
assign LUT_4[22932] = 32'b11111111111111111111011111111100;
assign LUT_4[22933] = 32'b11111111111111111000101011110100;
assign LUT_4[22934] = 32'b11111111111111111110111010100000;
assign LUT_4[22935] = 32'b11111111111111111000000110011000;
assign LUT_4[22936] = 32'b11111111111111111011101011110101;
assign LUT_4[22937] = 32'b11111111111111110100110111101101;
assign LUT_4[22938] = 32'b11111111111111111011000110011001;
assign LUT_4[22939] = 32'b11111111111111110100010010010001;
assign LUT_4[22940] = 32'b11111111111111111000101100010001;
assign LUT_4[22941] = 32'b11111111111111110001111000001001;
assign LUT_4[22942] = 32'b11111111111111111000000110110101;
assign LUT_4[22943] = 32'b11111111111111110001010010101101;
assign LUT_4[22944] = 32'b00000000000000000011001000111001;
assign LUT_4[22945] = 32'b11111111111111111100010100110001;
assign LUT_4[22946] = 32'b00000000000000000010100011011101;
assign LUT_4[22947] = 32'b11111111111111111011101111010101;
assign LUT_4[22948] = 32'b00000000000000000000001001010101;
assign LUT_4[22949] = 32'b11111111111111111001010101001101;
assign LUT_4[22950] = 32'b11111111111111111111100011111001;
assign LUT_4[22951] = 32'b11111111111111111000101111110001;
assign LUT_4[22952] = 32'b11111111111111111100010101001110;
assign LUT_4[22953] = 32'b11111111111111110101100001000110;
assign LUT_4[22954] = 32'b11111111111111111011101111110010;
assign LUT_4[22955] = 32'b11111111111111110100111011101010;
assign LUT_4[22956] = 32'b11111111111111111001010101101010;
assign LUT_4[22957] = 32'b11111111111111110010100001100010;
assign LUT_4[22958] = 32'b11111111111111111000110000001110;
assign LUT_4[22959] = 32'b11111111111111110001111100000110;
assign LUT_4[22960] = 32'b00000000000000000000111010100111;
assign LUT_4[22961] = 32'b11111111111111111010000110011111;
assign LUT_4[22962] = 32'b00000000000000000000010101001011;
assign LUT_4[22963] = 32'b11111111111111111001100001000011;
assign LUT_4[22964] = 32'b11111111111111111101111011000011;
assign LUT_4[22965] = 32'b11111111111111110111000110111011;
assign LUT_4[22966] = 32'b11111111111111111101010101100111;
assign LUT_4[22967] = 32'b11111111111111110110100001011111;
assign LUT_4[22968] = 32'b11111111111111111010000110111100;
assign LUT_4[22969] = 32'b11111111111111110011010010110100;
assign LUT_4[22970] = 32'b11111111111111111001100001100000;
assign LUT_4[22971] = 32'b11111111111111110010101101011000;
assign LUT_4[22972] = 32'b11111111111111110111000111011000;
assign LUT_4[22973] = 32'b11111111111111110000010011010000;
assign LUT_4[22974] = 32'b11111111111111110110100001111100;
assign LUT_4[22975] = 32'b11111111111111101111101101110100;
assign LUT_4[22976] = 32'b00000000000000000110000101000110;
assign LUT_4[22977] = 32'b11111111111111111111010000111110;
assign LUT_4[22978] = 32'b00000000000000000101011111101010;
assign LUT_4[22979] = 32'b11111111111111111110101011100010;
assign LUT_4[22980] = 32'b00000000000000000011000101100010;
assign LUT_4[22981] = 32'b11111111111111111100010001011010;
assign LUT_4[22982] = 32'b00000000000000000010100000000110;
assign LUT_4[22983] = 32'b11111111111111111011101011111110;
assign LUT_4[22984] = 32'b11111111111111111111010001011011;
assign LUT_4[22985] = 32'b11111111111111111000011101010011;
assign LUT_4[22986] = 32'b11111111111111111110101011111111;
assign LUT_4[22987] = 32'b11111111111111110111110111110111;
assign LUT_4[22988] = 32'b11111111111111111100010001110111;
assign LUT_4[22989] = 32'b11111111111111110101011101101111;
assign LUT_4[22990] = 32'b11111111111111111011101100011011;
assign LUT_4[22991] = 32'b11111111111111110100111000010011;
assign LUT_4[22992] = 32'b00000000000000000011110110110100;
assign LUT_4[22993] = 32'b11111111111111111101000010101100;
assign LUT_4[22994] = 32'b00000000000000000011010001011000;
assign LUT_4[22995] = 32'b11111111111111111100011101010000;
assign LUT_4[22996] = 32'b00000000000000000000110111010000;
assign LUT_4[22997] = 32'b11111111111111111010000011001000;
assign LUT_4[22998] = 32'b00000000000000000000010001110100;
assign LUT_4[22999] = 32'b11111111111111111001011101101100;
assign LUT_4[23000] = 32'b11111111111111111101000011001001;
assign LUT_4[23001] = 32'b11111111111111110110001111000001;
assign LUT_4[23002] = 32'b11111111111111111100011101101101;
assign LUT_4[23003] = 32'b11111111111111110101101001100101;
assign LUT_4[23004] = 32'b11111111111111111010000011100101;
assign LUT_4[23005] = 32'b11111111111111110011001111011101;
assign LUT_4[23006] = 32'b11111111111111111001011110001001;
assign LUT_4[23007] = 32'b11111111111111110010101010000001;
assign LUT_4[23008] = 32'b00000000000000000100100000001101;
assign LUT_4[23009] = 32'b11111111111111111101101100000101;
assign LUT_4[23010] = 32'b00000000000000000011111010110001;
assign LUT_4[23011] = 32'b11111111111111111101000110101001;
assign LUT_4[23012] = 32'b00000000000000000001100000101001;
assign LUT_4[23013] = 32'b11111111111111111010101100100001;
assign LUT_4[23014] = 32'b00000000000000000000111011001101;
assign LUT_4[23015] = 32'b11111111111111111010000111000101;
assign LUT_4[23016] = 32'b11111111111111111101101100100010;
assign LUT_4[23017] = 32'b11111111111111110110111000011010;
assign LUT_4[23018] = 32'b11111111111111111101000111000110;
assign LUT_4[23019] = 32'b11111111111111110110010010111110;
assign LUT_4[23020] = 32'b11111111111111111010101100111110;
assign LUT_4[23021] = 32'b11111111111111110011111000110110;
assign LUT_4[23022] = 32'b11111111111111111010000111100010;
assign LUT_4[23023] = 32'b11111111111111110011010011011010;
assign LUT_4[23024] = 32'b00000000000000000010010001111011;
assign LUT_4[23025] = 32'b11111111111111111011011101110011;
assign LUT_4[23026] = 32'b00000000000000000001101100011111;
assign LUT_4[23027] = 32'b11111111111111111010111000010111;
assign LUT_4[23028] = 32'b11111111111111111111010010010111;
assign LUT_4[23029] = 32'b11111111111111111000011110001111;
assign LUT_4[23030] = 32'b11111111111111111110101100111011;
assign LUT_4[23031] = 32'b11111111111111110111111000110011;
assign LUT_4[23032] = 32'b11111111111111111011011110010000;
assign LUT_4[23033] = 32'b11111111111111110100101010001000;
assign LUT_4[23034] = 32'b11111111111111111010111000110100;
assign LUT_4[23035] = 32'b11111111111111110100000100101100;
assign LUT_4[23036] = 32'b11111111111111111000011110101100;
assign LUT_4[23037] = 32'b11111111111111110001101010100100;
assign LUT_4[23038] = 32'b11111111111111110111111001010000;
assign LUT_4[23039] = 32'b11111111111111110001000101001000;
assign LUT_4[23040] = 32'b11111111111111111100010000001111;
assign LUT_4[23041] = 32'b11111111111111110101011100000111;
assign LUT_4[23042] = 32'b11111111111111111011101010110011;
assign LUT_4[23043] = 32'b11111111111111110100110110101011;
assign LUT_4[23044] = 32'b11111111111111111001010000101011;
assign LUT_4[23045] = 32'b11111111111111110010011100100011;
assign LUT_4[23046] = 32'b11111111111111111000101011001111;
assign LUT_4[23047] = 32'b11111111111111110001110111000111;
assign LUT_4[23048] = 32'b11111111111111110101011100100100;
assign LUT_4[23049] = 32'b11111111111111101110101000011100;
assign LUT_4[23050] = 32'b11111111111111110100110111001000;
assign LUT_4[23051] = 32'b11111111111111101110000011000000;
assign LUT_4[23052] = 32'b11111111111111110010011101000000;
assign LUT_4[23053] = 32'b11111111111111101011101000111000;
assign LUT_4[23054] = 32'b11111111111111110001110111100100;
assign LUT_4[23055] = 32'b11111111111111101011000011011100;
assign LUT_4[23056] = 32'b11111111111111111010000001111101;
assign LUT_4[23057] = 32'b11111111111111110011001101110101;
assign LUT_4[23058] = 32'b11111111111111111001011100100001;
assign LUT_4[23059] = 32'b11111111111111110010101000011001;
assign LUT_4[23060] = 32'b11111111111111110111000010011001;
assign LUT_4[23061] = 32'b11111111111111110000001110010001;
assign LUT_4[23062] = 32'b11111111111111110110011100111101;
assign LUT_4[23063] = 32'b11111111111111101111101000110101;
assign LUT_4[23064] = 32'b11111111111111110011001110010010;
assign LUT_4[23065] = 32'b11111111111111101100011010001010;
assign LUT_4[23066] = 32'b11111111111111110010101000110110;
assign LUT_4[23067] = 32'b11111111111111101011110100101110;
assign LUT_4[23068] = 32'b11111111111111110000001110101110;
assign LUT_4[23069] = 32'b11111111111111101001011010100110;
assign LUT_4[23070] = 32'b11111111111111101111101001010010;
assign LUT_4[23071] = 32'b11111111111111101000110101001010;
assign LUT_4[23072] = 32'b11111111111111111010101011010110;
assign LUT_4[23073] = 32'b11111111111111110011110111001110;
assign LUT_4[23074] = 32'b11111111111111111010000101111010;
assign LUT_4[23075] = 32'b11111111111111110011010001110010;
assign LUT_4[23076] = 32'b11111111111111110111101011110010;
assign LUT_4[23077] = 32'b11111111111111110000110111101010;
assign LUT_4[23078] = 32'b11111111111111110111000110010110;
assign LUT_4[23079] = 32'b11111111111111110000010010001110;
assign LUT_4[23080] = 32'b11111111111111110011110111101011;
assign LUT_4[23081] = 32'b11111111111111101101000011100011;
assign LUT_4[23082] = 32'b11111111111111110011010010001111;
assign LUT_4[23083] = 32'b11111111111111101100011110000111;
assign LUT_4[23084] = 32'b11111111111111110000111000000111;
assign LUT_4[23085] = 32'b11111111111111101010000011111111;
assign LUT_4[23086] = 32'b11111111111111110000010010101011;
assign LUT_4[23087] = 32'b11111111111111101001011110100011;
assign LUT_4[23088] = 32'b11111111111111111000011101000100;
assign LUT_4[23089] = 32'b11111111111111110001101000111100;
assign LUT_4[23090] = 32'b11111111111111110111110111101000;
assign LUT_4[23091] = 32'b11111111111111110001000011100000;
assign LUT_4[23092] = 32'b11111111111111110101011101100000;
assign LUT_4[23093] = 32'b11111111111111101110101001011000;
assign LUT_4[23094] = 32'b11111111111111110100111000000100;
assign LUT_4[23095] = 32'b11111111111111101110000011111100;
assign LUT_4[23096] = 32'b11111111111111110001101001011001;
assign LUT_4[23097] = 32'b11111111111111101010110101010001;
assign LUT_4[23098] = 32'b11111111111111110001000011111101;
assign LUT_4[23099] = 32'b11111111111111101010001111110101;
assign LUT_4[23100] = 32'b11111111111111101110101001110101;
assign LUT_4[23101] = 32'b11111111111111100111110101101101;
assign LUT_4[23102] = 32'b11111111111111101110000100011001;
assign LUT_4[23103] = 32'b11111111111111100111010000010001;
assign LUT_4[23104] = 32'b11111111111111111101100111100011;
assign LUT_4[23105] = 32'b11111111111111110110110011011011;
assign LUT_4[23106] = 32'b11111111111111111101000010000111;
assign LUT_4[23107] = 32'b11111111111111110110001101111111;
assign LUT_4[23108] = 32'b11111111111111111010100111111111;
assign LUT_4[23109] = 32'b11111111111111110011110011110111;
assign LUT_4[23110] = 32'b11111111111111111010000010100011;
assign LUT_4[23111] = 32'b11111111111111110011001110011011;
assign LUT_4[23112] = 32'b11111111111111110110110011111000;
assign LUT_4[23113] = 32'b11111111111111101111111111110000;
assign LUT_4[23114] = 32'b11111111111111110110001110011100;
assign LUT_4[23115] = 32'b11111111111111101111011010010100;
assign LUT_4[23116] = 32'b11111111111111110011110100010100;
assign LUT_4[23117] = 32'b11111111111111101101000000001100;
assign LUT_4[23118] = 32'b11111111111111110011001110111000;
assign LUT_4[23119] = 32'b11111111111111101100011010110000;
assign LUT_4[23120] = 32'b11111111111111111011011001010001;
assign LUT_4[23121] = 32'b11111111111111110100100101001001;
assign LUT_4[23122] = 32'b11111111111111111010110011110101;
assign LUT_4[23123] = 32'b11111111111111110011111111101101;
assign LUT_4[23124] = 32'b11111111111111111000011001101101;
assign LUT_4[23125] = 32'b11111111111111110001100101100101;
assign LUT_4[23126] = 32'b11111111111111110111110100010001;
assign LUT_4[23127] = 32'b11111111111111110001000000001001;
assign LUT_4[23128] = 32'b11111111111111110100100101100110;
assign LUT_4[23129] = 32'b11111111111111101101110001011110;
assign LUT_4[23130] = 32'b11111111111111110100000000001010;
assign LUT_4[23131] = 32'b11111111111111101101001100000010;
assign LUT_4[23132] = 32'b11111111111111110001100110000010;
assign LUT_4[23133] = 32'b11111111111111101010110001111010;
assign LUT_4[23134] = 32'b11111111111111110001000000100110;
assign LUT_4[23135] = 32'b11111111111111101010001100011110;
assign LUT_4[23136] = 32'b11111111111111111100000010101010;
assign LUT_4[23137] = 32'b11111111111111110101001110100010;
assign LUT_4[23138] = 32'b11111111111111111011011101001110;
assign LUT_4[23139] = 32'b11111111111111110100101001000110;
assign LUT_4[23140] = 32'b11111111111111111001000011000110;
assign LUT_4[23141] = 32'b11111111111111110010001110111110;
assign LUT_4[23142] = 32'b11111111111111111000011101101010;
assign LUT_4[23143] = 32'b11111111111111110001101001100010;
assign LUT_4[23144] = 32'b11111111111111110101001110111111;
assign LUT_4[23145] = 32'b11111111111111101110011010110111;
assign LUT_4[23146] = 32'b11111111111111110100101001100011;
assign LUT_4[23147] = 32'b11111111111111101101110101011011;
assign LUT_4[23148] = 32'b11111111111111110010001111011011;
assign LUT_4[23149] = 32'b11111111111111101011011011010011;
assign LUT_4[23150] = 32'b11111111111111110001101001111111;
assign LUT_4[23151] = 32'b11111111111111101010110101110111;
assign LUT_4[23152] = 32'b11111111111111111001110100011000;
assign LUT_4[23153] = 32'b11111111111111110011000000010000;
assign LUT_4[23154] = 32'b11111111111111111001001110111100;
assign LUT_4[23155] = 32'b11111111111111110010011010110100;
assign LUT_4[23156] = 32'b11111111111111110110110100110100;
assign LUT_4[23157] = 32'b11111111111111110000000000101100;
assign LUT_4[23158] = 32'b11111111111111110110001111011000;
assign LUT_4[23159] = 32'b11111111111111101111011011010000;
assign LUT_4[23160] = 32'b11111111111111110011000000101101;
assign LUT_4[23161] = 32'b11111111111111101100001100100101;
assign LUT_4[23162] = 32'b11111111111111110010011011010001;
assign LUT_4[23163] = 32'b11111111111111101011100111001001;
assign LUT_4[23164] = 32'b11111111111111110000000001001001;
assign LUT_4[23165] = 32'b11111111111111101001001101000001;
assign LUT_4[23166] = 32'b11111111111111101111011011101101;
assign LUT_4[23167] = 32'b11111111111111101000100111100101;
assign LUT_4[23168] = 32'b11111111111111111110110110010111;
assign LUT_4[23169] = 32'b11111111111111111000000010001111;
assign LUT_4[23170] = 32'b11111111111111111110010000111011;
assign LUT_4[23171] = 32'b11111111111111110111011100110011;
assign LUT_4[23172] = 32'b11111111111111111011110110110011;
assign LUT_4[23173] = 32'b11111111111111110101000010101011;
assign LUT_4[23174] = 32'b11111111111111111011010001010111;
assign LUT_4[23175] = 32'b11111111111111110100011101001111;
assign LUT_4[23176] = 32'b11111111111111111000000010101100;
assign LUT_4[23177] = 32'b11111111111111110001001110100100;
assign LUT_4[23178] = 32'b11111111111111110111011101010000;
assign LUT_4[23179] = 32'b11111111111111110000101001001000;
assign LUT_4[23180] = 32'b11111111111111110101000011001000;
assign LUT_4[23181] = 32'b11111111111111101110001111000000;
assign LUT_4[23182] = 32'b11111111111111110100011101101100;
assign LUT_4[23183] = 32'b11111111111111101101101001100100;
assign LUT_4[23184] = 32'b11111111111111111100101000000101;
assign LUT_4[23185] = 32'b11111111111111110101110011111101;
assign LUT_4[23186] = 32'b11111111111111111100000010101001;
assign LUT_4[23187] = 32'b11111111111111110101001110100001;
assign LUT_4[23188] = 32'b11111111111111111001101000100001;
assign LUT_4[23189] = 32'b11111111111111110010110100011001;
assign LUT_4[23190] = 32'b11111111111111111001000011000101;
assign LUT_4[23191] = 32'b11111111111111110010001110111101;
assign LUT_4[23192] = 32'b11111111111111110101110100011010;
assign LUT_4[23193] = 32'b11111111111111101111000000010010;
assign LUT_4[23194] = 32'b11111111111111110101001110111110;
assign LUT_4[23195] = 32'b11111111111111101110011010110110;
assign LUT_4[23196] = 32'b11111111111111110010110100110110;
assign LUT_4[23197] = 32'b11111111111111101100000000101110;
assign LUT_4[23198] = 32'b11111111111111110010001111011010;
assign LUT_4[23199] = 32'b11111111111111101011011011010010;
assign LUT_4[23200] = 32'b11111111111111111101010001011110;
assign LUT_4[23201] = 32'b11111111111111110110011101010110;
assign LUT_4[23202] = 32'b11111111111111111100101100000010;
assign LUT_4[23203] = 32'b11111111111111110101110111111010;
assign LUT_4[23204] = 32'b11111111111111111010010001111010;
assign LUT_4[23205] = 32'b11111111111111110011011101110010;
assign LUT_4[23206] = 32'b11111111111111111001101100011110;
assign LUT_4[23207] = 32'b11111111111111110010111000010110;
assign LUT_4[23208] = 32'b11111111111111110110011101110011;
assign LUT_4[23209] = 32'b11111111111111101111101001101011;
assign LUT_4[23210] = 32'b11111111111111110101111000010111;
assign LUT_4[23211] = 32'b11111111111111101111000100001111;
assign LUT_4[23212] = 32'b11111111111111110011011110001111;
assign LUT_4[23213] = 32'b11111111111111101100101010000111;
assign LUT_4[23214] = 32'b11111111111111110010111000110011;
assign LUT_4[23215] = 32'b11111111111111101100000100101011;
assign LUT_4[23216] = 32'b11111111111111111011000011001100;
assign LUT_4[23217] = 32'b11111111111111110100001111000100;
assign LUT_4[23218] = 32'b11111111111111111010011101110000;
assign LUT_4[23219] = 32'b11111111111111110011101001101000;
assign LUT_4[23220] = 32'b11111111111111111000000011101000;
assign LUT_4[23221] = 32'b11111111111111110001001111100000;
assign LUT_4[23222] = 32'b11111111111111110111011110001100;
assign LUT_4[23223] = 32'b11111111111111110000101010000100;
assign LUT_4[23224] = 32'b11111111111111110100001111100001;
assign LUT_4[23225] = 32'b11111111111111101101011011011001;
assign LUT_4[23226] = 32'b11111111111111110011101010000101;
assign LUT_4[23227] = 32'b11111111111111101100110101111101;
assign LUT_4[23228] = 32'b11111111111111110001001111111101;
assign LUT_4[23229] = 32'b11111111111111101010011011110101;
assign LUT_4[23230] = 32'b11111111111111110000101010100001;
assign LUT_4[23231] = 32'b11111111111111101001110110011001;
assign LUT_4[23232] = 32'b00000000000000000000001101101011;
assign LUT_4[23233] = 32'b11111111111111111001011001100011;
assign LUT_4[23234] = 32'b11111111111111111111101000001111;
assign LUT_4[23235] = 32'b11111111111111111000110100000111;
assign LUT_4[23236] = 32'b11111111111111111101001110000111;
assign LUT_4[23237] = 32'b11111111111111110110011001111111;
assign LUT_4[23238] = 32'b11111111111111111100101000101011;
assign LUT_4[23239] = 32'b11111111111111110101110100100011;
assign LUT_4[23240] = 32'b11111111111111111001011010000000;
assign LUT_4[23241] = 32'b11111111111111110010100101111000;
assign LUT_4[23242] = 32'b11111111111111111000110100100100;
assign LUT_4[23243] = 32'b11111111111111110010000000011100;
assign LUT_4[23244] = 32'b11111111111111110110011010011100;
assign LUT_4[23245] = 32'b11111111111111101111100110010100;
assign LUT_4[23246] = 32'b11111111111111110101110101000000;
assign LUT_4[23247] = 32'b11111111111111101111000000111000;
assign LUT_4[23248] = 32'b11111111111111111101111111011001;
assign LUT_4[23249] = 32'b11111111111111110111001011010001;
assign LUT_4[23250] = 32'b11111111111111111101011001111101;
assign LUT_4[23251] = 32'b11111111111111110110100101110101;
assign LUT_4[23252] = 32'b11111111111111111010111111110101;
assign LUT_4[23253] = 32'b11111111111111110100001011101101;
assign LUT_4[23254] = 32'b11111111111111111010011010011001;
assign LUT_4[23255] = 32'b11111111111111110011100110010001;
assign LUT_4[23256] = 32'b11111111111111110111001011101110;
assign LUT_4[23257] = 32'b11111111111111110000010111100110;
assign LUT_4[23258] = 32'b11111111111111110110100110010010;
assign LUT_4[23259] = 32'b11111111111111101111110010001010;
assign LUT_4[23260] = 32'b11111111111111110100001100001010;
assign LUT_4[23261] = 32'b11111111111111101101011000000010;
assign LUT_4[23262] = 32'b11111111111111110011100110101110;
assign LUT_4[23263] = 32'b11111111111111101100110010100110;
assign LUT_4[23264] = 32'b11111111111111111110101000110010;
assign LUT_4[23265] = 32'b11111111111111110111110100101010;
assign LUT_4[23266] = 32'b11111111111111111110000011010110;
assign LUT_4[23267] = 32'b11111111111111110111001111001110;
assign LUT_4[23268] = 32'b11111111111111111011101001001110;
assign LUT_4[23269] = 32'b11111111111111110100110101000110;
assign LUT_4[23270] = 32'b11111111111111111011000011110010;
assign LUT_4[23271] = 32'b11111111111111110100001111101010;
assign LUT_4[23272] = 32'b11111111111111110111110101000111;
assign LUT_4[23273] = 32'b11111111111111110001000000111111;
assign LUT_4[23274] = 32'b11111111111111110111001111101011;
assign LUT_4[23275] = 32'b11111111111111110000011011100011;
assign LUT_4[23276] = 32'b11111111111111110100110101100011;
assign LUT_4[23277] = 32'b11111111111111101110000001011011;
assign LUT_4[23278] = 32'b11111111111111110100010000000111;
assign LUT_4[23279] = 32'b11111111111111101101011011111111;
assign LUT_4[23280] = 32'b11111111111111111100011010100000;
assign LUT_4[23281] = 32'b11111111111111110101100110011000;
assign LUT_4[23282] = 32'b11111111111111111011110101000100;
assign LUT_4[23283] = 32'b11111111111111110101000000111100;
assign LUT_4[23284] = 32'b11111111111111111001011010111100;
assign LUT_4[23285] = 32'b11111111111111110010100110110100;
assign LUT_4[23286] = 32'b11111111111111111000110101100000;
assign LUT_4[23287] = 32'b11111111111111110010000001011000;
assign LUT_4[23288] = 32'b11111111111111110101100110110101;
assign LUT_4[23289] = 32'b11111111111111101110110010101101;
assign LUT_4[23290] = 32'b11111111111111110101000001011001;
assign LUT_4[23291] = 32'b11111111111111101110001101010001;
assign LUT_4[23292] = 32'b11111111111111110010100111010001;
assign LUT_4[23293] = 32'b11111111111111101011110011001001;
assign LUT_4[23294] = 32'b11111111111111110010000001110101;
assign LUT_4[23295] = 32'b11111111111111101011001101101101;
assign LUT_4[23296] = 32'b00000000000000000001001011110010;
assign LUT_4[23297] = 32'b11111111111111111010010111101010;
assign LUT_4[23298] = 32'b00000000000000000000100110010110;
assign LUT_4[23299] = 32'b11111111111111111001110010001110;
assign LUT_4[23300] = 32'b11111111111111111110001100001110;
assign LUT_4[23301] = 32'b11111111111111110111011000000110;
assign LUT_4[23302] = 32'b11111111111111111101100110110010;
assign LUT_4[23303] = 32'b11111111111111110110110010101010;
assign LUT_4[23304] = 32'b11111111111111111010011000000111;
assign LUT_4[23305] = 32'b11111111111111110011100011111111;
assign LUT_4[23306] = 32'b11111111111111111001110010101011;
assign LUT_4[23307] = 32'b11111111111111110010111110100011;
assign LUT_4[23308] = 32'b11111111111111110111011000100011;
assign LUT_4[23309] = 32'b11111111111111110000100100011011;
assign LUT_4[23310] = 32'b11111111111111110110110011000111;
assign LUT_4[23311] = 32'b11111111111111101111111110111111;
assign LUT_4[23312] = 32'b11111111111111111110111101100000;
assign LUT_4[23313] = 32'b11111111111111111000001001011000;
assign LUT_4[23314] = 32'b11111111111111111110011000000100;
assign LUT_4[23315] = 32'b11111111111111110111100011111100;
assign LUT_4[23316] = 32'b11111111111111111011111101111100;
assign LUT_4[23317] = 32'b11111111111111110101001001110100;
assign LUT_4[23318] = 32'b11111111111111111011011000100000;
assign LUT_4[23319] = 32'b11111111111111110100100100011000;
assign LUT_4[23320] = 32'b11111111111111111000001001110101;
assign LUT_4[23321] = 32'b11111111111111110001010101101101;
assign LUT_4[23322] = 32'b11111111111111110111100100011001;
assign LUT_4[23323] = 32'b11111111111111110000110000010001;
assign LUT_4[23324] = 32'b11111111111111110101001010010001;
assign LUT_4[23325] = 32'b11111111111111101110010110001001;
assign LUT_4[23326] = 32'b11111111111111110100100100110101;
assign LUT_4[23327] = 32'b11111111111111101101110000101101;
assign LUT_4[23328] = 32'b11111111111111111111100110111001;
assign LUT_4[23329] = 32'b11111111111111111000110010110001;
assign LUT_4[23330] = 32'b11111111111111111111000001011101;
assign LUT_4[23331] = 32'b11111111111111111000001101010101;
assign LUT_4[23332] = 32'b11111111111111111100100111010101;
assign LUT_4[23333] = 32'b11111111111111110101110011001101;
assign LUT_4[23334] = 32'b11111111111111111100000001111001;
assign LUT_4[23335] = 32'b11111111111111110101001101110001;
assign LUT_4[23336] = 32'b11111111111111111000110011001110;
assign LUT_4[23337] = 32'b11111111111111110001111111000110;
assign LUT_4[23338] = 32'b11111111111111111000001101110010;
assign LUT_4[23339] = 32'b11111111111111110001011001101010;
assign LUT_4[23340] = 32'b11111111111111110101110011101010;
assign LUT_4[23341] = 32'b11111111111111101110111111100010;
assign LUT_4[23342] = 32'b11111111111111110101001110001110;
assign LUT_4[23343] = 32'b11111111111111101110011010000110;
assign LUT_4[23344] = 32'b11111111111111111101011000100111;
assign LUT_4[23345] = 32'b11111111111111110110100100011111;
assign LUT_4[23346] = 32'b11111111111111111100110011001011;
assign LUT_4[23347] = 32'b11111111111111110101111111000011;
assign LUT_4[23348] = 32'b11111111111111111010011001000011;
assign LUT_4[23349] = 32'b11111111111111110011100100111011;
assign LUT_4[23350] = 32'b11111111111111111001110011100111;
assign LUT_4[23351] = 32'b11111111111111110010111111011111;
assign LUT_4[23352] = 32'b11111111111111110110100100111100;
assign LUT_4[23353] = 32'b11111111111111101111110000110100;
assign LUT_4[23354] = 32'b11111111111111110101111111100000;
assign LUT_4[23355] = 32'b11111111111111101111001011011000;
assign LUT_4[23356] = 32'b11111111111111110011100101011000;
assign LUT_4[23357] = 32'b11111111111111101100110001010000;
assign LUT_4[23358] = 32'b11111111111111110010111111111100;
assign LUT_4[23359] = 32'b11111111111111101100001011110100;
assign LUT_4[23360] = 32'b00000000000000000010100011000110;
assign LUT_4[23361] = 32'b11111111111111111011101110111110;
assign LUT_4[23362] = 32'b00000000000000000001111101101010;
assign LUT_4[23363] = 32'b11111111111111111011001001100010;
assign LUT_4[23364] = 32'b11111111111111111111100011100010;
assign LUT_4[23365] = 32'b11111111111111111000101111011010;
assign LUT_4[23366] = 32'b11111111111111111110111110000110;
assign LUT_4[23367] = 32'b11111111111111111000001001111110;
assign LUT_4[23368] = 32'b11111111111111111011101111011011;
assign LUT_4[23369] = 32'b11111111111111110100111011010011;
assign LUT_4[23370] = 32'b11111111111111111011001001111111;
assign LUT_4[23371] = 32'b11111111111111110100010101110111;
assign LUT_4[23372] = 32'b11111111111111111000101111110111;
assign LUT_4[23373] = 32'b11111111111111110001111011101111;
assign LUT_4[23374] = 32'b11111111111111111000001010011011;
assign LUT_4[23375] = 32'b11111111111111110001010110010011;
assign LUT_4[23376] = 32'b00000000000000000000010100110100;
assign LUT_4[23377] = 32'b11111111111111111001100000101100;
assign LUT_4[23378] = 32'b11111111111111111111101111011000;
assign LUT_4[23379] = 32'b11111111111111111000111011010000;
assign LUT_4[23380] = 32'b11111111111111111101010101010000;
assign LUT_4[23381] = 32'b11111111111111110110100001001000;
assign LUT_4[23382] = 32'b11111111111111111100101111110100;
assign LUT_4[23383] = 32'b11111111111111110101111011101100;
assign LUT_4[23384] = 32'b11111111111111111001100001001001;
assign LUT_4[23385] = 32'b11111111111111110010101101000001;
assign LUT_4[23386] = 32'b11111111111111111000111011101101;
assign LUT_4[23387] = 32'b11111111111111110010000111100101;
assign LUT_4[23388] = 32'b11111111111111110110100001100101;
assign LUT_4[23389] = 32'b11111111111111101111101101011101;
assign LUT_4[23390] = 32'b11111111111111110101111100001001;
assign LUT_4[23391] = 32'b11111111111111101111001000000001;
assign LUT_4[23392] = 32'b00000000000000000000111110001101;
assign LUT_4[23393] = 32'b11111111111111111010001010000101;
assign LUT_4[23394] = 32'b00000000000000000000011000110001;
assign LUT_4[23395] = 32'b11111111111111111001100100101001;
assign LUT_4[23396] = 32'b11111111111111111101111110101001;
assign LUT_4[23397] = 32'b11111111111111110111001010100001;
assign LUT_4[23398] = 32'b11111111111111111101011001001101;
assign LUT_4[23399] = 32'b11111111111111110110100101000101;
assign LUT_4[23400] = 32'b11111111111111111010001010100010;
assign LUT_4[23401] = 32'b11111111111111110011010110011010;
assign LUT_4[23402] = 32'b11111111111111111001100101000110;
assign LUT_4[23403] = 32'b11111111111111110010110000111110;
assign LUT_4[23404] = 32'b11111111111111110111001010111110;
assign LUT_4[23405] = 32'b11111111111111110000010110110110;
assign LUT_4[23406] = 32'b11111111111111110110100101100010;
assign LUT_4[23407] = 32'b11111111111111101111110001011010;
assign LUT_4[23408] = 32'b11111111111111111110101111111011;
assign LUT_4[23409] = 32'b11111111111111110111111011110011;
assign LUT_4[23410] = 32'b11111111111111111110001010011111;
assign LUT_4[23411] = 32'b11111111111111110111010110010111;
assign LUT_4[23412] = 32'b11111111111111111011110000010111;
assign LUT_4[23413] = 32'b11111111111111110100111100001111;
assign LUT_4[23414] = 32'b11111111111111111011001010111011;
assign LUT_4[23415] = 32'b11111111111111110100010110110011;
assign LUT_4[23416] = 32'b11111111111111110111111100010000;
assign LUT_4[23417] = 32'b11111111111111110001001000001000;
assign LUT_4[23418] = 32'b11111111111111110111010110110100;
assign LUT_4[23419] = 32'b11111111111111110000100010101100;
assign LUT_4[23420] = 32'b11111111111111110100111100101100;
assign LUT_4[23421] = 32'b11111111111111101110001000100100;
assign LUT_4[23422] = 32'b11111111111111110100010111010000;
assign LUT_4[23423] = 32'b11111111111111101101100011001000;
assign LUT_4[23424] = 32'b00000000000000000011110001111010;
assign LUT_4[23425] = 32'b11111111111111111100111101110010;
assign LUT_4[23426] = 32'b00000000000000000011001100011110;
assign LUT_4[23427] = 32'b11111111111111111100011000010110;
assign LUT_4[23428] = 32'b00000000000000000000110010010110;
assign LUT_4[23429] = 32'b11111111111111111001111110001110;
assign LUT_4[23430] = 32'b00000000000000000000001100111010;
assign LUT_4[23431] = 32'b11111111111111111001011000110010;
assign LUT_4[23432] = 32'b11111111111111111100111110001111;
assign LUT_4[23433] = 32'b11111111111111110110001010000111;
assign LUT_4[23434] = 32'b11111111111111111100011000110011;
assign LUT_4[23435] = 32'b11111111111111110101100100101011;
assign LUT_4[23436] = 32'b11111111111111111001111110101011;
assign LUT_4[23437] = 32'b11111111111111110011001010100011;
assign LUT_4[23438] = 32'b11111111111111111001011001001111;
assign LUT_4[23439] = 32'b11111111111111110010100101000111;
assign LUT_4[23440] = 32'b00000000000000000001100011101000;
assign LUT_4[23441] = 32'b11111111111111111010101111100000;
assign LUT_4[23442] = 32'b00000000000000000000111110001100;
assign LUT_4[23443] = 32'b11111111111111111010001010000100;
assign LUT_4[23444] = 32'b11111111111111111110100100000100;
assign LUT_4[23445] = 32'b11111111111111110111101111111100;
assign LUT_4[23446] = 32'b11111111111111111101111110101000;
assign LUT_4[23447] = 32'b11111111111111110111001010100000;
assign LUT_4[23448] = 32'b11111111111111111010101111111101;
assign LUT_4[23449] = 32'b11111111111111110011111011110101;
assign LUT_4[23450] = 32'b11111111111111111010001010100001;
assign LUT_4[23451] = 32'b11111111111111110011010110011001;
assign LUT_4[23452] = 32'b11111111111111110111110000011001;
assign LUT_4[23453] = 32'b11111111111111110000111100010001;
assign LUT_4[23454] = 32'b11111111111111110111001010111101;
assign LUT_4[23455] = 32'b11111111111111110000010110110101;
assign LUT_4[23456] = 32'b00000000000000000010001101000001;
assign LUT_4[23457] = 32'b11111111111111111011011000111001;
assign LUT_4[23458] = 32'b00000000000000000001100111100101;
assign LUT_4[23459] = 32'b11111111111111111010110011011101;
assign LUT_4[23460] = 32'b11111111111111111111001101011101;
assign LUT_4[23461] = 32'b11111111111111111000011001010101;
assign LUT_4[23462] = 32'b11111111111111111110101000000001;
assign LUT_4[23463] = 32'b11111111111111110111110011111001;
assign LUT_4[23464] = 32'b11111111111111111011011001010110;
assign LUT_4[23465] = 32'b11111111111111110100100101001110;
assign LUT_4[23466] = 32'b11111111111111111010110011111010;
assign LUT_4[23467] = 32'b11111111111111110011111111110010;
assign LUT_4[23468] = 32'b11111111111111111000011001110010;
assign LUT_4[23469] = 32'b11111111111111110001100101101010;
assign LUT_4[23470] = 32'b11111111111111110111110100010110;
assign LUT_4[23471] = 32'b11111111111111110001000000001110;
assign LUT_4[23472] = 32'b11111111111111111111111110101111;
assign LUT_4[23473] = 32'b11111111111111111001001010100111;
assign LUT_4[23474] = 32'b11111111111111111111011001010011;
assign LUT_4[23475] = 32'b11111111111111111000100101001011;
assign LUT_4[23476] = 32'b11111111111111111100111111001011;
assign LUT_4[23477] = 32'b11111111111111110110001011000011;
assign LUT_4[23478] = 32'b11111111111111111100011001101111;
assign LUT_4[23479] = 32'b11111111111111110101100101100111;
assign LUT_4[23480] = 32'b11111111111111111001001011000100;
assign LUT_4[23481] = 32'b11111111111111110010010110111100;
assign LUT_4[23482] = 32'b11111111111111111000100101101000;
assign LUT_4[23483] = 32'b11111111111111110001110001100000;
assign LUT_4[23484] = 32'b11111111111111110110001011100000;
assign LUT_4[23485] = 32'b11111111111111101111010111011000;
assign LUT_4[23486] = 32'b11111111111111110101100110000100;
assign LUT_4[23487] = 32'b11111111111111101110110001111100;
assign LUT_4[23488] = 32'b00000000000000000101001001001110;
assign LUT_4[23489] = 32'b11111111111111111110010101000110;
assign LUT_4[23490] = 32'b00000000000000000100100011110010;
assign LUT_4[23491] = 32'b11111111111111111101101111101010;
assign LUT_4[23492] = 32'b00000000000000000010001001101010;
assign LUT_4[23493] = 32'b11111111111111111011010101100010;
assign LUT_4[23494] = 32'b00000000000000000001100100001110;
assign LUT_4[23495] = 32'b11111111111111111010110000000110;
assign LUT_4[23496] = 32'b11111111111111111110010101100011;
assign LUT_4[23497] = 32'b11111111111111110111100001011011;
assign LUT_4[23498] = 32'b11111111111111111101110000000111;
assign LUT_4[23499] = 32'b11111111111111110110111011111111;
assign LUT_4[23500] = 32'b11111111111111111011010101111111;
assign LUT_4[23501] = 32'b11111111111111110100100001110111;
assign LUT_4[23502] = 32'b11111111111111111010110000100011;
assign LUT_4[23503] = 32'b11111111111111110011111100011011;
assign LUT_4[23504] = 32'b00000000000000000010111010111100;
assign LUT_4[23505] = 32'b11111111111111111100000110110100;
assign LUT_4[23506] = 32'b00000000000000000010010101100000;
assign LUT_4[23507] = 32'b11111111111111111011100001011000;
assign LUT_4[23508] = 32'b11111111111111111111111011011000;
assign LUT_4[23509] = 32'b11111111111111111001000111010000;
assign LUT_4[23510] = 32'b11111111111111111111010101111100;
assign LUT_4[23511] = 32'b11111111111111111000100001110100;
assign LUT_4[23512] = 32'b11111111111111111100000111010001;
assign LUT_4[23513] = 32'b11111111111111110101010011001001;
assign LUT_4[23514] = 32'b11111111111111111011100001110101;
assign LUT_4[23515] = 32'b11111111111111110100101101101101;
assign LUT_4[23516] = 32'b11111111111111111001000111101101;
assign LUT_4[23517] = 32'b11111111111111110010010011100101;
assign LUT_4[23518] = 32'b11111111111111111000100010010001;
assign LUT_4[23519] = 32'b11111111111111110001101110001001;
assign LUT_4[23520] = 32'b00000000000000000011100100010101;
assign LUT_4[23521] = 32'b11111111111111111100110000001101;
assign LUT_4[23522] = 32'b00000000000000000010111110111001;
assign LUT_4[23523] = 32'b11111111111111111100001010110001;
assign LUT_4[23524] = 32'b00000000000000000000100100110001;
assign LUT_4[23525] = 32'b11111111111111111001110000101001;
assign LUT_4[23526] = 32'b11111111111111111111111111010101;
assign LUT_4[23527] = 32'b11111111111111111001001011001101;
assign LUT_4[23528] = 32'b11111111111111111100110000101010;
assign LUT_4[23529] = 32'b11111111111111110101111100100010;
assign LUT_4[23530] = 32'b11111111111111111100001011001110;
assign LUT_4[23531] = 32'b11111111111111110101010111000110;
assign LUT_4[23532] = 32'b11111111111111111001110001000110;
assign LUT_4[23533] = 32'b11111111111111110010111100111110;
assign LUT_4[23534] = 32'b11111111111111111001001011101010;
assign LUT_4[23535] = 32'b11111111111111110010010111100010;
assign LUT_4[23536] = 32'b00000000000000000001010110000011;
assign LUT_4[23537] = 32'b11111111111111111010100001111011;
assign LUT_4[23538] = 32'b00000000000000000000110000100111;
assign LUT_4[23539] = 32'b11111111111111111001111100011111;
assign LUT_4[23540] = 32'b11111111111111111110010110011111;
assign LUT_4[23541] = 32'b11111111111111110111100010010111;
assign LUT_4[23542] = 32'b11111111111111111101110001000011;
assign LUT_4[23543] = 32'b11111111111111110110111100111011;
assign LUT_4[23544] = 32'b11111111111111111010100010011000;
assign LUT_4[23545] = 32'b11111111111111110011101110010000;
assign LUT_4[23546] = 32'b11111111111111111001111100111100;
assign LUT_4[23547] = 32'b11111111111111110011001000110100;
assign LUT_4[23548] = 32'b11111111111111110111100010110100;
assign LUT_4[23549] = 32'b11111111111111110000101110101100;
assign LUT_4[23550] = 32'b11111111111111110110111101011000;
assign LUT_4[23551] = 32'b11111111111111110000001001010000;
assign LUT_4[23552] = 32'b11111111111111111110110110100110;
assign LUT_4[23553] = 32'b11111111111111111000000010011110;
assign LUT_4[23554] = 32'b11111111111111111110010001001010;
assign LUT_4[23555] = 32'b11111111111111110111011101000010;
assign LUT_4[23556] = 32'b11111111111111111011110111000010;
assign LUT_4[23557] = 32'b11111111111111110101000010111010;
assign LUT_4[23558] = 32'b11111111111111111011010001100110;
assign LUT_4[23559] = 32'b11111111111111110100011101011110;
assign LUT_4[23560] = 32'b11111111111111111000000010111011;
assign LUT_4[23561] = 32'b11111111111111110001001110110011;
assign LUT_4[23562] = 32'b11111111111111110111011101011111;
assign LUT_4[23563] = 32'b11111111111111110000101001010111;
assign LUT_4[23564] = 32'b11111111111111110101000011010111;
assign LUT_4[23565] = 32'b11111111111111101110001111001111;
assign LUT_4[23566] = 32'b11111111111111110100011101111011;
assign LUT_4[23567] = 32'b11111111111111101101101001110011;
assign LUT_4[23568] = 32'b11111111111111111100101000010100;
assign LUT_4[23569] = 32'b11111111111111110101110100001100;
assign LUT_4[23570] = 32'b11111111111111111100000010111000;
assign LUT_4[23571] = 32'b11111111111111110101001110110000;
assign LUT_4[23572] = 32'b11111111111111111001101000110000;
assign LUT_4[23573] = 32'b11111111111111110010110100101000;
assign LUT_4[23574] = 32'b11111111111111111001000011010100;
assign LUT_4[23575] = 32'b11111111111111110010001111001100;
assign LUT_4[23576] = 32'b11111111111111110101110100101001;
assign LUT_4[23577] = 32'b11111111111111101111000000100001;
assign LUT_4[23578] = 32'b11111111111111110101001111001101;
assign LUT_4[23579] = 32'b11111111111111101110011011000101;
assign LUT_4[23580] = 32'b11111111111111110010110101000101;
assign LUT_4[23581] = 32'b11111111111111101100000000111101;
assign LUT_4[23582] = 32'b11111111111111110010001111101001;
assign LUT_4[23583] = 32'b11111111111111101011011011100001;
assign LUT_4[23584] = 32'b11111111111111111101010001101101;
assign LUT_4[23585] = 32'b11111111111111110110011101100101;
assign LUT_4[23586] = 32'b11111111111111111100101100010001;
assign LUT_4[23587] = 32'b11111111111111110101111000001001;
assign LUT_4[23588] = 32'b11111111111111111010010010001001;
assign LUT_4[23589] = 32'b11111111111111110011011110000001;
assign LUT_4[23590] = 32'b11111111111111111001101100101101;
assign LUT_4[23591] = 32'b11111111111111110010111000100101;
assign LUT_4[23592] = 32'b11111111111111110110011110000010;
assign LUT_4[23593] = 32'b11111111111111101111101001111010;
assign LUT_4[23594] = 32'b11111111111111110101111000100110;
assign LUT_4[23595] = 32'b11111111111111101111000100011110;
assign LUT_4[23596] = 32'b11111111111111110011011110011110;
assign LUT_4[23597] = 32'b11111111111111101100101010010110;
assign LUT_4[23598] = 32'b11111111111111110010111001000010;
assign LUT_4[23599] = 32'b11111111111111101100000100111010;
assign LUT_4[23600] = 32'b11111111111111111011000011011011;
assign LUT_4[23601] = 32'b11111111111111110100001111010011;
assign LUT_4[23602] = 32'b11111111111111111010011101111111;
assign LUT_4[23603] = 32'b11111111111111110011101001110111;
assign LUT_4[23604] = 32'b11111111111111111000000011110111;
assign LUT_4[23605] = 32'b11111111111111110001001111101111;
assign LUT_4[23606] = 32'b11111111111111110111011110011011;
assign LUT_4[23607] = 32'b11111111111111110000101010010011;
assign LUT_4[23608] = 32'b11111111111111110100001111110000;
assign LUT_4[23609] = 32'b11111111111111101101011011101000;
assign LUT_4[23610] = 32'b11111111111111110011101010010100;
assign LUT_4[23611] = 32'b11111111111111101100110110001100;
assign LUT_4[23612] = 32'b11111111111111110001010000001100;
assign LUT_4[23613] = 32'b11111111111111101010011100000100;
assign LUT_4[23614] = 32'b11111111111111110000101010110000;
assign LUT_4[23615] = 32'b11111111111111101001110110101000;
assign LUT_4[23616] = 32'b00000000000000000000001101111010;
assign LUT_4[23617] = 32'b11111111111111111001011001110010;
assign LUT_4[23618] = 32'b11111111111111111111101000011110;
assign LUT_4[23619] = 32'b11111111111111111000110100010110;
assign LUT_4[23620] = 32'b11111111111111111101001110010110;
assign LUT_4[23621] = 32'b11111111111111110110011010001110;
assign LUT_4[23622] = 32'b11111111111111111100101000111010;
assign LUT_4[23623] = 32'b11111111111111110101110100110010;
assign LUT_4[23624] = 32'b11111111111111111001011010001111;
assign LUT_4[23625] = 32'b11111111111111110010100110000111;
assign LUT_4[23626] = 32'b11111111111111111000110100110011;
assign LUT_4[23627] = 32'b11111111111111110010000000101011;
assign LUT_4[23628] = 32'b11111111111111110110011010101011;
assign LUT_4[23629] = 32'b11111111111111101111100110100011;
assign LUT_4[23630] = 32'b11111111111111110101110101001111;
assign LUT_4[23631] = 32'b11111111111111101111000001000111;
assign LUT_4[23632] = 32'b11111111111111111101111111101000;
assign LUT_4[23633] = 32'b11111111111111110111001011100000;
assign LUT_4[23634] = 32'b11111111111111111101011010001100;
assign LUT_4[23635] = 32'b11111111111111110110100110000100;
assign LUT_4[23636] = 32'b11111111111111111011000000000100;
assign LUT_4[23637] = 32'b11111111111111110100001011111100;
assign LUT_4[23638] = 32'b11111111111111111010011010101000;
assign LUT_4[23639] = 32'b11111111111111110011100110100000;
assign LUT_4[23640] = 32'b11111111111111110111001011111101;
assign LUT_4[23641] = 32'b11111111111111110000010111110101;
assign LUT_4[23642] = 32'b11111111111111110110100110100001;
assign LUT_4[23643] = 32'b11111111111111101111110010011001;
assign LUT_4[23644] = 32'b11111111111111110100001100011001;
assign LUT_4[23645] = 32'b11111111111111101101011000010001;
assign LUT_4[23646] = 32'b11111111111111110011100110111101;
assign LUT_4[23647] = 32'b11111111111111101100110010110101;
assign LUT_4[23648] = 32'b11111111111111111110101001000001;
assign LUT_4[23649] = 32'b11111111111111110111110100111001;
assign LUT_4[23650] = 32'b11111111111111111110000011100101;
assign LUT_4[23651] = 32'b11111111111111110111001111011101;
assign LUT_4[23652] = 32'b11111111111111111011101001011101;
assign LUT_4[23653] = 32'b11111111111111110100110101010101;
assign LUT_4[23654] = 32'b11111111111111111011000100000001;
assign LUT_4[23655] = 32'b11111111111111110100001111111001;
assign LUT_4[23656] = 32'b11111111111111110111110101010110;
assign LUT_4[23657] = 32'b11111111111111110001000001001110;
assign LUT_4[23658] = 32'b11111111111111110111001111111010;
assign LUT_4[23659] = 32'b11111111111111110000011011110010;
assign LUT_4[23660] = 32'b11111111111111110100110101110010;
assign LUT_4[23661] = 32'b11111111111111101110000001101010;
assign LUT_4[23662] = 32'b11111111111111110100010000010110;
assign LUT_4[23663] = 32'b11111111111111101101011100001110;
assign LUT_4[23664] = 32'b11111111111111111100011010101111;
assign LUT_4[23665] = 32'b11111111111111110101100110100111;
assign LUT_4[23666] = 32'b11111111111111111011110101010011;
assign LUT_4[23667] = 32'b11111111111111110101000001001011;
assign LUT_4[23668] = 32'b11111111111111111001011011001011;
assign LUT_4[23669] = 32'b11111111111111110010100111000011;
assign LUT_4[23670] = 32'b11111111111111111000110101101111;
assign LUT_4[23671] = 32'b11111111111111110010000001100111;
assign LUT_4[23672] = 32'b11111111111111110101100111000100;
assign LUT_4[23673] = 32'b11111111111111101110110010111100;
assign LUT_4[23674] = 32'b11111111111111110101000001101000;
assign LUT_4[23675] = 32'b11111111111111101110001101100000;
assign LUT_4[23676] = 32'b11111111111111110010100111100000;
assign LUT_4[23677] = 32'b11111111111111101011110011011000;
assign LUT_4[23678] = 32'b11111111111111110010000010000100;
assign LUT_4[23679] = 32'b11111111111111101011001101111100;
assign LUT_4[23680] = 32'b00000000000000000001011100101110;
assign LUT_4[23681] = 32'b11111111111111111010101000100110;
assign LUT_4[23682] = 32'b00000000000000000000110111010010;
assign LUT_4[23683] = 32'b11111111111111111010000011001010;
assign LUT_4[23684] = 32'b11111111111111111110011101001010;
assign LUT_4[23685] = 32'b11111111111111110111101001000010;
assign LUT_4[23686] = 32'b11111111111111111101110111101110;
assign LUT_4[23687] = 32'b11111111111111110111000011100110;
assign LUT_4[23688] = 32'b11111111111111111010101001000011;
assign LUT_4[23689] = 32'b11111111111111110011110100111011;
assign LUT_4[23690] = 32'b11111111111111111010000011100111;
assign LUT_4[23691] = 32'b11111111111111110011001111011111;
assign LUT_4[23692] = 32'b11111111111111110111101001011111;
assign LUT_4[23693] = 32'b11111111111111110000110101010111;
assign LUT_4[23694] = 32'b11111111111111110111000100000011;
assign LUT_4[23695] = 32'b11111111111111110000001111111011;
assign LUT_4[23696] = 32'b11111111111111111111001110011100;
assign LUT_4[23697] = 32'b11111111111111111000011010010100;
assign LUT_4[23698] = 32'b11111111111111111110101001000000;
assign LUT_4[23699] = 32'b11111111111111110111110100111000;
assign LUT_4[23700] = 32'b11111111111111111100001110111000;
assign LUT_4[23701] = 32'b11111111111111110101011010110000;
assign LUT_4[23702] = 32'b11111111111111111011101001011100;
assign LUT_4[23703] = 32'b11111111111111110100110101010100;
assign LUT_4[23704] = 32'b11111111111111111000011010110001;
assign LUT_4[23705] = 32'b11111111111111110001100110101001;
assign LUT_4[23706] = 32'b11111111111111110111110101010101;
assign LUT_4[23707] = 32'b11111111111111110001000001001101;
assign LUT_4[23708] = 32'b11111111111111110101011011001101;
assign LUT_4[23709] = 32'b11111111111111101110100111000101;
assign LUT_4[23710] = 32'b11111111111111110100110101110001;
assign LUT_4[23711] = 32'b11111111111111101110000001101001;
assign LUT_4[23712] = 32'b11111111111111111111110111110101;
assign LUT_4[23713] = 32'b11111111111111111001000011101101;
assign LUT_4[23714] = 32'b11111111111111111111010010011001;
assign LUT_4[23715] = 32'b11111111111111111000011110010001;
assign LUT_4[23716] = 32'b11111111111111111100111000010001;
assign LUT_4[23717] = 32'b11111111111111110110000100001001;
assign LUT_4[23718] = 32'b11111111111111111100010010110101;
assign LUT_4[23719] = 32'b11111111111111110101011110101101;
assign LUT_4[23720] = 32'b11111111111111111001000100001010;
assign LUT_4[23721] = 32'b11111111111111110010010000000010;
assign LUT_4[23722] = 32'b11111111111111111000011110101110;
assign LUT_4[23723] = 32'b11111111111111110001101010100110;
assign LUT_4[23724] = 32'b11111111111111110110000100100110;
assign LUT_4[23725] = 32'b11111111111111101111010000011110;
assign LUT_4[23726] = 32'b11111111111111110101011111001010;
assign LUT_4[23727] = 32'b11111111111111101110101011000010;
assign LUT_4[23728] = 32'b11111111111111111101101001100011;
assign LUT_4[23729] = 32'b11111111111111110110110101011011;
assign LUT_4[23730] = 32'b11111111111111111101000100000111;
assign LUT_4[23731] = 32'b11111111111111110110001111111111;
assign LUT_4[23732] = 32'b11111111111111111010101001111111;
assign LUT_4[23733] = 32'b11111111111111110011110101110111;
assign LUT_4[23734] = 32'b11111111111111111010000100100011;
assign LUT_4[23735] = 32'b11111111111111110011010000011011;
assign LUT_4[23736] = 32'b11111111111111110110110101111000;
assign LUT_4[23737] = 32'b11111111111111110000000001110000;
assign LUT_4[23738] = 32'b11111111111111110110010000011100;
assign LUT_4[23739] = 32'b11111111111111101111011100010100;
assign LUT_4[23740] = 32'b11111111111111110011110110010100;
assign LUT_4[23741] = 32'b11111111111111101101000010001100;
assign LUT_4[23742] = 32'b11111111111111110011010000111000;
assign LUT_4[23743] = 32'b11111111111111101100011100110000;
assign LUT_4[23744] = 32'b00000000000000000010110100000010;
assign LUT_4[23745] = 32'b11111111111111111011111111111010;
assign LUT_4[23746] = 32'b00000000000000000010001110100110;
assign LUT_4[23747] = 32'b11111111111111111011011010011110;
assign LUT_4[23748] = 32'b11111111111111111111110100011110;
assign LUT_4[23749] = 32'b11111111111111111001000000010110;
assign LUT_4[23750] = 32'b11111111111111111111001111000010;
assign LUT_4[23751] = 32'b11111111111111111000011010111010;
assign LUT_4[23752] = 32'b11111111111111111100000000010111;
assign LUT_4[23753] = 32'b11111111111111110101001100001111;
assign LUT_4[23754] = 32'b11111111111111111011011010111011;
assign LUT_4[23755] = 32'b11111111111111110100100110110011;
assign LUT_4[23756] = 32'b11111111111111111001000000110011;
assign LUT_4[23757] = 32'b11111111111111110010001100101011;
assign LUT_4[23758] = 32'b11111111111111111000011011010111;
assign LUT_4[23759] = 32'b11111111111111110001100111001111;
assign LUT_4[23760] = 32'b00000000000000000000100101110000;
assign LUT_4[23761] = 32'b11111111111111111001110001101000;
assign LUT_4[23762] = 32'b00000000000000000000000000010100;
assign LUT_4[23763] = 32'b11111111111111111001001100001100;
assign LUT_4[23764] = 32'b11111111111111111101100110001100;
assign LUT_4[23765] = 32'b11111111111111110110110010000100;
assign LUT_4[23766] = 32'b11111111111111111101000000110000;
assign LUT_4[23767] = 32'b11111111111111110110001100101000;
assign LUT_4[23768] = 32'b11111111111111111001110010000101;
assign LUT_4[23769] = 32'b11111111111111110010111101111101;
assign LUT_4[23770] = 32'b11111111111111111001001100101001;
assign LUT_4[23771] = 32'b11111111111111110010011000100001;
assign LUT_4[23772] = 32'b11111111111111110110110010100001;
assign LUT_4[23773] = 32'b11111111111111101111111110011001;
assign LUT_4[23774] = 32'b11111111111111110110001101000101;
assign LUT_4[23775] = 32'b11111111111111101111011000111101;
assign LUT_4[23776] = 32'b00000000000000000001001111001001;
assign LUT_4[23777] = 32'b11111111111111111010011011000001;
assign LUT_4[23778] = 32'b00000000000000000000101001101101;
assign LUT_4[23779] = 32'b11111111111111111001110101100101;
assign LUT_4[23780] = 32'b11111111111111111110001111100101;
assign LUT_4[23781] = 32'b11111111111111110111011011011101;
assign LUT_4[23782] = 32'b11111111111111111101101010001001;
assign LUT_4[23783] = 32'b11111111111111110110110110000001;
assign LUT_4[23784] = 32'b11111111111111111010011011011110;
assign LUT_4[23785] = 32'b11111111111111110011100111010110;
assign LUT_4[23786] = 32'b11111111111111111001110110000010;
assign LUT_4[23787] = 32'b11111111111111110011000001111010;
assign LUT_4[23788] = 32'b11111111111111110111011011111010;
assign LUT_4[23789] = 32'b11111111111111110000100111110010;
assign LUT_4[23790] = 32'b11111111111111110110110110011110;
assign LUT_4[23791] = 32'b11111111111111110000000010010110;
assign LUT_4[23792] = 32'b11111111111111111111000000110111;
assign LUT_4[23793] = 32'b11111111111111111000001100101111;
assign LUT_4[23794] = 32'b11111111111111111110011011011011;
assign LUT_4[23795] = 32'b11111111111111110111100111010011;
assign LUT_4[23796] = 32'b11111111111111111100000001010011;
assign LUT_4[23797] = 32'b11111111111111110101001101001011;
assign LUT_4[23798] = 32'b11111111111111111011011011110111;
assign LUT_4[23799] = 32'b11111111111111110100100111101111;
assign LUT_4[23800] = 32'b11111111111111111000001101001100;
assign LUT_4[23801] = 32'b11111111111111110001011001000100;
assign LUT_4[23802] = 32'b11111111111111110111100111110000;
assign LUT_4[23803] = 32'b11111111111111110000110011101000;
assign LUT_4[23804] = 32'b11111111111111110101001101101000;
assign LUT_4[23805] = 32'b11111111111111101110011001100000;
assign LUT_4[23806] = 32'b11111111111111110100101000001100;
assign LUT_4[23807] = 32'b11111111111111101101110100000100;
assign LUT_4[23808] = 32'b00000000000000000011110010001001;
assign LUT_4[23809] = 32'b11111111111111111100111110000001;
assign LUT_4[23810] = 32'b00000000000000000011001100101101;
assign LUT_4[23811] = 32'b11111111111111111100011000100101;
assign LUT_4[23812] = 32'b00000000000000000000110010100101;
assign LUT_4[23813] = 32'b11111111111111111001111110011101;
assign LUT_4[23814] = 32'b00000000000000000000001101001001;
assign LUT_4[23815] = 32'b11111111111111111001011001000001;
assign LUT_4[23816] = 32'b11111111111111111100111110011110;
assign LUT_4[23817] = 32'b11111111111111110110001010010110;
assign LUT_4[23818] = 32'b11111111111111111100011001000010;
assign LUT_4[23819] = 32'b11111111111111110101100100111010;
assign LUT_4[23820] = 32'b11111111111111111001111110111010;
assign LUT_4[23821] = 32'b11111111111111110011001010110010;
assign LUT_4[23822] = 32'b11111111111111111001011001011110;
assign LUT_4[23823] = 32'b11111111111111110010100101010110;
assign LUT_4[23824] = 32'b00000000000000000001100011110111;
assign LUT_4[23825] = 32'b11111111111111111010101111101111;
assign LUT_4[23826] = 32'b00000000000000000000111110011011;
assign LUT_4[23827] = 32'b11111111111111111010001010010011;
assign LUT_4[23828] = 32'b11111111111111111110100100010011;
assign LUT_4[23829] = 32'b11111111111111110111110000001011;
assign LUT_4[23830] = 32'b11111111111111111101111110110111;
assign LUT_4[23831] = 32'b11111111111111110111001010101111;
assign LUT_4[23832] = 32'b11111111111111111010110000001100;
assign LUT_4[23833] = 32'b11111111111111110011111100000100;
assign LUT_4[23834] = 32'b11111111111111111010001010110000;
assign LUT_4[23835] = 32'b11111111111111110011010110101000;
assign LUT_4[23836] = 32'b11111111111111110111110000101000;
assign LUT_4[23837] = 32'b11111111111111110000111100100000;
assign LUT_4[23838] = 32'b11111111111111110111001011001100;
assign LUT_4[23839] = 32'b11111111111111110000010111000100;
assign LUT_4[23840] = 32'b00000000000000000010001101010000;
assign LUT_4[23841] = 32'b11111111111111111011011001001000;
assign LUT_4[23842] = 32'b00000000000000000001100111110100;
assign LUT_4[23843] = 32'b11111111111111111010110011101100;
assign LUT_4[23844] = 32'b11111111111111111111001101101100;
assign LUT_4[23845] = 32'b11111111111111111000011001100100;
assign LUT_4[23846] = 32'b11111111111111111110101000010000;
assign LUT_4[23847] = 32'b11111111111111110111110100001000;
assign LUT_4[23848] = 32'b11111111111111111011011001100101;
assign LUT_4[23849] = 32'b11111111111111110100100101011101;
assign LUT_4[23850] = 32'b11111111111111111010110100001001;
assign LUT_4[23851] = 32'b11111111111111110100000000000001;
assign LUT_4[23852] = 32'b11111111111111111000011010000001;
assign LUT_4[23853] = 32'b11111111111111110001100101111001;
assign LUT_4[23854] = 32'b11111111111111110111110100100101;
assign LUT_4[23855] = 32'b11111111111111110001000000011101;
assign LUT_4[23856] = 32'b11111111111111111111111110111110;
assign LUT_4[23857] = 32'b11111111111111111001001010110110;
assign LUT_4[23858] = 32'b11111111111111111111011001100010;
assign LUT_4[23859] = 32'b11111111111111111000100101011010;
assign LUT_4[23860] = 32'b11111111111111111100111111011010;
assign LUT_4[23861] = 32'b11111111111111110110001011010010;
assign LUT_4[23862] = 32'b11111111111111111100011001111110;
assign LUT_4[23863] = 32'b11111111111111110101100101110110;
assign LUT_4[23864] = 32'b11111111111111111001001011010011;
assign LUT_4[23865] = 32'b11111111111111110010010111001011;
assign LUT_4[23866] = 32'b11111111111111111000100101110111;
assign LUT_4[23867] = 32'b11111111111111110001110001101111;
assign LUT_4[23868] = 32'b11111111111111110110001011101111;
assign LUT_4[23869] = 32'b11111111111111101111010111100111;
assign LUT_4[23870] = 32'b11111111111111110101100110010011;
assign LUT_4[23871] = 32'b11111111111111101110110010001011;
assign LUT_4[23872] = 32'b00000000000000000101001001011101;
assign LUT_4[23873] = 32'b11111111111111111110010101010101;
assign LUT_4[23874] = 32'b00000000000000000100100100000001;
assign LUT_4[23875] = 32'b11111111111111111101101111111001;
assign LUT_4[23876] = 32'b00000000000000000010001001111001;
assign LUT_4[23877] = 32'b11111111111111111011010101110001;
assign LUT_4[23878] = 32'b00000000000000000001100100011101;
assign LUT_4[23879] = 32'b11111111111111111010110000010101;
assign LUT_4[23880] = 32'b11111111111111111110010101110010;
assign LUT_4[23881] = 32'b11111111111111110111100001101010;
assign LUT_4[23882] = 32'b11111111111111111101110000010110;
assign LUT_4[23883] = 32'b11111111111111110110111100001110;
assign LUT_4[23884] = 32'b11111111111111111011010110001110;
assign LUT_4[23885] = 32'b11111111111111110100100010000110;
assign LUT_4[23886] = 32'b11111111111111111010110000110010;
assign LUT_4[23887] = 32'b11111111111111110011111100101010;
assign LUT_4[23888] = 32'b00000000000000000010111011001011;
assign LUT_4[23889] = 32'b11111111111111111100000111000011;
assign LUT_4[23890] = 32'b00000000000000000010010101101111;
assign LUT_4[23891] = 32'b11111111111111111011100001100111;
assign LUT_4[23892] = 32'b11111111111111111111111011100111;
assign LUT_4[23893] = 32'b11111111111111111001000111011111;
assign LUT_4[23894] = 32'b11111111111111111111010110001011;
assign LUT_4[23895] = 32'b11111111111111111000100010000011;
assign LUT_4[23896] = 32'b11111111111111111100000111100000;
assign LUT_4[23897] = 32'b11111111111111110101010011011000;
assign LUT_4[23898] = 32'b11111111111111111011100010000100;
assign LUT_4[23899] = 32'b11111111111111110100101101111100;
assign LUT_4[23900] = 32'b11111111111111111001000111111100;
assign LUT_4[23901] = 32'b11111111111111110010010011110100;
assign LUT_4[23902] = 32'b11111111111111111000100010100000;
assign LUT_4[23903] = 32'b11111111111111110001101110011000;
assign LUT_4[23904] = 32'b00000000000000000011100100100100;
assign LUT_4[23905] = 32'b11111111111111111100110000011100;
assign LUT_4[23906] = 32'b00000000000000000010111111001000;
assign LUT_4[23907] = 32'b11111111111111111100001011000000;
assign LUT_4[23908] = 32'b00000000000000000000100101000000;
assign LUT_4[23909] = 32'b11111111111111111001110000111000;
assign LUT_4[23910] = 32'b11111111111111111111111111100100;
assign LUT_4[23911] = 32'b11111111111111111001001011011100;
assign LUT_4[23912] = 32'b11111111111111111100110000111001;
assign LUT_4[23913] = 32'b11111111111111110101111100110001;
assign LUT_4[23914] = 32'b11111111111111111100001011011101;
assign LUT_4[23915] = 32'b11111111111111110101010111010101;
assign LUT_4[23916] = 32'b11111111111111111001110001010101;
assign LUT_4[23917] = 32'b11111111111111110010111101001101;
assign LUT_4[23918] = 32'b11111111111111111001001011111001;
assign LUT_4[23919] = 32'b11111111111111110010010111110001;
assign LUT_4[23920] = 32'b00000000000000000001010110010010;
assign LUT_4[23921] = 32'b11111111111111111010100010001010;
assign LUT_4[23922] = 32'b00000000000000000000110000110110;
assign LUT_4[23923] = 32'b11111111111111111001111100101110;
assign LUT_4[23924] = 32'b11111111111111111110010110101110;
assign LUT_4[23925] = 32'b11111111111111110111100010100110;
assign LUT_4[23926] = 32'b11111111111111111101110001010010;
assign LUT_4[23927] = 32'b11111111111111110110111101001010;
assign LUT_4[23928] = 32'b11111111111111111010100010100111;
assign LUT_4[23929] = 32'b11111111111111110011101110011111;
assign LUT_4[23930] = 32'b11111111111111111001111101001011;
assign LUT_4[23931] = 32'b11111111111111110011001001000011;
assign LUT_4[23932] = 32'b11111111111111110111100011000011;
assign LUT_4[23933] = 32'b11111111111111110000101110111011;
assign LUT_4[23934] = 32'b11111111111111110110111101100111;
assign LUT_4[23935] = 32'b11111111111111110000001001011111;
assign LUT_4[23936] = 32'b00000000000000000110011000010001;
assign LUT_4[23937] = 32'b11111111111111111111100100001001;
assign LUT_4[23938] = 32'b00000000000000000101110010110101;
assign LUT_4[23939] = 32'b11111111111111111110111110101101;
assign LUT_4[23940] = 32'b00000000000000000011011000101101;
assign LUT_4[23941] = 32'b11111111111111111100100100100101;
assign LUT_4[23942] = 32'b00000000000000000010110011010001;
assign LUT_4[23943] = 32'b11111111111111111011111111001001;
assign LUT_4[23944] = 32'b11111111111111111111100100100110;
assign LUT_4[23945] = 32'b11111111111111111000110000011110;
assign LUT_4[23946] = 32'b11111111111111111110111111001010;
assign LUT_4[23947] = 32'b11111111111111111000001011000010;
assign LUT_4[23948] = 32'b11111111111111111100100101000010;
assign LUT_4[23949] = 32'b11111111111111110101110000111010;
assign LUT_4[23950] = 32'b11111111111111111011111111100110;
assign LUT_4[23951] = 32'b11111111111111110101001011011110;
assign LUT_4[23952] = 32'b00000000000000000100001001111111;
assign LUT_4[23953] = 32'b11111111111111111101010101110111;
assign LUT_4[23954] = 32'b00000000000000000011100100100011;
assign LUT_4[23955] = 32'b11111111111111111100110000011011;
assign LUT_4[23956] = 32'b00000000000000000001001010011011;
assign LUT_4[23957] = 32'b11111111111111111010010110010011;
assign LUT_4[23958] = 32'b00000000000000000000100100111111;
assign LUT_4[23959] = 32'b11111111111111111001110000110111;
assign LUT_4[23960] = 32'b11111111111111111101010110010100;
assign LUT_4[23961] = 32'b11111111111111110110100010001100;
assign LUT_4[23962] = 32'b11111111111111111100110000111000;
assign LUT_4[23963] = 32'b11111111111111110101111100110000;
assign LUT_4[23964] = 32'b11111111111111111010010110110000;
assign LUT_4[23965] = 32'b11111111111111110011100010101000;
assign LUT_4[23966] = 32'b11111111111111111001110001010100;
assign LUT_4[23967] = 32'b11111111111111110010111101001100;
assign LUT_4[23968] = 32'b00000000000000000100110011011000;
assign LUT_4[23969] = 32'b11111111111111111101111111010000;
assign LUT_4[23970] = 32'b00000000000000000100001101111100;
assign LUT_4[23971] = 32'b11111111111111111101011001110100;
assign LUT_4[23972] = 32'b00000000000000000001110011110100;
assign LUT_4[23973] = 32'b11111111111111111010111111101100;
assign LUT_4[23974] = 32'b00000000000000000001001110011000;
assign LUT_4[23975] = 32'b11111111111111111010011010010000;
assign LUT_4[23976] = 32'b11111111111111111101111111101101;
assign LUT_4[23977] = 32'b11111111111111110111001011100101;
assign LUT_4[23978] = 32'b11111111111111111101011010010001;
assign LUT_4[23979] = 32'b11111111111111110110100110001001;
assign LUT_4[23980] = 32'b11111111111111111011000000001001;
assign LUT_4[23981] = 32'b11111111111111110100001100000001;
assign LUT_4[23982] = 32'b11111111111111111010011010101101;
assign LUT_4[23983] = 32'b11111111111111110011100110100101;
assign LUT_4[23984] = 32'b00000000000000000010100101000110;
assign LUT_4[23985] = 32'b11111111111111111011110000111110;
assign LUT_4[23986] = 32'b00000000000000000001111111101010;
assign LUT_4[23987] = 32'b11111111111111111011001011100010;
assign LUT_4[23988] = 32'b11111111111111111111100101100010;
assign LUT_4[23989] = 32'b11111111111111111000110001011010;
assign LUT_4[23990] = 32'b11111111111111111111000000000110;
assign LUT_4[23991] = 32'b11111111111111111000001011111110;
assign LUT_4[23992] = 32'b11111111111111111011110001011011;
assign LUT_4[23993] = 32'b11111111111111110100111101010011;
assign LUT_4[23994] = 32'b11111111111111111011001011111111;
assign LUT_4[23995] = 32'b11111111111111110100010111110111;
assign LUT_4[23996] = 32'b11111111111111111000110001110111;
assign LUT_4[23997] = 32'b11111111111111110001111101101111;
assign LUT_4[23998] = 32'b11111111111111111000001100011011;
assign LUT_4[23999] = 32'b11111111111111110001011000010011;
assign LUT_4[24000] = 32'b00000000000000000111101111100101;
assign LUT_4[24001] = 32'b00000000000000000000111011011101;
assign LUT_4[24002] = 32'b00000000000000000111001010001001;
assign LUT_4[24003] = 32'b00000000000000000000010110000001;
assign LUT_4[24004] = 32'b00000000000000000100110000000001;
assign LUT_4[24005] = 32'b11111111111111111101111011111001;
assign LUT_4[24006] = 32'b00000000000000000100001010100101;
assign LUT_4[24007] = 32'b11111111111111111101010110011101;
assign LUT_4[24008] = 32'b00000000000000000000111011111010;
assign LUT_4[24009] = 32'b11111111111111111010000111110010;
assign LUT_4[24010] = 32'b00000000000000000000010110011110;
assign LUT_4[24011] = 32'b11111111111111111001100010010110;
assign LUT_4[24012] = 32'b11111111111111111101111100010110;
assign LUT_4[24013] = 32'b11111111111111110111001000001110;
assign LUT_4[24014] = 32'b11111111111111111101010110111010;
assign LUT_4[24015] = 32'b11111111111111110110100010110010;
assign LUT_4[24016] = 32'b00000000000000000101100001010011;
assign LUT_4[24017] = 32'b11111111111111111110101101001011;
assign LUT_4[24018] = 32'b00000000000000000100111011110111;
assign LUT_4[24019] = 32'b11111111111111111110000111101111;
assign LUT_4[24020] = 32'b00000000000000000010100001101111;
assign LUT_4[24021] = 32'b11111111111111111011101101100111;
assign LUT_4[24022] = 32'b00000000000000000001111100010011;
assign LUT_4[24023] = 32'b11111111111111111011001000001011;
assign LUT_4[24024] = 32'b11111111111111111110101101101000;
assign LUT_4[24025] = 32'b11111111111111110111111001100000;
assign LUT_4[24026] = 32'b11111111111111111110001000001100;
assign LUT_4[24027] = 32'b11111111111111110111010100000100;
assign LUT_4[24028] = 32'b11111111111111111011101110000100;
assign LUT_4[24029] = 32'b11111111111111110100111001111100;
assign LUT_4[24030] = 32'b11111111111111111011001000101000;
assign LUT_4[24031] = 32'b11111111111111110100010100100000;
assign LUT_4[24032] = 32'b00000000000000000110001010101100;
assign LUT_4[24033] = 32'b11111111111111111111010110100100;
assign LUT_4[24034] = 32'b00000000000000000101100101010000;
assign LUT_4[24035] = 32'b11111111111111111110110001001000;
assign LUT_4[24036] = 32'b00000000000000000011001011001000;
assign LUT_4[24037] = 32'b11111111111111111100010111000000;
assign LUT_4[24038] = 32'b00000000000000000010100101101100;
assign LUT_4[24039] = 32'b11111111111111111011110001100100;
assign LUT_4[24040] = 32'b11111111111111111111010111000001;
assign LUT_4[24041] = 32'b11111111111111111000100010111001;
assign LUT_4[24042] = 32'b11111111111111111110110001100101;
assign LUT_4[24043] = 32'b11111111111111110111111101011101;
assign LUT_4[24044] = 32'b11111111111111111100010111011101;
assign LUT_4[24045] = 32'b11111111111111110101100011010101;
assign LUT_4[24046] = 32'b11111111111111111011110010000001;
assign LUT_4[24047] = 32'b11111111111111110100111101111001;
assign LUT_4[24048] = 32'b00000000000000000011111100011010;
assign LUT_4[24049] = 32'b11111111111111111101001000010010;
assign LUT_4[24050] = 32'b00000000000000000011010110111110;
assign LUT_4[24051] = 32'b11111111111111111100100010110110;
assign LUT_4[24052] = 32'b00000000000000000000111100110110;
assign LUT_4[24053] = 32'b11111111111111111010001000101110;
assign LUT_4[24054] = 32'b00000000000000000000010111011010;
assign LUT_4[24055] = 32'b11111111111111111001100011010010;
assign LUT_4[24056] = 32'b11111111111111111101001000101111;
assign LUT_4[24057] = 32'b11111111111111110110010100100111;
assign LUT_4[24058] = 32'b11111111111111111100100011010011;
assign LUT_4[24059] = 32'b11111111111111110101101111001011;
assign LUT_4[24060] = 32'b11111111111111111010001001001011;
assign LUT_4[24061] = 32'b11111111111111110011010101000011;
assign LUT_4[24062] = 32'b11111111111111111001100011101111;
assign LUT_4[24063] = 32'b11111111111111110010101111100111;
assign LUT_4[24064] = 32'b11111111111111111101111010101110;
assign LUT_4[24065] = 32'b11111111111111110111000110100110;
assign LUT_4[24066] = 32'b11111111111111111101010101010010;
assign LUT_4[24067] = 32'b11111111111111110110100001001010;
assign LUT_4[24068] = 32'b11111111111111111010111011001010;
assign LUT_4[24069] = 32'b11111111111111110100000111000010;
assign LUT_4[24070] = 32'b11111111111111111010010101101110;
assign LUT_4[24071] = 32'b11111111111111110011100001100110;
assign LUT_4[24072] = 32'b11111111111111110111000111000011;
assign LUT_4[24073] = 32'b11111111111111110000010010111011;
assign LUT_4[24074] = 32'b11111111111111110110100001100111;
assign LUT_4[24075] = 32'b11111111111111101111101101011111;
assign LUT_4[24076] = 32'b11111111111111110100000111011111;
assign LUT_4[24077] = 32'b11111111111111101101010011010111;
assign LUT_4[24078] = 32'b11111111111111110011100010000011;
assign LUT_4[24079] = 32'b11111111111111101100101101111011;
assign LUT_4[24080] = 32'b11111111111111111011101100011100;
assign LUT_4[24081] = 32'b11111111111111110100111000010100;
assign LUT_4[24082] = 32'b11111111111111111011000111000000;
assign LUT_4[24083] = 32'b11111111111111110100010010111000;
assign LUT_4[24084] = 32'b11111111111111111000101100111000;
assign LUT_4[24085] = 32'b11111111111111110001111000110000;
assign LUT_4[24086] = 32'b11111111111111111000000111011100;
assign LUT_4[24087] = 32'b11111111111111110001010011010100;
assign LUT_4[24088] = 32'b11111111111111110100111000110001;
assign LUT_4[24089] = 32'b11111111111111101110000100101001;
assign LUT_4[24090] = 32'b11111111111111110100010011010101;
assign LUT_4[24091] = 32'b11111111111111101101011111001101;
assign LUT_4[24092] = 32'b11111111111111110001111001001101;
assign LUT_4[24093] = 32'b11111111111111101011000101000101;
assign LUT_4[24094] = 32'b11111111111111110001010011110001;
assign LUT_4[24095] = 32'b11111111111111101010011111101001;
assign LUT_4[24096] = 32'b11111111111111111100010101110101;
assign LUT_4[24097] = 32'b11111111111111110101100001101101;
assign LUT_4[24098] = 32'b11111111111111111011110000011001;
assign LUT_4[24099] = 32'b11111111111111110100111100010001;
assign LUT_4[24100] = 32'b11111111111111111001010110010001;
assign LUT_4[24101] = 32'b11111111111111110010100010001001;
assign LUT_4[24102] = 32'b11111111111111111000110000110101;
assign LUT_4[24103] = 32'b11111111111111110001111100101101;
assign LUT_4[24104] = 32'b11111111111111110101100010001010;
assign LUT_4[24105] = 32'b11111111111111101110101110000010;
assign LUT_4[24106] = 32'b11111111111111110100111100101110;
assign LUT_4[24107] = 32'b11111111111111101110001000100110;
assign LUT_4[24108] = 32'b11111111111111110010100010100110;
assign LUT_4[24109] = 32'b11111111111111101011101110011110;
assign LUT_4[24110] = 32'b11111111111111110001111101001010;
assign LUT_4[24111] = 32'b11111111111111101011001001000010;
assign LUT_4[24112] = 32'b11111111111111111010000111100011;
assign LUT_4[24113] = 32'b11111111111111110011010011011011;
assign LUT_4[24114] = 32'b11111111111111111001100010000111;
assign LUT_4[24115] = 32'b11111111111111110010101101111111;
assign LUT_4[24116] = 32'b11111111111111110111000111111111;
assign LUT_4[24117] = 32'b11111111111111110000010011110111;
assign LUT_4[24118] = 32'b11111111111111110110100010100011;
assign LUT_4[24119] = 32'b11111111111111101111101110011011;
assign LUT_4[24120] = 32'b11111111111111110011010011111000;
assign LUT_4[24121] = 32'b11111111111111101100011111110000;
assign LUT_4[24122] = 32'b11111111111111110010101110011100;
assign LUT_4[24123] = 32'b11111111111111101011111010010100;
assign LUT_4[24124] = 32'b11111111111111110000010100010100;
assign LUT_4[24125] = 32'b11111111111111101001100000001100;
assign LUT_4[24126] = 32'b11111111111111101111101110111000;
assign LUT_4[24127] = 32'b11111111111111101000111010110000;
assign LUT_4[24128] = 32'b11111111111111111111010010000010;
assign LUT_4[24129] = 32'b11111111111111111000011101111010;
assign LUT_4[24130] = 32'b11111111111111111110101100100110;
assign LUT_4[24131] = 32'b11111111111111110111111000011110;
assign LUT_4[24132] = 32'b11111111111111111100010010011110;
assign LUT_4[24133] = 32'b11111111111111110101011110010110;
assign LUT_4[24134] = 32'b11111111111111111011101101000010;
assign LUT_4[24135] = 32'b11111111111111110100111000111010;
assign LUT_4[24136] = 32'b11111111111111111000011110010111;
assign LUT_4[24137] = 32'b11111111111111110001101010001111;
assign LUT_4[24138] = 32'b11111111111111110111111000111011;
assign LUT_4[24139] = 32'b11111111111111110001000100110011;
assign LUT_4[24140] = 32'b11111111111111110101011110110011;
assign LUT_4[24141] = 32'b11111111111111101110101010101011;
assign LUT_4[24142] = 32'b11111111111111110100111001010111;
assign LUT_4[24143] = 32'b11111111111111101110000101001111;
assign LUT_4[24144] = 32'b11111111111111111101000011110000;
assign LUT_4[24145] = 32'b11111111111111110110001111101000;
assign LUT_4[24146] = 32'b11111111111111111100011110010100;
assign LUT_4[24147] = 32'b11111111111111110101101010001100;
assign LUT_4[24148] = 32'b11111111111111111010000100001100;
assign LUT_4[24149] = 32'b11111111111111110011010000000100;
assign LUT_4[24150] = 32'b11111111111111111001011110110000;
assign LUT_4[24151] = 32'b11111111111111110010101010101000;
assign LUT_4[24152] = 32'b11111111111111110110010000000101;
assign LUT_4[24153] = 32'b11111111111111101111011011111101;
assign LUT_4[24154] = 32'b11111111111111110101101010101001;
assign LUT_4[24155] = 32'b11111111111111101110110110100001;
assign LUT_4[24156] = 32'b11111111111111110011010000100001;
assign LUT_4[24157] = 32'b11111111111111101100011100011001;
assign LUT_4[24158] = 32'b11111111111111110010101011000101;
assign LUT_4[24159] = 32'b11111111111111101011110110111101;
assign LUT_4[24160] = 32'b11111111111111111101101101001001;
assign LUT_4[24161] = 32'b11111111111111110110111001000001;
assign LUT_4[24162] = 32'b11111111111111111101000111101101;
assign LUT_4[24163] = 32'b11111111111111110110010011100101;
assign LUT_4[24164] = 32'b11111111111111111010101101100101;
assign LUT_4[24165] = 32'b11111111111111110011111001011101;
assign LUT_4[24166] = 32'b11111111111111111010001000001001;
assign LUT_4[24167] = 32'b11111111111111110011010100000001;
assign LUT_4[24168] = 32'b11111111111111110110111001011110;
assign LUT_4[24169] = 32'b11111111111111110000000101010110;
assign LUT_4[24170] = 32'b11111111111111110110010100000010;
assign LUT_4[24171] = 32'b11111111111111101111011111111010;
assign LUT_4[24172] = 32'b11111111111111110011111001111010;
assign LUT_4[24173] = 32'b11111111111111101101000101110010;
assign LUT_4[24174] = 32'b11111111111111110011010100011110;
assign LUT_4[24175] = 32'b11111111111111101100100000010110;
assign LUT_4[24176] = 32'b11111111111111111011011110110111;
assign LUT_4[24177] = 32'b11111111111111110100101010101111;
assign LUT_4[24178] = 32'b11111111111111111010111001011011;
assign LUT_4[24179] = 32'b11111111111111110100000101010011;
assign LUT_4[24180] = 32'b11111111111111111000011111010011;
assign LUT_4[24181] = 32'b11111111111111110001101011001011;
assign LUT_4[24182] = 32'b11111111111111110111111001110111;
assign LUT_4[24183] = 32'b11111111111111110001000101101111;
assign LUT_4[24184] = 32'b11111111111111110100101011001100;
assign LUT_4[24185] = 32'b11111111111111101101110111000100;
assign LUT_4[24186] = 32'b11111111111111110100000101110000;
assign LUT_4[24187] = 32'b11111111111111101101010001101000;
assign LUT_4[24188] = 32'b11111111111111110001101011101000;
assign LUT_4[24189] = 32'b11111111111111101010110111100000;
assign LUT_4[24190] = 32'b11111111111111110001000110001100;
assign LUT_4[24191] = 32'b11111111111111101010010010000100;
assign LUT_4[24192] = 32'b00000000000000000000100000110110;
assign LUT_4[24193] = 32'b11111111111111111001101100101110;
assign LUT_4[24194] = 32'b11111111111111111111111011011010;
assign LUT_4[24195] = 32'b11111111111111111001000111010010;
assign LUT_4[24196] = 32'b11111111111111111101100001010010;
assign LUT_4[24197] = 32'b11111111111111110110101101001010;
assign LUT_4[24198] = 32'b11111111111111111100111011110110;
assign LUT_4[24199] = 32'b11111111111111110110000111101110;
assign LUT_4[24200] = 32'b11111111111111111001101101001011;
assign LUT_4[24201] = 32'b11111111111111110010111001000011;
assign LUT_4[24202] = 32'b11111111111111111001000111101111;
assign LUT_4[24203] = 32'b11111111111111110010010011100111;
assign LUT_4[24204] = 32'b11111111111111110110101101100111;
assign LUT_4[24205] = 32'b11111111111111101111111001011111;
assign LUT_4[24206] = 32'b11111111111111110110001000001011;
assign LUT_4[24207] = 32'b11111111111111101111010100000011;
assign LUT_4[24208] = 32'b11111111111111111110010010100100;
assign LUT_4[24209] = 32'b11111111111111110111011110011100;
assign LUT_4[24210] = 32'b11111111111111111101101101001000;
assign LUT_4[24211] = 32'b11111111111111110110111001000000;
assign LUT_4[24212] = 32'b11111111111111111011010011000000;
assign LUT_4[24213] = 32'b11111111111111110100011110111000;
assign LUT_4[24214] = 32'b11111111111111111010101101100100;
assign LUT_4[24215] = 32'b11111111111111110011111001011100;
assign LUT_4[24216] = 32'b11111111111111110111011110111001;
assign LUT_4[24217] = 32'b11111111111111110000101010110001;
assign LUT_4[24218] = 32'b11111111111111110110111001011101;
assign LUT_4[24219] = 32'b11111111111111110000000101010101;
assign LUT_4[24220] = 32'b11111111111111110100011111010101;
assign LUT_4[24221] = 32'b11111111111111101101101011001101;
assign LUT_4[24222] = 32'b11111111111111110011111001111001;
assign LUT_4[24223] = 32'b11111111111111101101000101110001;
assign LUT_4[24224] = 32'b11111111111111111110111011111101;
assign LUT_4[24225] = 32'b11111111111111111000000111110101;
assign LUT_4[24226] = 32'b11111111111111111110010110100001;
assign LUT_4[24227] = 32'b11111111111111110111100010011001;
assign LUT_4[24228] = 32'b11111111111111111011111100011001;
assign LUT_4[24229] = 32'b11111111111111110101001000010001;
assign LUT_4[24230] = 32'b11111111111111111011010110111101;
assign LUT_4[24231] = 32'b11111111111111110100100010110101;
assign LUT_4[24232] = 32'b11111111111111111000001000010010;
assign LUT_4[24233] = 32'b11111111111111110001010100001010;
assign LUT_4[24234] = 32'b11111111111111110111100010110110;
assign LUT_4[24235] = 32'b11111111111111110000101110101110;
assign LUT_4[24236] = 32'b11111111111111110101001000101110;
assign LUT_4[24237] = 32'b11111111111111101110010100100110;
assign LUT_4[24238] = 32'b11111111111111110100100011010010;
assign LUT_4[24239] = 32'b11111111111111101101101111001010;
assign LUT_4[24240] = 32'b11111111111111111100101101101011;
assign LUT_4[24241] = 32'b11111111111111110101111001100011;
assign LUT_4[24242] = 32'b11111111111111111100001000001111;
assign LUT_4[24243] = 32'b11111111111111110101010100000111;
assign LUT_4[24244] = 32'b11111111111111111001101110000111;
assign LUT_4[24245] = 32'b11111111111111110010111001111111;
assign LUT_4[24246] = 32'b11111111111111111001001000101011;
assign LUT_4[24247] = 32'b11111111111111110010010100100011;
assign LUT_4[24248] = 32'b11111111111111110101111010000000;
assign LUT_4[24249] = 32'b11111111111111101111000101111000;
assign LUT_4[24250] = 32'b11111111111111110101010100100100;
assign LUT_4[24251] = 32'b11111111111111101110100000011100;
assign LUT_4[24252] = 32'b11111111111111110010111010011100;
assign LUT_4[24253] = 32'b11111111111111101100000110010100;
assign LUT_4[24254] = 32'b11111111111111110010010101000000;
assign LUT_4[24255] = 32'b11111111111111101011100000111000;
assign LUT_4[24256] = 32'b00000000000000000001111000001010;
assign LUT_4[24257] = 32'b11111111111111111011000100000010;
assign LUT_4[24258] = 32'b00000000000000000001010010101110;
assign LUT_4[24259] = 32'b11111111111111111010011110100110;
assign LUT_4[24260] = 32'b11111111111111111110111000100110;
assign LUT_4[24261] = 32'b11111111111111111000000100011110;
assign LUT_4[24262] = 32'b11111111111111111110010011001010;
assign LUT_4[24263] = 32'b11111111111111110111011111000010;
assign LUT_4[24264] = 32'b11111111111111111011000100011111;
assign LUT_4[24265] = 32'b11111111111111110100010000010111;
assign LUT_4[24266] = 32'b11111111111111111010011111000011;
assign LUT_4[24267] = 32'b11111111111111110011101010111011;
assign LUT_4[24268] = 32'b11111111111111111000000100111011;
assign LUT_4[24269] = 32'b11111111111111110001010000110011;
assign LUT_4[24270] = 32'b11111111111111110111011111011111;
assign LUT_4[24271] = 32'b11111111111111110000101011010111;
assign LUT_4[24272] = 32'b11111111111111111111101001111000;
assign LUT_4[24273] = 32'b11111111111111111000110101110000;
assign LUT_4[24274] = 32'b11111111111111111111000100011100;
assign LUT_4[24275] = 32'b11111111111111111000010000010100;
assign LUT_4[24276] = 32'b11111111111111111100101010010100;
assign LUT_4[24277] = 32'b11111111111111110101110110001100;
assign LUT_4[24278] = 32'b11111111111111111100000100111000;
assign LUT_4[24279] = 32'b11111111111111110101010000110000;
assign LUT_4[24280] = 32'b11111111111111111000110110001101;
assign LUT_4[24281] = 32'b11111111111111110010000010000101;
assign LUT_4[24282] = 32'b11111111111111111000010000110001;
assign LUT_4[24283] = 32'b11111111111111110001011100101001;
assign LUT_4[24284] = 32'b11111111111111110101110110101001;
assign LUT_4[24285] = 32'b11111111111111101111000010100001;
assign LUT_4[24286] = 32'b11111111111111110101010001001101;
assign LUT_4[24287] = 32'b11111111111111101110011101000101;
assign LUT_4[24288] = 32'b00000000000000000000010011010001;
assign LUT_4[24289] = 32'b11111111111111111001011111001001;
assign LUT_4[24290] = 32'b11111111111111111111101101110101;
assign LUT_4[24291] = 32'b11111111111111111000111001101101;
assign LUT_4[24292] = 32'b11111111111111111101010011101101;
assign LUT_4[24293] = 32'b11111111111111110110011111100101;
assign LUT_4[24294] = 32'b11111111111111111100101110010001;
assign LUT_4[24295] = 32'b11111111111111110101111010001001;
assign LUT_4[24296] = 32'b11111111111111111001011111100110;
assign LUT_4[24297] = 32'b11111111111111110010101011011110;
assign LUT_4[24298] = 32'b11111111111111111000111010001010;
assign LUT_4[24299] = 32'b11111111111111110010000110000010;
assign LUT_4[24300] = 32'b11111111111111110110100000000010;
assign LUT_4[24301] = 32'b11111111111111101111101011111010;
assign LUT_4[24302] = 32'b11111111111111110101111010100110;
assign LUT_4[24303] = 32'b11111111111111101111000110011110;
assign LUT_4[24304] = 32'b11111111111111111110000100111111;
assign LUT_4[24305] = 32'b11111111111111110111010000110111;
assign LUT_4[24306] = 32'b11111111111111111101011111100011;
assign LUT_4[24307] = 32'b11111111111111110110101011011011;
assign LUT_4[24308] = 32'b11111111111111111011000101011011;
assign LUT_4[24309] = 32'b11111111111111110100010001010011;
assign LUT_4[24310] = 32'b11111111111111111010011111111111;
assign LUT_4[24311] = 32'b11111111111111110011101011110111;
assign LUT_4[24312] = 32'b11111111111111110111010001010100;
assign LUT_4[24313] = 32'b11111111111111110000011101001100;
assign LUT_4[24314] = 32'b11111111111111110110101011111000;
assign LUT_4[24315] = 32'b11111111111111101111110111110000;
assign LUT_4[24316] = 32'b11111111111111110100010001110000;
assign LUT_4[24317] = 32'b11111111111111101101011101101000;
assign LUT_4[24318] = 32'b11111111111111110011101100010100;
assign LUT_4[24319] = 32'b11111111111111101100111000001100;
assign LUT_4[24320] = 32'b00000000000000000010110110010001;
assign LUT_4[24321] = 32'b11111111111111111100000010001001;
assign LUT_4[24322] = 32'b00000000000000000010010000110101;
assign LUT_4[24323] = 32'b11111111111111111011011100101101;
assign LUT_4[24324] = 32'b11111111111111111111110110101101;
assign LUT_4[24325] = 32'b11111111111111111001000010100101;
assign LUT_4[24326] = 32'b11111111111111111111010001010001;
assign LUT_4[24327] = 32'b11111111111111111000011101001001;
assign LUT_4[24328] = 32'b11111111111111111100000010100110;
assign LUT_4[24329] = 32'b11111111111111110101001110011110;
assign LUT_4[24330] = 32'b11111111111111111011011101001010;
assign LUT_4[24331] = 32'b11111111111111110100101001000010;
assign LUT_4[24332] = 32'b11111111111111111001000011000010;
assign LUT_4[24333] = 32'b11111111111111110010001110111010;
assign LUT_4[24334] = 32'b11111111111111111000011101100110;
assign LUT_4[24335] = 32'b11111111111111110001101001011110;
assign LUT_4[24336] = 32'b00000000000000000000100111111111;
assign LUT_4[24337] = 32'b11111111111111111001110011110111;
assign LUT_4[24338] = 32'b00000000000000000000000010100011;
assign LUT_4[24339] = 32'b11111111111111111001001110011011;
assign LUT_4[24340] = 32'b11111111111111111101101000011011;
assign LUT_4[24341] = 32'b11111111111111110110110100010011;
assign LUT_4[24342] = 32'b11111111111111111101000010111111;
assign LUT_4[24343] = 32'b11111111111111110110001110110111;
assign LUT_4[24344] = 32'b11111111111111111001110100010100;
assign LUT_4[24345] = 32'b11111111111111110011000000001100;
assign LUT_4[24346] = 32'b11111111111111111001001110111000;
assign LUT_4[24347] = 32'b11111111111111110010011010110000;
assign LUT_4[24348] = 32'b11111111111111110110110100110000;
assign LUT_4[24349] = 32'b11111111111111110000000000101000;
assign LUT_4[24350] = 32'b11111111111111110110001111010100;
assign LUT_4[24351] = 32'b11111111111111101111011011001100;
assign LUT_4[24352] = 32'b00000000000000000001010001011000;
assign LUT_4[24353] = 32'b11111111111111111010011101010000;
assign LUT_4[24354] = 32'b00000000000000000000101011111100;
assign LUT_4[24355] = 32'b11111111111111111001110111110100;
assign LUT_4[24356] = 32'b11111111111111111110010001110100;
assign LUT_4[24357] = 32'b11111111111111110111011101101100;
assign LUT_4[24358] = 32'b11111111111111111101101100011000;
assign LUT_4[24359] = 32'b11111111111111110110111000010000;
assign LUT_4[24360] = 32'b11111111111111111010011101101101;
assign LUT_4[24361] = 32'b11111111111111110011101001100101;
assign LUT_4[24362] = 32'b11111111111111111001111000010001;
assign LUT_4[24363] = 32'b11111111111111110011000100001001;
assign LUT_4[24364] = 32'b11111111111111110111011110001001;
assign LUT_4[24365] = 32'b11111111111111110000101010000001;
assign LUT_4[24366] = 32'b11111111111111110110111000101101;
assign LUT_4[24367] = 32'b11111111111111110000000100100101;
assign LUT_4[24368] = 32'b11111111111111111111000011000110;
assign LUT_4[24369] = 32'b11111111111111111000001110111110;
assign LUT_4[24370] = 32'b11111111111111111110011101101010;
assign LUT_4[24371] = 32'b11111111111111110111101001100010;
assign LUT_4[24372] = 32'b11111111111111111100000011100010;
assign LUT_4[24373] = 32'b11111111111111110101001111011010;
assign LUT_4[24374] = 32'b11111111111111111011011110000110;
assign LUT_4[24375] = 32'b11111111111111110100101001111110;
assign LUT_4[24376] = 32'b11111111111111111000001111011011;
assign LUT_4[24377] = 32'b11111111111111110001011011010011;
assign LUT_4[24378] = 32'b11111111111111110111101001111111;
assign LUT_4[24379] = 32'b11111111111111110000110101110111;
assign LUT_4[24380] = 32'b11111111111111110101001111110111;
assign LUT_4[24381] = 32'b11111111111111101110011011101111;
assign LUT_4[24382] = 32'b11111111111111110100101010011011;
assign LUT_4[24383] = 32'b11111111111111101101110110010011;
assign LUT_4[24384] = 32'b00000000000000000100001101100101;
assign LUT_4[24385] = 32'b11111111111111111101011001011101;
assign LUT_4[24386] = 32'b00000000000000000011101000001001;
assign LUT_4[24387] = 32'b11111111111111111100110100000001;
assign LUT_4[24388] = 32'b00000000000000000001001110000001;
assign LUT_4[24389] = 32'b11111111111111111010011001111001;
assign LUT_4[24390] = 32'b00000000000000000000101000100101;
assign LUT_4[24391] = 32'b11111111111111111001110100011101;
assign LUT_4[24392] = 32'b11111111111111111101011001111010;
assign LUT_4[24393] = 32'b11111111111111110110100101110010;
assign LUT_4[24394] = 32'b11111111111111111100110100011110;
assign LUT_4[24395] = 32'b11111111111111110110000000010110;
assign LUT_4[24396] = 32'b11111111111111111010011010010110;
assign LUT_4[24397] = 32'b11111111111111110011100110001110;
assign LUT_4[24398] = 32'b11111111111111111001110100111010;
assign LUT_4[24399] = 32'b11111111111111110011000000110010;
assign LUT_4[24400] = 32'b00000000000000000001111111010011;
assign LUT_4[24401] = 32'b11111111111111111011001011001011;
assign LUT_4[24402] = 32'b00000000000000000001011001110111;
assign LUT_4[24403] = 32'b11111111111111111010100101101111;
assign LUT_4[24404] = 32'b11111111111111111110111111101111;
assign LUT_4[24405] = 32'b11111111111111111000001011100111;
assign LUT_4[24406] = 32'b11111111111111111110011010010011;
assign LUT_4[24407] = 32'b11111111111111110111100110001011;
assign LUT_4[24408] = 32'b11111111111111111011001011101000;
assign LUT_4[24409] = 32'b11111111111111110100010111100000;
assign LUT_4[24410] = 32'b11111111111111111010100110001100;
assign LUT_4[24411] = 32'b11111111111111110011110010000100;
assign LUT_4[24412] = 32'b11111111111111111000001100000100;
assign LUT_4[24413] = 32'b11111111111111110001010111111100;
assign LUT_4[24414] = 32'b11111111111111110111100110101000;
assign LUT_4[24415] = 32'b11111111111111110000110010100000;
assign LUT_4[24416] = 32'b00000000000000000010101000101100;
assign LUT_4[24417] = 32'b11111111111111111011110100100100;
assign LUT_4[24418] = 32'b00000000000000000010000011010000;
assign LUT_4[24419] = 32'b11111111111111111011001111001000;
assign LUT_4[24420] = 32'b11111111111111111111101001001000;
assign LUT_4[24421] = 32'b11111111111111111000110101000000;
assign LUT_4[24422] = 32'b11111111111111111111000011101100;
assign LUT_4[24423] = 32'b11111111111111111000001111100100;
assign LUT_4[24424] = 32'b11111111111111111011110101000001;
assign LUT_4[24425] = 32'b11111111111111110101000000111001;
assign LUT_4[24426] = 32'b11111111111111111011001111100101;
assign LUT_4[24427] = 32'b11111111111111110100011011011101;
assign LUT_4[24428] = 32'b11111111111111111000110101011101;
assign LUT_4[24429] = 32'b11111111111111110010000001010101;
assign LUT_4[24430] = 32'b11111111111111111000010000000001;
assign LUT_4[24431] = 32'b11111111111111110001011011111001;
assign LUT_4[24432] = 32'b00000000000000000000011010011010;
assign LUT_4[24433] = 32'b11111111111111111001100110010010;
assign LUT_4[24434] = 32'b11111111111111111111110100111110;
assign LUT_4[24435] = 32'b11111111111111111001000000110110;
assign LUT_4[24436] = 32'b11111111111111111101011010110110;
assign LUT_4[24437] = 32'b11111111111111110110100110101110;
assign LUT_4[24438] = 32'b11111111111111111100110101011010;
assign LUT_4[24439] = 32'b11111111111111110110000001010010;
assign LUT_4[24440] = 32'b11111111111111111001100110101111;
assign LUT_4[24441] = 32'b11111111111111110010110010100111;
assign LUT_4[24442] = 32'b11111111111111111001000001010011;
assign LUT_4[24443] = 32'b11111111111111110010001101001011;
assign LUT_4[24444] = 32'b11111111111111110110100111001011;
assign LUT_4[24445] = 32'b11111111111111101111110011000011;
assign LUT_4[24446] = 32'b11111111111111110110000001101111;
assign LUT_4[24447] = 32'b11111111111111101111001101100111;
assign LUT_4[24448] = 32'b00000000000000000101011100011001;
assign LUT_4[24449] = 32'b11111111111111111110101000010001;
assign LUT_4[24450] = 32'b00000000000000000100110110111101;
assign LUT_4[24451] = 32'b11111111111111111110000010110101;
assign LUT_4[24452] = 32'b00000000000000000010011100110101;
assign LUT_4[24453] = 32'b11111111111111111011101000101101;
assign LUT_4[24454] = 32'b00000000000000000001110111011001;
assign LUT_4[24455] = 32'b11111111111111111011000011010001;
assign LUT_4[24456] = 32'b11111111111111111110101000101110;
assign LUT_4[24457] = 32'b11111111111111110111110100100110;
assign LUT_4[24458] = 32'b11111111111111111110000011010010;
assign LUT_4[24459] = 32'b11111111111111110111001111001010;
assign LUT_4[24460] = 32'b11111111111111111011101001001010;
assign LUT_4[24461] = 32'b11111111111111110100110101000010;
assign LUT_4[24462] = 32'b11111111111111111011000011101110;
assign LUT_4[24463] = 32'b11111111111111110100001111100110;
assign LUT_4[24464] = 32'b00000000000000000011001110000111;
assign LUT_4[24465] = 32'b11111111111111111100011001111111;
assign LUT_4[24466] = 32'b00000000000000000010101000101011;
assign LUT_4[24467] = 32'b11111111111111111011110100100011;
assign LUT_4[24468] = 32'b00000000000000000000001110100011;
assign LUT_4[24469] = 32'b11111111111111111001011010011011;
assign LUT_4[24470] = 32'b11111111111111111111101001000111;
assign LUT_4[24471] = 32'b11111111111111111000110100111111;
assign LUT_4[24472] = 32'b11111111111111111100011010011100;
assign LUT_4[24473] = 32'b11111111111111110101100110010100;
assign LUT_4[24474] = 32'b11111111111111111011110101000000;
assign LUT_4[24475] = 32'b11111111111111110101000000111000;
assign LUT_4[24476] = 32'b11111111111111111001011010111000;
assign LUT_4[24477] = 32'b11111111111111110010100110110000;
assign LUT_4[24478] = 32'b11111111111111111000110101011100;
assign LUT_4[24479] = 32'b11111111111111110010000001010100;
assign LUT_4[24480] = 32'b00000000000000000011110111100000;
assign LUT_4[24481] = 32'b11111111111111111101000011011000;
assign LUT_4[24482] = 32'b00000000000000000011010010000100;
assign LUT_4[24483] = 32'b11111111111111111100011101111100;
assign LUT_4[24484] = 32'b00000000000000000000110111111100;
assign LUT_4[24485] = 32'b11111111111111111010000011110100;
assign LUT_4[24486] = 32'b00000000000000000000010010100000;
assign LUT_4[24487] = 32'b11111111111111111001011110011000;
assign LUT_4[24488] = 32'b11111111111111111101000011110101;
assign LUT_4[24489] = 32'b11111111111111110110001111101101;
assign LUT_4[24490] = 32'b11111111111111111100011110011001;
assign LUT_4[24491] = 32'b11111111111111110101101010010001;
assign LUT_4[24492] = 32'b11111111111111111010000100010001;
assign LUT_4[24493] = 32'b11111111111111110011010000001001;
assign LUT_4[24494] = 32'b11111111111111111001011110110101;
assign LUT_4[24495] = 32'b11111111111111110010101010101101;
assign LUT_4[24496] = 32'b00000000000000000001101001001110;
assign LUT_4[24497] = 32'b11111111111111111010110101000110;
assign LUT_4[24498] = 32'b00000000000000000001000011110010;
assign LUT_4[24499] = 32'b11111111111111111010001111101010;
assign LUT_4[24500] = 32'b11111111111111111110101001101010;
assign LUT_4[24501] = 32'b11111111111111110111110101100010;
assign LUT_4[24502] = 32'b11111111111111111110000100001110;
assign LUT_4[24503] = 32'b11111111111111110111010000000110;
assign LUT_4[24504] = 32'b11111111111111111010110101100011;
assign LUT_4[24505] = 32'b11111111111111110100000001011011;
assign LUT_4[24506] = 32'b11111111111111111010010000000111;
assign LUT_4[24507] = 32'b11111111111111110011011011111111;
assign LUT_4[24508] = 32'b11111111111111110111110101111111;
assign LUT_4[24509] = 32'b11111111111111110001000001110111;
assign LUT_4[24510] = 32'b11111111111111110111010000100011;
assign LUT_4[24511] = 32'b11111111111111110000011100011011;
assign LUT_4[24512] = 32'b00000000000000000110110011101101;
assign LUT_4[24513] = 32'b11111111111111111111111111100101;
assign LUT_4[24514] = 32'b00000000000000000110001110010001;
assign LUT_4[24515] = 32'b11111111111111111111011010001001;
assign LUT_4[24516] = 32'b00000000000000000011110100001001;
assign LUT_4[24517] = 32'b11111111111111111101000000000001;
assign LUT_4[24518] = 32'b00000000000000000011001110101101;
assign LUT_4[24519] = 32'b11111111111111111100011010100101;
assign LUT_4[24520] = 32'b00000000000000000000000000000010;
assign LUT_4[24521] = 32'b11111111111111111001001011111010;
assign LUT_4[24522] = 32'b11111111111111111111011010100110;
assign LUT_4[24523] = 32'b11111111111111111000100110011110;
assign LUT_4[24524] = 32'b11111111111111111101000000011110;
assign LUT_4[24525] = 32'b11111111111111110110001100010110;
assign LUT_4[24526] = 32'b11111111111111111100011011000010;
assign LUT_4[24527] = 32'b11111111111111110101100110111010;
assign LUT_4[24528] = 32'b00000000000000000100100101011011;
assign LUT_4[24529] = 32'b11111111111111111101110001010011;
assign LUT_4[24530] = 32'b00000000000000000011111111111111;
assign LUT_4[24531] = 32'b11111111111111111101001011110111;
assign LUT_4[24532] = 32'b00000000000000000001100101110111;
assign LUT_4[24533] = 32'b11111111111111111010110001101111;
assign LUT_4[24534] = 32'b00000000000000000001000000011011;
assign LUT_4[24535] = 32'b11111111111111111010001100010011;
assign LUT_4[24536] = 32'b11111111111111111101110001110000;
assign LUT_4[24537] = 32'b11111111111111110110111101101000;
assign LUT_4[24538] = 32'b11111111111111111101001100010100;
assign LUT_4[24539] = 32'b11111111111111110110011000001100;
assign LUT_4[24540] = 32'b11111111111111111010110010001100;
assign LUT_4[24541] = 32'b11111111111111110011111110000100;
assign LUT_4[24542] = 32'b11111111111111111010001100110000;
assign LUT_4[24543] = 32'b11111111111111110011011000101000;
assign LUT_4[24544] = 32'b00000000000000000101001110110100;
assign LUT_4[24545] = 32'b11111111111111111110011010101100;
assign LUT_4[24546] = 32'b00000000000000000100101001011000;
assign LUT_4[24547] = 32'b11111111111111111101110101010000;
assign LUT_4[24548] = 32'b00000000000000000010001111010000;
assign LUT_4[24549] = 32'b11111111111111111011011011001000;
assign LUT_4[24550] = 32'b00000000000000000001101001110100;
assign LUT_4[24551] = 32'b11111111111111111010110101101100;
assign LUT_4[24552] = 32'b11111111111111111110011011001001;
assign LUT_4[24553] = 32'b11111111111111110111100111000001;
assign LUT_4[24554] = 32'b11111111111111111101110101101101;
assign LUT_4[24555] = 32'b11111111111111110111000001100101;
assign LUT_4[24556] = 32'b11111111111111111011011011100101;
assign LUT_4[24557] = 32'b11111111111111110100100111011101;
assign LUT_4[24558] = 32'b11111111111111111010110110001001;
assign LUT_4[24559] = 32'b11111111111111110100000010000001;
assign LUT_4[24560] = 32'b00000000000000000011000000100010;
assign LUT_4[24561] = 32'b11111111111111111100001100011010;
assign LUT_4[24562] = 32'b00000000000000000010011011000110;
assign LUT_4[24563] = 32'b11111111111111111011100110111110;
assign LUT_4[24564] = 32'b00000000000000000000000000111110;
assign LUT_4[24565] = 32'b11111111111111111001001100110110;
assign LUT_4[24566] = 32'b11111111111111111111011011100010;
assign LUT_4[24567] = 32'b11111111111111111000100111011010;
assign LUT_4[24568] = 32'b11111111111111111100001100110111;
assign LUT_4[24569] = 32'b11111111111111110101011000101111;
assign LUT_4[24570] = 32'b11111111111111111011100111011011;
assign LUT_4[24571] = 32'b11111111111111110100110011010011;
assign LUT_4[24572] = 32'b11111111111111111001001101010011;
assign LUT_4[24573] = 32'b11111111111111110010011001001011;
assign LUT_4[24574] = 32'b11111111111111111000100111110111;
assign LUT_4[24575] = 32'b11111111111111110001110011101111;
assign LUT_4[24576] = 32'b00000000000000001011101100011000;
assign LUT_4[24577] = 32'b00000000000000000100111000010000;
assign LUT_4[24578] = 32'b00000000000000001011000110111100;
assign LUT_4[24579] = 32'b00000000000000000100010010110100;
assign LUT_4[24580] = 32'b00000000000000001000101100110100;
assign LUT_4[24581] = 32'b00000000000000000001111000101100;
assign LUT_4[24582] = 32'b00000000000000001000000111011000;
assign LUT_4[24583] = 32'b00000000000000000001010011010000;
assign LUT_4[24584] = 32'b00000000000000000100111000101101;
assign LUT_4[24585] = 32'b11111111111111111110000100100101;
assign LUT_4[24586] = 32'b00000000000000000100010011010001;
assign LUT_4[24587] = 32'b11111111111111111101011111001001;
assign LUT_4[24588] = 32'b00000000000000000001111001001001;
assign LUT_4[24589] = 32'b11111111111111111011000101000001;
assign LUT_4[24590] = 32'b00000000000000000001010011101101;
assign LUT_4[24591] = 32'b11111111111111111010011111100101;
assign LUT_4[24592] = 32'b00000000000000001001011110000110;
assign LUT_4[24593] = 32'b00000000000000000010101001111110;
assign LUT_4[24594] = 32'b00000000000000001000111000101010;
assign LUT_4[24595] = 32'b00000000000000000010000100100010;
assign LUT_4[24596] = 32'b00000000000000000110011110100010;
assign LUT_4[24597] = 32'b11111111111111111111101010011010;
assign LUT_4[24598] = 32'b00000000000000000101111001000110;
assign LUT_4[24599] = 32'b11111111111111111111000100111110;
assign LUT_4[24600] = 32'b00000000000000000010101010011011;
assign LUT_4[24601] = 32'b11111111111111111011110110010011;
assign LUT_4[24602] = 32'b00000000000000000010000100111111;
assign LUT_4[24603] = 32'b11111111111111111011010000110111;
assign LUT_4[24604] = 32'b11111111111111111111101010110111;
assign LUT_4[24605] = 32'b11111111111111111000110110101111;
assign LUT_4[24606] = 32'b11111111111111111111000101011011;
assign LUT_4[24607] = 32'b11111111111111111000010001010011;
assign LUT_4[24608] = 32'b00000000000000001010000111011111;
assign LUT_4[24609] = 32'b00000000000000000011010011010111;
assign LUT_4[24610] = 32'b00000000000000001001100010000011;
assign LUT_4[24611] = 32'b00000000000000000010101101111011;
assign LUT_4[24612] = 32'b00000000000000000111000111111011;
assign LUT_4[24613] = 32'b00000000000000000000010011110011;
assign LUT_4[24614] = 32'b00000000000000000110100010011111;
assign LUT_4[24615] = 32'b11111111111111111111101110010111;
assign LUT_4[24616] = 32'b00000000000000000011010011110100;
assign LUT_4[24617] = 32'b11111111111111111100011111101100;
assign LUT_4[24618] = 32'b00000000000000000010101110011000;
assign LUT_4[24619] = 32'b11111111111111111011111010010000;
assign LUT_4[24620] = 32'b00000000000000000000010100010000;
assign LUT_4[24621] = 32'b11111111111111111001100000001000;
assign LUT_4[24622] = 32'b11111111111111111111101110110100;
assign LUT_4[24623] = 32'b11111111111111111000111010101100;
assign LUT_4[24624] = 32'b00000000000000000111111001001101;
assign LUT_4[24625] = 32'b00000000000000000001000101000101;
assign LUT_4[24626] = 32'b00000000000000000111010011110001;
assign LUT_4[24627] = 32'b00000000000000000000011111101001;
assign LUT_4[24628] = 32'b00000000000000000100111001101001;
assign LUT_4[24629] = 32'b11111111111111111110000101100001;
assign LUT_4[24630] = 32'b00000000000000000100010100001101;
assign LUT_4[24631] = 32'b11111111111111111101100000000101;
assign LUT_4[24632] = 32'b00000000000000000001000101100010;
assign LUT_4[24633] = 32'b11111111111111111010010001011010;
assign LUT_4[24634] = 32'b00000000000000000000100000000110;
assign LUT_4[24635] = 32'b11111111111111111001101011111110;
assign LUT_4[24636] = 32'b11111111111111111110000101111110;
assign LUT_4[24637] = 32'b11111111111111110111010001110110;
assign LUT_4[24638] = 32'b11111111111111111101100000100010;
assign LUT_4[24639] = 32'b11111111111111110110101100011010;
assign LUT_4[24640] = 32'b00000000000000001101000011101100;
assign LUT_4[24641] = 32'b00000000000000000110001111100100;
assign LUT_4[24642] = 32'b00000000000000001100011110010000;
assign LUT_4[24643] = 32'b00000000000000000101101010001000;
assign LUT_4[24644] = 32'b00000000000000001010000100001000;
assign LUT_4[24645] = 32'b00000000000000000011010000000000;
assign LUT_4[24646] = 32'b00000000000000001001011110101100;
assign LUT_4[24647] = 32'b00000000000000000010101010100100;
assign LUT_4[24648] = 32'b00000000000000000110010000000001;
assign LUT_4[24649] = 32'b11111111111111111111011011111001;
assign LUT_4[24650] = 32'b00000000000000000101101010100101;
assign LUT_4[24651] = 32'b11111111111111111110110110011101;
assign LUT_4[24652] = 32'b00000000000000000011010000011101;
assign LUT_4[24653] = 32'b11111111111111111100011100010101;
assign LUT_4[24654] = 32'b00000000000000000010101011000001;
assign LUT_4[24655] = 32'b11111111111111111011110110111001;
assign LUT_4[24656] = 32'b00000000000000001010110101011010;
assign LUT_4[24657] = 32'b00000000000000000100000001010010;
assign LUT_4[24658] = 32'b00000000000000001010001111111110;
assign LUT_4[24659] = 32'b00000000000000000011011011110110;
assign LUT_4[24660] = 32'b00000000000000000111110101110110;
assign LUT_4[24661] = 32'b00000000000000000001000001101110;
assign LUT_4[24662] = 32'b00000000000000000111010000011010;
assign LUT_4[24663] = 32'b00000000000000000000011100010010;
assign LUT_4[24664] = 32'b00000000000000000100000001101111;
assign LUT_4[24665] = 32'b11111111111111111101001101100111;
assign LUT_4[24666] = 32'b00000000000000000011011100010011;
assign LUT_4[24667] = 32'b11111111111111111100101000001011;
assign LUT_4[24668] = 32'b00000000000000000001000010001011;
assign LUT_4[24669] = 32'b11111111111111111010001110000011;
assign LUT_4[24670] = 32'b00000000000000000000011100101111;
assign LUT_4[24671] = 32'b11111111111111111001101000100111;
assign LUT_4[24672] = 32'b00000000000000001011011110110011;
assign LUT_4[24673] = 32'b00000000000000000100101010101011;
assign LUT_4[24674] = 32'b00000000000000001010111001010111;
assign LUT_4[24675] = 32'b00000000000000000100000101001111;
assign LUT_4[24676] = 32'b00000000000000001000011111001111;
assign LUT_4[24677] = 32'b00000000000000000001101011000111;
assign LUT_4[24678] = 32'b00000000000000000111111001110011;
assign LUT_4[24679] = 32'b00000000000000000001000101101011;
assign LUT_4[24680] = 32'b00000000000000000100101011001000;
assign LUT_4[24681] = 32'b11111111111111111101110111000000;
assign LUT_4[24682] = 32'b00000000000000000100000101101100;
assign LUT_4[24683] = 32'b11111111111111111101010001100100;
assign LUT_4[24684] = 32'b00000000000000000001101011100100;
assign LUT_4[24685] = 32'b11111111111111111010110111011100;
assign LUT_4[24686] = 32'b00000000000000000001000110001000;
assign LUT_4[24687] = 32'b11111111111111111010010010000000;
assign LUT_4[24688] = 32'b00000000000000001001010000100001;
assign LUT_4[24689] = 32'b00000000000000000010011100011001;
assign LUT_4[24690] = 32'b00000000000000001000101011000101;
assign LUT_4[24691] = 32'b00000000000000000001110110111101;
assign LUT_4[24692] = 32'b00000000000000000110010000111101;
assign LUT_4[24693] = 32'b11111111111111111111011100110101;
assign LUT_4[24694] = 32'b00000000000000000101101011100001;
assign LUT_4[24695] = 32'b11111111111111111110110111011001;
assign LUT_4[24696] = 32'b00000000000000000010011100110110;
assign LUT_4[24697] = 32'b11111111111111111011101000101110;
assign LUT_4[24698] = 32'b00000000000000000001110111011010;
assign LUT_4[24699] = 32'b11111111111111111011000011010010;
assign LUT_4[24700] = 32'b11111111111111111111011101010010;
assign LUT_4[24701] = 32'b11111111111111111000101001001010;
assign LUT_4[24702] = 32'b11111111111111111110110111110110;
assign LUT_4[24703] = 32'b11111111111111111000000011101110;
assign LUT_4[24704] = 32'b00000000000000001110010010100000;
assign LUT_4[24705] = 32'b00000000000000000111011110011000;
assign LUT_4[24706] = 32'b00000000000000001101101101000100;
assign LUT_4[24707] = 32'b00000000000000000110111000111100;
assign LUT_4[24708] = 32'b00000000000000001011010010111100;
assign LUT_4[24709] = 32'b00000000000000000100011110110100;
assign LUT_4[24710] = 32'b00000000000000001010101101100000;
assign LUT_4[24711] = 32'b00000000000000000011111001011000;
assign LUT_4[24712] = 32'b00000000000000000111011110110101;
assign LUT_4[24713] = 32'b00000000000000000000101010101101;
assign LUT_4[24714] = 32'b00000000000000000110111001011001;
assign LUT_4[24715] = 32'b00000000000000000000000101010001;
assign LUT_4[24716] = 32'b00000000000000000100011111010001;
assign LUT_4[24717] = 32'b11111111111111111101101011001001;
assign LUT_4[24718] = 32'b00000000000000000011111001110101;
assign LUT_4[24719] = 32'b11111111111111111101000101101101;
assign LUT_4[24720] = 32'b00000000000000001100000100001110;
assign LUT_4[24721] = 32'b00000000000000000101010000000110;
assign LUT_4[24722] = 32'b00000000000000001011011110110010;
assign LUT_4[24723] = 32'b00000000000000000100101010101010;
assign LUT_4[24724] = 32'b00000000000000001001000100101010;
assign LUT_4[24725] = 32'b00000000000000000010010000100010;
assign LUT_4[24726] = 32'b00000000000000001000011111001110;
assign LUT_4[24727] = 32'b00000000000000000001101011000110;
assign LUT_4[24728] = 32'b00000000000000000101010000100011;
assign LUT_4[24729] = 32'b11111111111111111110011100011011;
assign LUT_4[24730] = 32'b00000000000000000100101011000111;
assign LUT_4[24731] = 32'b11111111111111111101110110111111;
assign LUT_4[24732] = 32'b00000000000000000010010000111111;
assign LUT_4[24733] = 32'b11111111111111111011011100110111;
assign LUT_4[24734] = 32'b00000000000000000001101011100011;
assign LUT_4[24735] = 32'b11111111111111111010110111011011;
assign LUT_4[24736] = 32'b00000000000000001100101101100111;
assign LUT_4[24737] = 32'b00000000000000000101111001011111;
assign LUT_4[24738] = 32'b00000000000000001100001000001011;
assign LUT_4[24739] = 32'b00000000000000000101010100000011;
assign LUT_4[24740] = 32'b00000000000000001001101110000011;
assign LUT_4[24741] = 32'b00000000000000000010111001111011;
assign LUT_4[24742] = 32'b00000000000000001001001000100111;
assign LUT_4[24743] = 32'b00000000000000000010010100011111;
assign LUT_4[24744] = 32'b00000000000000000101111001111100;
assign LUT_4[24745] = 32'b11111111111111111111000101110100;
assign LUT_4[24746] = 32'b00000000000000000101010100100000;
assign LUT_4[24747] = 32'b11111111111111111110100000011000;
assign LUT_4[24748] = 32'b00000000000000000010111010011000;
assign LUT_4[24749] = 32'b11111111111111111100000110010000;
assign LUT_4[24750] = 32'b00000000000000000010010100111100;
assign LUT_4[24751] = 32'b11111111111111111011100000110100;
assign LUT_4[24752] = 32'b00000000000000001010011111010101;
assign LUT_4[24753] = 32'b00000000000000000011101011001101;
assign LUT_4[24754] = 32'b00000000000000001001111001111001;
assign LUT_4[24755] = 32'b00000000000000000011000101110001;
assign LUT_4[24756] = 32'b00000000000000000111011111110001;
assign LUT_4[24757] = 32'b00000000000000000000101011101001;
assign LUT_4[24758] = 32'b00000000000000000110111010010101;
assign LUT_4[24759] = 32'b00000000000000000000000110001101;
assign LUT_4[24760] = 32'b00000000000000000011101011101010;
assign LUT_4[24761] = 32'b11111111111111111100110111100010;
assign LUT_4[24762] = 32'b00000000000000000011000110001110;
assign LUT_4[24763] = 32'b11111111111111111100010010000110;
assign LUT_4[24764] = 32'b00000000000000000000101100000110;
assign LUT_4[24765] = 32'b11111111111111111001110111111110;
assign LUT_4[24766] = 32'b00000000000000000000000110101010;
assign LUT_4[24767] = 32'b11111111111111111001010010100010;
assign LUT_4[24768] = 32'b00000000000000001111101001110100;
assign LUT_4[24769] = 32'b00000000000000001000110101101100;
assign LUT_4[24770] = 32'b00000000000000001111000100011000;
assign LUT_4[24771] = 32'b00000000000000001000010000010000;
assign LUT_4[24772] = 32'b00000000000000001100101010010000;
assign LUT_4[24773] = 32'b00000000000000000101110110001000;
assign LUT_4[24774] = 32'b00000000000000001100000100110100;
assign LUT_4[24775] = 32'b00000000000000000101010000101100;
assign LUT_4[24776] = 32'b00000000000000001000110110001001;
assign LUT_4[24777] = 32'b00000000000000000010000010000001;
assign LUT_4[24778] = 32'b00000000000000001000010000101101;
assign LUT_4[24779] = 32'b00000000000000000001011100100101;
assign LUT_4[24780] = 32'b00000000000000000101110110100101;
assign LUT_4[24781] = 32'b11111111111111111111000010011101;
assign LUT_4[24782] = 32'b00000000000000000101010001001001;
assign LUT_4[24783] = 32'b11111111111111111110011101000001;
assign LUT_4[24784] = 32'b00000000000000001101011011100010;
assign LUT_4[24785] = 32'b00000000000000000110100111011010;
assign LUT_4[24786] = 32'b00000000000000001100110110000110;
assign LUT_4[24787] = 32'b00000000000000000110000001111110;
assign LUT_4[24788] = 32'b00000000000000001010011011111110;
assign LUT_4[24789] = 32'b00000000000000000011100111110110;
assign LUT_4[24790] = 32'b00000000000000001001110110100010;
assign LUT_4[24791] = 32'b00000000000000000011000010011010;
assign LUT_4[24792] = 32'b00000000000000000110100111110111;
assign LUT_4[24793] = 32'b11111111111111111111110011101111;
assign LUT_4[24794] = 32'b00000000000000000110000010011011;
assign LUT_4[24795] = 32'b11111111111111111111001110010011;
assign LUT_4[24796] = 32'b00000000000000000011101000010011;
assign LUT_4[24797] = 32'b11111111111111111100110100001011;
assign LUT_4[24798] = 32'b00000000000000000011000010110111;
assign LUT_4[24799] = 32'b11111111111111111100001110101111;
assign LUT_4[24800] = 32'b00000000000000001110000100111011;
assign LUT_4[24801] = 32'b00000000000000000111010000110011;
assign LUT_4[24802] = 32'b00000000000000001101011111011111;
assign LUT_4[24803] = 32'b00000000000000000110101011010111;
assign LUT_4[24804] = 32'b00000000000000001011000101010111;
assign LUT_4[24805] = 32'b00000000000000000100010001001111;
assign LUT_4[24806] = 32'b00000000000000001010011111111011;
assign LUT_4[24807] = 32'b00000000000000000011101011110011;
assign LUT_4[24808] = 32'b00000000000000000111010001010000;
assign LUT_4[24809] = 32'b00000000000000000000011101001000;
assign LUT_4[24810] = 32'b00000000000000000110101011110100;
assign LUT_4[24811] = 32'b11111111111111111111110111101100;
assign LUT_4[24812] = 32'b00000000000000000100010001101100;
assign LUT_4[24813] = 32'b11111111111111111101011101100100;
assign LUT_4[24814] = 32'b00000000000000000011101100010000;
assign LUT_4[24815] = 32'b11111111111111111100111000001000;
assign LUT_4[24816] = 32'b00000000000000001011110110101001;
assign LUT_4[24817] = 32'b00000000000000000101000010100001;
assign LUT_4[24818] = 32'b00000000000000001011010001001101;
assign LUT_4[24819] = 32'b00000000000000000100011101000101;
assign LUT_4[24820] = 32'b00000000000000001000110111000101;
assign LUT_4[24821] = 32'b00000000000000000010000010111101;
assign LUT_4[24822] = 32'b00000000000000001000010001101001;
assign LUT_4[24823] = 32'b00000000000000000001011101100001;
assign LUT_4[24824] = 32'b00000000000000000101000010111110;
assign LUT_4[24825] = 32'b11111111111111111110001110110110;
assign LUT_4[24826] = 32'b00000000000000000100011101100010;
assign LUT_4[24827] = 32'b11111111111111111101101001011010;
assign LUT_4[24828] = 32'b00000000000000000010000011011010;
assign LUT_4[24829] = 32'b11111111111111111011001111010010;
assign LUT_4[24830] = 32'b00000000000000000001011101111110;
assign LUT_4[24831] = 32'b11111111111111111010101001110110;
assign LUT_4[24832] = 32'b00000000000000010000100111111011;
assign LUT_4[24833] = 32'b00000000000000001001110011110011;
assign LUT_4[24834] = 32'b00000000000000010000000010011111;
assign LUT_4[24835] = 32'b00000000000000001001001110010111;
assign LUT_4[24836] = 32'b00000000000000001101101000010111;
assign LUT_4[24837] = 32'b00000000000000000110110100001111;
assign LUT_4[24838] = 32'b00000000000000001101000010111011;
assign LUT_4[24839] = 32'b00000000000000000110001110110011;
assign LUT_4[24840] = 32'b00000000000000001001110100010000;
assign LUT_4[24841] = 32'b00000000000000000011000000001000;
assign LUT_4[24842] = 32'b00000000000000001001001110110100;
assign LUT_4[24843] = 32'b00000000000000000010011010101100;
assign LUT_4[24844] = 32'b00000000000000000110110100101100;
assign LUT_4[24845] = 32'b00000000000000000000000000100100;
assign LUT_4[24846] = 32'b00000000000000000110001111010000;
assign LUT_4[24847] = 32'b11111111111111111111011011001000;
assign LUT_4[24848] = 32'b00000000000000001110011001101001;
assign LUT_4[24849] = 32'b00000000000000000111100101100001;
assign LUT_4[24850] = 32'b00000000000000001101110100001101;
assign LUT_4[24851] = 32'b00000000000000000111000000000101;
assign LUT_4[24852] = 32'b00000000000000001011011010000101;
assign LUT_4[24853] = 32'b00000000000000000100100101111101;
assign LUT_4[24854] = 32'b00000000000000001010110100101001;
assign LUT_4[24855] = 32'b00000000000000000100000000100001;
assign LUT_4[24856] = 32'b00000000000000000111100101111110;
assign LUT_4[24857] = 32'b00000000000000000000110001110110;
assign LUT_4[24858] = 32'b00000000000000000111000000100010;
assign LUT_4[24859] = 32'b00000000000000000000001100011010;
assign LUT_4[24860] = 32'b00000000000000000100100110011010;
assign LUT_4[24861] = 32'b11111111111111111101110010010010;
assign LUT_4[24862] = 32'b00000000000000000100000000111110;
assign LUT_4[24863] = 32'b11111111111111111101001100110110;
assign LUT_4[24864] = 32'b00000000000000001111000011000010;
assign LUT_4[24865] = 32'b00000000000000001000001110111010;
assign LUT_4[24866] = 32'b00000000000000001110011101100110;
assign LUT_4[24867] = 32'b00000000000000000111101001011110;
assign LUT_4[24868] = 32'b00000000000000001100000011011110;
assign LUT_4[24869] = 32'b00000000000000000101001111010110;
assign LUT_4[24870] = 32'b00000000000000001011011110000010;
assign LUT_4[24871] = 32'b00000000000000000100101001111010;
assign LUT_4[24872] = 32'b00000000000000001000001111010111;
assign LUT_4[24873] = 32'b00000000000000000001011011001111;
assign LUT_4[24874] = 32'b00000000000000000111101001111011;
assign LUT_4[24875] = 32'b00000000000000000000110101110011;
assign LUT_4[24876] = 32'b00000000000000000101001111110011;
assign LUT_4[24877] = 32'b11111111111111111110011011101011;
assign LUT_4[24878] = 32'b00000000000000000100101010010111;
assign LUT_4[24879] = 32'b11111111111111111101110110001111;
assign LUT_4[24880] = 32'b00000000000000001100110100110000;
assign LUT_4[24881] = 32'b00000000000000000110000000101000;
assign LUT_4[24882] = 32'b00000000000000001100001111010100;
assign LUT_4[24883] = 32'b00000000000000000101011011001100;
assign LUT_4[24884] = 32'b00000000000000001001110101001100;
assign LUT_4[24885] = 32'b00000000000000000011000001000100;
assign LUT_4[24886] = 32'b00000000000000001001001111110000;
assign LUT_4[24887] = 32'b00000000000000000010011011101000;
assign LUT_4[24888] = 32'b00000000000000000110000001000101;
assign LUT_4[24889] = 32'b11111111111111111111001100111101;
assign LUT_4[24890] = 32'b00000000000000000101011011101001;
assign LUT_4[24891] = 32'b11111111111111111110100111100001;
assign LUT_4[24892] = 32'b00000000000000000011000001100001;
assign LUT_4[24893] = 32'b11111111111111111100001101011001;
assign LUT_4[24894] = 32'b00000000000000000010011100000101;
assign LUT_4[24895] = 32'b11111111111111111011100111111101;
assign LUT_4[24896] = 32'b00000000000000010001111111001111;
assign LUT_4[24897] = 32'b00000000000000001011001011000111;
assign LUT_4[24898] = 32'b00000000000000010001011001110011;
assign LUT_4[24899] = 32'b00000000000000001010100101101011;
assign LUT_4[24900] = 32'b00000000000000001110111111101011;
assign LUT_4[24901] = 32'b00000000000000001000001011100011;
assign LUT_4[24902] = 32'b00000000000000001110011010001111;
assign LUT_4[24903] = 32'b00000000000000000111100110000111;
assign LUT_4[24904] = 32'b00000000000000001011001011100100;
assign LUT_4[24905] = 32'b00000000000000000100010111011100;
assign LUT_4[24906] = 32'b00000000000000001010100110001000;
assign LUT_4[24907] = 32'b00000000000000000011110010000000;
assign LUT_4[24908] = 32'b00000000000000001000001100000000;
assign LUT_4[24909] = 32'b00000000000000000001010111111000;
assign LUT_4[24910] = 32'b00000000000000000111100110100100;
assign LUT_4[24911] = 32'b00000000000000000000110010011100;
assign LUT_4[24912] = 32'b00000000000000001111110000111101;
assign LUT_4[24913] = 32'b00000000000000001000111100110101;
assign LUT_4[24914] = 32'b00000000000000001111001011100001;
assign LUT_4[24915] = 32'b00000000000000001000010111011001;
assign LUT_4[24916] = 32'b00000000000000001100110001011001;
assign LUT_4[24917] = 32'b00000000000000000101111101010001;
assign LUT_4[24918] = 32'b00000000000000001100001011111101;
assign LUT_4[24919] = 32'b00000000000000000101010111110101;
assign LUT_4[24920] = 32'b00000000000000001000111101010010;
assign LUT_4[24921] = 32'b00000000000000000010001001001010;
assign LUT_4[24922] = 32'b00000000000000001000010111110110;
assign LUT_4[24923] = 32'b00000000000000000001100011101110;
assign LUT_4[24924] = 32'b00000000000000000101111101101110;
assign LUT_4[24925] = 32'b11111111111111111111001001100110;
assign LUT_4[24926] = 32'b00000000000000000101011000010010;
assign LUT_4[24927] = 32'b11111111111111111110100100001010;
assign LUT_4[24928] = 32'b00000000000000010000011010010110;
assign LUT_4[24929] = 32'b00000000000000001001100110001110;
assign LUT_4[24930] = 32'b00000000000000001111110100111010;
assign LUT_4[24931] = 32'b00000000000000001001000000110010;
assign LUT_4[24932] = 32'b00000000000000001101011010110010;
assign LUT_4[24933] = 32'b00000000000000000110100110101010;
assign LUT_4[24934] = 32'b00000000000000001100110101010110;
assign LUT_4[24935] = 32'b00000000000000000110000001001110;
assign LUT_4[24936] = 32'b00000000000000001001100110101011;
assign LUT_4[24937] = 32'b00000000000000000010110010100011;
assign LUT_4[24938] = 32'b00000000000000001001000001001111;
assign LUT_4[24939] = 32'b00000000000000000010001101000111;
assign LUT_4[24940] = 32'b00000000000000000110100111000111;
assign LUT_4[24941] = 32'b11111111111111111111110010111111;
assign LUT_4[24942] = 32'b00000000000000000110000001101011;
assign LUT_4[24943] = 32'b11111111111111111111001101100011;
assign LUT_4[24944] = 32'b00000000000000001110001100000100;
assign LUT_4[24945] = 32'b00000000000000000111010111111100;
assign LUT_4[24946] = 32'b00000000000000001101100110101000;
assign LUT_4[24947] = 32'b00000000000000000110110010100000;
assign LUT_4[24948] = 32'b00000000000000001011001100100000;
assign LUT_4[24949] = 32'b00000000000000000100011000011000;
assign LUT_4[24950] = 32'b00000000000000001010100111000100;
assign LUT_4[24951] = 32'b00000000000000000011110010111100;
assign LUT_4[24952] = 32'b00000000000000000111011000011001;
assign LUT_4[24953] = 32'b00000000000000000000100100010001;
assign LUT_4[24954] = 32'b00000000000000000110110010111101;
assign LUT_4[24955] = 32'b11111111111111111111111110110101;
assign LUT_4[24956] = 32'b00000000000000000100011000110101;
assign LUT_4[24957] = 32'b11111111111111111101100100101101;
assign LUT_4[24958] = 32'b00000000000000000011110011011001;
assign LUT_4[24959] = 32'b11111111111111111100111111010001;
assign LUT_4[24960] = 32'b00000000000000010011001110000011;
assign LUT_4[24961] = 32'b00000000000000001100011001111011;
assign LUT_4[24962] = 32'b00000000000000010010101000100111;
assign LUT_4[24963] = 32'b00000000000000001011110100011111;
assign LUT_4[24964] = 32'b00000000000000010000001110011111;
assign LUT_4[24965] = 32'b00000000000000001001011010010111;
assign LUT_4[24966] = 32'b00000000000000001111101001000011;
assign LUT_4[24967] = 32'b00000000000000001000110100111011;
assign LUT_4[24968] = 32'b00000000000000001100011010011000;
assign LUT_4[24969] = 32'b00000000000000000101100110010000;
assign LUT_4[24970] = 32'b00000000000000001011110100111100;
assign LUT_4[24971] = 32'b00000000000000000101000000110100;
assign LUT_4[24972] = 32'b00000000000000001001011010110100;
assign LUT_4[24973] = 32'b00000000000000000010100110101100;
assign LUT_4[24974] = 32'b00000000000000001000110101011000;
assign LUT_4[24975] = 32'b00000000000000000010000001010000;
assign LUT_4[24976] = 32'b00000000000000010000111111110001;
assign LUT_4[24977] = 32'b00000000000000001010001011101001;
assign LUT_4[24978] = 32'b00000000000000010000011010010101;
assign LUT_4[24979] = 32'b00000000000000001001100110001101;
assign LUT_4[24980] = 32'b00000000000000001110000000001101;
assign LUT_4[24981] = 32'b00000000000000000111001100000101;
assign LUT_4[24982] = 32'b00000000000000001101011010110001;
assign LUT_4[24983] = 32'b00000000000000000110100110101001;
assign LUT_4[24984] = 32'b00000000000000001010001100000110;
assign LUT_4[24985] = 32'b00000000000000000011010111111110;
assign LUT_4[24986] = 32'b00000000000000001001100110101010;
assign LUT_4[24987] = 32'b00000000000000000010110010100010;
assign LUT_4[24988] = 32'b00000000000000000111001100100010;
assign LUT_4[24989] = 32'b00000000000000000000011000011010;
assign LUT_4[24990] = 32'b00000000000000000110100111000110;
assign LUT_4[24991] = 32'b11111111111111111111110010111110;
assign LUT_4[24992] = 32'b00000000000000010001101001001010;
assign LUT_4[24993] = 32'b00000000000000001010110101000010;
assign LUT_4[24994] = 32'b00000000000000010001000011101110;
assign LUT_4[24995] = 32'b00000000000000001010001111100110;
assign LUT_4[24996] = 32'b00000000000000001110101001100110;
assign LUT_4[24997] = 32'b00000000000000000111110101011110;
assign LUT_4[24998] = 32'b00000000000000001110000100001010;
assign LUT_4[24999] = 32'b00000000000000000111010000000010;
assign LUT_4[25000] = 32'b00000000000000001010110101011111;
assign LUT_4[25001] = 32'b00000000000000000100000001010111;
assign LUT_4[25002] = 32'b00000000000000001010010000000011;
assign LUT_4[25003] = 32'b00000000000000000011011011111011;
assign LUT_4[25004] = 32'b00000000000000000111110101111011;
assign LUT_4[25005] = 32'b00000000000000000001000001110011;
assign LUT_4[25006] = 32'b00000000000000000111010000011111;
assign LUT_4[25007] = 32'b00000000000000000000011100010111;
assign LUT_4[25008] = 32'b00000000000000001111011010111000;
assign LUT_4[25009] = 32'b00000000000000001000100110110000;
assign LUT_4[25010] = 32'b00000000000000001110110101011100;
assign LUT_4[25011] = 32'b00000000000000001000000001010100;
assign LUT_4[25012] = 32'b00000000000000001100011011010100;
assign LUT_4[25013] = 32'b00000000000000000101100111001100;
assign LUT_4[25014] = 32'b00000000000000001011110101111000;
assign LUT_4[25015] = 32'b00000000000000000101000001110000;
assign LUT_4[25016] = 32'b00000000000000001000100111001101;
assign LUT_4[25017] = 32'b00000000000000000001110011000101;
assign LUT_4[25018] = 32'b00000000000000001000000001110001;
assign LUT_4[25019] = 32'b00000000000000000001001101101001;
assign LUT_4[25020] = 32'b00000000000000000101100111101001;
assign LUT_4[25021] = 32'b11111111111111111110110011100001;
assign LUT_4[25022] = 32'b00000000000000000101000010001101;
assign LUT_4[25023] = 32'b11111111111111111110001110000101;
assign LUT_4[25024] = 32'b00000000000000010100100101010111;
assign LUT_4[25025] = 32'b00000000000000001101110001001111;
assign LUT_4[25026] = 32'b00000000000000010011111111111011;
assign LUT_4[25027] = 32'b00000000000000001101001011110011;
assign LUT_4[25028] = 32'b00000000000000010001100101110011;
assign LUT_4[25029] = 32'b00000000000000001010110001101011;
assign LUT_4[25030] = 32'b00000000000000010001000000010111;
assign LUT_4[25031] = 32'b00000000000000001010001100001111;
assign LUT_4[25032] = 32'b00000000000000001101110001101100;
assign LUT_4[25033] = 32'b00000000000000000110111101100100;
assign LUT_4[25034] = 32'b00000000000000001101001100010000;
assign LUT_4[25035] = 32'b00000000000000000110011000001000;
assign LUT_4[25036] = 32'b00000000000000001010110010001000;
assign LUT_4[25037] = 32'b00000000000000000011111110000000;
assign LUT_4[25038] = 32'b00000000000000001010001100101100;
assign LUT_4[25039] = 32'b00000000000000000011011000100100;
assign LUT_4[25040] = 32'b00000000000000010010010111000101;
assign LUT_4[25041] = 32'b00000000000000001011100010111101;
assign LUT_4[25042] = 32'b00000000000000010001110001101001;
assign LUT_4[25043] = 32'b00000000000000001010111101100001;
assign LUT_4[25044] = 32'b00000000000000001111010111100001;
assign LUT_4[25045] = 32'b00000000000000001000100011011001;
assign LUT_4[25046] = 32'b00000000000000001110110010000101;
assign LUT_4[25047] = 32'b00000000000000000111111101111101;
assign LUT_4[25048] = 32'b00000000000000001011100011011010;
assign LUT_4[25049] = 32'b00000000000000000100101111010010;
assign LUT_4[25050] = 32'b00000000000000001010111101111110;
assign LUT_4[25051] = 32'b00000000000000000100001001110110;
assign LUT_4[25052] = 32'b00000000000000001000100011110110;
assign LUT_4[25053] = 32'b00000000000000000001101111101110;
assign LUT_4[25054] = 32'b00000000000000000111111110011010;
assign LUT_4[25055] = 32'b00000000000000000001001010010010;
assign LUT_4[25056] = 32'b00000000000000010011000000011110;
assign LUT_4[25057] = 32'b00000000000000001100001100010110;
assign LUT_4[25058] = 32'b00000000000000010010011011000010;
assign LUT_4[25059] = 32'b00000000000000001011100110111010;
assign LUT_4[25060] = 32'b00000000000000010000000000111010;
assign LUT_4[25061] = 32'b00000000000000001001001100110010;
assign LUT_4[25062] = 32'b00000000000000001111011011011110;
assign LUT_4[25063] = 32'b00000000000000001000100111010110;
assign LUT_4[25064] = 32'b00000000000000001100001100110011;
assign LUT_4[25065] = 32'b00000000000000000101011000101011;
assign LUT_4[25066] = 32'b00000000000000001011100111010111;
assign LUT_4[25067] = 32'b00000000000000000100110011001111;
assign LUT_4[25068] = 32'b00000000000000001001001101001111;
assign LUT_4[25069] = 32'b00000000000000000010011001000111;
assign LUT_4[25070] = 32'b00000000000000001000100111110011;
assign LUT_4[25071] = 32'b00000000000000000001110011101011;
assign LUT_4[25072] = 32'b00000000000000010000110010001100;
assign LUT_4[25073] = 32'b00000000000000001001111110000100;
assign LUT_4[25074] = 32'b00000000000000010000001100110000;
assign LUT_4[25075] = 32'b00000000000000001001011000101000;
assign LUT_4[25076] = 32'b00000000000000001101110010101000;
assign LUT_4[25077] = 32'b00000000000000000110111110100000;
assign LUT_4[25078] = 32'b00000000000000001101001101001100;
assign LUT_4[25079] = 32'b00000000000000000110011001000100;
assign LUT_4[25080] = 32'b00000000000000001001111110100001;
assign LUT_4[25081] = 32'b00000000000000000011001010011001;
assign LUT_4[25082] = 32'b00000000000000001001011001000101;
assign LUT_4[25083] = 32'b00000000000000000010100100111101;
assign LUT_4[25084] = 32'b00000000000000000110111110111101;
assign LUT_4[25085] = 32'b00000000000000000000001010110101;
assign LUT_4[25086] = 32'b00000000000000000110011001100001;
assign LUT_4[25087] = 32'b11111111111111111111100101011001;
assign LUT_4[25088] = 32'b00000000000000001010110000100000;
assign LUT_4[25089] = 32'b00000000000000000011111100011000;
assign LUT_4[25090] = 32'b00000000000000001010001011000100;
assign LUT_4[25091] = 32'b00000000000000000011010110111100;
assign LUT_4[25092] = 32'b00000000000000000111110000111100;
assign LUT_4[25093] = 32'b00000000000000000000111100110100;
assign LUT_4[25094] = 32'b00000000000000000111001011100000;
assign LUT_4[25095] = 32'b00000000000000000000010111011000;
assign LUT_4[25096] = 32'b00000000000000000011111100110101;
assign LUT_4[25097] = 32'b11111111111111111101001000101101;
assign LUT_4[25098] = 32'b00000000000000000011010111011001;
assign LUT_4[25099] = 32'b11111111111111111100100011010001;
assign LUT_4[25100] = 32'b00000000000000000000111101010001;
assign LUT_4[25101] = 32'b11111111111111111010001001001001;
assign LUT_4[25102] = 32'b00000000000000000000010111110101;
assign LUT_4[25103] = 32'b11111111111111111001100011101101;
assign LUT_4[25104] = 32'b00000000000000001000100010001110;
assign LUT_4[25105] = 32'b00000000000000000001101110000110;
assign LUT_4[25106] = 32'b00000000000000000111111100110010;
assign LUT_4[25107] = 32'b00000000000000000001001000101010;
assign LUT_4[25108] = 32'b00000000000000000101100010101010;
assign LUT_4[25109] = 32'b11111111111111111110101110100010;
assign LUT_4[25110] = 32'b00000000000000000100111101001110;
assign LUT_4[25111] = 32'b11111111111111111110001001000110;
assign LUT_4[25112] = 32'b00000000000000000001101110100011;
assign LUT_4[25113] = 32'b11111111111111111010111010011011;
assign LUT_4[25114] = 32'b00000000000000000001001001000111;
assign LUT_4[25115] = 32'b11111111111111111010010100111111;
assign LUT_4[25116] = 32'b11111111111111111110101110111111;
assign LUT_4[25117] = 32'b11111111111111110111111010110111;
assign LUT_4[25118] = 32'b11111111111111111110001001100011;
assign LUT_4[25119] = 32'b11111111111111110111010101011011;
assign LUT_4[25120] = 32'b00000000000000001001001011100111;
assign LUT_4[25121] = 32'b00000000000000000010010111011111;
assign LUT_4[25122] = 32'b00000000000000001000100110001011;
assign LUT_4[25123] = 32'b00000000000000000001110010000011;
assign LUT_4[25124] = 32'b00000000000000000110001100000011;
assign LUT_4[25125] = 32'b11111111111111111111010111111011;
assign LUT_4[25126] = 32'b00000000000000000101100110100111;
assign LUT_4[25127] = 32'b11111111111111111110110010011111;
assign LUT_4[25128] = 32'b00000000000000000010010111111100;
assign LUT_4[25129] = 32'b11111111111111111011100011110100;
assign LUT_4[25130] = 32'b00000000000000000001110010100000;
assign LUT_4[25131] = 32'b11111111111111111010111110011000;
assign LUT_4[25132] = 32'b11111111111111111111011000011000;
assign LUT_4[25133] = 32'b11111111111111111000100100010000;
assign LUT_4[25134] = 32'b11111111111111111110110010111100;
assign LUT_4[25135] = 32'b11111111111111110111111110110100;
assign LUT_4[25136] = 32'b00000000000000000110111101010101;
assign LUT_4[25137] = 32'b00000000000000000000001001001101;
assign LUT_4[25138] = 32'b00000000000000000110010111111001;
assign LUT_4[25139] = 32'b11111111111111111111100011110001;
assign LUT_4[25140] = 32'b00000000000000000011111101110001;
assign LUT_4[25141] = 32'b11111111111111111101001001101001;
assign LUT_4[25142] = 32'b00000000000000000011011000010101;
assign LUT_4[25143] = 32'b11111111111111111100100100001101;
assign LUT_4[25144] = 32'b00000000000000000000001001101010;
assign LUT_4[25145] = 32'b11111111111111111001010101100010;
assign LUT_4[25146] = 32'b11111111111111111111100100001110;
assign LUT_4[25147] = 32'b11111111111111111000110000000110;
assign LUT_4[25148] = 32'b11111111111111111101001010000110;
assign LUT_4[25149] = 32'b11111111111111110110010101111110;
assign LUT_4[25150] = 32'b11111111111111111100100100101010;
assign LUT_4[25151] = 32'b11111111111111110101110000100010;
assign LUT_4[25152] = 32'b00000000000000001100000111110100;
assign LUT_4[25153] = 32'b00000000000000000101010011101100;
assign LUT_4[25154] = 32'b00000000000000001011100010011000;
assign LUT_4[25155] = 32'b00000000000000000100101110010000;
assign LUT_4[25156] = 32'b00000000000000001001001000010000;
assign LUT_4[25157] = 32'b00000000000000000010010100001000;
assign LUT_4[25158] = 32'b00000000000000001000100010110100;
assign LUT_4[25159] = 32'b00000000000000000001101110101100;
assign LUT_4[25160] = 32'b00000000000000000101010100001001;
assign LUT_4[25161] = 32'b11111111111111111110100000000001;
assign LUT_4[25162] = 32'b00000000000000000100101110101101;
assign LUT_4[25163] = 32'b11111111111111111101111010100101;
assign LUT_4[25164] = 32'b00000000000000000010010100100101;
assign LUT_4[25165] = 32'b11111111111111111011100000011101;
assign LUT_4[25166] = 32'b00000000000000000001101111001001;
assign LUT_4[25167] = 32'b11111111111111111010111011000001;
assign LUT_4[25168] = 32'b00000000000000001001111001100010;
assign LUT_4[25169] = 32'b00000000000000000011000101011010;
assign LUT_4[25170] = 32'b00000000000000001001010100000110;
assign LUT_4[25171] = 32'b00000000000000000010011111111110;
assign LUT_4[25172] = 32'b00000000000000000110111001111110;
assign LUT_4[25173] = 32'b00000000000000000000000101110110;
assign LUT_4[25174] = 32'b00000000000000000110010100100010;
assign LUT_4[25175] = 32'b11111111111111111111100000011010;
assign LUT_4[25176] = 32'b00000000000000000011000101110111;
assign LUT_4[25177] = 32'b11111111111111111100010001101111;
assign LUT_4[25178] = 32'b00000000000000000010100000011011;
assign LUT_4[25179] = 32'b11111111111111111011101100010011;
assign LUT_4[25180] = 32'b00000000000000000000000110010011;
assign LUT_4[25181] = 32'b11111111111111111001010010001011;
assign LUT_4[25182] = 32'b11111111111111111111100000110111;
assign LUT_4[25183] = 32'b11111111111111111000101100101111;
assign LUT_4[25184] = 32'b00000000000000001010100010111011;
assign LUT_4[25185] = 32'b00000000000000000011101110110011;
assign LUT_4[25186] = 32'b00000000000000001001111101011111;
assign LUT_4[25187] = 32'b00000000000000000011001001010111;
assign LUT_4[25188] = 32'b00000000000000000111100011010111;
assign LUT_4[25189] = 32'b00000000000000000000101111001111;
assign LUT_4[25190] = 32'b00000000000000000110111101111011;
assign LUT_4[25191] = 32'b00000000000000000000001001110011;
assign LUT_4[25192] = 32'b00000000000000000011101111010000;
assign LUT_4[25193] = 32'b11111111111111111100111011001000;
assign LUT_4[25194] = 32'b00000000000000000011001001110100;
assign LUT_4[25195] = 32'b11111111111111111100010101101100;
assign LUT_4[25196] = 32'b00000000000000000000101111101100;
assign LUT_4[25197] = 32'b11111111111111111001111011100100;
assign LUT_4[25198] = 32'b00000000000000000000001010010000;
assign LUT_4[25199] = 32'b11111111111111111001010110001000;
assign LUT_4[25200] = 32'b00000000000000001000010100101001;
assign LUT_4[25201] = 32'b00000000000000000001100000100001;
assign LUT_4[25202] = 32'b00000000000000000111101111001101;
assign LUT_4[25203] = 32'b00000000000000000000111011000101;
assign LUT_4[25204] = 32'b00000000000000000101010101000101;
assign LUT_4[25205] = 32'b11111111111111111110100000111101;
assign LUT_4[25206] = 32'b00000000000000000100101111101001;
assign LUT_4[25207] = 32'b11111111111111111101111011100001;
assign LUT_4[25208] = 32'b00000000000000000001100000111110;
assign LUT_4[25209] = 32'b11111111111111111010101100110110;
assign LUT_4[25210] = 32'b00000000000000000000111011100010;
assign LUT_4[25211] = 32'b11111111111111111010000111011010;
assign LUT_4[25212] = 32'b11111111111111111110100001011010;
assign LUT_4[25213] = 32'b11111111111111110111101101010010;
assign LUT_4[25214] = 32'b11111111111111111101111011111110;
assign LUT_4[25215] = 32'b11111111111111110111000111110110;
assign LUT_4[25216] = 32'b00000000000000001101010110101000;
assign LUT_4[25217] = 32'b00000000000000000110100010100000;
assign LUT_4[25218] = 32'b00000000000000001100110001001100;
assign LUT_4[25219] = 32'b00000000000000000101111101000100;
assign LUT_4[25220] = 32'b00000000000000001010010111000100;
assign LUT_4[25221] = 32'b00000000000000000011100010111100;
assign LUT_4[25222] = 32'b00000000000000001001110001101000;
assign LUT_4[25223] = 32'b00000000000000000010111101100000;
assign LUT_4[25224] = 32'b00000000000000000110100010111101;
assign LUT_4[25225] = 32'b11111111111111111111101110110101;
assign LUT_4[25226] = 32'b00000000000000000101111101100001;
assign LUT_4[25227] = 32'b11111111111111111111001001011001;
assign LUT_4[25228] = 32'b00000000000000000011100011011001;
assign LUT_4[25229] = 32'b11111111111111111100101111010001;
assign LUT_4[25230] = 32'b00000000000000000010111101111101;
assign LUT_4[25231] = 32'b11111111111111111100001001110101;
assign LUT_4[25232] = 32'b00000000000000001011001000010110;
assign LUT_4[25233] = 32'b00000000000000000100010100001110;
assign LUT_4[25234] = 32'b00000000000000001010100010111010;
assign LUT_4[25235] = 32'b00000000000000000011101110110010;
assign LUT_4[25236] = 32'b00000000000000001000001000110010;
assign LUT_4[25237] = 32'b00000000000000000001010100101010;
assign LUT_4[25238] = 32'b00000000000000000111100011010110;
assign LUT_4[25239] = 32'b00000000000000000000101111001110;
assign LUT_4[25240] = 32'b00000000000000000100010100101011;
assign LUT_4[25241] = 32'b11111111111111111101100000100011;
assign LUT_4[25242] = 32'b00000000000000000011101111001111;
assign LUT_4[25243] = 32'b11111111111111111100111011000111;
assign LUT_4[25244] = 32'b00000000000000000001010101000111;
assign LUT_4[25245] = 32'b11111111111111111010100000111111;
assign LUT_4[25246] = 32'b00000000000000000000101111101011;
assign LUT_4[25247] = 32'b11111111111111111001111011100011;
assign LUT_4[25248] = 32'b00000000000000001011110001101111;
assign LUT_4[25249] = 32'b00000000000000000100111101100111;
assign LUT_4[25250] = 32'b00000000000000001011001100010011;
assign LUT_4[25251] = 32'b00000000000000000100011000001011;
assign LUT_4[25252] = 32'b00000000000000001000110010001011;
assign LUT_4[25253] = 32'b00000000000000000001111110000011;
assign LUT_4[25254] = 32'b00000000000000001000001100101111;
assign LUT_4[25255] = 32'b00000000000000000001011000100111;
assign LUT_4[25256] = 32'b00000000000000000100111110000100;
assign LUT_4[25257] = 32'b11111111111111111110001001111100;
assign LUT_4[25258] = 32'b00000000000000000100011000101000;
assign LUT_4[25259] = 32'b11111111111111111101100100100000;
assign LUT_4[25260] = 32'b00000000000000000001111110100000;
assign LUT_4[25261] = 32'b11111111111111111011001010011000;
assign LUT_4[25262] = 32'b00000000000000000001011001000100;
assign LUT_4[25263] = 32'b11111111111111111010100100111100;
assign LUT_4[25264] = 32'b00000000000000001001100011011101;
assign LUT_4[25265] = 32'b00000000000000000010101111010101;
assign LUT_4[25266] = 32'b00000000000000001000111110000001;
assign LUT_4[25267] = 32'b00000000000000000010001001111001;
assign LUT_4[25268] = 32'b00000000000000000110100011111001;
assign LUT_4[25269] = 32'b11111111111111111111101111110001;
assign LUT_4[25270] = 32'b00000000000000000101111110011101;
assign LUT_4[25271] = 32'b11111111111111111111001010010101;
assign LUT_4[25272] = 32'b00000000000000000010101111110010;
assign LUT_4[25273] = 32'b11111111111111111011111011101010;
assign LUT_4[25274] = 32'b00000000000000000010001010010110;
assign LUT_4[25275] = 32'b11111111111111111011010110001110;
assign LUT_4[25276] = 32'b11111111111111111111110000001110;
assign LUT_4[25277] = 32'b11111111111111111000111100000110;
assign LUT_4[25278] = 32'b11111111111111111111001010110010;
assign LUT_4[25279] = 32'b11111111111111111000010110101010;
assign LUT_4[25280] = 32'b00000000000000001110101101111100;
assign LUT_4[25281] = 32'b00000000000000000111111001110100;
assign LUT_4[25282] = 32'b00000000000000001110001000100000;
assign LUT_4[25283] = 32'b00000000000000000111010100011000;
assign LUT_4[25284] = 32'b00000000000000001011101110011000;
assign LUT_4[25285] = 32'b00000000000000000100111010010000;
assign LUT_4[25286] = 32'b00000000000000001011001000111100;
assign LUT_4[25287] = 32'b00000000000000000100010100110100;
assign LUT_4[25288] = 32'b00000000000000000111111010010001;
assign LUT_4[25289] = 32'b00000000000000000001000110001001;
assign LUT_4[25290] = 32'b00000000000000000111010100110101;
assign LUT_4[25291] = 32'b00000000000000000000100000101101;
assign LUT_4[25292] = 32'b00000000000000000100111010101101;
assign LUT_4[25293] = 32'b11111111111111111110000110100101;
assign LUT_4[25294] = 32'b00000000000000000100010101010001;
assign LUT_4[25295] = 32'b11111111111111111101100001001001;
assign LUT_4[25296] = 32'b00000000000000001100011111101010;
assign LUT_4[25297] = 32'b00000000000000000101101011100010;
assign LUT_4[25298] = 32'b00000000000000001011111010001110;
assign LUT_4[25299] = 32'b00000000000000000101000110000110;
assign LUT_4[25300] = 32'b00000000000000001001100000000110;
assign LUT_4[25301] = 32'b00000000000000000010101011111110;
assign LUT_4[25302] = 32'b00000000000000001000111010101010;
assign LUT_4[25303] = 32'b00000000000000000010000110100010;
assign LUT_4[25304] = 32'b00000000000000000101101011111111;
assign LUT_4[25305] = 32'b11111111111111111110110111110111;
assign LUT_4[25306] = 32'b00000000000000000101000110100011;
assign LUT_4[25307] = 32'b11111111111111111110010010011011;
assign LUT_4[25308] = 32'b00000000000000000010101100011011;
assign LUT_4[25309] = 32'b11111111111111111011111000010011;
assign LUT_4[25310] = 32'b00000000000000000010000110111111;
assign LUT_4[25311] = 32'b11111111111111111011010010110111;
assign LUT_4[25312] = 32'b00000000000000001101001001000011;
assign LUT_4[25313] = 32'b00000000000000000110010100111011;
assign LUT_4[25314] = 32'b00000000000000001100100011100111;
assign LUT_4[25315] = 32'b00000000000000000101101111011111;
assign LUT_4[25316] = 32'b00000000000000001010001001011111;
assign LUT_4[25317] = 32'b00000000000000000011010101010111;
assign LUT_4[25318] = 32'b00000000000000001001100100000011;
assign LUT_4[25319] = 32'b00000000000000000010101111111011;
assign LUT_4[25320] = 32'b00000000000000000110010101011000;
assign LUT_4[25321] = 32'b11111111111111111111100001010000;
assign LUT_4[25322] = 32'b00000000000000000101101111111100;
assign LUT_4[25323] = 32'b11111111111111111110111011110100;
assign LUT_4[25324] = 32'b00000000000000000011010101110100;
assign LUT_4[25325] = 32'b11111111111111111100100001101100;
assign LUT_4[25326] = 32'b00000000000000000010110000011000;
assign LUT_4[25327] = 32'b11111111111111111011111100010000;
assign LUT_4[25328] = 32'b00000000000000001010111010110001;
assign LUT_4[25329] = 32'b00000000000000000100000110101001;
assign LUT_4[25330] = 32'b00000000000000001010010101010101;
assign LUT_4[25331] = 32'b00000000000000000011100001001101;
assign LUT_4[25332] = 32'b00000000000000000111111011001101;
assign LUT_4[25333] = 32'b00000000000000000001000111000101;
assign LUT_4[25334] = 32'b00000000000000000111010101110001;
assign LUT_4[25335] = 32'b00000000000000000000100001101001;
assign LUT_4[25336] = 32'b00000000000000000100000111000110;
assign LUT_4[25337] = 32'b11111111111111111101010010111110;
assign LUT_4[25338] = 32'b00000000000000000011100001101010;
assign LUT_4[25339] = 32'b11111111111111111100101101100010;
assign LUT_4[25340] = 32'b00000000000000000001000111100010;
assign LUT_4[25341] = 32'b11111111111111111010010011011010;
assign LUT_4[25342] = 32'b00000000000000000000100010000110;
assign LUT_4[25343] = 32'b11111111111111111001101101111110;
assign LUT_4[25344] = 32'b00000000000000001111101100000011;
assign LUT_4[25345] = 32'b00000000000000001000110111111011;
assign LUT_4[25346] = 32'b00000000000000001111000110100111;
assign LUT_4[25347] = 32'b00000000000000001000010010011111;
assign LUT_4[25348] = 32'b00000000000000001100101100011111;
assign LUT_4[25349] = 32'b00000000000000000101111000010111;
assign LUT_4[25350] = 32'b00000000000000001100000111000011;
assign LUT_4[25351] = 32'b00000000000000000101010010111011;
assign LUT_4[25352] = 32'b00000000000000001000111000011000;
assign LUT_4[25353] = 32'b00000000000000000010000100010000;
assign LUT_4[25354] = 32'b00000000000000001000010010111100;
assign LUT_4[25355] = 32'b00000000000000000001011110110100;
assign LUT_4[25356] = 32'b00000000000000000101111000110100;
assign LUT_4[25357] = 32'b11111111111111111111000100101100;
assign LUT_4[25358] = 32'b00000000000000000101010011011000;
assign LUT_4[25359] = 32'b11111111111111111110011111010000;
assign LUT_4[25360] = 32'b00000000000000001101011101110001;
assign LUT_4[25361] = 32'b00000000000000000110101001101001;
assign LUT_4[25362] = 32'b00000000000000001100111000010101;
assign LUT_4[25363] = 32'b00000000000000000110000100001101;
assign LUT_4[25364] = 32'b00000000000000001010011110001101;
assign LUT_4[25365] = 32'b00000000000000000011101010000101;
assign LUT_4[25366] = 32'b00000000000000001001111000110001;
assign LUT_4[25367] = 32'b00000000000000000011000100101001;
assign LUT_4[25368] = 32'b00000000000000000110101010000110;
assign LUT_4[25369] = 32'b11111111111111111111110101111110;
assign LUT_4[25370] = 32'b00000000000000000110000100101010;
assign LUT_4[25371] = 32'b11111111111111111111010000100010;
assign LUT_4[25372] = 32'b00000000000000000011101010100010;
assign LUT_4[25373] = 32'b11111111111111111100110110011010;
assign LUT_4[25374] = 32'b00000000000000000011000101000110;
assign LUT_4[25375] = 32'b11111111111111111100010000111110;
assign LUT_4[25376] = 32'b00000000000000001110000111001010;
assign LUT_4[25377] = 32'b00000000000000000111010011000010;
assign LUT_4[25378] = 32'b00000000000000001101100001101110;
assign LUT_4[25379] = 32'b00000000000000000110101101100110;
assign LUT_4[25380] = 32'b00000000000000001011000111100110;
assign LUT_4[25381] = 32'b00000000000000000100010011011110;
assign LUT_4[25382] = 32'b00000000000000001010100010001010;
assign LUT_4[25383] = 32'b00000000000000000011101110000010;
assign LUT_4[25384] = 32'b00000000000000000111010011011111;
assign LUT_4[25385] = 32'b00000000000000000000011111010111;
assign LUT_4[25386] = 32'b00000000000000000110101110000011;
assign LUT_4[25387] = 32'b11111111111111111111111001111011;
assign LUT_4[25388] = 32'b00000000000000000100010011111011;
assign LUT_4[25389] = 32'b11111111111111111101011111110011;
assign LUT_4[25390] = 32'b00000000000000000011101110011111;
assign LUT_4[25391] = 32'b11111111111111111100111010010111;
assign LUT_4[25392] = 32'b00000000000000001011111000111000;
assign LUT_4[25393] = 32'b00000000000000000101000100110000;
assign LUT_4[25394] = 32'b00000000000000001011010011011100;
assign LUT_4[25395] = 32'b00000000000000000100011111010100;
assign LUT_4[25396] = 32'b00000000000000001000111001010100;
assign LUT_4[25397] = 32'b00000000000000000010000101001100;
assign LUT_4[25398] = 32'b00000000000000001000010011111000;
assign LUT_4[25399] = 32'b00000000000000000001011111110000;
assign LUT_4[25400] = 32'b00000000000000000101000101001101;
assign LUT_4[25401] = 32'b11111111111111111110010001000101;
assign LUT_4[25402] = 32'b00000000000000000100011111110001;
assign LUT_4[25403] = 32'b11111111111111111101101011101001;
assign LUT_4[25404] = 32'b00000000000000000010000101101001;
assign LUT_4[25405] = 32'b11111111111111111011010001100001;
assign LUT_4[25406] = 32'b00000000000000000001100000001101;
assign LUT_4[25407] = 32'b11111111111111111010101100000101;
assign LUT_4[25408] = 32'b00000000000000010001000011010111;
assign LUT_4[25409] = 32'b00000000000000001010001111001111;
assign LUT_4[25410] = 32'b00000000000000010000011101111011;
assign LUT_4[25411] = 32'b00000000000000001001101001110011;
assign LUT_4[25412] = 32'b00000000000000001110000011110011;
assign LUT_4[25413] = 32'b00000000000000000111001111101011;
assign LUT_4[25414] = 32'b00000000000000001101011110010111;
assign LUT_4[25415] = 32'b00000000000000000110101010001111;
assign LUT_4[25416] = 32'b00000000000000001010001111101100;
assign LUT_4[25417] = 32'b00000000000000000011011011100100;
assign LUT_4[25418] = 32'b00000000000000001001101010010000;
assign LUT_4[25419] = 32'b00000000000000000010110110001000;
assign LUT_4[25420] = 32'b00000000000000000111010000001000;
assign LUT_4[25421] = 32'b00000000000000000000011100000000;
assign LUT_4[25422] = 32'b00000000000000000110101010101100;
assign LUT_4[25423] = 32'b11111111111111111111110110100100;
assign LUT_4[25424] = 32'b00000000000000001110110101000101;
assign LUT_4[25425] = 32'b00000000000000001000000000111101;
assign LUT_4[25426] = 32'b00000000000000001110001111101001;
assign LUT_4[25427] = 32'b00000000000000000111011011100001;
assign LUT_4[25428] = 32'b00000000000000001011110101100001;
assign LUT_4[25429] = 32'b00000000000000000101000001011001;
assign LUT_4[25430] = 32'b00000000000000001011010000000101;
assign LUT_4[25431] = 32'b00000000000000000100011011111101;
assign LUT_4[25432] = 32'b00000000000000001000000001011010;
assign LUT_4[25433] = 32'b00000000000000000001001101010010;
assign LUT_4[25434] = 32'b00000000000000000111011011111110;
assign LUT_4[25435] = 32'b00000000000000000000100111110110;
assign LUT_4[25436] = 32'b00000000000000000101000001110110;
assign LUT_4[25437] = 32'b11111111111111111110001101101110;
assign LUT_4[25438] = 32'b00000000000000000100011100011010;
assign LUT_4[25439] = 32'b11111111111111111101101000010010;
assign LUT_4[25440] = 32'b00000000000000001111011110011110;
assign LUT_4[25441] = 32'b00000000000000001000101010010110;
assign LUT_4[25442] = 32'b00000000000000001110111001000010;
assign LUT_4[25443] = 32'b00000000000000001000000100111010;
assign LUT_4[25444] = 32'b00000000000000001100011110111010;
assign LUT_4[25445] = 32'b00000000000000000101101010110010;
assign LUT_4[25446] = 32'b00000000000000001011111001011110;
assign LUT_4[25447] = 32'b00000000000000000101000101010110;
assign LUT_4[25448] = 32'b00000000000000001000101010110011;
assign LUT_4[25449] = 32'b00000000000000000001110110101011;
assign LUT_4[25450] = 32'b00000000000000001000000101010111;
assign LUT_4[25451] = 32'b00000000000000000001010001001111;
assign LUT_4[25452] = 32'b00000000000000000101101011001111;
assign LUT_4[25453] = 32'b11111111111111111110110111000111;
assign LUT_4[25454] = 32'b00000000000000000101000101110011;
assign LUT_4[25455] = 32'b11111111111111111110010001101011;
assign LUT_4[25456] = 32'b00000000000000001101010000001100;
assign LUT_4[25457] = 32'b00000000000000000110011100000100;
assign LUT_4[25458] = 32'b00000000000000001100101010110000;
assign LUT_4[25459] = 32'b00000000000000000101110110101000;
assign LUT_4[25460] = 32'b00000000000000001010010000101000;
assign LUT_4[25461] = 32'b00000000000000000011011100100000;
assign LUT_4[25462] = 32'b00000000000000001001101011001100;
assign LUT_4[25463] = 32'b00000000000000000010110111000100;
assign LUT_4[25464] = 32'b00000000000000000110011100100001;
assign LUT_4[25465] = 32'b11111111111111111111101000011001;
assign LUT_4[25466] = 32'b00000000000000000101110111000101;
assign LUT_4[25467] = 32'b11111111111111111111000010111101;
assign LUT_4[25468] = 32'b00000000000000000011011100111101;
assign LUT_4[25469] = 32'b11111111111111111100101000110101;
assign LUT_4[25470] = 32'b00000000000000000010110111100001;
assign LUT_4[25471] = 32'b11111111111111111100000011011001;
assign LUT_4[25472] = 32'b00000000000000010010010010001011;
assign LUT_4[25473] = 32'b00000000000000001011011110000011;
assign LUT_4[25474] = 32'b00000000000000010001101100101111;
assign LUT_4[25475] = 32'b00000000000000001010111000100111;
assign LUT_4[25476] = 32'b00000000000000001111010010100111;
assign LUT_4[25477] = 32'b00000000000000001000011110011111;
assign LUT_4[25478] = 32'b00000000000000001110101101001011;
assign LUT_4[25479] = 32'b00000000000000000111111001000011;
assign LUT_4[25480] = 32'b00000000000000001011011110100000;
assign LUT_4[25481] = 32'b00000000000000000100101010011000;
assign LUT_4[25482] = 32'b00000000000000001010111001000100;
assign LUT_4[25483] = 32'b00000000000000000100000100111100;
assign LUT_4[25484] = 32'b00000000000000001000011110111100;
assign LUT_4[25485] = 32'b00000000000000000001101010110100;
assign LUT_4[25486] = 32'b00000000000000000111111001100000;
assign LUT_4[25487] = 32'b00000000000000000001000101011000;
assign LUT_4[25488] = 32'b00000000000000010000000011111001;
assign LUT_4[25489] = 32'b00000000000000001001001111110001;
assign LUT_4[25490] = 32'b00000000000000001111011110011101;
assign LUT_4[25491] = 32'b00000000000000001000101010010101;
assign LUT_4[25492] = 32'b00000000000000001101000100010101;
assign LUT_4[25493] = 32'b00000000000000000110010000001101;
assign LUT_4[25494] = 32'b00000000000000001100011110111001;
assign LUT_4[25495] = 32'b00000000000000000101101010110001;
assign LUT_4[25496] = 32'b00000000000000001001010000001110;
assign LUT_4[25497] = 32'b00000000000000000010011100000110;
assign LUT_4[25498] = 32'b00000000000000001000101010110010;
assign LUT_4[25499] = 32'b00000000000000000001110110101010;
assign LUT_4[25500] = 32'b00000000000000000110010000101010;
assign LUT_4[25501] = 32'b11111111111111111111011100100010;
assign LUT_4[25502] = 32'b00000000000000000101101011001110;
assign LUT_4[25503] = 32'b11111111111111111110110111000110;
assign LUT_4[25504] = 32'b00000000000000010000101101010010;
assign LUT_4[25505] = 32'b00000000000000001001111001001010;
assign LUT_4[25506] = 32'b00000000000000010000000111110110;
assign LUT_4[25507] = 32'b00000000000000001001010011101110;
assign LUT_4[25508] = 32'b00000000000000001101101101101110;
assign LUT_4[25509] = 32'b00000000000000000110111001100110;
assign LUT_4[25510] = 32'b00000000000000001101001000010010;
assign LUT_4[25511] = 32'b00000000000000000110010100001010;
assign LUT_4[25512] = 32'b00000000000000001001111001100111;
assign LUT_4[25513] = 32'b00000000000000000011000101011111;
assign LUT_4[25514] = 32'b00000000000000001001010100001011;
assign LUT_4[25515] = 32'b00000000000000000010100000000011;
assign LUT_4[25516] = 32'b00000000000000000110111010000011;
assign LUT_4[25517] = 32'b00000000000000000000000101111011;
assign LUT_4[25518] = 32'b00000000000000000110010100100111;
assign LUT_4[25519] = 32'b11111111111111111111100000011111;
assign LUT_4[25520] = 32'b00000000000000001110011111000000;
assign LUT_4[25521] = 32'b00000000000000000111101010111000;
assign LUT_4[25522] = 32'b00000000000000001101111001100100;
assign LUT_4[25523] = 32'b00000000000000000111000101011100;
assign LUT_4[25524] = 32'b00000000000000001011011111011100;
assign LUT_4[25525] = 32'b00000000000000000100101011010100;
assign LUT_4[25526] = 32'b00000000000000001010111010000000;
assign LUT_4[25527] = 32'b00000000000000000100000101111000;
assign LUT_4[25528] = 32'b00000000000000000111101011010101;
assign LUT_4[25529] = 32'b00000000000000000000110111001101;
assign LUT_4[25530] = 32'b00000000000000000111000101111001;
assign LUT_4[25531] = 32'b00000000000000000000010001110001;
assign LUT_4[25532] = 32'b00000000000000000100101011110001;
assign LUT_4[25533] = 32'b11111111111111111101110111101001;
assign LUT_4[25534] = 32'b00000000000000000100000110010101;
assign LUT_4[25535] = 32'b11111111111111111101010010001101;
assign LUT_4[25536] = 32'b00000000000000010011101001011111;
assign LUT_4[25537] = 32'b00000000000000001100110101010111;
assign LUT_4[25538] = 32'b00000000000000010011000100000011;
assign LUT_4[25539] = 32'b00000000000000001100001111111011;
assign LUT_4[25540] = 32'b00000000000000010000101001111011;
assign LUT_4[25541] = 32'b00000000000000001001110101110011;
assign LUT_4[25542] = 32'b00000000000000010000000100011111;
assign LUT_4[25543] = 32'b00000000000000001001010000010111;
assign LUT_4[25544] = 32'b00000000000000001100110101110100;
assign LUT_4[25545] = 32'b00000000000000000110000001101100;
assign LUT_4[25546] = 32'b00000000000000001100010000011000;
assign LUT_4[25547] = 32'b00000000000000000101011100010000;
assign LUT_4[25548] = 32'b00000000000000001001110110010000;
assign LUT_4[25549] = 32'b00000000000000000011000010001000;
assign LUT_4[25550] = 32'b00000000000000001001010000110100;
assign LUT_4[25551] = 32'b00000000000000000010011100101100;
assign LUT_4[25552] = 32'b00000000000000010001011011001101;
assign LUT_4[25553] = 32'b00000000000000001010100111000101;
assign LUT_4[25554] = 32'b00000000000000010000110101110001;
assign LUT_4[25555] = 32'b00000000000000001010000001101001;
assign LUT_4[25556] = 32'b00000000000000001110011011101001;
assign LUT_4[25557] = 32'b00000000000000000111100111100001;
assign LUT_4[25558] = 32'b00000000000000001101110110001101;
assign LUT_4[25559] = 32'b00000000000000000111000010000101;
assign LUT_4[25560] = 32'b00000000000000001010100111100010;
assign LUT_4[25561] = 32'b00000000000000000011110011011010;
assign LUT_4[25562] = 32'b00000000000000001010000010000110;
assign LUT_4[25563] = 32'b00000000000000000011001101111110;
assign LUT_4[25564] = 32'b00000000000000000111100111111110;
assign LUT_4[25565] = 32'b00000000000000000000110011110110;
assign LUT_4[25566] = 32'b00000000000000000111000010100010;
assign LUT_4[25567] = 32'b00000000000000000000001110011010;
assign LUT_4[25568] = 32'b00000000000000010010000100100110;
assign LUT_4[25569] = 32'b00000000000000001011010000011110;
assign LUT_4[25570] = 32'b00000000000000010001011111001010;
assign LUT_4[25571] = 32'b00000000000000001010101011000010;
assign LUT_4[25572] = 32'b00000000000000001111000101000010;
assign LUT_4[25573] = 32'b00000000000000001000010000111010;
assign LUT_4[25574] = 32'b00000000000000001110011111100110;
assign LUT_4[25575] = 32'b00000000000000000111101011011110;
assign LUT_4[25576] = 32'b00000000000000001011010000111011;
assign LUT_4[25577] = 32'b00000000000000000100011100110011;
assign LUT_4[25578] = 32'b00000000000000001010101011011111;
assign LUT_4[25579] = 32'b00000000000000000011110111010111;
assign LUT_4[25580] = 32'b00000000000000001000010001010111;
assign LUT_4[25581] = 32'b00000000000000000001011101001111;
assign LUT_4[25582] = 32'b00000000000000000111101011111011;
assign LUT_4[25583] = 32'b00000000000000000000110111110011;
assign LUT_4[25584] = 32'b00000000000000001111110110010100;
assign LUT_4[25585] = 32'b00000000000000001001000010001100;
assign LUT_4[25586] = 32'b00000000000000001111010000111000;
assign LUT_4[25587] = 32'b00000000000000001000011100110000;
assign LUT_4[25588] = 32'b00000000000000001100110110110000;
assign LUT_4[25589] = 32'b00000000000000000110000010101000;
assign LUT_4[25590] = 32'b00000000000000001100010001010100;
assign LUT_4[25591] = 32'b00000000000000000101011101001100;
assign LUT_4[25592] = 32'b00000000000000001001000010101001;
assign LUT_4[25593] = 32'b00000000000000000010001110100001;
assign LUT_4[25594] = 32'b00000000000000001000011101001101;
assign LUT_4[25595] = 32'b00000000000000000001101001000101;
assign LUT_4[25596] = 32'b00000000000000000110000011000101;
assign LUT_4[25597] = 32'b11111111111111111111001110111101;
assign LUT_4[25598] = 32'b00000000000000000101011101101001;
assign LUT_4[25599] = 32'b11111111111111111110101001100001;
assign LUT_4[25600] = 32'b00000000000000001101010110110111;
assign LUT_4[25601] = 32'b00000000000000000110100010101111;
assign LUT_4[25602] = 32'b00000000000000001100110001011011;
assign LUT_4[25603] = 32'b00000000000000000101111101010011;
assign LUT_4[25604] = 32'b00000000000000001010010111010011;
assign LUT_4[25605] = 32'b00000000000000000011100011001011;
assign LUT_4[25606] = 32'b00000000000000001001110001110111;
assign LUT_4[25607] = 32'b00000000000000000010111101101111;
assign LUT_4[25608] = 32'b00000000000000000110100011001100;
assign LUT_4[25609] = 32'b11111111111111111111101111000100;
assign LUT_4[25610] = 32'b00000000000000000101111101110000;
assign LUT_4[25611] = 32'b11111111111111111111001001101000;
assign LUT_4[25612] = 32'b00000000000000000011100011101000;
assign LUT_4[25613] = 32'b11111111111111111100101111100000;
assign LUT_4[25614] = 32'b00000000000000000010111110001100;
assign LUT_4[25615] = 32'b11111111111111111100001010000100;
assign LUT_4[25616] = 32'b00000000000000001011001000100101;
assign LUT_4[25617] = 32'b00000000000000000100010100011101;
assign LUT_4[25618] = 32'b00000000000000001010100011001001;
assign LUT_4[25619] = 32'b00000000000000000011101111000001;
assign LUT_4[25620] = 32'b00000000000000001000001001000001;
assign LUT_4[25621] = 32'b00000000000000000001010100111001;
assign LUT_4[25622] = 32'b00000000000000000111100011100101;
assign LUT_4[25623] = 32'b00000000000000000000101111011101;
assign LUT_4[25624] = 32'b00000000000000000100010100111010;
assign LUT_4[25625] = 32'b11111111111111111101100000110010;
assign LUT_4[25626] = 32'b00000000000000000011101111011110;
assign LUT_4[25627] = 32'b11111111111111111100111011010110;
assign LUT_4[25628] = 32'b00000000000000000001010101010110;
assign LUT_4[25629] = 32'b11111111111111111010100001001110;
assign LUT_4[25630] = 32'b00000000000000000000101111111010;
assign LUT_4[25631] = 32'b11111111111111111001111011110010;
assign LUT_4[25632] = 32'b00000000000000001011110001111110;
assign LUT_4[25633] = 32'b00000000000000000100111101110110;
assign LUT_4[25634] = 32'b00000000000000001011001100100010;
assign LUT_4[25635] = 32'b00000000000000000100011000011010;
assign LUT_4[25636] = 32'b00000000000000001000110010011010;
assign LUT_4[25637] = 32'b00000000000000000001111110010010;
assign LUT_4[25638] = 32'b00000000000000001000001100111110;
assign LUT_4[25639] = 32'b00000000000000000001011000110110;
assign LUT_4[25640] = 32'b00000000000000000100111110010011;
assign LUT_4[25641] = 32'b11111111111111111110001010001011;
assign LUT_4[25642] = 32'b00000000000000000100011000110111;
assign LUT_4[25643] = 32'b11111111111111111101100100101111;
assign LUT_4[25644] = 32'b00000000000000000001111110101111;
assign LUT_4[25645] = 32'b11111111111111111011001010100111;
assign LUT_4[25646] = 32'b00000000000000000001011001010011;
assign LUT_4[25647] = 32'b11111111111111111010100101001011;
assign LUT_4[25648] = 32'b00000000000000001001100011101100;
assign LUT_4[25649] = 32'b00000000000000000010101111100100;
assign LUT_4[25650] = 32'b00000000000000001000111110010000;
assign LUT_4[25651] = 32'b00000000000000000010001010001000;
assign LUT_4[25652] = 32'b00000000000000000110100100001000;
assign LUT_4[25653] = 32'b11111111111111111111110000000000;
assign LUT_4[25654] = 32'b00000000000000000101111110101100;
assign LUT_4[25655] = 32'b11111111111111111111001010100100;
assign LUT_4[25656] = 32'b00000000000000000010110000000001;
assign LUT_4[25657] = 32'b11111111111111111011111011111001;
assign LUT_4[25658] = 32'b00000000000000000010001010100101;
assign LUT_4[25659] = 32'b11111111111111111011010110011101;
assign LUT_4[25660] = 32'b11111111111111111111110000011101;
assign LUT_4[25661] = 32'b11111111111111111000111100010101;
assign LUT_4[25662] = 32'b11111111111111111111001011000001;
assign LUT_4[25663] = 32'b11111111111111111000010110111001;
assign LUT_4[25664] = 32'b00000000000000001110101110001011;
assign LUT_4[25665] = 32'b00000000000000000111111010000011;
assign LUT_4[25666] = 32'b00000000000000001110001000101111;
assign LUT_4[25667] = 32'b00000000000000000111010100100111;
assign LUT_4[25668] = 32'b00000000000000001011101110100111;
assign LUT_4[25669] = 32'b00000000000000000100111010011111;
assign LUT_4[25670] = 32'b00000000000000001011001001001011;
assign LUT_4[25671] = 32'b00000000000000000100010101000011;
assign LUT_4[25672] = 32'b00000000000000000111111010100000;
assign LUT_4[25673] = 32'b00000000000000000001000110011000;
assign LUT_4[25674] = 32'b00000000000000000111010101000100;
assign LUT_4[25675] = 32'b00000000000000000000100000111100;
assign LUT_4[25676] = 32'b00000000000000000100111010111100;
assign LUT_4[25677] = 32'b11111111111111111110000110110100;
assign LUT_4[25678] = 32'b00000000000000000100010101100000;
assign LUT_4[25679] = 32'b11111111111111111101100001011000;
assign LUT_4[25680] = 32'b00000000000000001100011111111001;
assign LUT_4[25681] = 32'b00000000000000000101101011110001;
assign LUT_4[25682] = 32'b00000000000000001011111010011101;
assign LUT_4[25683] = 32'b00000000000000000101000110010101;
assign LUT_4[25684] = 32'b00000000000000001001100000010101;
assign LUT_4[25685] = 32'b00000000000000000010101100001101;
assign LUT_4[25686] = 32'b00000000000000001000111010111001;
assign LUT_4[25687] = 32'b00000000000000000010000110110001;
assign LUT_4[25688] = 32'b00000000000000000101101100001110;
assign LUT_4[25689] = 32'b11111111111111111110111000000110;
assign LUT_4[25690] = 32'b00000000000000000101000110110010;
assign LUT_4[25691] = 32'b11111111111111111110010010101010;
assign LUT_4[25692] = 32'b00000000000000000010101100101010;
assign LUT_4[25693] = 32'b11111111111111111011111000100010;
assign LUT_4[25694] = 32'b00000000000000000010000111001110;
assign LUT_4[25695] = 32'b11111111111111111011010011000110;
assign LUT_4[25696] = 32'b00000000000000001101001001010010;
assign LUT_4[25697] = 32'b00000000000000000110010101001010;
assign LUT_4[25698] = 32'b00000000000000001100100011110110;
assign LUT_4[25699] = 32'b00000000000000000101101111101110;
assign LUT_4[25700] = 32'b00000000000000001010001001101110;
assign LUT_4[25701] = 32'b00000000000000000011010101100110;
assign LUT_4[25702] = 32'b00000000000000001001100100010010;
assign LUT_4[25703] = 32'b00000000000000000010110000001010;
assign LUT_4[25704] = 32'b00000000000000000110010101100111;
assign LUT_4[25705] = 32'b11111111111111111111100001011111;
assign LUT_4[25706] = 32'b00000000000000000101110000001011;
assign LUT_4[25707] = 32'b11111111111111111110111100000011;
assign LUT_4[25708] = 32'b00000000000000000011010110000011;
assign LUT_4[25709] = 32'b11111111111111111100100001111011;
assign LUT_4[25710] = 32'b00000000000000000010110000100111;
assign LUT_4[25711] = 32'b11111111111111111011111100011111;
assign LUT_4[25712] = 32'b00000000000000001010111011000000;
assign LUT_4[25713] = 32'b00000000000000000100000110111000;
assign LUT_4[25714] = 32'b00000000000000001010010101100100;
assign LUT_4[25715] = 32'b00000000000000000011100001011100;
assign LUT_4[25716] = 32'b00000000000000000111111011011100;
assign LUT_4[25717] = 32'b00000000000000000001000111010100;
assign LUT_4[25718] = 32'b00000000000000000111010110000000;
assign LUT_4[25719] = 32'b00000000000000000000100001111000;
assign LUT_4[25720] = 32'b00000000000000000100000111010101;
assign LUT_4[25721] = 32'b11111111111111111101010011001101;
assign LUT_4[25722] = 32'b00000000000000000011100001111001;
assign LUT_4[25723] = 32'b11111111111111111100101101110001;
assign LUT_4[25724] = 32'b00000000000000000001000111110001;
assign LUT_4[25725] = 32'b11111111111111111010010011101001;
assign LUT_4[25726] = 32'b00000000000000000000100010010101;
assign LUT_4[25727] = 32'b11111111111111111001101110001101;
assign LUT_4[25728] = 32'b00000000000000001111111100111111;
assign LUT_4[25729] = 32'b00000000000000001001001000110111;
assign LUT_4[25730] = 32'b00000000000000001111010111100011;
assign LUT_4[25731] = 32'b00000000000000001000100011011011;
assign LUT_4[25732] = 32'b00000000000000001100111101011011;
assign LUT_4[25733] = 32'b00000000000000000110001001010011;
assign LUT_4[25734] = 32'b00000000000000001100010111111111;
assign LUT_4[25735] = 32'b00000000000000000101100011110111;
assign LUT_4[25736] = 32'b00000000000000001001001001010100;
assign LUT_4[25737] = 32'b00000000000000000010010101001100;
assign LUT_4[25738] = 32'b00000000000000001000100011111000;
assign LUT_4[25739] = 32'b00000000000000000001101111110000;
assign LUT_4[25740] = 32'b00000000000000000110001001110000;
assign LUT_4[25741] = 32'b11111111111111111111010101101000;
assign LUT_4[25742] = 32'b00000000000000000101100100010100;
assign LUT_4[25743] = 32'b11111111111111111110110000001100;
assign LUT_4[25744] = 32'b00000000000000001101101110101101;
assign LUT_4[25745] = 32'b00000000000000000110111010100101;
assign LUT_4[25746] = 32'b00000000000000001101001001010001;
assign LUT_4[25747] = 32'b00000000000000000110010101001001;
assign LUT_4[25748] = 32'b00000000000000001010101111001001;
assign LUT_4[25749] = 32'b00000000000000000011111011000001;
assign LUT_4[25750] = 32'b00000000000000001010001001101101;
assign LUT_4[25751] = 32'b00000000000000000011010101100101;
assign LUT_4[25752] = 32'b00000000000000000110111011000010;
assign LUT_4[25753] = 32'b00000000000000000000000110111010;
assign LUT_4[25754] = 32'b00000000000000000110010101100110;
assign LUT_4[25755] = 32'b11111111111111111111100001011110;
assign LUT_4[25756] = 32'b00000000000000000011111011011110;
assign LUT_4[25757] = 32'b11111111111111111101000111010110;
assign LUT_4[25758] = 32'b00000000000000000011010110000010;
assign LUT_4[25759] = 32'b11111111111111111100100001111010;
assign LUT_4[25760] = 32'b00000000000000001110011000000110;
assign LUT_4[25761] = 32'b00000000000000000111100011111110;
assign LUT_4[25762] = 32'b00000000000000001101110010101010;
assign LUT_4[25763] = 32'b00000000000000000110111110100010;
assign LUT_4[25764] = 32'b00000000000000001011011000100010;
assign LUT_4[25765] = 32'b00000000000000000100100100011010;
assign LUT_4[25766] = 32'b00000000000000001010110011000110;
assign LUT_4[25767] = 32'b00000000000000000011111110111110;
assign LUT_4[25768] = 32'b00000000000000000111100100011011;
assign LUT_4[25769] = 32'b00000000000000000000110000010011;
assign LUT_4[25770] = 32'b00000000000000000110111110111111;
assign LUT_4[25771] = 32'b00000000000000000000001010110111;
assign LUT_4[25772] = 32'b00000000000000000100100100110111;
assign LUT_4[25773] = 32'b11111111111111111101110000101111;
assign LUT_4[25774] = 32'b00000000000000000011111111011011;
assign LUT_4[25775] = 32'b11111111111111111101001011010011;
assign LUT_4[25776] = 32'b00000000000000001100001001110100;
assign LUT_4[25777] = 32'b00000000000000000101010101101100;
assign LUT_4[25778] = 32'b00000000000000001011100100011000;
assign LUT_4[25779] = 32'b00000000000000000100110000010000;
assign LUT_4[25780] = 32'b00000000000000001001001010010000;
assign LUT_4[25781] = 32'b00000000000000000010010110001000;
assign LUT_4[25782] = 32'b00000000000000001000100100110100;
assign LUT_4[25783] = 32'b00000000000000000001110000101100;
assign LUT_4[25784] = 32'b00000000000000000101010110001001;
assign LUT_4[25785] = 32'b11111111111111111110100010000001;
assign LUT_4[25786] = 32'b00000000000000000100110000101101;
assign LUT_4[25787] = 32'b11111111111111111101111100100101;
assign LUT_4[25788] = 32'b00000000000000000010010110100101;
assign LUT_4[25789] = 32'b11111111111111111011100010011101;
assign LUT_4[25790] = 32'b00000000000000000001110001001001;
assign LUT_4[25791] = 32'b11111111111111111010111101000001;
assign LUT_4[25792] = 32'b00000000000000010001010100010011;
assign LUT_4[25793] = 32'b00000000000000001010100000001011;
assign LUT_4[25794] = 32'b00000000000000010000101110110111;
assign LUT_4[25795] = 32'b00000000000000001001111010101111;
assign LUT_4[25796] = 32'b00000000000000001110010100101111;
assign LUT_4[25797] = 32'b00000000000000000111100000100111;
assign LUT_4[25798] = 32'b00000000000000001101101111010011;
assign LUT_4[25799] = 32'b00000000000000000110111011001011;
assign LUT_4[25800] = 32'b00000000000000001010100000101000;
assign LUT_4[25801] = 32'b00000000000000000011101100100000;
assign LUT_4[25802] = 32'b00000000000000001001111011001100;
assign LUT_4[25803] = 32'b00000000000000000011000111000100;
assign LUT_4[25804] = 32'b00000000000000000111100001000100;
assign LUT_4[25805] = 32'b00000000000000000000101100111100;
assign LUT_4[25806] = 32'b00000000000000000110111011101000;
assign LUT_4[25807] = 32'b00000000000000000000000111100000;
assign LUT_4[25808] = 32'b00000000000000001111000110000001;
assign LUT_4[25809] = 32'b00000000000000001000010001111001;
assign LUT_4[25810] = 32'b00000000000000001110100000100101;
assign LUT_4[25811] = 32'b00000000000000000111101100011101;
assign LUT_4[25812] = 32'b00000000000000001100000110011101;
assign LUT_4[25813] = 32'b00000000000000000101010010010101;
assign LUT_4[25814] = 32'b00000000000000001011100001000001;
assign LUT_4[25815] = 32'b00000000000000000100101100111001;
assign LUT_4[25816] = 32'b00000000000000001000010010010110;
assign LUT_4[25817] = 32'b00000000000000000001011110001110;
assign LUT_4[25818] = 32'b00000000000000000111101100111010;
assign LUT_4[25819] = 32'b00000000000000000000111000110010;
assign LUT_4[25820] = 32'b00000000000000000101010010110010;
assign LUT_4[25821] = 32'b11111111111111111110011110101010;
assign LUT_4[25822] = 32'b00000000000000000100101101010110;
assign LUT_4[25823] = 32'b11111111111111111101111001001110;
assign LUT_4[25824] = 32'b00000000000000001111101111011010;
assign LUT_4[25825] = 32'b00000000000000001000111011010010;
assign LUT_4[25826] = 32'b00000000000000001111001001111110;
assign LUT_4[25827] = 32'b00000000000000001000010101110110;
assign LUT_4[25828] = 32'b00000000000000001100101111110110;
assign LUT_4[25829] = 32'b00000000000000000101111011101110;
assign LUT_4[25830] = 32'b00000000000000001100001010011010;
assign LUT_4[25831] = 32'b00000000000000000101010110010010;
assign LUT_4[25832] = 32'b00000000000000001000111011101111;
assign LUT_4[25833] = 32'b00000000000000000010000111100111;
assign LUT_4[25834] = 32'b00000000000000001000010110010011;
assign LUT_4[25835] = 32'b00000000000000000001100010001011;
assign LUT_4[25836] = 32'b00000000000000000101111100001011;
assign LUT_4[25837] = 32'b11111111111111111111001000000011;
assign LUT_4[25838] = 32'b00000000000000000101010110101111;
assign LUT_4[25839] = 32'b11111111111111111110100010100111;
assign LUT_4[25840] = 32'b00000000000000001101100001001000;
assign LUT_4[25841] = 32'b00000000000000000110101101000000;
assign LUT_4[25842] = 32'b00000000000000001100111011101100;
assign LUT_4[25843] = 32'b00000000000000000110000111100100;
assign LUT_4[25844] = 32'b00000000000000001010100001100100;
assign LUT_4[25845] = 32'b00000000000000000011101101011100;
assign LUT_4[25846] = 32'b00000000000000001001111100001000;
assign LUT_4[25847] = 32'b00000000000000000011001000000000;
assign LUT_4[25848] = 32'b00000000000000000110101101011101;
assign LUT_4[25849] = 32'b11111111111111111111111001010101;
assign LUT_4[25850] = 32'b00000000000000000110001000000001;
assign LUT_4[25851] = 32'b11111111111111111111010011111001;
assign LUT_4[25852] = 32'b00000000000000000011101101111001;
assign LUT_4[25853] = 32'b11111111111111111100111001110001;
assign LUT_4[25854] = 32'b00000000000000000011001000011101;
assign LUT_4[25855] = 32'b11111111111111111100010100010101;
assign LUT_4[25856] = 32'b00000000000000010010010010011010;
assign LUT_4[25857] = 32'b00000000000000001011011110010010;
assign LUT_4[25858] = 32'b00000000000000010001101100111110;
assign LUT_4[25859] = 32'b00000000000000001010111000110110;
assign LUT_4[25860] = 32'b00000000000000001111010010110110;
assign LUT_4[25861] = 32'b00000000000000001000011110101110;
assign LUT_4[25862] = 32'b00000000000000001110101101011010;
assign LUT_4[25863] = 32'b00000000000000000111111001010010;
assign LUT_4[25864] = 32'b00000000000000001011011110101111;
assign LUT_4[25865] = 32'b00000000000000000100101010100111;
assign LUT_4[25866] = 32'b00000000000000001010111001010011;
assign LUT_4[25867] = 32'b00000000000000000100000101001011;
assign LUT_4[25868] = 32'b00000000000000001000011111001011;
assign LUT_4[25869] = 32'b00000000000000000001101011000011;
assign LUT_4[25870] = 32'b00000000000000000111111001101111;
assign LUT_4[25871] = 32'b00000000000000000001000101100111;
assign LUT_4[25872] = 32'b00000000000000010000000100001000;
assign LUT_4[25873] = 32'b00000000000000001001010000000000;
assign LUT_4[25874] = 32'b00000000000000001111011110101100;
assign LUT_4[25875] = 32'b00000000000000001000101010100100;
assign LUT_4[25876] = 32'b00000000000000001101000100100100;
assign LUT_4[25877] = 32'b00000000000000000110010000011100;
assign LUT_4[25878] = 32'b00000000000000001100011111001000;
assign LUT_4[25879] = 32'b00000000000000000101101011000000;
assign LUT_4[25880] = 32'b00000000000000001001010000011101;
assign LUT_4[25881] = 32'b00000000000000000010011100010101;
assign LUT_4[25882] = 32'b00000000000000001000101011000001;
assign LUT_4[25883] = 32'b00000000000000000001110110111001;
assign LUT_4[25884] = 32'b00000000000000000110010000111001;
assign LUT_4[25885] = 32'b11111111111111111111011100110001;
assign LUT_4[25886] = 32'b00000000000000000101101011011101;
assign LUT_4[25887] = 32'b11111111111111111110110111010101;
assign LUT_4[25888] = 32'b00000000000000010000101101100001;
assign LUT_4[25889] = 32'b00000000000000001001111001011001;
assign LUT_4[25890] = 32'b00000000000000010000001000000101;
assign LUT_4[25891] = 32'b00000000000000001001010011111101;
assign LUT_4[25892] = 32'b00000000000000001101101101111101;
assign LUT_4[25893] = 32'b00000000000000000110111001110101;
assign LUT_4[25894] = 32'b00000000000000001101001000100001;
assign LUT_4[25895] = 32'b00000000000000000110010100011001;
assign LUT_4[25896] = 32'b00000000000000001001111001110110;
assign LUT_4[25897] = 32'b00000000000000000011000101101110;
assign LUT_4[25898] = 32'b00000000000000001001010100011010;
assign LUT_4[25899] = 32'b00000000000000000010100000010010;
assign LUT_4[25900] = 32'b00000000000000000110111010010010;
assign LUT_4[25901] = 32'b00000000000000000000000110001010;
assign LUT_4[25902] = 32'b00000000000000000110010100110110;
assign LUT_4[25903] = 32'b11111111111111111111100000101110;
assign LUT_4[25904] = 32'b00000000000000001110011111001111;
assign LUT_4[25905] = 32'b00000000000000000111101011000111;
assign LUT_4[25906] = 32'b00000000000000001101111001110011;
assign LUT_4[25907] = 32'b00000000000000000111000101101011;
assign LUT_4[25908] = 32'b00000000000000001011011111101011;
assign LUT_4[25909] = 32'b00000000000000000100101011100011;
assign LUT_4[25910] = 32'b00000000000000001010111010001111;
assign LUT_4[25911] = 32'b00000000000000000100000110000111;
assign LUT_4[25912] = 32'b00000000000000000111101011100100;
assign LUT_4[25913] = 32'b00000000000000000000110111011100;
assign LUT_4[25914] = 32'b00000000000000000111000110001000;
assign LUT_4[25915] = 32'b00000000000000000000010010000000;
assign LUT_4[25916] = 32'b00000000000000000100101100000000;
assign LUT_4[25917] = 32'b11111111111111111101110111111000;
assign LUT_4[25918] = 32'b00000000000000000100000110100100;
assign LUT_4[25919] = 32'b11111111111111111101010010011100;
assign LUT_4[25920] = 32'b00000000000000010011101001101110;
assign LUT_4[25921] = 32'b00000000000000001100110101100110;
assign LUT_4[25922] = 32'b00000000000000010011000100010010;
assign LUT_4[25923] = 32'b00000000000000001100010000001010;
assign LUT_4[25924] = 32'b00000000000000010000101010001010;
assign LUT_4[25925] = 32'b00000000000000001001110110000010;
assign LUT_4[25926] = 32'b00000000000000010000000100101110;
assign LUT_4[25927] = 32'b00000000000000001001010000100110;
assign LUT_4[25928] = 32'b00000000000000001100110110000011;
assign LUT_4[25929] = 32'b00000000000000000110000001111011;
assign LUT_4[25930] = 32'b00000000000000001100010000100111;
assign LUT_4[25931] = 32'b00000000000000000101011100011111;
assign LUT_4[25932] = 32'b00000000000000001001110110011111;
assign LUT_4[25933] = 32'b00000000000000000011000010010111;
assign LUT_4[25934] = 32'b00000000000000001001010001000011;
assign LUT_4[25935] = 32'b00000000000000000010011100111011;
assign LUT_4[25936] = 32'b00000000000000010001011011011100;
assign LUT_4[25937] = 32'b00000000000000001010100111010100;
assign LUT_4[25938] = 32'b00000000000000010000110110000000;
assign LUT_4[25939] = 32'b00000000000000001010000001111000;
assign LUT_4[25940] = 32'b00000000000000001110011011111000;
assign LUT_4[25941] = 32'b00000000000000000111100111110000;
assign LUT_4[25942] = 32'b00000000000000001101110110011100;
assign LUT_4[25943] = 32'b00000000000000000111000010010100;
assign LUT_4[25944] = 32'b00000000000000001010100111110001;
assign LUT_4[25945] = 32'b00000000000000000011110011101001;
assign LUT_4[25946] = 32'b00000000000000001010000010010101;
assign LUT_4[25947] = 32'b00000000000000000011001110001101;
assign LUT_4[25948] = 32'b00000000000000000111101000001101;
assign LUT_4[25949] = 32'b00000000000000000000110100000101;
assign LUT_4[25950] = 32'b00000000000000000111000010110001;
assign LUT_4[25951] = 32'b00000000000000000000001110101001;
assign LUT_4[25952] = 32'b00000000000000010010000100110101;
assign LUT_4[25953] = 32'b00000000000000001011010000101101;
assign LUT_4[25954] = 32'b00000000000000010001011111011001;
assign LUT_4[25955] = 32'b00000000000000001010101011010001;
assign LUT_4[25956] = 32'b00000000000000001111000101010001;
assign LUT_4[25957] = 32'b00000000000000001000010001001001;
assign LUT_4[25958] = 32'b00000000000000001110011111110101;
assign LUT_4[25959] = 32'b00000000000000000111101011101101;
assign LUT_4[25960] = 32'b00000000000000001011010001001010;
assign LUT_4[25961] = 32'b00000000000000000100011101000010;
assign LUT_4[25962] = 32'b00000000000000001010101011101110;
assign LUT_4[25963] = 32'b00000000000000000011110111100110;
assign LUT_4[25964] = 32'b00000000000000001000010001100110;
assign LUT_4[25965] = 32'b00000000000000000001011101011110;
assign LUT_4[25966] = 32'b00000000000000000111101100001010;
assign LUT_4[25967] = 32'b00000000000000000000111000000010;
assign LUT_4[25968] = 32'b00000000000000001111110110100011;
assign LUT_4[25969] = 32'b00000000000000001001000010011011;
assign LUT_4[25970] = 32'b00000000000000001111010001000111;
assign LUT_4[25971] = 32'b00000000000000001000011100111111;
assign LUT_4[25972] = 32'b00000000000000001100110110111111;
assign LUT_4[25973] = 32'b00000000000000000110000010110111;
assign LUT_4[25974] = 32'b00000000000000001100010001100011;
assign LUT_4[25975] = 32'b00000000000000000101011101011011;
assign LUT_4[25976] = 32'b00000000000000001001000010111000;
assign LUT_4[25977] = 32'b00000000000000000010001110110000;
assign LUT_4[25978] = 32'b00000000000000001000011101011100;
assign LUT_4[25979] = 32'b00000000000000000001101001010100;
assign LUT_4[25980] = 32'b00000000000000000110000011010100;
assign LUT_4[25981] = 32'b11111111111111111111001111001100;
assign LUT_4[25982] = 32'b00000000000000000101011101111000;
assign LUT_4[25983] = 32'b11111111111111111110101001110000;
assign LUT_4[25984] = 32'b00000000000000010100111000100010;
assign LUT_4[25985] = 32'b00000000000000001110000100011010;
assign LUT_4[25986] = 32'b00000000000000010100010011000110;
assign LUT_4[25987] = 32'b00000000000000001101011110111110;
assign LUT_4[25988] = 32'b00000000000000010001111000111110;
assign LUT_4[25989] = 32'b00000000000000001011000100110110;
assign LUT_4[25990] = 32'b00000000000000010001010011100010;
assign LUT_4[25991] = 32'b00000000000000001010011111011010;
assign LUT_4[25992] = 32'b00000000000000001110000100110111;
assign LUT_4[25993] = 32'b00000000000000000111010000101111;
assign LUT_4[25994] = 32'b00000000000000001101011111011011;
assign LUT_4[25995] = 32'b00000000000000000110101011010011;
assign LUT_4[25996] = 32'b00000000000000001011000101010011;
assign LUT_4[25997] = 32'b00000000000000000100010001001011;
assign LUT_4[25998] = 32'b00000000000000001010011111110111;
assign LUT_4[25999] = 32'b00000000000000000011101011101111;
assign LUT_4[26000] = 32'b00000000000000010010101010010000;
assign LUT_4[26001] = 32'b00000000000000001011110110001000;
assign LUT_4[26002] = 32'b00000000000000010010000100110100;
assign LUT_4[26003] = 32'b00000000000000001011010000101100;
assign LUT_4[26004] = 32'b00000000000000001111101010101100;
assign LUT_4[26005] = 32'b00000000000000001000110110100100;
assign LUT_4[26006] = 32'b00000000000000001111000101010000;
assign LUT_4[26007] = 32'b00000000000000001000010001001000;
assign LUT_4[26008] = 32'b00000000000000001011110110100101;
assign LUT_4[26009] = 32'b00000000000000000101000010011101;
assign LUT_4[26010] = 32'b00000000000000001011010001001001;
assign LUT_4[26011] = 32'b00000000000000000100011101000001;
assign LUT_4[26012] = 32'b00000000000000001000110111000001;
assign LUT_4[26013] = 32'b00000000000000000010000010111001;
assign LUT_4[26014] = 32'b00000000000000001000010001100101;
assign LUT_4[26015] = 32'b00000000000000000001011101011101;
assign LUT_4[26016] = 32'b00000000000000010011010011101001;
assign LUT_4[26017] = 32'b00000000000000001100011111100001;
assign LUT_4[26018] = 32'b00000000000000010010101110001101;
assign LUT_4[26019] = 32'b00000000000000001011111010000101;
assign LUT_4[26020] = 32'b00000000000000010000010100000101;
assign LUT_4[26021] = 32'b00000000000000001001011111111101;
assign LUT_4[26022] = 32'b00000000000000001111101110101001;
assign LUT_4[26023] = 32'b00000000000000001000111010100001;
assign LUT_4[26024] = 32'b00000000000000001100011111111110;
assign LUT_4[26025] = 32'b00000000000000000101101011110110;
assign LUT_4[26026] = 32'b00000000000000001011111010100010;
assign LUT_4[26027] = 32'b00000000000000000101000110011010;
assign LUT_4[26028] = 32'b00000000000000001001100000011010;
assign LUT_4[26029] = 32'b00000000000000000010101100010010;
assign LUT_4[26030] = 32'b00000000000000001000111010111110;
assign LUT_4[26031] = 32'b00000000000000000010000110110110;
assign LUT_4[26032] = 32'b00000000000000010001000101010111;
assign LUT_4[26033] = 32'b00000000000000001010010001001111;
assign LUT_4[26034] = 32'b00000000000000010000011111111011;
assign LUT_4[26035] = 32'b00000000000000001001101011110011;
assign LUT_4[26036] = 32'b00000000000000001110000101110011;
assign LUT_4[26037] = 32'b00000000000000000111010001101011;
assign LUT_4[26038] = 32'b00000000000000001101100000010111;
assign LUT_4[26039] = 32'b00000000000000000110101100001111;
assign LUT_4[26040] = 32'b00000000000000001010010001101100;
assign LUT_4[26041] = 32'b00000000000000000011011101100100;
assign LUT_4[26042] = 32'b00000000000000001001101100010000;
assign LUT_4[26043] = 32'b00000000000000000010111000001000;
assign LUT_4[26044] = 32'b00000000000000000111010010001000;
assign LUT_4[26045] = 32'b00000000000000000000011110000000;
assign LUT_4[26046] = 32'b00000000000000000110101100101100;
assign LUT_4[26047] = 32'b11111111111111111111111000100100;
assign LUT_4[26048] = 32'b00000000000000010110001111110110;
assign LUT_4[26049] = 32'b00000000000000001111011011101110;
assign LUT_4[26050] = 32'b00000000000000010101101010011010;
assign LUT_4[26051] = 32'b00000000000000001110110110010010;
assign LUT_4[26052] = 32'b00000000000000010011010000010010;
assign LUT_4[26053] = 32'b00000000000000001100011100001010;
assign LUT_4[26054] = 32'b00000000000000010010101010110110;
assign LUT_4[26055] = 32'b00000000000000001011110110101110;
assign LUT_4[26056] = 32'b00000000000000001111011100001011;
assign LUT_4[26057] = 32'b00000000000000001000101000000011;
assign LUT_4[26058] = 32'b00000000000000001110110110101111;
assign LUT_4[26059] = 32'b00000000000000001000000010100111;
assign LUT_4[26060] = 32'b00000000000000001100011100100111;
assign LUT_4[26061] = 32'b00000000000000000101101000011111;
assign LUT_4[26062] = 32'b00000000000000001011110111001011;
assign LUT_4[26063] = 32'b00000000000000000101000011000011;
assign LUT_4[26064] = 32'b00000000000000010100000001100100;
assign LUT_4[26065] = 32'b00000000000000001101001101011100;
assign LUT_4[26066] = 32'b00000000000000010011011100001000;
assign LUT_4[26067] = 32'b00000000000000001100101000000000;
assign LUT_4[26068] = 32'b00000000000000010001000010000000;
assign LUT_4[26069] = 32'b00000000000000001010001101111000;
assign LUT_4[26070] = 32'b00000000000000010000011100100100;
assign LUT_4[26071] = 32'b00000000000000001001101000011100;
assign LUT_4[26072] = 32'b00000000000000001101001101111001;
assign LUT_4[26073] = 32'b00000000000000000110011001110001;
assign LUT_4[26074] = 32'b00000000000000001100101000011101;
assign LUT_4[26075] = 32'b00000000000000000101110100010101;
assign LUT_4[26076] = 32'b00000000000000001010001110010101;
assign LUT_4[26077] = 32'b00000000000000000011011010001101;
assign LUT_4[26078] = 32'b00000000000000001001101000111001;
assign LUT_4[26079] = 32'b00000000000000000010110100110001;
assign LUT_4[26080] = 32'b00000000000000010100101010111101;
assign LUT_4[26081] = 32'b00000000000000001101110110110101;
assign LUT_4[26082] = 32'b00000000000000010100000101100001;
assign LUT_4[26083] = 32'b00000000000000001101010001011001;
assign LUT_4[26084] = 32'b00000000000000010001101011011001;
assign LUT_4[26085] = 32'b00000000000000001010110111010001;
assign LUT_4[26086] = 32'b00000000000000010001000101111101;
assign LUT_4[26087] = 32'b00000000000000001010010001110101;
assign LUT_4[26088] = 32'b00000000000000001101110111010010;
assign LUT_4[26089] = 32'b00000000000000000111000011001010;
assign LUT_4[26090] = 32'b00000000000000001101010001110110;
assign LUT_4[26091] = 32'b00000000000000000110011101101110;
assign LUT_4[26092] = 32'b00000000000000001010110111101110;
assign LUT_4[26093] = 32'b00000000000000000100000011100110;
assign LUT_4[26094] = 32'b00000000000000001010010010010010;
assign LUT_4[26095] = 32'b00000000000000000011011110001010;
assign LUT_4[26096] = 32'b00000000000000010010011100101011;
assign LUT_4[26097] = 32'b00000000000000001011101000100011;
assign LUT_4[26098] = 32'b00000000000000010001110111001111;
assign LUT_4[26099] = 32'b00000000000000001011000011000111;
assign LUT_4[26100] = 32'b00000000000000001111011101000111;
assign LUT_4[26101] = 32'b00000000000000001000101000111111;
assign LUT_4[26102] = 32'b00000000000000001110110111101011;
assign LUT_4[26103] = 32'b00000000000000001000000011100011;
assign LUT_4[26104] = 32'b00000000000000001011101001000000;
assign LUT_4[26105] = 32'b00000000000000000100110100111000;
assign LUT_4[26106] = 32'b00000000000000001011000011100100;
assign LUT_4[26107] = 32'b00000000000000000100001111011100;
assign LUT_4[26108] = 32'b00000000000000001000101001011100;
assign LUT_4[26109] = 32'b00000000000000000001110101010100;
assign LUT_4[26110] = 32'b00000000000000001000000100000000;
assign LUT_4[26111] = 32'b00000000000000000001001111111000;
assign LUT_4[26112] = 32'b00000000000000001100011010111111;
assign LUT_4[26113] = 32'b00000000000000000101100110110111;
assign LUT_4[26114] = 32'b00000000000000001011110101100011;
assign LUT_4[26115] = 32'b00000000000000000101000001011011;
assign LUT_4[26116] = 32'b00000000000000001001011011011011;
assign LUT_4[26117] = 32'b00000000000000000010100111010011;
assign LUT_4[26118] = 32'b00000000000000001000110101111111;
assign LUT_4[26119] = 32'b00000000000000000010000001110111;
assign LUT_4[26120] = 32'b00000000000000000101100111010100;
assign LUT_4[26121] = 32'b11111111111111111110110011001100;
assign LUT_4[26122] = 32'b00000000000000000101000001111000;
assign LUT_4[26123] = 32'b11111111111111111110001101110000;
assign LUT_4[26124] = 32'b00000000000000000010100111110000;
assign LUT_4[26125] = 32'b11111111111111111011110011101000;
assign LUT_4[26126] = 32'b00000000000000000010000010010100;
assign LUT_4[26127] = 32'b11111111111111111011001110001100;
assign LUT_4[26128] = 32'b00000000000000001010001100101101;
assign LUT_4[26129] = 32'b00000000000000000011011000100101;
assign LUT_4[26130] = 32'b00000000000000001001100111010001;
assign LUT_4[26131] = 32'b00000000000000000010110011001001;
assign LUT_4[26132] = 32'b00000000000000000111001101001001;
assign LUT_4[26133] = 32'b00000000000000000000011001000001;
assign LUT_4[26134] = 32'b00000000000000000110100111101101;
assign LUT_4[26135] = 32'b11111111111111111111110011100101;
assign LUT_4[26136] = 32'b00000000000000000011011001000010;
assign LUT_4[26137] = 32'b11111111111111111100100100111010;
assign LUT_4[26138] = 32'b00000000000000000010110011100110;
assign LUT_4[26139] = 32'b11111111111111111011111111011110;
assign LUT_4[26140] = 32'b00000000000000000000011001011110;
assign LUT_4[26141] = 32'b11111111111111111001100101010110;
assign LUT_4[26142] = 32'b11111111111111111111110100000010;
assign LUT_4[26143] = 32'b11111111111111111000111111111010;
assign LUT_4[26144] = 32'b00000000000000001010110110000110;
assign LUT_4[26145] = 32'b00000000000000000100000001111110;
assign LUT_4[26146] = 32'b00000000000000001010010000101010;
assign LUT_4[26147] = 32'b00000000000000000011011100100010;
assign LUT_4[26148] = 32'b00000000000000000111110110100010;
assign LUT_4[26149] = 32'b00000000000000000001000010011010;
assign LUT_4[26150] = 32'b00000000000000000111010001000110;
assign LUT_4[26151] = 32'b00000000000000000000011100111110;
assign LUT_4[26152] = 32'b00000000000000000100000010011011;
assign LUT_4[26153] = 32'b11111111111111111101001110010011;
assign LUT_4[26154] = 32'b00000000000000000011011100111111;
assign LUT_4[26155] = 32'b11111111111111111100101000110111;
assign LUT_4[26156] = 32'b00000000000000000001000010110111;
assign LUT_4[26157] = 32'b11111111111111111010001110101111;
assign LUT_4[26158] = 32'b00000000000000000000011101011011;
assign LUT_4[26159] = 32'b11111111111111111001101001010011;
assign LUT_4[26160] = 32'b00000000000000001000100111110100;
assign LUT_4[26161] = 32'b00000000000000000001110011101100;
assign LUT_4[26162] = 32'b00000000000000001000000010011000;
assign LUT_4[26163] = 32'b00000000000000000001001110010000;
assign LUT_4[26164] = 32'b00000000000000000101101000010000;
assign LUT_4[26165] = 32'b11111111111111111110110100001000;
assign LUT_4[26166] = 32'b00000000000000000101000010110100;
assign LUT_4[26167] = 32'b11111111111111111110001110101100;
assign LUT_4[26168] = 32'b00000000000000000001110100001001;
assign LUT_4[26169] = 32'b11111111111111111011000000000001;
assign LUT_4[26170] = 32'b00000000000000000001001110101101;
assign LUT_4[26171] = 32'b11111111111111111010011010100101;
assign LUT_4[26172] = 32'b11111111111111111110110100100101;
assign LUT_4[26173] = 32'b11111111111111111000000000011101;
assign LUT_4[26174] = 32'b11111111111111111110001111001001;
assign LUT_4[26175] = 32'b11111111111111110111011011000001;
assign LUT_4[26176] = 32'b00000000000000001101110010010011;
assign LUT_4[26177] = 32'b00000000000000000110111110001011;
assign LUT_4[26178] = 32'b00000000000000001101001100110111;
assign LUT_4[26179] = 32'b00000000000000000110011000101111;
assign LUT_4[26180] = 32'b00000000000000001010110010101111;
assign LUT_4[26181] = 32'b00000000000000000011111110100111;
assign LUT_4[26182] = 32'b00000000000000001010001101010011;
assign LUT_4[26183] = 32'b00000000000000000011011001001011;
assign LUT_4[26184] = 32'b00000000000000000110111110101000;
assign LUT_4[26185] = 32'b00000000000000000000001010100000;
assign LUT_4[26186] = 32'b00000000000000000110011001001100;
assign LUT_4[26187] = 32'b11111111111111111111100101000100;
assign LUT_4[26188] = 32'b00000000000000000011111111000100;
assign LUT_4[26189] = 32'b11111111111111111101001010111100;
assign LUT_4[26190] = 32'b00000000000000000011011001101000;
assign LUT_4[26191] = 32'b11111111111111111100100101100000;
assign LUT_4[26192] = 32'b00000000000000001011100100000001;
assign LUT_4[26193] = 32'b00000000000000000100101111111001;
assign LUT_4[26194] = 32'b00000000000000001010111110100101;
assign LUT_4[26195] = 32'b00000000000000000100001010011101;
assign LUT_4[26196] = 32'b00000000000000001000100100011101;
assign LUT_4[26197] = 32'b00000000000000000001110000010101;
assign LUT_4[26198] = 32'b00000000000000000111111111000001;
assign LUT_4[26199] = 32'b00000000000000000001001010111001;
assign LUT_4[26200] = 32'b00000000000000000100110000010110;
assign LUT_4[26201] = 32'b11111111111111111101111100001110;
assign LUT_4[26202] = 32'b00000000000000000100001010111010;
assign LUT_4[26203] = 32'b11111111111111111101010110110010;
assign LUT_4[26204] = 32'b00000000000000000001110000110010;
assign LUT_4[26205] = 32'b11111111111111111010111100101010;
assign LUT_4[26206] = 32'b00000000000000000001001011010110;
assign LUT_4[26207] = 32'b11111111111111111010010111001110;
assign LUT_4[26208] = 32'b00000000000000001100001101011010;
assign LUT_4[26209] = 32'b00000000000000000101011001010010;
assign LUT_4[26210] = 32'b00000000000000001011100111111110;
assign LUT_4[26211] = 32'b00000000000000000100110011110110;
assign LUT_4[26212] = 32'b00000000000000001001001101110110;
assign LUT_4[26213] = 32'b00000000000000000010011001101110;
assign LUT_4[26214] = 32'b00000000000000001000101000011010;
assign LUT_4[26215] = 32'b00000000000000000001110100010010;
assign LUT_4[26216] = 32'b00000000000000000101011001101111;
assign LUT_4[26217] = 32'b11111111111111111110100101100111;
assign LUT_4[26218] = 32'b00000000000000000100110100010011;
assign LUT_4[26219] = 32'b11111111111111111110000000001011;
assign LUT_4[26220] = 32'b00000000000000000010011010001011;
assign LUT_4[26221] = 32'b11111111111111111011100110000011;
assign LUT_4[26222] = 32'b00000000000000000001110100101111;
assign LUT_4[26223] = 32'b11111111111111111011000000100111;
assign LUT_4[26224] = 32'b00000000000000001001111111001000;
assign LUT_4[26225] = 32'b00000000000000000011001011000000;
assign LUT_4[26226] = 32'b00000000000000001001011001101100;
assign LUT_4[26227] = 32'b00000000000000000010100101100100;
assign LUT_4[26228] = 32'b00000000000000000110111111100100;
assign LUT_4[26229] = 32'b00000000000000000000001011011100;
assign LUT_4[26230] = 32'b00000000000000000110011010001000;
assign LUT_4[26231] = 32'b11111111111111111111100110000000;
assign LUT_4[26232] = 32'b00000000000000000011001011011101;
assign LUT_4[26233] = 32'b11111111111111111100010111010101;
assign LUT_4[26234] = 32'b00000000000000000010100110000001;
assign LUT_4[26235] = 32'b11111111111111111011110001111001;
assign LUT_4[26236] = 32'b00000000000000000000001011111001;
assign LUT_4[26237] = 32'b11111111111111111001010111110001;
assign LUT_4[26238] = 32'b11111111111111111111100110011101;
assign LUT_4[26239] = 32'b11111111111111111000110010010101;
assign LUT_4[26240] = 32'b00000000000000001111000001000111;
assign LUT_4[26241] = 32'b00000000000000001000001100111111;
assign LUT_4[26242] = 32'b00000000000000001110011011101011;
assign LUT_4[26243] = 32'b00000000000000000111100111100011;
assign LUT_4[26244] = 32'b00000000000000001100000001100011;
assign LUT_4[26245] = 32'b00000000000000000101001101011011;
assign LUT_4[26246] = 32'b00000000000000001011011100000111;
assign LUT_4[26247] = 32'b00000000000000000100100111111111;
assign LUT_4[26248] = 32'b00000000000000001000001101011100;
assign LUT_4[26249] = 32'b00000000000000000001011001010100;
assign LUT_4[26250] = 32'b00000000000000000111101000000000;
assign LUT_4[26251] = 32'b00000000000000000000110011111000;
assign LUT_4[26252] = 32'b00000000000000000101001101111000;
assign LUT_4[26253] = 32'b11111111111111111110011001110000;
assign LUT_4[26254] = 32'b00000000000000000100101000011100;
assign LUT_4[26255] = 32'b11111111111111111101110100010100;
assign LUT_4[26256] = 32'b00000000000000001100110010110101;
assign LUT_4[26257] = 32'b00000000000000000101111110101101;
assign LUT_4[26258] = 32'b00000000000000001100001101011001;
assign LUT_4[26259] = 32'b00000000000000000101011001010001;
assign LUT_4[26260] = 32'b00000000000000001001110011010001;
assign LUT_4[26261] = 32'b00000000000000000010111111001001;
assign LUT_4[26262] = 32'b00000000000000001001001101110101;
assign LUT_4[26263] = 32'b00000000000000000010011001101101;
assign LUT_4[26264] = 32'b00000000000000000101111111001010;
assign LUT_4[26265] = 32'b11111111111111111111001011000010;
assign LUT_4[26266] = 32'b00000000000000000101011001101110;
assign LUT_4[26267] = 32'b11111111111111111110100101100110;
assign LUT_4[26268] = 32'b00000000000000000010111111100110;
assign LUT_4[26269] = 32'b11111111111111111100001011011110;
assign LUT_4[26270] = 32'b00000000000000000010011010001010;
assign LUT_4[26271] = 32'b11111111111111111011100110000010;
assign LUT_4[26272] = 32'b00000000000000001101011100001110;
assign LUT_4[26273] = 32'b00000000000000000110101000000110;
assign LUT_4[26274] = 32'b00000000000000001100110110110010;
assign LUT_4[26275] = 32'b00000000000000000110000010101010;
assign LUT_4[26276] = 32'b00000000000000001010011100101010;
assign LUT_4[26277] = 32'b00000000000000000011101000100010;
assign LUT_4[26278] = 32'b00000000000000001001110111001110;
assign LUT_4[26279] = 32'b00000000000000000011000011000110;
assign LUT_4[26280] = 32'b00000000000000000110101000100011;
assign LUT_4[26281] = 32'b11111111111111111111110100011011;
assign LUT_4[26282] = 32'b00000000000000000110000011000111;
assign LUT_4[26283] = 32'b11111111111111111111001110111111;
assign LUT_4[26284] = 32'b00000000000000000011101000111111;
assign LUT_4[26285] = 32'b11111111111111111100110100110111;
assign LUT_4[26286] = 32'b00000000000000000011000011100011;
assign LUT_4[26287] = 32'b11111111111111111100001111011011;
assign LUT_4[26288] = 32'b00000000000000001011001101111100;
assign LUT_4[26289] = 32'b00000000000000000100011001110100;
assign LUT_4[26290] = 32'b00000000000000001010101000100000;
assign LUT_4[26291] = 32'b00000000000000000011110100011000;
assign LUT_4[26292] = 32'b00000000000000001000001110011000;
assign LUT_4[26293] = 32'b00000000000000000001011010010000;
assign LUT_4[26294] = 32'b00000000000000000111101000111100;
assign LUT_4[26295] = 32'b00000000000000000000110100110100;
assign LUT_4[26296] = 32'b00000000000000000100011010010001;
assign LUT_4[26297] = 32'b11111111111111111101100110001001;
assign LUT_4[26298] = 32'b00000000000000000011110100110101;
assign LUT_4[26299] = 32'b11111111111111111101000000101101;
assign LUT_4[26300] = 32'b00000000000000000001011010101101;
assign LUT_4[26301] = 32'b11111111111111111010100110100101;
assign LUT_4[26302] = 32'b00000000000000000000110101010001;
assign LUT_4[26303] = 32'b11111111111111111010000001001001;
assign LUT_4[26304] = 32'b00000000000000010000011000011011;
assign LUT_4[26305] = 32'b00000000000000001001100100010011;
assign LUT_4[26306] = 32'b00000000000000001111110010111111;
assign LUT_4[26307] = 32'b00000000000000001000111110110111;
assign LUT_4[26308] = 32'b00000000000000001101011000110111;
assign LUT_4[26309] = 32'b00000000000000000110100100101111;
assign LUT_4[26310] = 32'b00000000000000001100110011011011;
assign LUT_4[26311] = 32'b00000000000000000101111111010011;
assign LUT_4[26312] = 32'b00000000000000001001100100110000;
assign LUT_4[26313] = 32'b00000000000000000010110000101000;
assign LUT_4[26314] = 32'b00000000000000001000111111010100;
assign LUT_4[26315] = 32'b00000000000000000010001011001100;
assign LUT_4[26316] = 32'b00000000000000000110100101001100;
assign LUT_4[26317] = 32'b11111111111111111111110001000100;
assign LUT_4[26318] = 32'b00000000000000000101111111110000;
assign LUT_4[26319] = 32'b11111111111111111111001011101000;
assign LUT_4[26320] = 32'b00000000000000001110001010001001;
assign LUT_4[26321] = 32'b00000000000000000111010110000001;
assign LUT_4[26322] = 32'b00000000000000001101100100101101;
assign LUT_4[26323] = 32'b00000000000000000110110000100101;
assign LUT_4[26324] = 32'b00000000000000001011001010100101;
assign LUT_4[26325] = 32'b00000000000000000100010110011101;
assign LUT_4[26326] = 32'b00000000000000001010100101001001;
assign LUT_4[26327] = 32'b00000000000000000011110001000001;
assign LUT_4[26328] = 32'b00000000000000000111010110011110;
assign LUT_4[26329] = 32'b00000000000000000000100010010110;
assign LUT_4[26330] = 32'b00000000000000000110110001000010;
assign LUT_4[26331] = 32'b11111111111111111111111100111010;
assign LUT_4[26332] = 32'b00000000000000000100010110111010;
assign LUT_4[26333] = 32'b11111111111111111101100010110010;
assign LUT_4[26334] = 32'b00000000000000000011110001011110;
assign LUT_4[26335] = 32'b11111111111111111100111101010110;
assign LUT_4[26336] = 32'b00000000000000001110110011100010;
assign LUT_4[26337] = 32'b00000000000000000111111111011010;
assign LUT_4[26338] = 32'b00000000000000001110001110000110;
assign LUT_4[26339] = 32'b00000000000000000111011001111110;
assign LUT_4[26340] = 32'b00000000000000001011110011111110;
assign LUT_4[26341] = 32'b00000000000000000100111111110110;
assign LUT_4[26342] = 32'b00000000000000001011001110100010;
assign LUT_4[26343] = 32'b00000000000000000100011010011010;
assign LUT_4[26344] = 32'b00000000000000000111111111110111;
assign LUT_4[26345] = 32'b00000000000000000001001011101111;
assign LUT_4[26346] = 32'b00000000000000000111011010011011;
assign LUT_4[26347] = 32'b00000000000000000000100110010011;
assign LUT_4[26348] = 32'b00000000000000000101000000010011;
assign LUT_4[26349] = 32'b11111111111111111110001100001011;
assign LUT_4[26350] = 32'b00000000000000000100011010110111;
assign LUT_4[26351] = 32'b11111111111111111101100110101111;
assign LUT_4[26352] = 32'b00000000000000001100100101010000;
assign LUT_4[26353] = 32'b00000000000000000101110001001000;
assign LUT_4[26354] = 32'b00000000000000001011111111110100;
assign LUT_4[26355] = 32'b00000000000000000101001011101100;
assign LUT_4[26356] = 32'b00000000000000001001100101101100;
assign LUT_4[26357] = 32'b00000000000000000010110001100100;
assign LUT_4[26358] = 32'b00000000000000001001000000010000;
assign LUT_4[26359] = 32'b00000000000000000010001100001000;
assign LUT_4[26360] = 32'b00000000000000000101110001100101;
assign LUT_4[26361] = 32'b11111111111111111110111101011101;
assign LUT_4[26362] = 32'b00000000000000000101001100001001;
assign LUT_4[26363] = 32'b11111111111111111110011000000001;
assign LUT_4[26364] = 32'b00000000000000000010110010000001;
assign LUT_4[26365] = 32'b11111111111111111011111101111001;
assign LUT_4[26366] = 32'b00000000000000000010001100100101;
assign LUT_4[26367] = 32'b11111111111111111011011000011101;
assign LUT_4[26368] = 32'b00000000000000010001010110100010;
assign LUT_4[26369] = 32'b00000000000000001010100010011010;
assign LUT_4[26370] = 32'b00000000000000010000110001000110;
assign LUT_4[26371] = 32'b00000000000000001001111100111110;
assign LUT_4[26372] = 32'b00000000000000001110010110111110;
assign LUT_4[26373] = 32'b00000000000000000111100010110110;
assign LUT_4[26374] = 32'b00000000000000001101110001100010;
assign LUT_4[26375] = 32'b00000000000000000110111101011010;
assign LUT_4[26376] = 32'b00000000000000001010100010110111;
assign LUT_4[26377] = 32'b00000000000000000011101110101111;
assign LUT_4[26378] = 32'b00000000000000001001111101011011;
assign LUT_4[26379] = 32'b00000000000000000011001001010011;
assign LUT_4[26380] = 32'b00000000000000000111100011010011;
assign LUT_4[26381] = 32'b00000000000000000000101111001011;
assign LUT_4[26382] = 32'b00000000000000000110111101110111;
assign LUT_4[26383] = 32'b00000000000000000000001001101111;
assign LUT_4[26384] = 32'b00000000000000001111001000010000;
assign LUT_4[26385] = 32'b00000000000000001000010100001000;
assign LUT_4[26386] = 32'b00000000000000001110100010110100;
assign LUT_4[26387] = 32'b00000000000000000111101110101100;
assign LUT_4[26388] = 32'b00000000000000001100001000101100;
assign LUT_4[26389] = 32'b00000000000000000101010100100100;
assign LUT_4[26390] = 32'b00000000000000001011100011010000;
assign LUT_4[26391] = 32'b00000000000000000100101111001000;
assign LUT_4[26392] = 32'b00000000000000001000010100100101;
assign LUT_4[26393] = 32'b00000000000000000001100000011101;
assign LUT_4[26394] = 32'b00000000000000000111101111001001;
assign LUT_4[26395] = 32'b00000000000000000000111011000001;
assign LUT_4[26396] = 32'b00000000000000000101010101000001;
assign LUT_4[26397] = 32'b11111111111111111110100000111001;
assign LUT_4[26398] = 32'b00000000000000000100101111100101;
assign LUT_4[26399] = 32'b11111111111111111101111011011101;
assign LUT_4[26400] = 32'b00000000000000001111110001101001;
assign LUT_4[26401] = 32'b00000000000000001000111101100001;
assign LUT_4[26402] = 32'b00000000000000001111001100001101;
assign LUT_4[26403] = 32'b00000000000000001000011000000101;
assign LUT_4[26404] = 32'b00000000000000001100110010000101;
assign LUT_4[26405] = 32'b00000000000000000101111101111101;
assign LUT_4[26406] = 32'b00000000000000001100001100101001;
assign LUT_4[26407] = 32'b00000000000000000101011000100001;
assign LUT_4[26408] = 32'b00000000000000001000111101111110;
assign LUT_4[26409] = 32'b00000000000000000010001001110110;
assign LUT_4[26410] = 32'b00000000000000001000011000100010;
assign LUT_4[26411] = 32'b00000000000000000001100100011010;
assign LUT_4[26412] = 32'b00000000000000000101111110011010;
assign LUT_4[26413] = 32'b11111111111111111111001010010010;
assign LUT_4[26414] = 32'b00000000000000000101011000111110;
assign LUT_4[26415] = 32'b11111111111111111110100100110110;
assign LUT_4[26416] = 32'b00000000000000001101100011010111;
assign LUT_4[26417] = 32'b00000000000000000110101111001111;
assign LUT_4[26418] = 32'b00000000000000001100111101111011;
assign LUT_4[26419] = 32'b00000000000000000110001001110011;
assign LUT_4[26420] = 32'b00000000000000001010100011110011;
assign LUT_4[26421] = 32'b00000000000000000011101111101011;
assign LUT_4[26422] = 32'b00000000000000001001111110010111;
assign LUT_4[26423] = 32'b00000000000000000011001010001111;
assign LUT_4[26424] = 32'b00000000000000000110101111101100;
assign LUT_4[26425] = 32'b11111111111111111111111011100100;
assign LUT_4[26426] = 32'b00000000000000000110001010010000;
assign LUT_4[26427] = 32'b11111111111111111111010110001000;
assign LUT_4[26428] = 32'b00000000000000000011110000001000;
assign LUT_4[26429] = 32'b11111111111111111100111100000000;
assign LUT_4[26430] = 32'b00000000000000000011001010101100;
assign LUT_4[26431] = 32'b11111111111111111100010110100100;
assign LUT_4[26432] = 32'b00000000000000010010101101110110;
assign LUT_4[26433] = 32'b00000000000000001011111001101110;
assign LUT_4[26434] = 32'b00000000000000010010001000011010;
assign LUT_4[26435] = 32'b00000000000000001011010100010010;
assign LUT_4[26436] = 32'b00000000000000001111101110010010;
assign LUT_4[26437] = 32'b00000000000000001000111010001010;
assign LUT_4[26438] = 32'b00000000000000001111001000110110;
assign LUT_4[26439] = 32'b00000000000000001000010100101110;
assign LUT_4[26440] = 32'b00000000000000001011111010001011;
assign LUT_4[26441] = 32'b00000000000000000101000110000011;
assign LUT_4[26442] = 32'b00000000000000001011010100101111;
assign LUT_4[26443] = 32'b00000000000000000100100000100111;
assign LUT_4[26444] = 32'b00000000000000001000111010100111;
assign LUT_4[26445] = 32'b00000000000000000010000110011111;
assign LUT_4[26446] = 32'b00000000000000001000010101001011;
assign LUT_4[26447] = 32'b00000000000000000001100001000011;
assign LUT_4[26448] = 32'b00000000000000010000011111100100;
assign LUT_4[26449] = 32'b00000000000000001001101011011100;
assign LUT_4[26450] = 32'b00000000000000001111111010001000;
assign LUT_4[26451] = 32'b00000000000000001001000110000000;
assign LUT_4[26452] = 32'b00000000000000001101100000000000;
assign LUT_4[26453] = 32'b00000000000000000110101011111000;
assign LUT_4[26454] = 32'b00000000000000001100111010100100;
assign LUT_4[26455] = 32'b00000000000000000110000110011100;
assign LUT_4[26456] = 32'b00000000000000001001101011111001;
assign LUT_4[26457] = 32'b00000000000000000010110111110001;
assign LUT_4[26458] = 32'b00000000000000001001000110011101;
assign LUT_4[26459] = 32'b00000000000000000010010010010101;
assign LUT_4[26460] = 32'b00000000000000000110101100010101;
assign LUT_4[26461] = 32'b11111111111111111111111000001101;
assign LUT_4[26462] = 32'b00000000000000000110000110111001;
assign LUT_4[26463] = 32'b11111111111111111111010010110001;
assign LUT_4[26464] = 32'b00000000000000010001001000111101;
assign LUT_4[26465] = 32'b00000000000000001010010100110101;
assign LUT_4[26466] = 32'b00000000000000010000100011100001;
assign LUT_4[26467] = 32'b00000000000000001001101111011001;
assign LUT_4[26468] = 32'b00000000000000001110001001011001;
assign LUT_4[26469] = 32'b00000000000000000111010101010001;
assign LUT_4[26470] = 32'b00000000000000001101100011111101;
assign LUT_4[26471] = 32'b00000000000000000110101111110101;
assign LUT_4[26472] = 32'b00000000000000001010010101010010;
assign LUT_4[26473] = 32'b00000000000000000011100001001010;
assign LUT_4[26474] = 32'b00000000000000001001101111110110;
assign LUT_4[26475] = 32'b00000000000000000010111011101110;
assign LUT_4[26476] = 32'b00000000000000000111010101101110;
assign LUT_4[26477] = 32'b00000000000000000000100001100110;
assign LUT_4[26478] = 32'b00000000000000000110110000010010;
assign LUT_4[26479] = 32'b11111111111111111111111100001010;
assign LUT_4[26480] = 32'b00000000000000001110111010101011;
assign LUT_4[26481] = 32'b00000000000000001000000110100011;
assign LUT_4[26482] = 32'b00000000000000001110010101001111;
assign LUT_4[26483] = 32'b00000000000000000111100001000111;
assign LUT_4[26484] = 32'b00000000000000001011111011000111;
assign LUT_4[26485] = 32'b00000000000000000101000110111111;
assign LUT_4[26486] = 32'b00000000000000001011010101101011;
assign LUT_4[26487] = 32'b00000000000000000100100001100011;
assign LUT_4[26488] = 32'b00000000000000001000000111000000;
assign LUT_4[26489] = 32'b00000000000000000001010010111000;
assign LUT_4[26490] = 32'b00000000000000000111100001100100;
assign LUT_4[26491] = 32'b00000000000000000000101101011100;
assign LUT_4[26492] = 32'b00000000000000000101000111011100;
assign LUT_4[26493] = 32'b11111111111111111110010011010100;
assign LUT_4[26494] = 32'b00000000000000000100100010000000;
assign LUT_4[26495] = 32'b11111111111111111101101101111000;
assign LUT_4[26496] = 32'b00000000000000010011111100101010;
assign LUT_4[26497] = 32'b00000000000000001101001000100010;
assign LUT_4[26498] = 32'b00000000000000010011010111001110;
assign LUT_4[26499] = 32'b00000000000000001100100011000110;
assign LUT_4[26500] = 32'b00000000000000010000111101000110;
assign LUT_4[26501] = 32'b00000000000000001010001000111110;
assign LUT_4[26502] = 32'b00000000000000010000010111101010;
assign LUT_4[26503] = 32'b00000000000000001001100011100010;
assign LUT_4[26504] = 32'b00000000000000001101001000111111;
assign LUT_4[26505] = 32'b00000000000000000110010100110111;
assign LUT_4[26506] = 32'b00000000000000001100100011100011;
assign LUT_4[26507] = 32'b00000000000000000101101111011011;
assign LUT_4[26508] = 32'b00000000000000001010001001011011;
assign LUT_4[26509] = 32'b00000000000000000011010101010011;
assign LUT_4[26510] = 32'b00000000000000001001100011111111;
assign LUT_4[26511] = 32'b00000000000000000010101111110111;
assign LUT_4[26512] = 32'b00000000000000010001101110011000;
assign LUT_4[26513] = 32'b00000000000000001010111010010000;
assign LUT_4[26514] = 32'b00000000000000010001001000111100;
assign LUT_4[26515] = 32'b00000000000000001010010100110100;
assign LUT_4[26516] = 32'b00000000000000001110101110110100;
assign LUT_4[26517] = 32'b00000000000000000111111010101100;
assign LUT_4[26518] = 32'b00000000000000001110001001011000;
assign LUT_4[26519] = 32'b00000000000000000111010101010000;
assign LUT_4[26520] = 32'b00000000000000001010111010101101;
assign LUT_4[26521] = 32'b00000000000000000100000110100101;
assign LUT_4[26522] = 32'b00000000000000001010010101010001;
assign LUT_4[26523] = 32'b00000000000000000011100001001001;
assign LUT_4[26524] = 32'b00000000000000000111111011001001;
assign LUT_4[26525] = 32'b00000000000000000001000111000001;
assign LUT_4[26526] = 32'b00000000000000000111010101101101;
assign LUT_4[26527] = 32'b00000000000000000000100001100101;
assign LUT_4[26528] = 32'b00000000000000010010010111110001;
assign LUT_4[26529] = 32'b00000000000000001011100011101001;
assign LUT_4[26530] = 32'b00000000000000010001110010010101;
assign LUT_4[26531] = 32'b00000000000000001010111110001101;
assign LUT_4[26532] = 32'b00000000000000001111011000001101;
assign LUT_4[26533] = 32'b00000000000000001000100100000101;
assign LUT_4[26534] = 32'b00000000000000001110110010110001;
assign LUT_4[26535] = 32'b00000000000000000111111110101001;
assign LUT_4[26536] = 32'b00000000000000001011100100000110;
assign LUT_4[26537] = 32'b00000000000000000100101111111110;
assign LUT_4[26538] = 32'b00000000000000001010111110101010;
assign LUT_4[26539] = 32'b00000000000000000100001010100010;
assign LUT_4[26540] = 32'b00000000000000001000100100100010;
assign LUT_4[26541] = 32'b00000000000000000001110000011010;
assign LUT_4[26542] = 32'b00000000000000000111111111000110;
assign LUT_4[26543] = 32'b00000000000000000001001010111110;
assign LUT_4[26544] = 32'b00000000000000010000001001011111;
assign LUT_4[26545] = 32'b00000000000000001001010101010111;
assign LUT_4[26546] = 32'b00000000000000001111100100000011;
assign LUT_4[26547] = 32'b00000000000000001000101111111011;
assign LUT_4[26548] = 32'b00000000000000001101001001111011;
assign LUT_4[26549] = 32'b00000000000000000110010101110011;
assign LUT_4[26550] = 32'b00000000000000001100100100011111;
assign LUT_4[26551] = 32'b00000000000000000101110000010111;
assign LUT_4[26552] = 32'b00000000000000001001010101110100;
assign LUT_4[26553] = 32'b00000000000000000010100001101100;
assign LUT_4[26554] = 32'b00000000000000001000110000011000;
assign LUT_4[26555] = 32'b00000000000000000001111100010000;
assign LUT_4[26556] = 32'b00000000000000000110010110010000;
assign LUT_4[26557] = 32'b11111111111111111111100010001000;
assign LUT_4[26558] = 32'b00000000000000000101110000110100;
assign LUT_4[26559] = 32'b11111111111111111110111100101100;
assign LUT_4[26560] = 32'b00000000000000010101010011111110;
assign LUT_4[26561] = 32'b00000000000000001110011111110110;
assign LUT_4[26562] = 32'b00000000000000010100101110100010;
assign LUT_4[26563] = 32'b00000000000000001101111010011010;
assign LUT_4[26564] = 32'b00000000000000010010010100011010;
assign LUT_4[26565] = 32'b00000000000000001011100000010010;
assign LUT_4[26566] = 32'b00000000000000010001101110111110;
assign LUT_4[26567] = 32'b00000000000000001010111010110110;
assign LUT_4[26568] = 32'b00000000000000001110100000010011;
assign LUT_4[26569] = 32'b00000000000000000111101100001011;
assign LUT_4[26570] = 32'b00000000000000001101111010110111;
assign LUT_4[26571] = 32'b00000000000000000111000110101111;
assign LUT_4[26572] = 32'b00000000000000001011100000101111;
assign LUT_4[26573] = 32'b00000000000000000100101100100111;
assign LUT_4[26574] = 32'b00000000000000001010111011010011;
assign LUT_4[26575] = 32'b00000000000000000100000111001011;
assign LUT_4[26576] = 32'b00000000000000010011000101101100;
assign LUT_4[26577] = 32'b00000000000000001100010001100100;
assign LUT_4[26578] = 32'b00000000000000010010100000010000;
assign LUT_4[26579] = 32'b00000000000000001011101100001000;
assign LUT_4[26580] = 32'b00000000000000010000000110001000;
assign LUT_4[26581] = 32'b00000000000000001001010010000000;
assign LUT_4[26582] = 32'b00000000000000001111100000101100;
assign LUT_4[26583] = 32'b00000000000000001000101100100100;
assign LUT_4[26584] = 32'b00000000000000001100010010000001;
assign LUT_4[26585] = 32'b00000000000000000101011101111001;
assign LUT_4[26586] = 32'b00000000000000001011101100100101;
assign LUT_4[26587] = 32'b00000000000000000100111000011101;
assign LUT_4[26588] = 32'b00000000000000001001010010011101;
assign LUT_4[26589] = 32'b00000000000000000010011110010101;
assign LUT_4[26590] = 32'b00000000000000001000101101000001;
assign LUT_4[26591] = 32'b00000000000000000001111000111001;
assign LUT_4[26592] = 32'b00000000000000010011101111000101;
assign LUT_4[26593] = 32'b00000000000000001100111010111101;
assign LUT_4[26594] = 32'b00000000000000010011001001101001;
assign LUT_4[26595] = 32'b00000000000000001100010101100001;
assign LUT_4[26596] = 32'b00000000000000010000101111100001;
assign LUT_4[26597] = 32'b00000000000000001001111011011001;
assign LUT_4[26598] = 32'b00000000000000010000001010000101;
assign LUT_4[26599] = 32'b00000000000000001001010101111101;
assign LUT_4[26600] = 32'b00000000000000001100111011011010;
assign LUT_4[26601] = 32'b00000000000000000110000111010010;
assign LUT_4[26602] = 32'b00000000000000001100010101111110;
assign LUT_4[26603] = 32'b00000000000000000101100001110110;
assign LUT_4[26604] = 32'b00000000000000001001111011110110;
assign LUT_4[26605] = 32'b00000000000000000011000111101110;
assign LUT_4[26606] = 32'b00000000000000001001010110011010;
assign LUT_4[26607] = 32'b00000000000000000010100010010010;
assign LUT_4[26608] = 32'b00000000000000010001100000110011;
assign LUT_4[26609] = 32'b00000000000000001010101100101011;
assign LUT_4[26610] = 32'b00000000000000010000111011010111;
assign LUT_4[26611] = 32'b00000000000000001010000111001111;
assign LUT_4[26612] = 32'b00000000000000001110100001001111;
assign LUT_4[26613] = 32'b00000000000000000111101101000111;
assign LUT_4[26614] = 32'b00000000000000001101111011110011;
assign LUT_4[26615] = 32'b00000000000000000111000111101011;
assign LUT_4[26616] = 32'b00000000000000001010101101001000;
assign LUT_4[26617] = 32'b00000000000000000011111001000000;
assign LUT_4[26618] = 32'b00000000000000001010000111101100;
assign LUT_4[26619] = 32'b00000000000000000011010011100100;
assign LUT_4[26620] = 32'b00000000000000000111101101100100;
assign LUT_4[26621] = 32'b00000000000000000000111001011100;
assign LUT_4[26622] = 32'b00000000000000000111001000001000;
assign LUT_4[26623] = 32'b00000000000000000000010100000000;
assign LUT_4[26624] = 32'b00000000000000000111001011100010;
assign LUT_4[26625] = 32'b00000000000000000000010111011010;
assign LUT_4[26626] = 32'b00000000000000000110100110000110;
assign LUT_4[26627] = 32'b11111111111111111111110001111110;
assign LUT_4[26628] = 32'b00000000000000000100001011111110;
assign LUT_4[26629] = 32'b11111111111111111101010111110110;
assign LUT_4[26630] = 32'b00000000000000000011100110100010;
assign LUT_4[26631] = 32'b11111111111111111100110010011010;
assign LUT_4[26632] = 32'b00000000000000000000010111110111;
assign LUT_4[26633] = 32'b11111111111111111001100011101111;
assign LUT_4[26634] = 32'b11111111111111111111110010011011;
assign LUT_4[26635] = 32'b11111111111111111000111110010011;
assign LUT_4[26636] = 32'b11111111111111111101011000010011;
assign LUT_4[26637] = 32'b11111111111111110110100100001011;
assign LUT_4[26638] = 32'b11111111111111111100110010110111;
assign LUT_4[26639] = 32'b11111111111111110101111110101111;
assign LUT_4[26640] = 32'b00000000000000000100111101010000;
assign LUT_4[26641] = 32'b11111111111111111110001001001000;
assign LUT_4[26642] = 32'b00000000000000000100010111110100;
assign LUT_4[26643] = 32'b11111111111111111101100011101100;
assign LUT_4[26644] = 32'b00000000000000000001111101101100;
assign LUT_4[26645] = 32'b11111111111111111011001001100100;
assign LUT_4[26646] = 32'b00000000000000000001011000010000;
assign LUT_4[26647] = 32'b11111111111111111010100100001000;
assign LUT_4[26648] = 32'b11111111111111111110001001100101;
assign LUT_4[26649] = 32'b11111111111111110111010101011101;
assign LUT_4[26650] = 32'b11111111111111111101100100001001;
assign LUT_4[26651] = 32'b11111111111111110110110000000001;
assign LUT_4[26652] = 32'b11111111111111111011001010000001;
assign LUT_4[26653] = 32'b11111111111111110100010101111001;
assign LUT_4[26654] = 32'b11111111111111111010100100100101;
assign LUT_4[26655] = 32'b11111111111111110011110000011101;
assign LUT_4[26656] = 32'b00000000000000000101100110101001;
assign LUT_4[26657] = 32'b11111111111111111110110010100001;
assign LUT_4[26658] = 32'b00000000000000000101000001001101;
assign LUT_4[26659] = 32'b11111111111111111110001101000101;
assign LUT_4[26660] = 32'b00000000000000000010100111000101;
assign LUT_4[26661] = 32'b11111111111111111011110010111101;
assign LUT_4[26662] = 32'b00000000000000000010000001101001;
assign LUT_4[26663] = 32'b11111111111111111011001101100001;
assign LUT_4[26664] = 32'b11111111111111111110110010111110;
assign LUT_4[26665] = 32'b11111111111111110111111110110110;
assign LUT_4[26666] = 32'b11111111111111111110001101100010;
assign LUT_4[26667] = 32'b11111111111111110111011001011010;
assign LUT_4[26668] = 32'b11111111111111111011110011011010;
assign LUT_4[26669] = 32'b11111111111111110100111111010010;
assign LUT_4[26670] = 32'b11111111111111111011001101111110;
assign LUT_4[26671] = 32'b11111111111111110100011001110110;
assign LUT_4[26672] = 32'b00000000000000000011011000010111;
assign LUT_4[26673] = 32'b11111111111111111100100100001111;
assign LUT_4[26674] = 32'b00000000000000000010110010111011;
assign LUT_4[26675] = 32'b11111111111111111011111110110011;
assign LUT_4[26676] = 32'b00000000000000000000011000110011;
assign LUT_4[26677] = 32'b11111111111111111001100100101011;
assign LUT_4[26678] = 32'b11111111111111111111110011010111;
assign LUT_4[26679] = 32'b11111111111111111000111111001111;
assign LUT_4[26680] = 32'b11111111111111111100100100101100;
assign LUT_4[26681] = 32'b11111111111111110101110000100100;
assign LUT_4[26682] = 32'b11111111111111111011111111010000;
assign LUT_4[26683] = 32'b11111111111111110101001011001000;
assign LUT_4[26684] = 32'b11111111111111111001100101001000;
assign LUT_4[26685] = 32'b11111111111111110010110001000000;
assign LUT_4[26686] = 32'b11111111111111111000111111101100;
assign LUT_4[26687] = 32'b11111111111111110010001011100100;
assign LUT_4[26688] = 32'b00000000000000001000100010110110;
assign LUT_4[26689] = 32'b00000000000000000001101110101110;
assign LUT_4[26690] = 32'b00000000000000000111111101011010;
assign LUT_4[26691] = 32'b00000000000000000001001001010010;
assign LUT_4[26692] = 32'b00000000000000000101100011010010;
assign LUT_4[26693] = 32'b11111111111111111110101111001010;
assign LUT_4[26694] = 32'b00000000000000000100111101110110;
assign LUT_4[26695] = 32'b11111111111111111110001001101110;
assign LUT_4[26696] = 32'b00000000000000000001101111001011;
assign LUT_4[26697] = 32'b11111111111111111010111011000011;
assign LUT_4[26698] = 32'b00000000000000000001001001101111;
assign LUT_4[26699] = 32'b11111111111111111010010101100111;
assign LUT_4[26700] = 32'b11111111111111111110101111100111;
assign LUT_4[26701] = 32'b11111111111111110111111011011111;
assign LUT_4[26702] = 32'b11111111111111111110001010001011;
assign LUT_4[26703] = 32'b11111111111111110111010110000011;
assign LUT_4[26704] = 32'b00000000000000000110010100100100;
assign LUT_4[26705] = 32'b11111111111111111111100000011100;
assign LUT_4[26706] = 32'b00000000000000000101101111001000;
assign LUT_4[26707] = 32'b11111111111111111110111011000000;
assign LUT_4[26708] = 32'b00000000000000000011010101000000;
assign LUT_4[26709] = 32'b11111111111111111100100000111000;
assign LUT_4[26710] = 32'b00000000000000000010101111100100;
assign LUT_4[26711] = 32'b11111111111111111011111011011100;
assign LUT_4[26712] = 32'b11111111111111111111100000111001;
assign LUT_4[26713] = 32'b11111111111111111000101100110001;
assign LUT_4[26714] = 32'b11111111111111111110111011011101;
assign LUT_4[26715] = 32'b11111111111111111000000111010101;
assign LUT_4[26716] = 32'b11111111111111111100100001010101;
assign LUT_4[26717] = 32'b11111111111111110101101101001101;
assign LUT_4[26718] = 32'b11111111111111111011111011111001;
assign LUT_4[26719] = 32'b11111111111111110101000111110001;
assign LUT_4[26720] = 32'b00000000000000000110111101111101;
assign LUT_4[26721] = 32'b00000000000000000000001001110101;
assign LUT_4[26722] = 32'b00000000000000000110011000100001;
assign LUT_4[26723] = 32'b11111111111111111111100100011001;
assign LUT_4[26724] = 32'b00000000000000000011111110011001;
assign LUT_4[26725] = 32'b11111111111111111101001010010001;
assign LUT_4[26726] = 32'b00000000000000000011011000111101;
assign LUT_4[26727] = 32'b11111111111111111100100100110101;
assign LUT_4[26728] = 32'b00000000000000000000001010010010;
assign LUT_4[26729] = 32'b11111111111111111001010110001010;
assign LUT_4[26730] = 32'b11111111111111111111100100110110;
assign LUT_4[26731] = 32'b11111111111111111000110000101110;
assign LUT_4[26732] = 32'b11111111111111111101001010101110;
assign LUT_4[26733] = 32'b11111111111111110110010110100110;
assign LUT_4[26734] = 32'b11111111111111111100100101010010;
assign LUT_4[26735] = 32'b11111111111111110101110001001010;
assign LUT_4[26736] = 32'b00000000000000000100101111101011;
assign LUT_4[26737] = 32'b11111111111111111101111011100011;
assign LUT_4[26738] = 32'b00000000000000000100001010001111;
assign LUT_4[26739] = 32'b11111111111111111101010110000111;
assign LUT_4[26740] = 32'b00000000000000000001110000000111;
assign LUT_4[26741] = 32'b11111111111111111010111011111111;
assign LUT_4[26742] = 32'b00000000000000000001001010101011;
assign LUT_4[26743] = 32'b11111111111111111010010110100011;
assign LUT_4[26744] = 32'b11111111111111111101111100000000;
assign LUT_4[26745] = 32'b11111111111111110111000111111000;
assign LUT_4[26746] = 32'b11111111111111111101010110100100;
assign LUT_4[26747] = 32'b11111111111111110110100010011100;
assign LUT_4[26748] = 32'b11111111111111111010111100011100;
assign LUT_4[26749] = 32'b11111111111111110100001000010100;
assign LUT_4[26750] = 32'b11111111111111111010010111000000;
assign LUT_4[26751] = 32'b11111111111111110011100010111000;
assign LUT_4[26752] = 32'b00000000000000001001110001101010;
assign LUT_4[26753] = 32'b00000000000000000010111101100010;
assign LUT_4[26754] = 32'b00000000000000001001001100001110;
assign LUT_4[26755] = 32'b00000000000000000010011000000110;
assign LUT_4[26756] = 32'b00000000000000000110110010000110;
assign LUT_4[26757] = 32'b11111111111111111111111101111110;
assign LUT_4[26758] = 32'b00000000000000000110001100101010;
assign LUT_4[26759] = 32'b11111111111111111111011000100010;
assign LUT_4[26760] = 32'b00000000000000000010111101111111;
assign LUT_4[26761] = 32'b11111111111111111100001001110111;
assign LUT_4[26762] = 32'b00000000000000000010011000100011;
assign LUT_4[26763] = 32'b11111111111111111011100100011011;
assign LUT_4[26764] = 32'b11111111111111111111111110011011;
assign LUT_4[26765] = 32'b11111111111111111001001010010011;
assign LUT_4[26766] = 32'b11111111111111111111011000111111;
assign LUT_4[26767] = 32'b11111111111111111000100100110111;
assign LUT_4[26768] = 32'b00000000000000000111100011011000;
assign LUT_4[26769] = 32'b00000000000000000000101111010000;
assign LUT_4[26770] = 32'b00000000000000000110111101111100;
assign LUT_4[26771] = 32'b00000000000000000000001001110100;
assign LUT_4[26772] = 32'b00000000000000000100100011110100;
assign LUT_4[26773] = 32'b11111111111111111101101111101100;
assign LUT_4[26774] = 32'b00000000000000000011111110011000;
assign LUT_4[26775] = 32'b11111111111111111101001010010000;
assign LUT_4[26776] = 32'b00000000000000000000101111101101;
assign LUT_4[26777] = 32'b11111111111111111001111011100101;
assign LUT_4[26778] = 32'b00000000000000000000001010010001;
assign LUT_4[26779] = 32'b11111111111111111001010110001001;
assign LUT_4[26780] = 32'b11111111111111111101110000001001;
assign LUT_4[26781] = 32'b11111111111111110110111100000001;
assign LUT_4[26782] = 32'b11111111111111111101001010101101;
assign LUT_4[26783] = 32'b11111111111111110110010110100101;
assign LUT_4[26784] = 32'b00000000000000001000001100110001;
assign LUT_4[26785] = 32'b00000000000000000001011000101001;
assign LUT_4[26786] = 32'b00000000000000000111100111010101;
assign LUT_4[26787] = 32'b00000000000000000000110011001101;
assign LUT_4[26788] = 32'b00000000000000000101001101001101;
assign LUT_4[26789] = 32'b11111111111111111110011001000101;
assign LUT_4[26790] = 32'b00000000000000000100100111110001;
assign LUT_4[26791] = 32'b11111111111111111101110011101001;
assign LUT_4[26792] = 32'b00000000000000000001011001000110;
assign LUT_4[26793] = 32'b11111111111111111010100100111110;
assign LUT_4[26794] = 32'b00000000000000000000110011101010;
assign LUT_4[26795] = 32'b11111111111111111001111111100010;
assign LUT_4[26796] = 32'b11111111111111111110011001100010;
assign LUT_4[26797] = 32'b11111111111111110111100101011010;
assign LUT_4[26798] = 32'b11111111111111111101110100000110;
assign LUT_4[26799] = 32'b11111111111111110110111111111110;
assign LUT_4[26800] = 32'b00000000000000000101111110011111;
assign LUT_4[26801] = 32'b11111111111111111111001010010111;
assign LUT_4[26802] = 32'b00000000000000000101011001000011;
assign LUT_4[26803] = 32'b11111111111111111110100100111011;
assign LUT_4[26804] = 32'b00000000000000000010111110111011;
assign LUT_4[26805] = 32'b11111111111111111100001010110011;
assign LUT_4[26806] = 32'b00000000000000000010011001011111;
assign LUT_4[26807] = 32'b11111111111111111011100101010111;
assign LUT_4[26808] = 32'b11111111111111111111001010110100;
assign LUT_4[26809] = 32'b11111111111111111000010110101100;
assign LUT_4[26810] = 32'b11111111111111111110100101011000;
assign LUT_4[26811] = 32'b11111111111111110111110001010000;
assign LUT_4[26812] = 32'b11111111111111111100001011010000;
assign LUT_4[26813] = 32'b11111111111111110101010111001000;
assign LUT_4[26814] = 32'b11111111111111111011100101110100;
assign LUT_4[26815] = 32'b11111111111111110100110001101100;
assign LUT_4[26816] = 32'b00000000000000001011001000111110;
assign LUT_4[26817] = 32'b00000000000000000100010100110110;
assign LUT_4[26818] = 32'b00000000000000001010100011100010;
assign LUT_4[26819] = 32'b00000000000000000011101111011010;
assign LUT_4[26820] = 32'b00000000000000001000001001011010;
assign LUT_4[26821] = 32'b00000000000000000001010101010010;
assign LUT_4[26822] = 32'b00000000000000000111100011111110;
assign LUT_4[26823] = 32'b00000000000000000000101111110110;
assign LUT_4[26824] = 32'b00000000000000000100010101010011;
assign LUT_4[26825] = 32'b11111111111111111101100001001011;
assign LUT_4[26826] = 32'b00000000000000000011101111110111;
assign LUT_4[26827] = 32'b11111111111111111100111011101111;
assign LUT_4[26828] = 32'b00000000000000000001010101101111;
assign LUT_4[26829] = 32'b11111111111111111010100001100111;
assign LUT_4[26830] = 32'b00000000000000000000110000010011;
assign LUT_4[26831] = 32'b11111111111111111001111100001011;
assign LUT_4[26832] = 32'b00000000000000001000111010101100;
assign LUT_4[26833] = 32'b00000000000000000010000110100100;
assign LUT_4[26834] = 32'b00000000000000001000010101010000;
assign LUT_4[26835] = 32'b00000000000000000001100001001000;
assign LUT_4[26836] = 32'b00000000000000000101111011001000;
assign LUT_4[26837] = 32'b11111111111111111111000111000000;
assign LUT_4[26838] = 32'b00000000000000000101010101101100;
assign LUT_4[26839] = 32'b11111111111111111110100001100100;
assign LUT_4[26840] = 32'b00000000000000000010000111000001;
assign LUT_4[26841] = 32'b11111111111111111011010010111001;
assign LUT_4[26842] = 32'b00000000000000000001100001100101;
assign LUT_4[26843] = 32'b11111111111111111010101101011101;
assign LUT_4[26844] = 32'b11111111111111111111000111011101;
assign LUT_4[26845] = 32'b11111111111111111000010011010101;
assign LUT_4[26846] = 32'b11111111111111111110100010000001;
assign LUT_4[26847] = 32'b11111111111111110111101101111001;
assign LUT_4[26848] = 32'b00000000000000001001100100000101;
assign LUT_4[26849] = 32'b00000000000000000010101111111101;
assign LUT_4[26850] = 32'b00000000000000001000111110101001;
assign LUT_4[26851] = 32'b00000000000000000010001010100001;
assign LUT_4[26852] = 32'b00000000000000000110100100100001;
assign LUT_4[26853] = 32'b11111111111111111111110000011001;
assign LUT_4[26854] = 32'b00000000000000000101111111000101;
assign LUT_4[26855] = 32'b11111111111111111111001010111101;
assign LUT_4[26856] = 32'b00000000000000000010110000011010;
assign LUT_4[26857] = 32'b11111111111111111011111100010010;
assign LUT_4[26858] = 32'b00000000000000000010001010111110;
assign LUT_4[26859] = 32'b11111111111111111011010110110110;
assign LUT_4[26860] = 32'b11111111111111111111110000110110;
assign LUT_4[26861] = 32'b11111111111111111000111100101110;
assign LUT_4[26862] = 32'b11111111111111111111001011011010;
assign LUT_4[26863] = 32'b11111111111111111000010111010010;
assign LUT_4[26864] = 32'b00000000000000000111010101110011;
assign LUT_4[26865] = 32'b00000000000000000000100001101011;
assign LUT_4[26866] = 32'b00000000000000000110110000010111;
assign LUT_4[26867] = 32'b11111111111111111111111100001111;
assign LUT_4[26868] = 32'b00000000000000000100010110001111;
assign LUT_4[26869] = 32'b11111111111111111101100010000111;
assign LUT_4[26870] = 32'b00000000000000000011110000110011;
assign LUT_4[26871] = 32'b11111111111111111100111100101011;
assign LUT_4[26872] = 32'b00000000000000000000100010001000;
assign LUT_4[26873] = 32'b11111111111111111001101110000000;
assign LUT_4[26874] = 32'b11111111111111111111111100101100;
assign LUT_4[26875] = 32'b11111111111111111001001000100100;
assign LUT_4[26876] = 32'b11111111111111111101100010100100;
assign LUT_4[26877] = 32'b11111111111111110110101110011100;
assign LUT_4[26878] = 32'b11111111111111111100111101001000;
assign LUT_4[26879] = 32'b11111111111111110110001001000000;
assign LUT_4[26880] = 32'b00000000000000001100000111000101;
assign LUT_4[26881] = 32'b00000000000000000101010010111101;
assign LUT_4[26882] = 32'b00000000000000001011100001101001;
assign LUT_4[26883] = 32'b00000000000000000100101101100001;
assign LUT_4[26884] = 32'b00000000000000001001000111100001;
assign LUT_4[26885] = 32'b00000000000000000010010011011001;
assign LUT_4[26886] = 32'b00000000000000001000100010000101;
assign LUT_4[26887] = 32'b00000000000000000001101101111101;
assign LUT_4[26888] = 32'b00000000000000000101010011011010;
assign LUT_4[26889] = 32'b11111111111111111110011111010010;
assign LUT_4[26890] = 32'b00000000000000000100101101111110;
assign LUT_4[26891] = 32'b11111111111111111101111001110110;
assign LUT_4[26892] = 32'b00000000000000000010010011110110;
assign LUT_4[26893] = 32'b11111111111111111011011111101110;
assign LUT_4[26894] = 32'b00000000000000000001101110011010;
assign LUT_4[26895] = 32'b11111111111111111010111010010010;
assign LUT_4[26896] = 32'b00000000000000001001111000110011;
assign LUT_4[26897] = 32'b00000000000000000011000100101011;
assign LUT_4[26898] = 32'b00000000000000001001010011010111;
assign LUT_4[26899] = 32'b00000000000000000010011111001111;
assign LUT_4[26900] = 32'b00000000000000000110111001001111;
assign LUT_4[26901] = 32'b00000000000000000000000101000111;
assign LUT_4[26902] = 32'b00000000000000000110010011110011;
assign LUT_4[26903] = 32'b11111111111111111111011111101011;
assign LUT_4[26904] = 32'b00000000000000000011000101001000;
assign LUT_4[26905] = 32'b11111111111111111100010001000000;
assign LUT_4[26906] = 32'b00000000000000000010011111101100;
assign LUT_4[26907] = 32'b11111111111111111011101011100100;
assign LUT_4[26908] = 32'b00000000000000000000000101100100;
assign LUT_4[26909] = 32'b11111111111111111001010001011100;
assign LUT_4[26910] = 32'b11111111111111111111100000001000;
assign LUT_4[26911] = 32'b11111111111111111000101100000000;
assign LUT_4[26912] = 32'b00000000000000001010100010001100;
assign LUT_4[26913] = 32'b00000000000000000011101110000100;
assign LUT_4[26914] = 32'b00000000000000001001111100110000;
assign LUT_4[26915] = 32'b00000000000000000011001000101000;
assign LUT_4[26916] = 32'b00000000000000000111100010101000;
assign LUT_4[26917] = 32'b00000000000000000000101110100000;
assign LUT_4[26918] = 32'b00000000000000000110111101001100;
assign LUT_4[26919] = 32'b00000000000000000000001001000100;
assign LUT_4[26920] = 32'b00000000000000000011101110100001;
assign LUT_4[26921] = 32'b11111111111111111100111010011001;
assign LUT_4[26922] = 32'b00000000000000000011001001000101;
assign LUT_4[26923] = 32'b11111111111111111100010100111101;
assign LUT_4[26924] = 32'b00000000000000000000101110111101;
assign LUT_4[26925] = 32'b11111111111111111001111010110101;
assign LUT_4[26926] = 32'b00000000000000000000001001100001;
assign LUT_4[26927] = 32'b11111111111111111001010101011001;
assign LUT_4[26928] = 32'b00000000000000001000010011111010;
assign LUT_4[26929] = 32'b00000000000000000001011111110010;
assign LUT_4[26930] = 32'b00000000000000000111101110011110;
assign LUT_4[26931] = 32'b00000000000000000000111010010110;
assign LUT_4[26932] = 32'b00000000000000000101010100010110;
assign LUT_4[26933] = 32'b11111111111111111110100000001110;
assign LUT_4[26934] = 32'b00000000000000000100101110111010;
assign LUT_4[26935] = 32'b11111111111111111101111010110010;
assign LUT_4[26936] = 32'b00000000000000000001100000001111;
assign LUT_4[26937] = 32'b11111111111111111010101100000111;
assign LUT_4[26938] = 32'b00000000000000000000111010110011;
assign LUT_4[26939] = 32'b11111111111111111010000110101011;
assign LUT_4[26940] = 32'b11111111111111111110100000101011;
assign LUT_4[26941] = 32'b11111111111111110111101100100011;
assign LUT_4[26942] = 32'b11111111111111111101111011001111;
assign LUT_4[26943] = 32'b11111111111111110111000111000111;
assign LUT_4[26944] = 32'b00000000000000001101011110011001;
assign LUT_4[26945] = 32'b00000000000000000110101010010001;
assign LUT_4[26946] = 32'b00000000000000001100111000111101;
assign LUT_4[26947] = 32'b00000000000000000110000100110101;
assign LUT_4[26948] = 32'b00000000000000001010011110110101;
assign LUT_4[26949] = 32'b00000000000000000011101010101101;
assign LUT_4[26950] = 32'b00000000000000001001111001011001;
assign LUT_4[26951] = 32'b00000000000000000011000101010001;
assign LUT_4[26952] = 32'b00000000000000000110101010101110;
assign LUT_4[26953] = 32'b11111111111111111111110110100110;
assign LUT_4[26954] = 32'b00000000000000000110000101010010;
assign LUT_4[26955] = 32'b11111111111111111111010001001010;
assign LUT_4[26956] = 32'b00000000000000000011101011001010;
assign LUT_4[26957] = 32'b11111111111111111100110111000010;
assign LUT_4[26958] = 32'b00000000000000000011000101101110;
assign LUT_4[26959] = 32'b11111111111111111100010001100110;
assign LUT_4[26960] = 32'b00000000000000001011010000000111;
assign LUT_4[26961] = 32'b00000000000000000100011011111111;
assign LUT_4[26962] = 32'b00000000000000001010101010101011;
assign LUT_4[26963] = 32'b00000000000000000011110110100011;
assign LUT_4[26964] = 32'b00000000000000001000010000100011;
assign LUT_4[26965] = 32'b00000000000000000001011100011011;
assign LUT_4[26966] = 32'b00000000000000000111101011000111;
assign LUT_4[26967] = 32'b00000000000000000000110110111111;
assign LUT_4[26968] = 32'b00000000000000000100011100011100;
assign LUT_4[26969] = 32'b11111111111111111101101000010100;
assign LUT_4[26970] = 32'b00000000000000000011110111000000;
assign LUT_4[26971] = 32'b11111111111111111101000010111000;
assign LUT_4[26972] = 32'b00000000000000000001011100111000;
assign LUT_4[26973] = 32'b11111111111111111010101000110000;
assign LUT_4[26974] = 32'b00000000000000000000110111011100;
assign LUT_4[26975] = 32'b11111111111111111010000011010100;
assign LUT_4[26976] = 32'b00000000000000001011111001100000;
assign LUT_4[26977] = 32'b00000000000000000101000101011000;
assign LUT_4[26978] = 32'b00000000000000001011010100000100;
assign LUT_4[26979] = 32'b00000000000000000100011111111100;
assign LUT_4[26980] = 32'b00000000000000001000111001111100;
assign LUT_4[26981] = 32'b00000000000000000010000101110100;
assign LUT_4[26982] = 32'b00000000000000001000010100100000;
assign LUT_4[26983] = 32'b00000000000000000001100000011000;
assign LUT_4[26984] = 32'b00000000000000000101000101110101;
assign LUT_4[26985] = 32'b11111111111111111110010001101101;
assign LUT_4[26986] = 32'b00000000000000000100100000011001;
assign LUT_4[26987] = 32'b11111111111111111101101100010001;
assign LUT_4[26988] = 32'b00000000000000000010000110010001;
assign LUT_4[26989] = 32'b11111111111111111011010010001001;
assign LUT_4[26990] = 32'b00000000000000000001100000110101;
assign LUT_4[26991] = 32'b11111111111111111010101100101101;
assign LUT_4[26992] = 32'b00000000000000001001101011001110;
assign LUT_4[26993] = 32'b00000000000000000010110111000110;
assign LUT_4[26994] = 32'b00000000000000001001000101110010;
assign LUT_4[26995] = 32'b00000000000000000010010001101010;
assign LUT_4[26996] = 32'b00000000000000000110101011101010;
assign LUT_4[26997] = 32'b11111111111111111111110111100010;
assign LUT_4[26998] = 32'b00000000000000000110000110001110;
assign LUT_4[26999] = 32'b11111111111111111111010010000110;
assign LUT_4[27000] = 32'b00000000000000000010110111100011;
assign LUT_4[27001] = 32'b11111111111111111100000011011011;
assign LUT_4[27002] = 32'b00000000000000000010010010000111;
assign LUT_4[27003] = 32'b11111111111111111011011101111111;
assign LUT_4[27004] = 32'b11111111111111111111110111111111;
assign LUT_4[27005] = 32'b11111111111111111001000011110111;
assign LUT_4[27006] = 32'b11111111111111111111010010100011;
assign LUT_4[27007] = 32'b11111111111111111000011110011011;
assign LUT_4[27008] = 32'b00000000000000001110101101001101;
assign LUT_4[27009] = 32'b00000000000000000111111001000101;
assign LUT_4[27010] = 32'b00000000000000001110000111110001;
assign LUT_4[27011] = 32'b00000000000000000111010011101001;
assign LUT_4[27012] = 32'b00000000000000001011101101101001;
assign LUT_4[27013] = 32'b00000000000000000100111001100001;
assign LUT_4[27014] = 32'b00000000000000001011001000001101;
assign LUT_4[27015] = 32'b00000000000000000100010100000101;
assign LUT_4[27016] = 32'b00000000000000000111111001100010;
assign LUT_4[27017] = 32'b00000000000000000001000101011010;
assign LUT_4[27018] = 32'b00000000000000000111010100000110;
assign LUT_4[27019] = 32'b00000000000000000000011111111110;
assign LUT_4[27020] = 32'b00000000000000000100111001111110;
assign LUT_4[27021] = 32'b11111111111111111110000101110110;
assign LUT_4[27022] = 32'b00000000000000000100010100100010;
assign LUT_4[27023] = 32'b11111111111111111101100000011010;
assign LUT_4[27024] = 32'b00000000000000001100011110111011;
assign LUT_4[27025] = 32'b00000000000000000101101010110011;
assign LUT_4[27026] = 32'b00000000000000001011111001011111;
assign LUT_4[27027] = 32'b00000000000000000101000101010111;
assign LUT_4[27028] = 32'b00000000000000001001011111010111;
assign LUT_4[27029] = 32'b00000000000000000010101011001111;
assign LUT_4[27030] = 32'b00000000000000001000111001111011;
assign LUT_4[27031] = 32'b00000000000000000010000101110011;
assign LUT_4[27032] = 32'b00000000000000000101101011010000;
assign LUT_4[27033] = 32'b11111111111111111110110111001000;
assign LUT_4[27034] = 32'b00000000000000000101000101110100;
assign LUT_4[27035] = 32'b11111111111111111110010001101100;
assign LUT_4[27036] = 32'b00000000000000000010101011101100;
assign LUT_4[27037] = 32'b11111111111111111011110111100100;
assign LUT_4[27038] = 32'b00000000000000000010000110010000;
assign LUT_4[27039] = 32'b11111111111111111011010010001000;
assign LUT_4[27040] = 32'b00000000000000001101001000010100;
assign LUT_4[27041] = 32'b00000000000000000110010100001100;
assign LUT_4[27042] = 32'b00000000000000001100100010111000;
assign LUT_4[27043] = 32'b00000000000000000101101110110000;
assign LUT_4[27044] = 32'b00000000000000001010001000110000;
assign LUT_4[27045] = 32'b00000000000000000011010100101000;
assign LUT_4[27046] = 32'b00000000000000001001100011010100;
assign LUT_4[27047] = 32'b00000000000000000010101111001100;
assign LUT_4[27048] = 32'b00000000000000000110010100101001;
assign LUT_4[27049] = 32'b11111111111111111111100000100001;
assign LUT_4[27050] = 32'b00000000000000000101101111001101;
assign LUT_4[27051] = 32'b11111111111111111110111011000101;
assign LUT_4[27052] = 32'b00000000000000000011010101000101;
assign LUT_4[27053] = 32'b11111111111111111100100000111101;
assign LUT_4[27054] = 32'b00000000000000000010101111101001;
assign LUT_4[27055] = 32'b11111111111111111011111011100001;
assign LUT_4[27056] = 32'b00000000000000001010111010000010;
assign LUT_4[27057] = 32'b00000000000000000100000101111010;
assign LUT_4[27058] = 32'b00000000000000001010010100100110;
assign LUT_4[27059] = 32'b00000000000000000011100000011110;
assign LUT_4[27060] = 32'b00000000000000000111111010011110;
assign LUT_4[27061] = 32'b00000000000000000001000110010110;
assign LUT_4[27062] = 32'b00000000000000000111010101000010;
assign LUT_4[27063] = 32'b00000000000000000000100000111010;
assign LUT_4[27064] = 32'b00000000000000000100000110010111;
assign LUT_4[27065] = 32'b11111111111111111101010010001111;
assign LUT_4[27066] = 32'b00000000000000000011100000111011;
assign LUT_4[27067] = 32'b11111111111111111100101100110011;
assign LUT_4[27068] = 32'b00000000000000000001000110110011;
assign LUT_4[27069] = 32'b11111111111111111010010010101011;
assign LUT_4[27070] = 32'b00000000000000000000100001010111;
assign LUT_4[27071] = 32'b11111111111111111001101101001111;
assign LUT_4[27072] = 32'b00000000000000010000000100100001;
assign LUT_4[27073] = 32'b00000000000000001001010000011001;
assign LUT_4[27074] = 32'b00000000000000001111011111000101;
assign LUT_4[27075] = 32'b00000000000000001000101010111101;
assign LUT_4[27076] = 32'b00000000000000001101000100111101;
assign LUT_4[27077] = 32'b00000000000000000110010000110101;
assign LUT_4[27078] = 32'b00000000000000001100011111100001;
assign LUT_4[27079] = 32'b00000000000000000101101011011001;
assign LUT_4[27080] = 32'b00000000000000001001010000110110;
assign LUT_4[27081] = 32'b00000000000000000010011100101110;
assign LUT_4[27082] = 32'b00000000000000001000101011011010;
assign LUT_4[27083] = 32'b00000000000000000001110111010010;
assign LUT_4[27084] = 32'b00000000000000000110010001010010;
assign LUT_4[27085] = 32'b11111111111111111111011101001010;
assign LUT_4[27086] = 32'b00000000000000000101101011110110;
assign LUT_4[27087] = 32'b11111111111111111110110111101110;
assign LUT_4[27088] = 32'b00000000000000001101110110001111;
assign LUT_4[27089] = 32'b00000000000000000111000010000111;
assign LUT_4[27090] = 32'b00000000000000001101010000110011;
assign LUT_4[27091] = 32'b00000000000000000110011100101011;
assign LUT_4[27092] = 32'b00000000000000001010110110101011;
assign LUT_4[27093] = 32'b00000000000000000100000010100011;
assign LUT_4[27094] = 32'b00000000000000001010010001001111;
assign LUT_4[27095] = 32'b00000000000000000011011101000111;
assign LUT_4[27096] = 32'b00000000000000000111000010100100;
assign LUT_4[27097] = 32'b00000000000000000000001110011100;
assign LUT_4[27098] = 32'b00000000000000000110011101001000;
assign LUT_4[27099] = 32'b11111111111111111111101001000000;
assign LUT_4[27100] = 32'b00000000000000000100000011000000;
assign LUT_4[27101] = 32'b11111111111111111101001110111000;
assign LUT_4[27102] = 32'b00000000000000000011011101100100;
assign LUT_4[27103] = 32'b11111111111111111100101001011100;
assign LUT_4[27104] = 32'b00000000000000001110011111101000;
assign LUT_4[27105] = 32'b00000000000000000111101011100000;
assign LUT_4[27106] = 32'b00000000000000001101111010001100;
assign LUT_4[27107] = 32'b00000000000000000111000110000100;
assign LUT_4[27108] = 32'b00000000000000001011100000000100;
assign LUT_4[27109] = 32'b00000000000000000100101011111100;
assign LUT_4[27110] = 32'b00000000000000001010111010101000;
assign LUT_4[27111] = 32'b00000000000000000100000110100000;
assign LUT_4[27112] = 32'b00000000000000000111101011111101;
assign LUT_4[27113] = 32'b00000000000000000000110111110101;
assign LUT_4[27114] = 32'b00000000000000000111000110100001;
assign LUT_4[27115] = 32'b00000000000000000000010010011001;
assign LUT_4[27116] = 32'b00000000000000000100101100011001;
assign LUT_4[27117] = 32'b11111111111111111101111000010001;
assign LUT_4[27118] = 32'b00000000000000000100000110111101;
assign LUT_4[27119] = 32'b11111111111111111101010010110101;
assign LUT_4[27120] = 32'b00000000000000001100010001010110;
assign LUT_4[27121] = 32'b00000000000000000101011101001110;
assign LUT_4[27122] = 32'b00000000000000001011101011111010;
assign LUT_4[27123] = 32'b00000000000000000100110111110010;
assign LUT_4[27124] = 32'b00000000000000001001010001110010;
assign LUT_4[27125] = 32'b00000000000000000010011101101010;
assign LUT_4[27126] = 32'b00000000000000001000101100010110;
assign LUT_4[27127] = 32'b00000000000000000001111000001110;
assign LUT_4[27128] = 32'b00000000000000000101011101101011;
assign LUT_4[27129] = 32'b11111111111111111110101001100011;
assign LUT_4[27130] = 32'b00000000000000000100111000001111;
assign LUT_4[27131] = 32'b11111111111111111110000100000111;
assign LUT_4[27132] = 32'b00000000000000000010011110000111;
assign LUT_4[27133] = 32'b11111111111111111011101001111111;
assign LUT_4[27134] = 32'b00000000000000000001111000101011;
assign LUT_4[27135] = 32'b11111111111111111011000100100011;
assign LUT_4[27136] = 32'b00000000000000000110001111101010;
assign LUT_4[27137] = 32'b11111111111111111111011011100010;
assign LUT_4[27138] = 32'b00000000000000000101101010001110;
assign LUT_4[27139] = 32'b11111111111111111110110110000110;
assign LUT_4[27140] = 32'b00000000000000000011010000000110;
assign LUT_4[27141] = 32'b11111111111111111100011011111110;
assign LUT_4[27142] = 32'b00000000000000000010101010101010;
assign LUT_4[27143] = 32'b11111111111111111011110110100010;
assign LUT_4[27144] = 32'b11111111111111111111011011111111;
assign LUT_4[27145] = 32'b11111111111111111000100111110111;
assign LUT_4[27146] = 32'b11111111111111111110110110100011;
assign LUT_4[27147] = 32'b11111111111111111000000010011011;
assign LUT_4[27148] = 32'b11111111111111111100011100011011;
assign LUT_4[27149] = 32'b11111111111111110101101000010011;
assign LUT_4[27150] = 32'b11111111111111111011110110111111;
assign LUT_4[27151] = 32'b11111111111111110101000010110111;
assign LUT_4[27152] = 32'b00000000000000000100000001011000;
assign LUT_4[27153] = 32'b11111111111111111101001101010000;
assign LUT_4[27154] = 32'b00000000000000000011011011111100;
assign LUT_4[27155] = 32'b11111111111111111100100111110100;
assign LUT_4[27156] = 32'b00000000000000000001000001110100;
assign LUT_4[27157] = 32'b11111111111111111010001101101100;
assign LUT_4[27158] = 32'b00000000000000000000011100011000;
assign LUT_4[27159] = 32'b11111111111111111001101000010000;
assign LUT_4[27160] = 32'b11111111111111111101001101101101;
assign LUT_4[27161] = 32'b11111111111111110110011001100101;
assign LUT_4[27162] = 32'b11111111111111111100101000010001;
assign LUT_4[27163] = 32'b11111111111111110101110100001001;
assign LUT_4[27164] = 32'b11111111111111111010001110001001;
assign LUT_4[27165] = 32'b11111111111111110011011010000001;
assign LUT_4[27166] = 32'b11111111111111111001101000101101;
assign LUT_4[27167] = 32'b11111111111111110010110100100101;
assign LUT_4[27168] = 32'b00000000000000000100101010110001;
assign LUT_4[27169] = 32'b11111111111111111101110110101001;
assign LUT_4[27170] = 32'b00000000000000000100000101010101;
assign LUT_4[27171] = 32'b11111111111111111101010001001101;
assign LUT_4[27172] = 32'b00000000000000000001101011001101;
assign LUT_4[27173] = 32'b11111111111111111010110111000101;
assign LUT_4[27174] = 32'b00000000000000000001000101110001;
assign LUT_4[27175] = 32'b11111111111111111010010001101001;
assign LUT_4[27176] = 32'b11111111111111111101110111000110;
assign LUT_4[27177] = 32'b11111111111111110111000010111110;
assign LUT_4[27178] = 32'b11111111111111111101010001101010;
assign LUT_4[27179] = 32'b11111111111111110110011101100010;
assign LUT_4[27180] = 32'b11111111111111111010110111100010;
assign LUT_4[27181] = 32'b11111111111111110100000011011010;
assign LUT_4[27182] = 32'b11111111111111111010010010000110;
assign LUT_4[27183] = 32'b11111111111111110011011101111110;
assign LUT_4[27184] = 32'b00000000000000000010011100011111;
assign LUT_4[27185] = 32'b11111111111111111011101000010111;
assign LUT_4[27186] = 32'b00000000000000000001110111000011;
assign LUT_4[27187] = 32'b11111111111111111011000010111011;
assign LUT_4[27188] = 32'b11111111111111111111011100111011;
assign LUT_4[27189] = 32'b11111111111111111000101000110011;
assign LUT_4[27190] = 32'b11111111111111111110110111011111;
assign LUT_4[27191] = 32'b11111111111111111000000011010111;
assign LUT_4[27192] = 32'b11111111111111111011101000110100;
assign LUT_4[27193] = 32'b11111111111111110100110100101100;
assign LUT_4[27194] = 32'b11111111111111111011000011011000;
assign LUT_4[27195] = 32'b11111111111111110100001111010000;
assign LUT_4[27196] = 32'b11111111111111111000101001010000;
assign LUT_4[27197] = 32'b11111111111111110001110101001000;
assign LUT_4[27198] = 32'b11111111111111111000000011110100;
assign LUT_4[27199] = 32'b11111111111111110001001111101100;
assign LUT_4[27200] = 32'b00000000000000000111100110111110;
assign LUT_4[27201] = 32'b00000000000000000000110010110110;
assign LUT_4[27202] = 32'b00000000000000000111000001100010;
assign LUT_4[27203] = 32'b00000000000000000000001101011010;
assign LUT_4[27204] = 32'b00000000000000000100100111011010;
assign LUT_4[27205] = 32'b11111111111111111101110011010010;
assign LUT_4[27206] = 32'b00000000000000000100000001111110;
assign LUT_4[27207] = 32'b11111111111111111101001101110110;
assign LUT_4[27208] = 32'b00000000000000000000110011010011;
assign LUT_4[27209] = 32'b11111111111111111001111111001011;
assign LUT_4[27210] = 32'b00000000000000000000001101110111;
assign LUT_4[27211] = 32'b11111111111111111001011001101111;
assign LUT_4[27212] = 32'b11111111111111111101110011101111;
assign LUT_4[27213] = 32'b11111111111111110110111111100111;
assign LUT_4[27214] = 32'b11111111111111111101001110010011;
assign LUT_4[27215] = 32'b11111111111111110110011010001011;
assign LUT_4[27216] = 32'b00000000000000000101011000101100;
assign LUT_4[27217] = 32'b11111111111111111110100100100100;
assign LUT_4[27218] = 32'b00000000000000000100110011010000;
assign LUT_4[27219] = 32'b11111111111111111101111111001000;
assign LUT_4[27220] = 32'b00000000000000000010011001001000;
assign LUT_4[27221] = 32'b11111111111111111011100101000000;
assign LUT_4[27222] = 32'b00000000000000000001110011101100;
assign LUT_4[27223] = 32'b11111111111111111010111111100100;
assign LUT_4[27224] = 32'b11111111111111111110100101000001;
assign LUT_4[27225] = 32'b11111111111111110111110000111001;
assign LUT_4[27226] = 32'b11111111111111111101111111100101;
assign LUT_4[27227] = 32'b11111111111111110111001011011101;
assign LUT_4[27228] = 32'b11111111111111111011100101011101;
assign LUT_4[27229] = 32'b11111111111111110100110001010101;
assign LUT_4[27230] = 32'b11111111111111111011000000000001;
assign LUT_4[27231] = 32'b11111111111111110100001011111001;
assign LUT_4[27232] = 32'b00000000000000000110000010000101;
assign LUT_4[27233] = 32'b11111111111111111111001101111101;
assign LUT_4[27234] = 32'b00000000000000000101011100101001;
assign LUT_4[27235] = 32'b11111111111111111110101000100001;
assign LUT_4[27236] = 32'b00000000000000000011000010100001;
assign LUT_4[27237] = 32'b11111111111111111100001110011001;
assign LUT_4[27238] = 32'b00000000000000000010011101000101;
assign LUT_4[27239] = 32'b11111111111111111011101000111101;
assign LUT_4[27240] = 32'b11111111111111111111001110011010;
assign LUT_4[27241] = 32'b11111111111111111000011010010010;
assign LUT_4[27242] = 32'b11111111111111111110101000111110;
assign LUT_4[27243] = 32'b11111111111111110111110100110110;
assign LUT_4[27244] = 32'b11111111111111111100001110110110;
assign LUT_4[27245] = 32'b11111111111111110101011010101110;
assign LUT_4[27246] = 32'b11111111111111111011101001011010;
assign LUT_4[27247] = 32'b11111111111111110100110101010010;
assign LUT_4[27248] = 32'b00000000000000000011110011110011;
assign LUT_4[27249] = 32'b11111111111111111100111111101011;
assign LUT_4[27250] = 32'b00000000000000000011001110010111;
assign LUT_4[27251] = 32'b11111111111111111100011010001111;
assign LUT_4[27252] = 32'b00000000000000000000110100001111;
assign LUT_4[27253] = 32'b11111111111111111010000000000111;
assign LUT_4[27254] = 32'b00000000000000000000001110110011;
assign LUT_4[27255] = 32'b11111111111111111001011010101011;
assign LUT_4[27256] = 32'b11111111111111111101000000001000;
assign LUT_4[27257] = 32'b11111111111111110110001100000000;
assign LUT_4[27258] = 32'b11111111111111111100011010101100;
assign LUT_4[27259] = 32'b11111111111111110101100110100100;
assign LUT_4[27260] = 32'b11111111111111111010000000100100;
assign LUT_4[27261] = 32'b11111111111111110011001100011100;
assign LUT_4[27262] = 32'b11111111111111111001011011001000;
assign LUT_4[27263] = 32'b11111111111111110010100111000000;
assign LUT_4[27264] = 32'b00000000000000001000110101110010;
assign LUT_4[27265] = 32'b00000000000000000010000001101010;
assign LUT_4[27266] = 32'b00000000000000001000010000010110;
assign LUT_4[27267] = 32'b00000000000000000001011100001110;
assign LUT_4[27268] = 32'b00000000000000000101110110001110;
assign LUT_4[27269] = 32'b11111111111111111111000010000110;
assign LUT_4[27270] = 32'b00000000000000000101010000110010;
assign LUT_4[27271] = 32'b11111111111111111110011100101010;
assign LUT_4[27272] = 32'b00000000000000000010000010000111;
assign LUT_4[27273] = 32'b11111111111111111011001101111111;
assign LUT_4[27274] = 32'b00000000000000000001011100101011;
assign LUT_4[27275] = 32'b11111111111111111010101000100011;
assign LUT_4[27276] = 32'b11111111111111111111000010100011;
assign LUT_4[27277] = 32'b11111111111111111000001110011011;
assign LUT_4[27278] = 32'b11111111111111111110011101000111;
assign LUT_4[27279] = 32'b11111111111111110111101000111111;
assign LUT_4[27280] = 32'b00000000000000000110100111100000;
assign LUT_4[27281] = 32'b11111111111111111111110011011000;
assign LUT_4[27282] = 32'b00000000000000000110000010000100;
assign LUT_4[27283] = 32'b11111111111111111111001101111100;
assign LUT_4[27284] = 32'b00000000000000000011100111111100;
assign LUT_4[27285] = 32'b11111111111111111100110011110100;
assign LUT_4[27286] = 32'b00000000000000000011000010100000;
assign LUT_4[27287] = 32'b11111111111111111100001110011000;
assign LUT_4[27288] = 32'b11111111111111111111110011110101;
assign LUT_4[27289] = 32'b11111111111111111000111111101101;
assign LUT_4[27290] = 32'b11111111111111111111001110011001;
assign LUT_4[27291] = 32'b11111111111111111000011010010001;
assign LUT_4[27292] = 32'b11111111111111111100110100010001;
assign LUT_4[27293] = 32'b11111111111111110110000000001001;
assign LUT_4[27294] = 32'b11111111111111111100001110110101;
assign LUT_4[27295] = 32'b11111111111111110101011010101101;
assign LUT_4[27296] = 32'b00000000000000000111010000111001;
assign LUT_4[27297] = 32'b00000000000000000000011100110001;
assign LUT_4[27298] = 32'b00000000000000000110101011011101;
assign LUT_4[27299] = 32'b11111111111111111111110111010101;
assign LUT_4[27300] = 32'b00000000000000000100010001010101;
assign LUT_4[27301] = 32'b11111111111111111101011101001101;
assign LUT_4[27302] = 32'b00000000000000000011101011111001;
assign LUT_4[27303] = 32'b11111111111111111100110111110001;
assign LUT_4[27304] = 32'b00000000000000000000011101001110;
assign LUT_4[27305] = 32'b11111111111111111001101001000110;
assign LUT_4[27306] = 32'b11111111111111111111110111110010;
assign LUT_4[27307] = 32'b11111111111111111001000011101010;
assign LUT_4[27308] = 32'b11111111111111111101011101101010;
assign LUT_4[27309] = 32'b11111111111111110110101001100010;
assign LUT_4[27310] = 32'b11111111111111111100111000001110;
assign LUT_4[27311] = 32'b11111111111111110110000100000110;
assign LUT_4[27312] = 32'b00000000000000000101000010100111;
assign LUT_4[27313] = 32'b11111111111111111110001110011111;
assign LUT_4[27314] = 32'b00000000000000000100011101001011;
assign LUT_4[27315] = 32'b11111111111111111101101001000011;
assign LUT_4[27316] = 32'b00000000000000000010000011000011;
assign LUT_4[27317] = 32'b11111111111111111011001110111011;
assign LUT_4[27318] = 32'b00000000000000000001011101100111;
assign LUT_4[27319] = 32'b11111111111111111010101001011111;
assign LUT_4[27320] = 32'b11111111111111111110001110111100;
assign LUT_4[27321] = 32'b11111111111111110111011010110100;
assign LUT_4[27322] = 32'b11111111111111111101101001100000;
assign LUT_4[27323] = 32'b11111111111111110110110101011000;
assign LUT_4[27324] = 32'b11111111111111111011001111011000;
assign LUT_4[27325] = 32'b11111111111111110100011011010000;
assign LUT_4[27326] = 32'b11111111111111111010101001111100;
assign LUT_4[27327] = 32'b11111111111111110011110101110100;
assign LUT_4[27328] = 32'b00000000000000001010001101000110;
assign LUT_4[27329] = 32'b00000000000000000011011000111110;
assign LUT_4[27330] = 32'b00000000000000001001100111101010;
assign LUT_4[27331] = 32'b00000000000000000010110011100010;
assign LUT_4[27332] = 32'b00000000000000000111001101100010;
assign LUT_4[27333] = 32'b00000000000000000000011001011010;
assign LUT_4[27334] = 32'b00000000000000000110101000000110;
assign LUT_4[27335] = 32'b11111111111111111111110011111110;
assign LUT_4[27336] = 32'b00000000000000000011011001011011;
assign LUT_4[27337] = 32'b11111111111111111100100101010011;
assign LUT_4[27338] = 32'b00000000000000000010110011111111;
assign LUT_4[27339] = 32'b11111111111111111011111111110111;
assign LUT_4[27340] = 32'b00000000000000000000011001110111;
assign LUT_4[27341] = 32'b11111111111111111001100101101111;
assign LUT_4[27342] = 32'b11111111111111111111110100011011;
assign LUT_4[27343] = 32'b11111111111111111001000000010011;
assign LUT_4[27344] = 32'b00000000000000000111111110110100;
assign LUT_4[27345] = 32'b00000000000000000001001010101100;
assign LUT_4[27346] = 32'b00000000000000000111011001011000;
assign LUT_4[27347] = 32'b00000000000000000000100101010000;
assign LUT_4[27348] = 32'b00000000000000000100111111010000;
assign LUT_4[27349] = 32'b11111111111111111110001011001000;
assign LUT_4[27350] = 32'b00000000000000000100011001110100;
assign LUT_4[27351] = 32'b11111111111111111101100101101100;
assign LUT_4[27352] = 32'b00000000000000000001001011001001;
assign LUT_4[27353] = 32'b11111111111111111010010111000001;
assign LUT_4[27354] = 32'b00000000000000000000100101101101;
assign LUT_4[27355] = 32'b11111111111111111001110001100101;
assign LUT_4[27356] = 32'b11111111111111111110001011100101;
assign LUT_4[27357] = 32'b11111111111111110111010111011101;
assign LUT_4[27358] = 32'b11111111111111111101100110001001;
assign LUT_4[27359] = 32'b11111111111111110110110010000001;
assign LUT_4[27360] = 32'b00000000000000001000101000001101;
assign LUT_4[27361] = 32'b00000000000000000001110100000101;
assign LUT_4[27362] = 32'b00000000000000001000000010110001;
assign LUT_4[27363] = 32'b00000000000000000001001110101001;
assign LUT_4[27364] = 32'b00000000000000000101101000101001;
assign LUT_4[27365] = 32'b11111111111111111110110100100001;
assign LUT_4[27366] = 32'b00000000000000000101000011001101;
assign LUT_4[27367] = 32'b11111111111111111110001111000101;
assign LUT_4[27368] = 32'b00000000000000000001110100100010;
assign LUT_4[27369] = 32'b11111111111111111011000000011010;
assign LUT_4[27370] = 32'b00000000000000000001001111000110;
assign LUT_4[27371] = 32'b11111111111111111010011010111110;
assign LUT_4[27372] = 32'b11111111111111111110110100111110;
assign LUT_4[27373] = 32'b11111111111111111000000000110110;
assign LUT_4[27374] = 32'b11111111111111111110001111100010;
assign LUT_4[27375] = 32'b11111111111111110111011011011010;
assign LUT_4[27376] = 32'b00000000000000000110011001111011;
assign LUT_4[27377] = 32'b11111111111111111111100101110011;
assign LUT_4[27378] = 32'b00000000000000000101110100011111;
assign LUT_4[27379] = 32'b11111111111111111111000000010111;
assign LUT_4[27380] = 32'b00000000000000000011011010010111;
assign LUT_4[27381] = 32'b11111111111111111100100110001111;
assign LUT_4[27382] = 32'b00000000000000000010110100111011;
assign LUT_4[27383] = 32'b11111111111111111100000000110011;
assign LUT_4[27384] = 32'b11111111111111111111100110010000;
assign LUT_4[27385] = 32'b11111111111111111000110010001000;
assign LUT_4[27386] = 32'b11111111111111111111000000110100;
assign LUT_4[27387] = 32'b11111111111111111000001100101100;
assign LUT_4[27388] = 32'b11111111111111111100100110101100;
assign LUT_4[27389] = 32'b11111111111111110101110010100100;
assign LUT_4[27390] = 32'b11111111111111111100000001010000;
assign LUT_4[27391] = 32'b11111111111111110101001101001000;
assign LUT_4[27392] = 32'b00000000000000001011001011001101;
assign LUT_4[27393] = 32'b00000000000000000100010111000101;
assign LUT_4[27394] = 32'b00000000000000001010100101110001;
assign LUT_4[27395] = 32'b00000000000000000011110001101001;
assign LUT_4[27396] = 32'b00000000000000001000001011101001;
assign LUT_4[27397] = 32'b00000000000000000001010111100001;
assign LUT_4[27398] = 32'b00000000000000000111100110001101;
assign LUT_4[27399] = 32'b00000000000000000000110010000101;
assign LUT_4[27400] = 32'b00000000000000000100010111100010;
assign LUT_4[27401] = 32'b11111111111111111101100011011010;
assign LUT_4[27402] = 32'b00000000000000000011110010000110;
assign LUT_4[27403] = 32'b11111111111111111100111101111110;
assign LUT_4[27404] = 32'b00000000000000000001010111111110;
assign LUT_4[27405] = 32'b11111111111111111010100011110110;
assign LUT_4[27406] = 32'b00000000000000000000110010100010;
assign LUT_4[27407] = 32'b11111111111111111001111110011010;
assign LUT_4[27408] = 32'b00000000000000001000111100111011;
assign LUT_4[27409] = 32'b00000000000000000010001000110011;
assign LUT_4[27410] = 32'b00000000000000001000010111011111;
assign LUT_4[27411] = 32'b00000000000000000001100011010111;
assign LUT_4[27412] = 32'b00000000000000000101111101010111;
assign LUT_4[27413] = 32'b11111111111111111111001001001111;
assign LUT_4[27414] = 32'b00000000000000000101010111111011;
assign LUT_4[27415] = 32'b11111111111111111110100011110011;
assign LUT_4[27416] = 32'b00000000000000000010001001010000;
assign LUT_4[27417] = 32'b11111111111111111011010101001000;
assign LUT_4[27418] = 32'b00000000000000000001100011110100;
assign LUT_4[27419] = 32'b11111111111111111010101111101100;
assign LUT_4[27420] = 32'b11111111111111111111001001101100;
assign LUT_4[27421] = 32'b11111111111111111000010101100100;
assign LUT_4[27422] = 32'b11111111111111111110100100010000;
assign LUT_4[27423] = 32'b11111111111111110111110000001000;
assign LUT_4[27424] = 32'b00000000000000001001100110010100;
assign LUT_4[27425] = 32'b00000000000000000010110010001100;
assign LUT_4[27426] = 32'b00000000000000001001000000111000;
assign LUT_4[27427] = 32'b00000000000000000010001100110000;
assign LUT_4[27428] = 32'b00000000000000000110100110110000;
assign LUT_4[27429] = 32'b11111111111111111111110010101000;
assign LUT_4[27430] = 32'b00000000000000000110000001010100;
assign LUT_4[27431] = 32'b11111111111111111111001101001100;
assign LUT_4[27432] = 32'b00000000000000000010110010101001;
assign LUT_4[27433] = 32'b11111111111111111011111110100001;
assign LUT_4[27434] = 32'b00000000000000000010001101001101;
assign LUT_4[27435] = 32'b11111111111111111011011001000101;
assign LUT_4[27436] = 32'b11111111111111111111110011000101;
assign LUT_4[27437] = 32'b11111111111111111000111110111101;
assign LUT_4[27438] = 32'b11111111111111111111001101101001;
assign LUT_4[27439] = 32'b11111111111111111000011001100001;
assign LUT_4[27440] = 32'b00000000000000000111011000000010;
assign LUT_4[27441] = 32'b00000000000000000000100011111010;
assign LUT_4[27442] = 32'b00000000000000000110110010100110;
assign LUT_4[27443] = 32'b11111111111111111111111110011110;
assign LUT_4[27444] = 32'b00000000000000000100011000011110;
assign LUT_4[27445] = 32'b11111111111111111101100100010110;
assign LUT_4[27446] = 32'b00000000000000000011110011000010;
assign LUT_4[27447] = 32'b11111111111111111100111110111010;
assign LUT_4[27448] = 32'b00000000000000000000100100010111;
assign LUT_4[27449] = 32'b11111111111111111001110000001111;
assign LUT_4[27450] = 32'b11111111111111111111111110111011;
assign LUT_4[27451] = 32'b11111111111111111001001010110011;
assign LUT_4[27452] = 32'b11111111111111111101100100110011;
assign LUT_4[27453] = 32'b11111111111111110110110000101011;
assign LUT_4[27454] = 32'b11111111111111111100111111010111;
assign LUT_4[27455] = 32'b11111111111111110110001011001111;
assign LUT_4[27456] = 32'b00000000000000001100100010100001;
assign LUT_4[27457] = 32'b00000000000000000101101110011001;
assign LUT_4[27458] = 32'b00000000000000001011111101000101;
assign LUT_4[27459] = 32'b00000000000000000101001000111101;
assign LUT_4[27460] = 32'b00000000000000001001100010111101;
assign LUT_4[27461] = 32'b00000000000000000010101110110101;
assign LUT_4[27462] = 32'b00000000000000001000111101100001;
assign LUT_4[27463] = 32'b00000000000000000010001001011001;
assign LUT_4[27464] = 32'b00000000000000000101101110110110;
assign LUT_4[27465] = 32'b11111111111111111110111010101110;
assign LUT_4[27466] = 32'b00000000000000000101001001011010;
assign LUT_4[27467] = 32'b11111111111111111110010101010010;
assign LUT_4[27468] = 32'b00000000000000000010101111010010;
assign LUT_4[27469] = 32'b11111111111111111011111011001010;
assign LUT_4[27470] = 32'b00000000000000000010001001110110;
assign LUT_4[27471] = 32'b11111111111111111011010101101110;
assign LUT_4[27472] = 32'b00000000000000001010010100001111;
assign LUT_4[27473] = 32'b00000000000000000011100000000111;
assign LUT_4[27474] = 32'b00000000000000001001101110110011;
assign LUT_4[27475] = 32'b00000000000000000010111010101011;
assign LUT_4[27476] = 32'b00000000000000000111010100101011;
assign LUT_4[27477] = 32'b00000000000000000000100000100011;
assign LUT_4[27478] = 32'b00000000000000000110101111001111;
assign LUT_4[27479] = 32'b11111111111111111111111011000111;
assign LUT_4[27480] = 32'b00000000000000000011100000100100;
assign LUT_4[27481] = 32'b11111111111111111100101100011100;
assign LUT_4[27482] = 32'b00000000000000000010111011001000;
assign LUT_4[27483] = 32'b11111111111111111100000111000000;
assign LUT_4[27484] = 32'b00000000000000000000100001000000;
assign LUT_4[27485] = 32'b11111111111111111001101100111000;
assign LUT_4[27486] = 32'b11111111111111111111111011100100;
assign LUT_4[27487] = 32'b11111111111111111001000111011100;
assign LUT_4[27488] = 32'b00000000000000001010111101101000;
assign LUT_4[27489] = 32'b00000000000000000100001001100000;
assign LUT_4[27490] = 32'b00000000000000001010011000001100;
assign LUT_4[27491] = 32'b00000000000000000011100100000100;
assign LUT_4[27492] = 32'b00000000000000000111111110000100;
assign LUT_4[27493] = 32'b00000000000000000001001001111100;
assign LUT_4[27494] = 32'b00000000000000000111011000101000;
assign LUT_4[27495] = 32'b00000000000000000000100100100000;
assign LUT_4[27496] = 32'b00000000000000000100001001111101;
assign LUT_4[27497] = 32'b11111111111111111101010101110101;
assign LUT_4[27498] = 32'b00000000000000000011100100100001;
assign LUT_4[27499] = 32'b11111111111111111100110000011001;
assign LUT_4[27500] = 32'b00000000000000000001001010011001;
assign LUT_4[27501] = 32'b11111111111111111010010110010001;
assign LUT_4[27502] = 32'b00000000000000000000100100111101;
assign LUT_4[27503] = 32'b11111111111111111001110000110101;
assign LUT_4[27504] = 32'b00000000000000001000101111010110;
assign LUT_4[27505] = 32'b00000000000000000001111011001110;
assign LUT_4[27506] = 32'b00000000000000001000001001111010;
assign LUT_4[27507] = 32'b00000000000000000001010101110010;
assign LUT_4[27508] = 32'b00000000000000000101101111110010;
assign LUT_4[27509] = 32'b11111111111111111110111011101010;
assign LUT_4[27510] = 32'b00000000000000000101001010010110;
assign LUT_4[27511] = 32'b11111111111111111110010110001110;
assign LUT_4[27512] = 32'b00000000000000000001111011101011;
assign LUT_4[27513] = 32'b11111111111111111011000111100011;
assign LUT_4[27514] = 32'b00000000000000000001010110001111;
assign LUT_4[27515] = 32'b11111111111111111010100010000111;
assign LUT_4[27516] = 32'b11111111111111111110111100000111;
assign LUT_4[27517] = 32'b11111111111111111000000111111111;
assign LUT_4[27518] = 32'b11111111111111111110010110101011;
assign LUT_4[27519] = 32'b11111111111111110111100010100011;
assign LUT_4[27520] = 32'b00000000000000001101110001010101;
assign LUT_4[27521] = 32'b00000000000000000110111101001101;
assign LUT_4[27522] = 32'b00000000000000001101001011111001;
assign LUT_4[27523] = 32'b00000000000000000110010111110001;
assign LUT_4[27524] = 32'b00000000000000001010110001110001;
assign LUT_4[27525] = 32'b00000000000000000011111101101001;
assign LUT_4[27526] = 32'b00000000000000001010001100010101;
assign LUT_4[27527] = 32'b00000000000000000011011000001101;
assign LUT_4[27528] = 32'b00000000000000000110111101101010;
assign LUT_4[27529] = 32'b00000000000000000000001001100010;
assign LUT_4[27530] = 32'b00000000000000000110011000001110;
assign LUT_4[27531] = 32'b11111111111111111111100100000110;
assign LUT_4[27532] = 32'b00000000000000000011111110000110;
assign LUT_4[27533] = 32'b11111111111111111101001001111110;
assign LUT_4[27534] = 32'b00000000000000000011011000101010;
assign LUT_4[27535] = 32'b11111111111111111100100100100010;
assign LUT_4[27536] = 32'b00000000000000001011100011000011;
assign LUT_4[27537] = 32'b00000000000000000100101110111011;
assign LUT_4[27538] = 32'b00000000000000001010111101100111;
assign LUT_4[27539] = 32'b00000000000000000100001001011111;
assign LUT_4[27540] = 32'b00000000000000001000100011011111;
assign LUT_4[27541] = 32'b00000000000000000001101111010111;
assign LUT_4[27542] = 32'b00000000000000000111111110000011;
assign LUT_4[27543] = 32'b00000000000000000001001001111011;
assign LUT_4[27544] = 32'b00000000000000000100101111011000;
assign LUT_4[27545] = 32'b11111111111111111101111011010000;
assign LUT_4[27546] = 32'b00000000000000000100001001111100;
assign LUT_4[27547] = 32'b11111111111111111101010101110100;
assign LUT_4[27548] = 32'b00000000000000000001101111110100;
assign LUT_4[27549] = 32'b11111111111111111010111011101100;
assign LUT_4[27550] = 32'b00000000000000000001001010011000;
assign LUT_4[27551] = 32'b11111111111111111010010110010000;
assign LUT_4[27552] = 32'b00000000000000001100001100011100;
assign LUT_4[27553] = 32'b00000000000000000101011000010100;
assign LUT_4[27554] = 32'b00000000000000001011100111000000;
assign LUT_4[27555] = 32'b00000000000000000100110010111000;
assign LUT_4[27556] = 32'b00000000000000001001001100111000;
assign LUT_4[27557] = 32'b00000000000000000010011000110000;
assign LUT_4[27558] = 32'b00000000000000001000100111011100;
assign LUT_4[27559] = 32'b00000000000000000001110011010100;
assign LUT_4[27560] = 32'b00000000000000000101011000110001;
assign LUT_4[27561] = 32'b11111111111111111110100100101001;
assign LUT_4[27562] = 32'b00000000000000000100110011010101;
assign LUT_4[27563] = 32'b11111111111111111101111111001101;
assign LUT_4[27564] = 32'b00000000000000000010011001001101;
assign LUT_4[27565] = 32'b11111111111111111011100101000101;
assign LUT_4[27566] = 32'b00000000000000000001110011110001;
assign LUT_4[27567] = 32'b11111111111111111010111111101001;
assign LUT_4[27568] = 32'b00000000000000001001111110001010;
assign LUT_4[27569] = 32'b00000000000000000011001010000010;
assign LUT_4[27570] = 32'b00000000000000001001011000101110;
assign LUT_4[27571] = 32'b00000000000000000010100100100110;
assign LUT_4[27572] = 32'b00000000000000000110111110100110;
assign LUT_4[27573] = 32'b00000000000000000000001010011110;
assign LUT_4[27574] = 32'b00000000000000000110011001001010;
assign LUT_4[27575] = 32'b11111111111111111111100101000010;
assign LUT_4[27576] = 32'b00000000000000000011001010011111;
assign LUT_4[27577] = 32'b11111111111111111100010110010111;
assign LUT_4[27578] = 32'b00000000000000000010100101000011;
assign LUT_4[27579] = 32'b11111111111111111011110000111011;
assign LUT_4[27580] = 32'b00000000000000000000001010111011;
assign LUT_4[27581] = 32'b11111111111111111001010110110011;
assign LUT_4[27582] = 32'b11111111111111111111100101011111;
assign LUT_4[27583] = 32'b11111111111111111000110001010111;
assign LUT_4[27584] = 32'b00000000000000001111001000101001;
assign LUT_4[27585] = 32'b00000000000000001000010100100001;
assign LUT_4[27586] = 32'b00000000000000001110100011001101;
assign LUT_4[27587] = 32'b00000000000000000111101111000101;
assign LUT_4[27588] = 32'b00000000000000001100001001000101;
assign LUT_4[27589] = 32'b00000000000000000101010100111101;
assign LUT_4[27590] = 32'b00000000000000001011100011101001;
assign LUT_4[27591] = 32'b00000000000000000100101111100001;
assign LUT_4[27592] = 32'b00000000000000001000010100111110;
assign LUT_4[27593] = 32'b00000000000000000001100000110110;
assign LUT_4[27594] = 32'b00000000000000000111101111100010;
assign LUT_4[27595] = 32'b00000000000000000000111011011010;
assign LUT_4[27596] = 32'b00000000000000000101010101011010;
assign LUT_4[27597] = 32'b11111111111111111110100001010010;
assign LUT_4[27598] = 32'b00000000000000000100101111111110;
assign LUT_4[27599] = 32'b11111111111111111101111011110110;
assign LUT_4[27600] = 32'b00000000000000001100111010010111;
assign LUT_4[27601] = 32'b00000000000000000110000110001111;
assign LUT_4[27602] = 32'b00000000000000001100010100111011;
assign LUT_4[27603] = 32'b00000000000000000101100000110011;
assign LUT_4[27604] = 32'b00000000000000001001111010110011;
assign LUT_4[27605] = 32'b00000000000000000011000110101011;
assign LUT_4[27606] = 32'b00000000000000001001010101010111;
assign LUT_4[27607] = 32'b00000000000000000010100001001111;
assign LUT_4[27608] = 32'b00000000000000000110000110101100;
assign LUT_4[27609] = 32'b11111111111111111111010010100100;
assign LUT_4[27610] = 32'b00000000000000000101100001010000;
assign LUT_4[27611] = 32'b11111111111111111110101101001000;
assign LUT_4[27612] = 32'b00000000000000000011000111001000;
assign LUT_4[27613] = 32'b11111111111111111100010011000000;
assign LUT_4[27614] = 32'b00000000000000000010100001101100;
assign LUT_4[27615] = 32'b11111111111111111011101101100100;
assign LUT_4[27616] = 32'b00000000000000001101100011110000;
assign LUT_4[27617] = 32'b00000000000000000110101111101000;
assign LUT_4[27618] = 32'b00000000000000001100111110010100;
assign LUT_4[27619] = 32'b00000000000000000110001010001100;
assign LUT_4[27620] = 32'b00000000000000001010100100001100;
assign LUT_4[27621] = 32'b00000000000000000011110000000100;
assign LUT_4[27622] = 32'b00000000000000001001111110110000;
assign LUT_4[27623] = 32'b00000000000000000011001010101000;
assign LUT_4[27624] = 32'b00000000000000000110110000000101;
assign LUT_4[27625] = 32'b11111111111111111111111011111101;
assign LUT_4[27626] = 32'b00000000000000000110001010101001;
assign LUT_4[27627] = 32'b11111111111111111111010110100001;
assign LUT_4[27628] = 32'b00000000000000000011110000100001;
assign LUT_4[27629] = 32'b11111111111111111100111100011001;
assign LUT_4[27630] = 32'b00000000000000000011001011000101;
assign LUT_4[27631] = 32'b11111111111111111100010110111101;
assign LUT_4[27632] = 32'b00000000000000001011010101011110;
assign LUT_4[27633] = 32'b00000000000000000100100001010110;
assign LUT_4[27634] = 32'b00000000000000001010110000000010;
assign LUT_4[27635] = 32'b00000000000000000011111011111010;
assign LUT_4[27636] = 32'b00000000000000001000010101111010;
assign LUT_4[27637] = 32'b00000000000000000001100001110010;
assign LUT_4[27638] = 32'b00000000000000000111110000011110;
assign LUT_4[27639] = 32'b00000000000000000000111100010110;
assign LUT_4[27640] = 32'b00000000000000000100100001110011;
assign LUT_4[27641] = 32'b11111111111111111101101101101011;
assign LUT_4[27642] = 32'b00000000000000000011111100010111;
assign LUT_4[27643] = 32'b11111111111111111101001000001111;
assign LUT_4[27644] = 32'b00000000000000000001100010001111;
assign LUT_4[27645] = 32'b11111111111111111010101110000111;
assign LUT_4[27646] = 32'b00000000000000000000111100110011;
assign LUT_4[27647] = 32'b11111111111111111010001000101011;
assign LUT_4[27648] = 32'b00000000000000001000110110000001;
assign LUT_4[27649] = 32'b00000000000000000010000001111001;
assign LUT_4[27650] = 32'b00000000000000001000010000100101;
assign LUT_4[27651] = 32'b00000000000000000001011100011101;
assign LUT_4[27652] = 32'b00000000000000000101110110011101;
assign LUT_4[27653] = 32'b11111111111111111111000010010101;
assign LUT_4[27654] = 32'b00000000000000000101010001000001;
assign LUT_4[27655] = 32'b11111111111111111110011100111001;
assign LUT_4[27656] = 32'b00000000000000000010000010010110;
assign LUT_4[27657] = 32'b11111111111111111011001110001110;
assign LUT_4[27658] = 32'b00000000000000000001011100111010;
assign LUT_4[27659] = 32'b11111111111111111010101000110010;
assign LUT_4[27660] = 32'b11111111111111111111000010110010;
assign LUT_4[27661] = 32'b11111111111111111000001110101010;
assign LUT_4[27662] = 32'b11111111111111111110011101010110;
assign LUT_4[27663] = 32'b11111111111111110111101001001110;
assign LUT_4[27664] = 32'b00000000000000000110100111101111;
assign LUT_4[27665] = 32'b11111111111111111111110011100111;
assign LUT_4[27666] = 32'b00000000000000000110000010010011;
assign LUT_4[27667] = 32'b11111111111111111111001110001011;
assign LUT_4[27668] = 32'b00000000000000000011101000001011;
assign LUT_4[27669] = 32'b11111111111111111100110100000011;
assign LUT_4[27670] = 32'b00000000000000000011000010101111;
assign LUT_4[27671] = 32'b11111111111111111100001110100111;
assign LUT_4[27672] = 32'b11111111111111111111110100000100;
assign LUT_4[27673] = 32'b11111111111111111000111111111100;
assign LUT_4[27674] = 32'b11111111111111111111001110101000;
assign LUT_4[27675] = 32'b11111111111111111000011010100000;
assign LUT_4[27676] = 32'b11111111111111111100110100100000;
assign LUT_4[27677] = 32'b11111111111111110110000000011000;
assign LUT_4[27678] = 32'b11111111111111111100001111000100;
assign LUT_4[27679] = 32'b11111111111111110101011010111100;
assign LUT_4[27680] = 32'b00000000000000000111010001001000;
assign LUT_4[27681] = 32'b00000000000000000000011101000000;
assign LUT_4[27682] = 32'b00000000000000000110101011101100;
assign LUT_4[27683] = 32'b11111111111111111111110111100100;
assign LUT_4[27684] = 32'b00000000000000000100010001100100;
assign LUT_4[27685] = 32'b11111111111111111101011101011100;
assign LUT_4[27686] = 32'b00000000000000000011101100001000;
assign LUT_4[27687] = 32'b11111111111111111100111000000000;
assign LUT_4[27688] = 32'b00000000000000000000011101011101;
assign LUT_4[27689] = 32'b11111111111111111001101001010101;
assign LUT_4[27690] = 32'b11111111111111111111111000000001;
assign LUT_4[27691] = 32'b11111111111111111001000011111001;
assign LUT_4[27692] = 32'b11111111111111111101011101111001;
assign LUT_4[27693] = 32'b11111111111111110110101001110001;
assign LUT_4[27694] = 32'b11111111111111111100111000011101;
assign LUT_4[27695] = 32'b11111111111111110110000100010101;
assign LUT_4[27696] = 32'b00000000000000000101000010110110;
assign LUT_4[27697] = 32'b11111111111111111110001110101110;
assign LUT_4[27698] = 32'b00000000000000000100011101011010;
assign LUT_4[27699] = 32'b11111111111111111101101001010010;
assign LUT_4[27700] = 32'b00000000000000000010000011010010;
assign LUT_4[27701] = 32'b11111111111111111011001111001010;
assign LUT_4[27702] = 32'b00000000000000000001011101110110;
assign LUT_4[27703] = 32'b11111111111111111010101001101110;
assign LUT_4[27704] = 32'b11111111111111111110001111001011;
assign LUT_4[27705] = 32'b11111111111111110111011011000011;
assign LUT_4[27706] = 32'b11111111111111111101101001101111;
assign LUT_4[27707] = 32'b11111111111111110110110101100111;
assign LUT_4[27708] = 32'b11111111111111111011001111100111;
assign LUT_4[27709] = 32'b11111111111111110100011011011111;
assign LUT_4[27710] = 32'b11111111111111111010101010001011;
assign LUT_4[27711] = 32'b11111111111111110011110110000011;
assign LUT_4[27712] = 32'b00000000000000001010001101010101;
assign LUT_4[27713] = 32'b00000000000000000011011001001101;
assign LUT_4[27714] = 32'b00000000000000001001100111111001;
assign LUT_4[27715] = 32'b00000000000000000010110011110001;
assign LUT_4[27716] = 32'b00000000000000000111001101110001;
assign LUT_4[27717] = 32'b00000000000000000000011001101001;
assign LUT_4[27718] = 32'b00000000000000000110101000010101;
assign LUT_4[27719] = 32'b11111111111111111111110100001101;
assign LUT_4[27720] = 32'b00000000000000000011011001101010;
assign LUT_4[27721] = 32'b11111111111111111100100101100010;
assign LUT_4[27722] = 32'b00000000000000000010110100001110;
assign LUT_4[27723] = 32'b11111111111111111100000000000110;
assign LUT_4[27724] = 32'b00000000000000000000011010000110;
assign LUT_4[27725] = 32'b11111111111111111001100101111110;
assign LUT_4[27726] = 32'b11111111111111111111110100101010;
assign LUT_4[27727] = 32'b11111111111111111001000000100010;
assign LUT_4[27728] = 32'b00000000000000000111111111000011;
assign LUT_4[27729] = 32'b00000000000000000001001010111011;
assign LUT_4[27730] = 32'b00000000000000000111011001100111;
assign LUT_4[27731] = 32'b00000000000000000000100101011111;
assign LUT_4[27732] = 32'b00000000000000000100111111011111;
assign LUT_4[27733] = 32'b11111111111111111110001011010111;
assign LUT_4[27734] = 32'b00000000000000000100011010000011;
assign LUT_4[27735] = 32'b11111111111111111101100101111011;
assign LUT_4[27736] = 32'b00000000000000000001001011011000;
assign LUT_4[27737] = 32'b11111111111111111010010111010000;
assign LUT_4[27738] = 32'b00000000000000000000100101111100;
assign LUT_4[27739] = 32'b11111111111111111001110001110100;
assign LUT_4[27740] = 32'b11111111111111111110001011110100;
assign LUT_4[27741] = 32'b11111111111111110111010111101100;
assign LUT_4[27742] = 32'b11111111111111111101100110011000;
assign LUT_4[27743] = 32'b11111111111111110110110010010000;
assign LUT_4[27744] = 32'b00000000000000001000101000011100;
assign LUT_4[27745] = 32'b00000000000000000001110100010100;
assign LUT_4[27746] = 32'b00000000000000001000000011000000;
assign LUT_4[27747] = 32'b00000000000000000001001110111000;
assign LUT_4[27748] = 32'b00000000000000000101101000111000;
assign LUT_4[27749] = 32'b11111111111111111110110100110000;
assign LUT_4[27750] = 32'b00000000000000000101000011011100;
assign LUT_4[27751] = 32'b11111111111111111110001111010100;
assign LUT_4[27752] = 32'b00000000000000000001110100110001;
assign LUT_4[27753] = 32'b11111111111111111011000000101001;
assign LUT_4[27754] = 32'b00000000000000000001001111010101;
assign LUT_4[27755] = 32'b11111111111111111010011011001101;
assign LUT_4[27756] = 32'b11111111111111111110110101001101;
assign LUT_4[27757] = 32'b11111111111111111000000001000101;
assign LUT_4[27758] = 32'b11111111111111111110001111110001;
assign LUT_4[27759] = 32'b11111111111111110111011011101001;
assign LUT_4[27760] = 32'b00000000000000000110011010001010;
assign LUT_4[27761] = 32'b11111111111111111111100110000010;
assign LUT_4[27762] = 32'b00000000000000000101110100101110;
assign LUT_4[27763] = 32'b11111111111111111111000000100110;
assign LUT_4[27764] = 32'b00000000000000000011011010100110;
assign LUT_4[27765] = 32'b11111111111111111100100110011110;
assign LUT_4[27766] = 32'b00000000000000000010110101001010;
assign LUT_4[27767] = 32'b11111111111111111100000001000010;
assign LUT_4[27768] = 32'b11111111111111111111100110011111;
assign LUT_4[27769] = 32'b11111111111111111000110010010111;
assign LUT_4[27770] = 32'b11111111111111111111000001000011;
assign LUT_4[27771] = 32'b11111111111111111000001100111011;
assign LUT_4[27772] = 32'b11111111111111111100100110111011;
assign LUT_4[27773] = 32'b11111111111111110101110010110011;
assign LUT_4[27774] = 32'b11111111111111111100000001011111;
assign LUT_4[27775] = 32'b11111111111111110101001101010111;
assign LUT_4[27776] = 32'b00000000000000001011011100001001;
assign LUT_4[27777] = 32'b00000000000000000100101000000001;
assign LUT_4[27778] = 32'b00000000000000001010110110101101;
assign LUT_4[27779] = 32'b00000000000000000100000010100101;
assign LUT_4[27780] = 32'b00000000000000001000011100100101;
assign LUT_4[27781] = 32'b00000000000000000001101000011101;
assign LUT_4[27782] = 32'b00000000000000000111110111001001;
assign LUT_4[27783] = 32'b00000000000000000001000011000001;
assign LUT_4[27784] = 32'b00000000000000000100101000011110;
assign LUT_4[27785] = 32'b11111111111111111101110100010110;
assign LUT_4[27786] = 32'b00000000000000000100000011000010;
assign LUT_4[27787] = 32'b11111111111111111101001110111010;
assign LUT_4[27788] = 32'b00000000000000000001101000111010;
assign LUT_4[27789] = 32'b11111111111111111010110100110010;
assign LUT_4[27790] = 32'b00000000000000000001000011011110;
assign LUT_4[27791] = 32'b11111111111111111010001111010110;
assign LUT_4[27792] = 32'b00000000000000001001001101110111;
assign LUT_4[27793] = 32'b00000000000000000010011001101111;
assign LUT_4[27794] = 32'b00000000000000001000101000011011;
assign LUT_4[27795] = 32'b00000000000000000001110100010011;
assign LUT_4[27796] = 32'b00000000000000000110001110010011;
assign LUT_4[27797] = 32'b11111111111111111111011010001011;
assign LUT_4[27798] = 32'b00000000000000000101101000110111;
assign LUT_4[27799] = 32'b11111111111111111110110100101111;
assign LUT_4[27800] = 32'b00000000000000000010011010001100;
assign LUT_4[27801] = 32'b11111111111111111011100110000100;
assign LUT_4[27802] = 32'b00000000000000000001110100110000;
assign LUT_4[27803] = 32'b11111111111111111011000000101000;
assign LUT_4[27804] = 32'b11111111111111111111011010101000;
assign LUT_4[27805] = 32'b11111111111111111000100110100000;
assign LUT_4[27806] = 32'b11111111111111111110110101001100;
assign LUT_4[27807] = 32'b11111111111111111000000001000100;
assign LUT_4[27808] = 32'b00000000000000001001110111010000;
assign LUT_4[27809] = 32'b00000000000000000011000011001000;
assign LUT_4[27810] = 32'b00000000000000001001010001110100;
assign LUT_4[27811] = 32'b00000000000000000010011101101100;
assign LUT_4[27812] = 32'b00000000000000000110110111101100;
assign LUT_4[27813] = 32'b00000000000000000000000011100100;
assign LUT_4[27814] = 32'b00000000000000000110010010010000;
assign LUT_4[27815] = 32'b11111111111111111111011110001000;
assign LUT_4[27816] = 32'b00000000000000000011000011100101;
assign LUT_4[27817] = 32'b11111111111111111100001111011101;
assign LUT_4[27818] = 32'b00000000000000000010011110001001;
assign LUT_4[27819] = 32'b11111111111111111011101010000001;
assign LUT_4[27820] = 32'b00000000000000000000000100000001;
assign LUT_4[27821] = 32'b11111111111111111001001111111001;
assign LUT_4[27822] = 32'b11111111111111111111011110100101;
assign LUT_4[27823] = 32'b11111111111111111000101010011101;
assign LUT_4[27824] = 32'b00000000000000000111101000111110;
assign LUT_4[27825] = 32'b00000000000000000000110100110110;
assign LUT_4[27826] = 32'b00000000000000000111000011100010;
assign LUT_4[27827] = 32'b00000000000000000000001111011010;
assign LUT_4[27828] = 32'b00000000000000000100101001011010;
assign LUT_4[27829] = 32'b11111111111111111101110101010010;
assign LUT_4[27830] = 32'b00000000000000000100000011111110;
assign LUT_4[27831] = 32'b11111111111111111101001111110110;
assign LUT_4[27832] = 32'b00000000000000000000110101010011;
assign LUT_4[27833] = 32'b11111111111111111010000001001011;
assign LUT_4[27834] = 32'b00000000000000000000001111110111;
assign LUT_4[27835] = 32'b11111111111111111001011011101111;
assign LUT_4[27836] = 32'b11111111111111111101110101101111;
assign LUT_4[27837] = 32'b11111111111111110111000001100111;
assign LUT_4[27838] = 32'b11111111111111111101010000010011;
assign LUT_4[27839] = 32'b11111111111111110110011100001011;
assign LUT_4[27840] = 32'b00000000000000001100110011011101;
assign LUT_4[27841] = 32'b00000000000000000101111111010101;
assign LUT_4[27842] = 32'b00000000000000001100001110000001;
assign LUT_4[27843] = 32'b00000000000000000101011001111001;
assign LUT_4[27844] = 32'b00000000000000001001110011111001;
assign LUT_4[27845] = 32'b00000000000000000010111111110001;
assign LUT_4[27846] = 32'b00000000000000001001001110011101;
assign LUT_4[27847] = 32'b00000000000000000010011010010101;
assign LUT_4[27848] = 32'b00000000000000000101111111110010;
assign LUT_4[27849] = 32'b11111111111111111111001011101010;
assign LUT_4[27850] = 32'b00000000000000000101011010010110;
assign LUT_4[27851] = 32'b11111111111111111110100110001110;
assign LUT_4[27852] = 32'b00000000000000000011000000001110;
assign LUT_4[27853] = 32'b11111111111111111100001100000110;
assign LUT_4[27854] = 32'b00000000000000000010011010110010;
assign LUT_4[27855] = 32'b11111111111111111011100110101010;
assign LUT_4[27856] = 32'b00000000000000001010100101001011;
assign LUT_4[27857] = 32'b00000000000000000011110001000011;
assign LUT_4[27858] = 32'b00000000000000001001111111101111;
assign LUT_4[27859] = 32'b00000000000000000011001011100111;
assign LUT_4[27860] = 32'b00000000000000000111100101100111;
assign LUT_4[27861] = 32'b00000000000000000000110001011111;
assign LUT_4[27862] = 32'b00000000000000000111000000001011;
assign LUT_4[27863] = 32'b00000000000000000000001100000011;
assign LUT_4[27864] = 32'b00000000000000000011110001100000;
assign LUT_4[27865] = 32'b11111111111111111100111101011000;
assign LUT_4[27866] = 32'b00000000000000000011001100000100;
assign LUT_4[27867] = 32'b11111111111111111100010111111100;
assign LUT_4[27868] = 32'b00000000000000000000110001111100;
assign LUT_4[27869] = 32'b11111111111111111001111101110100;
assign LUT_4[27870] = 32'b00000000000000000000001100100000;
assign LUT_4[27871] = 32'b11111111111111111001011000011000;
assign LUT_4[27872] = 32'b00000000000000001011001110100100;
assign LUT_4[27873] = 32'b00000000000000000100011010011100;
assign LUT_4[27874] = 32'b00000000000000001010101001001000;
assign LUT_4[27875] = 32'b00000000000000000011110101000000;
assign LUT_4[27876] = 32'b00000000000000001000001111000000;
assign LUT_4[27877] = 32'b00000000000000000001011010111000;
assign LUT_4[27878] = 32'b00000000000000000111101001100100;
assign LUT_4[27879] = 32'b00000000000000000000110101011100;
assign LUT_4[27880] = 32'b00000000000000000100011010111001;
assign LUT_4[27881] = 32'b11111111111111111101100110110001;
assign LUT_4[27882] = 32'b00000000000000000011110101011101;
assign LUT_4[27883] = 32'b11111111111111111101000001010101;
assign LUT_4[27884] = 32'b00000000000000000001011011010101;
assign LUT_4[27885] = 32'b11111111111111111010100111001101;
assign LUT_4[27886] = 32'b00000000000000000000110101111001;
assign LUT_4[27887] = 32'b11111111111111111010000001110001;
assign LUT_4[27888] = 32'b00000000000000001001000000010010;
assign LUT_4[27889] = 32'b00000000000000000010001100001010;
assign LUT_4[27890] = 32'b00000000000000001000011010110110;
assign LUT_4[27891] = 32'b00000000000000000001100110101110;
assign LUT_4[27892] = 32'b00000000000000000110000000101110;
assign LUT_4[27893] = 32'b11111111111111111111001100100110;
assign LUT_4[27894] = 32'b00000000000000000101011011010010;
assign LUT_4[27895] = 32'b11111111111111111110100111001010;
assign LUT_4[27896] = 32'b00000000000000000010001100100111;
assign LUT_4[27897] = 32'b11111111111111111011011000011111;
assign LUT_4[27898] = 32'b00000000000000000001100111001011;
assign LUT_4[27899] = 32'b11111111111111111010110011000011;
assign LUT_4[27900] = 32'b11111111111111111111001101000011;
assign LUT_4[27901] = 32'b11111111111111111000011000111011;
assign LUT_4[27902] = 32'b11111111111111111110100111100111;
assign LUT_4[27903] = 32'b11111111111111110111110011011111;
assign LUT_4[27904] = 32'b00000000000000001101110001100100;
assign LUT_4[27905] = 32'b00000000000000000110111101011100;
assign LUT_4[27906] = 32'b00000000000000001101001100001000;
assign LUT_4[27907] = 32'b00000000000000000110011000000000;
assign LUT_4[27908] = 32'b00000000000000001010110010000000;
assign LUT_4[27909] = 32'b00000000000000000011111101111000;
assign LUT_4[27910] = 32'b00000000000000001010001100100100;
assign LUT_4[27911] = 32'b00000000000000000011011000011100;
assign LUT_4[27912] = 32'b00000000000000000110111101111001;
assign LUT_4[27913] = 32'b00000000000000000000001001110001;
assign LUT_4[27914] = 32'b00000000000000000110011000011101;
assign LUT_4[27915] = 32'b11111111111111111111100100010101;
assign LUT_4[27916] = 32'b00000000000000000011111110010101;
assign LUT_4[27917] = 32'b11111111111111111101001010001101;
assign LUT_4[27918] = 32'b00000000000000000011011000111001;
assign LUT_4[27919] = 32'b11111111111111111100100100110001;
assign LUT_4[27920] = 32'b00000000000000001011100011010010;
assign LUT_4[27921] = 32'b00000000000000000100101111001010;
assign LUT_4[27922] = 32'b00000000000000001010111101110110;
assign LUT_4[27923] = 32'b00000000000000000100001001101110;
assign LUT_4[27924] = 32'b00000000000000001000100011101110;
assign LUT_4[27925] = 32'b00000000000000000001101111100110;
assign LUT_4[27926] = 32'b00000000000000000111111110010010;
assign LUT_4[27927] = 32'b00000000000000000001001010001010;
assign LUT_4[27928] = 32'b00000000000000000100101111100111;
assign LUT_4[27929] = 32'b11111111111111111101111011011111;
assign LUT_4[27930] = 32'b00000000000000000100001010001011;
assign LUT_4[27931] = 32'b11111111111111111101010110000011;
assign LUT_4[27932] = 32'b00000000000000000001110000000011;
assign LUT_4[27933] = 32'b11111111111111111010111011111011;
assign LUT_4[27934] = 32'b00000000000000000001001010100111;
assign LUT_4[27935] = 32'b11111111111111111010010110011111;
assign LUT_4[27936] = 32'b00000000000000001100001100101011;
assign LUT_4[27937] = 32'b00000000000000000101011000100011;
assign LUT_4[27938] = 32'b00000000000000001011100111001111;
assign LUT_4[27939] = 32'b00000000000000000100110011000111;
assign LUT_4[27940] = 32'b00000000000000001001001101000111;
assign LUT_4[27941] = 32'b00000000000000000010011000111111;
assign LUT_4[27942] = 32'b00000000000000001000100111101011;
assign LUT_4[27943] = 32'b00000000000000000001110011100011;
assign LUT_4[27944] = 32'b00000000000000000101011001000000;
assign LUT_4[27945] = 32'b11111111111111111110100100111000;
assign LUT_4[27946] = 32'b00000000000000000100110011100100;
assign LUT_4[27947] = 32'b11111111111111111101111111011100;
assign LUT_4[27948] = 32'b00000000000000000010011001011100;
assign LUT_4[27949] = 32'b11111111111111111011100101010100;
assign LUT_4[27950] = 32'b00000000000000000001110100000000;
assign LUT_4[27951] = 32'b11111111111111111010111111111000;
assign LUT_4[27952] = 32'b00000000000000001001111110011001;
assign LUT_4[27953] = 32'b00000000000000000011001010010001;
assign LUT_4[27954] = 32'b00000000000000001001011000111101;
assign LUT_4[27955] = 32'b00000000000000000010100100110101;
assign LUT_4[27956] = 32'b00000000000000000110111110110101;
assign LUT_4[27957] = 32'b00000000000000000000001010101101;
assign LUT_4[27958] = 32'b00000000000000000110011001011001;
assign LUT_4[27959] = 32'b11111111111111111111100101010001;
assign LUT_4[27960] = 32'b00000000000000000011001010101110;
assign LUT_4[27961] = 32'b11111111111111111100010110100110;
assign LUT_4[27962] = 32'b00000000000000000010100101010010;
assign LUT_4[27963] = 32'b11111111111111111011110001001010;
assign LUT_4[27964] = 32'b00000000000000000000001011001010;
assign LUT_4[27965] = 32'b11111111111111111001010111000010;
assign LUT_4[27966] = 32'b11111111111111111111100101101110;
assign LUT_4[27967] = 32'b11111111111111111000110001100110;
assign LUT_4[27968] = 32'b00000000000000001111001000111000;
assign LUT_4[27969] = 32'b00000000000000001000010100110000;
assign LUT_4[27970] = 32'b00000000000000001110100011011100;
assign LUT_4[27971] = 32'b00000000000000000111101111010100;
assign LUT_4[27972] = 32'b00000000000000001100001001010100;
assign LUT_4[27973] = 32'b00000000000000000101010101001100;
assign LUT_4[27974] = 32'b00000000000000001011100011111000;
assign LUT_4[27975] = 32'b00000000000000000100101111110000;
assign LUT_4[27976] = 32'b00000000000000001000010101001101;
assign LUT_4[27977] = 32'b00000000000000000001100001000101;
assign LUT_4[27978] = 32'b00000000000000000111101111110001;
assign LUT_4[27979] = 32'b00000000000000000000111011101001;
assign LUT_4[27980] = 32'b00000000000000000101010101101001;
assign LUT_4[27981] = 32'b11111111111111111110100001100001;
assign LUT_4[27982] = 32'b00000000000000000100110000001101;
assign LUT_4[27983] = 32'b11111111111111111101111100000101;
assign LUT_4[27984] = 32'b00000000000000001100111010100110;
assign LUT_4[27985] = 32'b00000000000000000110000110011110;
assign LUT_4[27986] = 32'b00000000000000001100010101001010;
assign LUT_4[27987] = 32'b00000000000000000101100001000010;
assign LUT_4[27988] = 32'b00000000000000001001111011000010;
assign LUT_4[27989] = 32'b00000000000000000011000110111010;
assign LUT_4[27990] = 32'b00000000000000001001010101100110;
assign LUT_4[27991] = 32'b00000000000000000010100001011110;
assign LUT_4[27992] = 32'b00000000000000000110000110111011;
assign LUT_4[27993] = 32'b11111111111111111111010010110011;
assign LUT_4[27994] = 32'b00000000000000000101100001011111;
assign LUT_4[27995] = 32'b11111111111111111110101101010111;
assign LUT_4[27996] = 32'b00000000000000000011000111010111;
assign LUT_4[27997] = 32'b11111111111111111100010011001111;
assign LUT_4[27998] = 32'b00000000000000000010100001111011;
assign LUT_4[27999] = 32'b11111111111111111011101101110011;
assign LUT_4[28000] = 32'b00000000000000001101100011111111;
assign LUT_4[28001] = 32'b00000000000000000110101111110111;
assign LUT_4[28002] = 32'b00000000000000001100111110100011;
assign LUT_4[28003] = 32'b00000000000000000110001010011011;
assign LUT_4[28004] = 32'b00000000000000001010100100011011;
assign LUT_4[28005] = 32'b00000000000000000011110000010011;
assign LUT_4[28006] = 32'b00000000000000001001111110111111;
assign LUT_4[28007] = 32'b00000000000000000011001010110111;
assign LUT_4[28008] = 32'b00000000000000000110110000010100;
assign LUT_4[28009] = 32'b11111111111111111111111100001100;
assign LUT_4[28010] = 32'b00000000000000000110001010111000;
assign LUT_4[28011] = 32'b11111111111111111111010110110000;
assign LUT_4[28012] = 32'b00000000000000000011110000110000;
assign LUT_4[28013] = 32'b11111111111111111100111100101000;
assign LUT_4[28014] = 32'b00000000000000000011001011010100;
assign LUT_4[28015] = 32'b11111111111111111100010111001100;
assign LUT_4[28016] = 32'b00000000000000001011010101101101;
assign LUT_4[28017] = 32'b00000000000000000100100001100101;
assign LUT_4[28018] = 32'b00000000000000001010110000010001;
assign LUT_4[28019] = 32'b00000000000000000011111100001001;
assign LUT_4[28020] = 32'b00000000000000001000010110001001;
assign LUT_4[28021] = 32'b00000000000000000001100010000001;
assign LUT_4[28022] = 32'b00000000000000000111110000101101;
assign LUT_4[28023] = 32'b00000000000000000000111100100101;
assign LUT_4[28024] = 32'b00000000000000000100100010000010;
assign LUT_4[28025] = 32'b11111111111111111101101101111010;
assign LUT_4[28026] = 32'b00000000000000000011111100100110;
assign LUT_4[28027] = 32'b11111111111111111101001000011110;
assign LUT_4[28028] = 32'b00000000000000000001100010011110;
assign LUT_4[28029] = 32'b11111111111111111010101110010110;
assign LUT_4[28030] = 32'b00000000000000000000111101000010;
assign LUT_4[28031] = 32'b11111111111111111010001000111010;
assign LUT_4[28032] = 32'b00000000000000010000010111101100;
assign LUT_4[28033] = 32'b00000000000000001001100011100100;
assign LUT_4[28034] = 32'b00000000000000001111110010010000;
assign LUT_4[28035] = 32'b00000000000000001000111110001000;
assign LUT_4[28036] = 32'b00000000000000001101011000001000;
assign LUT_4[28037] = 32'b00000000000000000110100100000000;
assign LUT_4[28038] = 32'b00000000000000001100110010101100;
assign LUT_4[28039] = 32'b00000000000000000101111110100100;
assign LUT_4[28040] = 32'b00000000000000001001100100000001;
assign LUT_4[28041] = 32'b00000000000000000010101111111001;
assign LUT_4[28042] = 32'b00000000000000001000111110100101;
assign LUT_4[28043] = 32'b00000000000000000010001010011101;
assign LUT_4[28044] = 32'b00000000000000000110100100011101;
assign LUT_4[28045] = 32'b11111111111111111111110000010101;
assign LUT_4[28046] = 32'b00000000000000000101111111000001;
assign LUT_4[28047] = 32'b11111111111111111111001010111001;
assign LUT_4[28048] = 32'b00000000000000001110001001011010;
assign LUT_4[28049] = 32'b00000000000000000111010101010010;
assign LUT_4[28050] = 32'b00000000000000001101100011111110;
assign LUT_4[28051] = 32'b00000000000000000110101111110110;
assign LUT_4[28052] = 32'b00000000000000001011001001110110;
assign LUT_4[28053] = 32'b00000000000000000100010101101110;
assign LUT_4[28054] = 32'b00000000000000001010100100011010;
assign LUT_4[28055] = 32'b00000000000000000011110000010010;
assign LUT_4[28056] = 32'b00000000000000000111010101101111;
assign LUT_4[28057] = 32'b00000000000000000000100001100111;
assign LUT_4[28058] = 32'b00000000000000000110110000010011;
assign LUT_4[28059] = 32'b11111111111111111111111100001011;
assign LUT_4[28060] = 32'b00000000000000000100010110001011;
assign LUT_4[28061] = 32'b11111111111111111101100010000011;
assign LUT_4[28062] = 32'b00000000000000000011110000101111;
assign LUT_4[28063] = 32'b11111111111111111100111100100111;
assign LUT_4[28064] = 32'b00000000000000001110110010110011;
assign LUT_4[28065] = 32'b00000000000000000111111110101011;
assign LUT_4[28066] = 32'b00000000000000001110001101010111;
assign LUT_4[28067] = 32'b00000000000000000111011001001111;
assign LUT_4[28068] = 32'b00000000000000001011110011001111;
assign LUT_4[28069] = 32'b00000000000000000100111111000111;
assign LUT_4[28070] = 32'b00000000000000001011001101110011;
assign LUT_4[28071] = 32'b00000000000000000100011001101011;
assign LUT_4[28072] = 32'b00000000000000000111111111001000;
assign LUT_4[28073] = 32'b00000000000000000001001011000000;
assign LUT_4[28074] = 32'b00000000000000000111011001101100;
assign LUT_4[28075] = 32'b00000000000000000000100101100100;
assign LUT_4[28076] = 32'b00000000000000000100111111100100;
assign LUT_4[28077] = 32'b11111111111111111110001011011100;
assign LUT_4[28078] = 32'b00000000000000000100011010001000;
assign LUT_4[28079] = 32'b11111111111111111101100110000000;
assign LUT_4[28080] = 32'b00000000000000001100100100100001;
assign LUT_4[28081] = 32'b00000000000000000101110000011001;
assign LUT_4[28082] = 32'b00000000000000001011111111000101;
assign LUT_4[28083] = 32'b00000000000000000101001010111101;
assign LUT_4[28084] = 32'b00000000000000001001100100111101;
assign LUT_4[28085] = 32'b00000000000000000010110000110101;
assign LUT_4[28086] = 32'b00000000000000001000111111100001;
assign LUT_4[28087] = 32'b00000000000000000010001011011001;
assign LUT_4[28088] = 32'b00000000000000000101110000110110;
assign LUT_4[28089] = 32'b11111111111111111110111100101110;
assign LUT_4[28090] = 32'b00000000000000000101001011011010;
assign LUT_4[28091] = 32'b11111111111111111110010111010010;
assign LUT_4[28092] = 32'b00000000000000000010110001010010;
assign LUT_4[28093] = 32'b11111111111111111011111101001010;
assign LUT_4[28094] = 32'b00000000000000000010001011110110;
assign LUT_4[28095] = 32'b11111111111111111011010111101110;
assign LUT_4[28096] = 32'b00000000000000010001101111000000;
assign LUT_4[28097] = 32'b00000000000000001010111010111000;
assign LUT_4[28098] = 32'b00000000000000010001001001100100;
assign LUT_4[28099] = 32'b00000000000000001010010101011100;
assign LUT_4[28100] = 32'b00000000000000001110101111011100;
assign LUT_4[28101] = 32'b00000000000000000111111011010100;
assign LUT_4[28102] = 32'b00000000000000001110001010000000;
assign LUT_4[28103] = 32'b00000000000000000111010101111000;
assign LUT_4[28104] = 32'b00000000000000001010111011010101;
assign LUT_4[28105] = 32'b00000000000000000100000111001101;
assign LUT_4[28106] = 32'b00000000000000001010010101111001;
assign LUT_4[28107] = 32'b00000000000000000011100001110001;
assign LUT_4[28108] = 32'b00000000000000000111111011110001;
assign LUT_4[28109] = 32'b00000000000000000001000111101001;
assign LUT_4[28110] = 32'b00000000000000000111010110010101;
assign LUT_4[28111] = 32'b00000000000000000000100010001101;
assign LUT_4[28112] = 32'b00000000000000001111100000101110;
assign LUT_4[28113] = 32'b00000000000000001000101100100110;
assign LUT_4[28114] = 32'b00000000000000001110111011010010;
assign LUT_4[28115] = 32'b00000000000000001000000111001010;
assign LUT_4[28116] = 32'b00000000000000001100100001001010;
assign LUT_4[28117] = 32'b00000000000000000101101101000010;
assign LUT_4[28118] = 32'b00000000000000001011111011101110;
assign LUT_4[28119] = 32'b00000000000000000101000111100110;
assign LUT_4[28120] = 32'b00000000000000001000101101000011;
assign LUT_4[28121] = 32'b00000000000000000001111000111011;
assign LUT_4[28122] = 32'b00000000000000001000000111100111;
assign LUT_4[28123] = 32'b00000000000000000001010011011111;
assign LUT_4[28124] = 32'b00000000000000000101101101011111;
assign LUT_4[28125] = 32'b11111111111111111110111001010111;
assign LUT_4[28126] = 32'b00000000000000000101001000000011;
assign LUT_4[28127] = 32'b11111111111111111110010011111011;
assign LUT_4[28128] = 32'b00000000000000010000001010000111;
assign LUT_4[28129] = 32'b00000000000000001001010101111111;
assign LUT_4[28130] = 32'b00000000000000001111100100101011;
assign LUT_4[28131] = 32'b00000000000000001000110000100011;
assign LUT_4[28132] = 32'b00000000000000001101001010100011;
assign LUT_4[28133] = 32'b00000000000000000110010110011011;
assign LUT_4[28134] = 32'b00000000000000001100100101000111;
assign LUT_4[28135] = 32'b00000000000000000101110000111111;
assign LUT_4[28136] = 32'b00000000000000001001010110011100;
assign LUT_4[28137] = 32'b00000000000000000010100010010100;
assign LUT_4[28138] = 32'b00000000000000001000110001000000;
assign LUT_4[28139] = 32'b00000000000000000001111100111000;
assign LUT_4[28140] = 32'b00000000000000000110010110111000;
assign LUT_4[28141] = 32'b11111111111111111111100010110000;
assign LUT_4[28142] = 32'b00000000000000000101110001011100;
assign LUT_4[28143] = 32'b11111111111111111110111101010100;
assign LUT_4[28144] = 32'b00000000000000001101111011110101;
assign LUT_4[28145] = 32'b00000000000000000111000111101101;
assign LUT_4[28146] = 32'b00000000000000001101010110011001;
assign LUT_4[28147] = 32'b00000000000000000110100010010001;
assign LUT_4[28148] = 32'b00000000000000001010111100010001;
assign LUT_4[28149] = 32'b00000000000000000100001000001001;
assign LUT_4[28150] = 32'b00000000000000001010010110110101;
assign LUT_4[28151] = 32'b00000000000000000011100010101101;
assign LUT_4[28152] = 32'b00000000000000000111001000001010;
assign LUT_4[28153] = 32'b00000000000000000000010100000010;
assign LUT_4[28154] = 32'b00000000000000000110100010101110;
assign LUT_4[28155] = 32'b11111111111111111111101110100110;
assign LUT_4[28156] = 32'b00000000000000000100001000100110;
assign LUT_4[28157] = 32'b11111111111111111101010100011110;
assign LUT_4[28158] = 32'b00000000000000000011100011001010;
assign LUT_4[28159] = 32'b11111111111111111100101111000010;
assign LUT_4[28160] = 32'b00000000000000000111111010001001;
assign LUT_4[28161] = 32'b00000000000000000001000110000001;
assign LUT_4[28162] = 32'b00000000000000000111010100101101;
assign LUT_4[28163] = 32'b00000000000000000000100000100101;
assign LUT_4[28164] = 32'b00000000000000000100111010100101;
assign LUT_4[28165] = 32'b11111111111111111110000110011101;
assign LUT_4[28166] = 32'b00000000000000000100010101001001;
assign LUT_4[28167] = 32'b11111111111111111101100001000001;
assign LUT_4[28168] = 32'b00000000000000000001000110011110;
assign LUT_4[28169] = 32'b11111111111111111010010010010110;
assign LUT_4[28170] = 32'b00000000000000000000100001000010;
assign LUT_4[28171] = 32'b11111111111111111001101100111010;
assign LUT_4[28172] = 32'b11111111111111111110000110111010;
assign LUT_4[28173] = 32'b11111111111111110111010010110010;
assign LUT_4[28174] = 32'b11111111111111111101100001011110;
assign LUT_4[28175] = 32'b11111111111111110110101101010110;
assign LUT_4[28176] = 32'b00000000000000000101101011110111;
assign LUT_4[28177] = 32'b11111111111111111110110111101111;
assign LUT_4[28178] = 32'b00000000000000000101000110011011;
assign LUT_4[28179] = 32'b11111111111111111110010010010011;
assign LUT_4[28180] = 32'b00000000000000000010101100010011;
assign LUT_4[28181] = 32'b11111111111111111011111000001011;
assign LUT_4[28182] = 32'b00000000000000000010000110110111;
assign LUT_4[28183] = 32'b11111111111111111011010010101111;
assign LUT_4[28184] = 32'b11111111111111111110111000001100;
assign LUT_4[28185] = 32'b11111111111111111000000100000100;
assign LUT_4[28186] = 32'b11111111111111111110010010110000;
assign LUT_4[28187] = 32'b11111111111111110111011110101000;
assign LUT_4[28188] = 32'b11111111111111111011111000101000;
assign LUT_4[28189] = 32'b11111111111111110101000100100000;
assign LUT_4[28190] = 32'b11111111111111111011010011001100;
assign LUT_4[28191] = 32'b11111111111111110100011111000100;
assign LUT_4[28192] = 32'b00000000000000000110010101010000;
assign LUT_4[28193] = 32'b11111111111111111111100001001000;
assign LUT_4[28194] = 32'b00000000000000000101101111110100;
assign LUT_4[28195] = 32'b11111111111111111110111011101100;
assign LUT_4[28196] = 32'b00000000000000000011010101101100;
assign LUT_4[28197] = 32'b11111111111111111100100001100100;
assign LUT_4[28198] = 32'b00000000000000000010110000010000;
assign LUT_4[28199] = 32'b11111111111111111011111100001000;
assign LUT_4[28200] = 32'b11111111111111111111100001100101;
assign LUT_4[28201] = 32'b11111111111111111000101101011101;
assign LUT_4[28202] = 32'b11111111111111111110111100001001;
assign LUT_4[28203] = 32'b11111111111111111000001000000001;
assign LUT_4[28204] = 32'b11111111111111111100100010000001;
assign LUT_4[28205] = 32'b11111111111111110101101101111001;
assign LUT_4[28206] = 32'b11111111111111111011111100100101;
assign LUT_4[28207] = 32'b11111111111111110101001000011101;
assign LUT_4[28208] = 32'b00000000000000000100000110111110;
assign LUT_4[28209] = 32'b11111111111111111101010010110110;
assign LUT_4[28210] = 32'b00000000000000000011100001100010;
assign LUT_4[28211] = 32'b11111111111111111100101101011010;
assign LUT_4[28212] = 32'b00000000000000000001000111011010;
assign LUT_4[28213] = 32'b11111111111111111010010011010010;
assign LUT_4[28214] = 32'b00000000000000000000100001111110;
assign LUT_4[28215] = 32'b11111111111111111001101101110110;
assign LUT_4[28216] = 32'b11111111111111111101010011010011;
assign LUT_4[28217] = 32'b11111111111111110110011111001011;
assign LUT_4[28218] = 32'b11111111111111111100101101110111;
assign LUT_4[28219] = 32'b11111111111111110101111001101111;
assign LUT_4[28220] = 32'b11111111111111111010010011101111;
assign LUT_4[28221] = 32'b11111111111111110011011111100111;
assign LUT_4[28222] = 32'b11111111111111111001101110010011;
assign LUT_4[28223] = 32'b11111111111111110010111010001011;
assign LUT_4[28224] = 32'b00000000000000001001010001011101;
assign LUT_4[28225] = 32'b00000000000000000010011101010101;
assign LUT_4[28226] = 32'b00000000000000001000101100000001;
assign LUT_4[28227] = 32'b00000000000000000001110111111001;
assign LUT_4[28228] = 32'b00000000000000000110010001111001;
assign LUT_4[28229] = 32'b11111111111111111111011101110001;
assign LUT_4[28230] = 32'b00000000000000000101101100011101;
assign LUT_4[28231] = 32'b11111111111111111110111000010101;
assign LUT_4[28232] = 32'b00000000000000000010011101110010;
assign LUT_4[28233] = 32'b11111111111111111011101001101010;
assign LUT_4[28234] = 32'b00000000000000000001111000010110;
assign LUT_4[28235] = 32'b11111111111111111011000100001110;
assign LUT_4[28236] = 32'b11111111111111111111011110001110;
assign LUT_4[28237] = 32'b11111111111111111000101010000110;
assign LUT_4[28238] = 32'b11111111111111111110111000110010;
assign LUT_4[28239] = 32'b11111111111111111000000100101010;
assign LUT_4[28240] = 32'b00000000000000000111000011001011;
assign LUT_4[28241] = 32'b00000000000000000000001111000011;
assign LUT_4[28242] = 32'b00000000000000000110011101101111;
assign LUT_4[28243] = 32'b11111111111111111111101001100111;
assign LUT_4[28244] = 32'b00000000000000000100000011100111;
assign LUT_4[28245] = 32'b11111111111111111101001111011111;
assign LUT_4[28246] = 32'b00000000000000000011011110001011;
assign LUT_4[28247] = 32'b11111111111111111100101010000011;
assign LUT_4[28248] = 32'b00000000000000000000001111100000;
assign LUT_4[28249] = 32'b11111111111111111001011011011000;
assign LUT_4[28250] = 32'b11111111111111111111101010000100;
assign LUT_4[28251] = 32'b11111111111111111000110101111100;
assign LUT_4[28252] = 32'b11111111111111111101001111111100;
assign LUT_4[28253] = 32'b11111111111111110110011011110100;
assign LUT_4[28254] = 32'b11111111111111111100101010100000;
assign LUT_4[28255] = 32'b11111111111111110101110110011000;
assign LUT_4[28256] = 32'b00000000000000000111101100100100;
assign LUT_4[28257] = 32'b00000000000000000000111000011100;
assign LUT_4[28258] = 32'b00000000000000000111000111001000;
assign LUT_4[28259] = 32'b00000000000000000000010011000000;
assign LUT_4[28260] = 32'b00000000000000000100101101000000;
assign LUT_4[28261] = 32'b11111111111111111101111000111000;
assign LUT_4[28262] = 32'b00000000000000000100000111100100;
assign LUT_4[28263] = 32'b11111111111111111101010011011100;
assign LUT_4[28264] = 32'b00000000000000000000111000111001;
assign LUT_4[28265] = 32'b11111111111111111010000100110001;
assign LUT_4[28266] = 32'b00000000000000000000010011011101;
assign LUT_4[28267] = 32'b11111111111111111001011111010101;
assign LUT_4[28268] = 32'b11111111111111111101111001010101;
assign LUT_4[28269] = 32'b11111111111111110111000101001101;
assign LUT_4[28270] = 32'b11111111111111111101010011111001;
assign LUT_4[28271] = 32'b11111111111111110110011111110001;
assign LUT_4[28272] = 32'b00000000000000000101011110010010;
assign LUT_4[28273] = 32'b11111111111111111110101010001010;
assign LUT_4[28274] = 32'b00000000000000000100111000110110;
assign LUT_4[28275] = 32'b11111111111111111110000100101110;
assign LUT_4[28276] = 32'b00000000000000000010011110101110;
assign LUT_4[28277] = 32'b11111111111111111011101010100110;
assign LUT_4[28278] = 32'b00000000000000000001111001010010;
assign LUT_4[28279] = 32'b11111111111111111011000101001010;
assign LUT_4[28280] = 32'b11111111111111111110101010100111;
assign LUT_4[28281] = 32'b11111111111111110111110110011111;
assign LUT_4[28282] = 32'b11111111111111111110000101001011;
assign LUT_4[28283] = 32'b11111111111111110111010001000011;
assign LUT_4[28284] = 32'b11111111111111111011101011000011;
assign LUT_4[28285] = 32'b11111111111111110100110110111011;
assign LUT_4[28286] = 32'b11111111111111111011000101100111;
assign LUT_4[28287] = 32'b11111111111111110100010001011111;
assign LUT_4[28288] = 32'b00000000000000001010100000010001;
assign LUT_4[28289] = 32'b00000000000000000011101100001001;
assign LUT_4[28290] = 32'b00000000000000001001111010110101;
assign LUT_4[28291] = 32'b00000000000000000011000110101101;
assign LUT_4[28292] = 32'b00000000000000000111100000101101;
assign LUT_4[28293] = 32'b00000000000000000000101100100101;
assign LUT_4[28294] = 32'b00000000000000000110111011010001;
assign LUT_4[28295] = 32'b00000000000000000000000111001001;
assign LUT_4[28296] = 32'b00000000000000000011101100100110;
assign LUT_4[28297] = 32'b11111111111111111100111000011110;
assign LUT_4[28298] = 32'b00000000000000000011000111001010;
assign LUT_4[28299] = 32'b11111111111111111100010011000010;
assign LUT_4[28300] = 32'b00000000000000000000101101000010;
assign LUT_4[28301] = 32'b11111111111111111001111000111010;
assign LUT_4[28302] = 32'b00000000000000000000000111100110;
assign LUT_4[28303] = 32'b11111111111111111001010011011110;
assign LUT_4[28304] = 32'b00000000000000001000010001111111;
assign LUT_4[28305] = 32'b00000000000000000001011101110111;
assign LUT_4[28306] = 32'b00000000000000000111101100100011;
assign LUT_4[28307] = 32'b00000000000000000000111000011011;
assign LUT_4[28308] = 32'b00000000000000000101010010011011;
assign LUT_4[28309] = 32'b11111111111111111110011110010011;
assign LUT_4[28310] = 32'b00000000000000000100101100111111;
assign LUT_4[28311] = 32'b11111111111111111101111000110111;
assign LUT_4[28312] = 32'b00000000000000000001011110010100;
assign LUT_4[28313] = 32'b11111111111111111010101010001100;
assign LUT_4[28314] = 32'b00000000000000000000111000111000;
assign LUT_4[28315] = 32'b11111111111111111010000100110000;
assign LUT_4[28316] = 32'b11111111111111111110011110110000;
assign LUT_4[28317] = 32'b11111111111111110111101010101000;
assign LUT_4[28318] = 32'b11111111111111111101111001010100;
assign LUT_4[28319] = 32'b11111111111111110111000101001100;
assign LUT_4[28320] = 32'b00000000000000001000111011011000;
assign LUT_4[28321] = 32'b00000000000000000010000111010000;
assign LUT_4[28322] = 32'b00000000000000001000010101111100;
assign LUT_4[28323] = 32'b00000000000000000001100001110100;
assign LUT_4[28324] = 32'b00000000000000000101111011110100;
assign LUT_4[28325] = 32'b11111111111111111111000111101100;
assign LUT_4[28326] = 32'b00000000000000000101010110011000;
assign LUT_4[28327] = 32'b11111111111111111110100010010000;
assign LUT_4[28328] = 32'b00000000000000000010000111101101;
assign LUT_4[28329] = 32'b11111111111111111011010011100101;
assign LUT_4[28330] = 32'b00000000000000000001100010010001;
assign LUT_4[28331] = 32'b11111111111111111010101110001001;
assign LUT_4[28332] = 32'b11111111111111111111001000001001;
assign LUT_4[28333] = 32'b11111111111111111000010100000001;
assign LUT_4[28334] = 32'b11111111111111111110100010101101;
assign LUT_4[28335] = 32'b11111111111111110111101110100101;
assign LUT_4[28336] = 32'b00000000000000000110101101000110;
assign LUT_4[28337] = 32'b11111111111111111111111000111110;
assign LUT_4[28338] = 32'b00000000000000000110000111101010;
assign LUT_4[28339] = 32'b11111111111111111111010011100010;
assign LUT_4[28340] = 32'b00000000000000000011101101100010;
assign LUT_4[28341] = 32'b11111111111111111100111001011010;
assign LUT_4[28342] = 32'b00000000000000000011001000000110;
assign LUT_4[28343] = 32'b11111111111111111100010011111110;
assign LUT_4[28344] = 32'b11111111111111111111111001011011;
assign LUT_4[28345] = 32'b11111111111111111001000101010011;
assign LUT_4[28346] = 32'b11111111111111111111010011111111;
assign LUT_4[28347] = 32'b11111111111111111000011111110111;
assign LUT_4[28348] = 32'b11111111111111111100111001110111;
assign LUT_4[28349] = 32'b11111111111111110110000101101111;
assign LUT_4[28350] = 32'b11111111111111111100010100011011;
assign LUT_4[28351] = 32'b11111111111111110101100000010011;
assign LUT_4[28352] = 32'b00000000000000001011110111100101;
assign LUT_4[28353] = 32'b00000000000000000101000011011101;
assign LUT_4[28354] = 32'b00000000000000001011010010001001;
assign LUT_4[28355] = 32'b00000000000000000100011110000001;
assign LUT_4[28356] = 32'b00000000000000001000111000000001;
assign LUT_4[28357] = 32'b00000000000000000010000011111001;
assign LUT_4[28358] = 32'b00000000000000001000010010100101;
assign LUT_4[28359] = 32'b00000000000000000001011110011101;
assign LUT_4[28360] = 32'b00000000000000000101000011111010;
assign LUT_4[28361] = 32'b11111111111111111110001111110010;
assign LUT_4[28362] = 32'b00000000000000000100011110011110;
assign LUT_4[28363] = 32'b11111111111111111101101010010110;
assign LUT_4[28364] = 32'b00000000000000000010000100010110;
assign LUT_4[28365] = 32'b11111111111111111011010000001110;
assign LUT_4[28366] = 32'b00000000000000000001011110111010;
assign LUT_4[28367] = 32'b11111111111111111010101010110010;
assign LUT_4[28368] = 32'b00000000000000001001101001010011;
assign LUT_4[28369] = 32'b00000000000000000010110101001011;
assign LUT_4[28370] = 32'b00000000000000001001000011110111;
assign LUT_4[28371] = 32'b00000000000000000010001111101111;
assign LUT_4[28372] = 32'b00000000000000000110101001101111;
assign LUT_4[28373] = 32'b11111111111111111111110101100111;
assign LUT_4[28374] = 32'b00000000000000000110000100010011;
assign LUT_4[28375] = 32'b11111111111111111111010000001011;
assign LUT_4[28376] = 32'b00000000000000000010110101101000;
assign LUT_4[28377] = 32'b11111111111111111100000001100000;
assign LUT_4[28378] = 32'b00000000000000000010010000001100;
assign LUT_4[28379] = 32'b11111111111111111011011100000100;
assign LUT_4[28380] = 32'b11111111111111111111110110000100;
assign LUT_4[28381] = 32'b11111111111111111001000001111100;
assign LUT_4[28382] = 32'b11111111111111111111010000101000;
assign LUT_4[28383] = 32'b11111111111111111000011100100000;
assign LUT_4[28384] = 32'b00000000000000001010010010101100;
assign LUT_4[28385] = 32'b00000000000000000011011110100100;
assign LUT_4[28386] = 32'b00000000000000001001101101010000;
assign LUT_4[28387] = 32'b00000000000000000010111001001000;
assign LUT_4[28388] = 32'b00000000000000000111010011001000;
assign LUT_4[28389] = 32'b00000000000000000000011111000000;
assign LUT_4[28390] = 32'b00000000000000000110101101101100;
assign LUT_4[28391] = 32'b11111111111111111111111001100100;
assign LUT_4[28392] = 32'b00000000000000000011011111000001;
assign LUT_4[28393] = 32'b11111111111111111100101010111001;
assign LUT_4[28394] = 32'b00000000000000000010111001100101;
assign LUT_4[28395] = 32'b11111111111111111100000101011101;
assign LUT_4[28396] = 32'b00000000000000000000011111011101;
assign LUT_4[28397] = 32'b11111111111111111001101011010101;
assign LUT_4[28398] = 32'b11111111111111111111111010000001;
assign LUT_4[28399] = 32'b11111111111111111001000101111001;
assign LUT_4[28400] = 32'b00000000000000001000000100011010;
assign LUT_4[28401] = 32'b00000000000000000001010000010010;
assign LUT_4[28402] = 32'b00000000000000000111011110111110;
assign LUT_4[28403] = 32'b00000000000000000000101010110110;
assign LUT_4[28404] = 32'b00000000000000000101000100110110;
assign LUT_4[28405] = 32'b11111111111111111110010000101110;
assign LUT_4[28406] = 32'b00000000000000000100011111011010;
assign LUT_4[28407] = 32'b11111111111111111101101011010010;
assign LUT_4[28408] = 32'b00000000000000000001010000101111;
assign LUT_4[28409] = 32'b11111111111111111010011100100111;
assign LUT_4[28410] = 32'b00000000000000000000101011010011;
assign LUT_4[28411] = 32'b11111111111111111001110111001011;
assign LUT_4[28412] = 32'b11111111111111111110010001001011;
assign LUT_4[28413] = 32'b11111111111111110111011101000011;
assign LUT_4[28414] = 32'b11111111111111111101101011101111;
assign LUT_4[28415] = 32'b11111111111111110110110111100111;
assign LUT_4[28416] = 32'b00000000000000001100110101101100;
assign LUT_4[28417] = 32'b00000000000000000110000001100100;
assign LUT_4[28418] = 32'b00000000000000001100010000010000;
assign LUT_4[28419] = 32'b00000000000000000101011100001000;
assign LUT_4[28420] = 32'b00000000000000001001110110001000;
assign LUT_4[28421] = 32'b00000000000000000011000010000000;
assign LUT_4[28422] = 32'b00000000000000001001010000101100;
assign LUT_4[28423] = 32'b00000000000000000010011100100100;
assign LUT_4[28424] = 32'b00000000000000000110000010000001;
assign LUT_4[28425] = 32'b11111111111111111111001101111001;
assign LUT_4[28426] = 32'b00000000000000000101011100100101;
assign LUT_4[28427] = 32'b11111111111111111110101000011101;
assign LUT_4[28428] = 32'b00000000000000000011000010011101;
assign LUT_4[28429] = 32'b11111111111111111100001110010101;
assign LUT_4[28430] = 32'b00000000000000000010011101000001;
assign LUT_4[28431] = 32'b11111111111111111011101000111001;
assign LUT_4[28432] = 32'b00000000000000001010100111011010;
assign LUT_4[28433] = 32'b00000000000000000011110011010010;
assign LUT_4[28434] = 32'b00000000000000001010000001111110;
assign LUT_4[28435] = 32'b00000000000000000011001101110110;
assign LUT_4[28436] = 32'b00000000000000000111100111110110;
assign LUT_4[28437] = 32'b00000000000000000000110011101110;
assign LUT_4[28438] = 32'b00000000000000000111000010011010;
assign LUT_4[28439] = 32'b00000000000000000000001110010010;
assign LUT_4[28440] = 32'b00000000000000000011110011101111;
assign LUT_4[28441] = 32'b11111111111111111100111111100111;
assign LUT_4[28442] = 32'b00000000000000000011001110010011;
assign LUT_4[28443] = 32'b11111111111111111100011010001011;
assign LUT_4[28444] = 32'b00000000000000000000110100001011;
assign LUT_4[28445] = 32'b11111111111111111010000000000011;
assign LUT_4[28446] = 32'b00000000000000000000001110101111;
assign LUT_4[28447] = 32'b11111111111111111001011010100111;
assign LUT_4[28448] = 32'b00000000000000001011010000110011;
assign LUT_4[28449] = 32'b00000000000000000100011100101011;
assign LUT_4[28450] = 32'b00000000000000001010101011010111;
assign LUT_4[28451] = 32'b00000000000000000011110111001111;
assign LUT_4[28452] = 32'b00000000000000001000010001001111;
assign LUT_4[28453] = 32'b00000000000000000001011101000111;
assign LUT_4[28454] = 32'b00000000000000000111101011110011;
assign LUT_4[28455] = 32'b00000000000000000000110111101011;
assign LUT_4[28456] = 32'b00000000000000000100011101001000;
assign LUT_4[28457] = 32'b11111111111111111101101001000000;
assign LUT_4[28458] = 32'b00000000000000000011110111101100;
assign LUT_4[28459] = 32'b11111111111111111101000011100100;
assign LUT_4[28460] = 32'b00000000000000000001011101100100;
assign LUT_4[28461] = 32'b11111111111111111010101001011100;
assign LUT_4[28462] = 32'b00000000000000000000111000001000;
assign LUT_4[28463] = 32'b11111111111111111010000100000000;
assign LUT_4[28464] = 32'b00000000000000001001000010100001;
assign LUT_4[28465] = 32'b00000000000000000010001110011001;
assign LUT_4[28466] = 32'b00000000000000001000011101000101;
assign LUT_4[28467] = 32'b00000000000000000001101000111101;
assign LUT_4[28468] = 32'b00000000000000000110000010111101;
assign LUT_4[28469] = 32'b11111111111111111111001110110101;
assign LUT_4[28470] = 32'b00000000000000000101011101100001;
assign LUT_4[28471] = 32'b11111111111111111110101001011001;
assign LUT_4[28472] = 32'b00000000000000000010001110110110;
assign LUT_4[28473] = 32'b11111111111111111011011010101110;
assign LUT_4[28474] = 32'b00000000000000000001101001011010;
assign LUT_4[28475] = 32'b11111111111111111010110101010010;
assign LUT_4[28476] = 32'b11111111111111111111001111010010;
assign LUT_4[28477] = 32'b11111111111111111000011011001010;
assign LUT_4[28478] = 32'b11111111111111111110101001110110;
assign LUT_4[28479] = 32'b11111111111111110111110101101110;
assign LUT_4[28480] = 32'b00000000000000001110001101000000;
assign LUT_4[28481] = 32'b00000000000000000111011000111000;
assign LUT_4[28482] = 32'b00000000000000001101100111100100;
assign LUT_4[28483] = 32'b00000000000000000110110011011100;
assign LUT_4[28484] = 32'b00000000000000001011001101011100;
assign LUT_4[28485] = 32'b00000000000000000100011001010100;
assign LUT_4[28486] = 32'b00000000000000001010101000000000;
assign LUT_4[28487] = 32'b00000000000000000011110011111000;
assign LUT_4[28488] = 32'b00000000000000000111011001010101;
assign LUT_4[28489] = 32'b00000000000000000000100101001101;
assign LUT_4[28490] = 32'b00000000000000000110110011111001;
assign LUT_4[28491] = 32'b11111111111111111111111111110001;
assign LUT_4[28492] = 32'b00000000000000000100011001110001;
assign LUT_4[28493] = 32'b11111111111111111101100101101001;
assign LUT_4[28494] = 32'b00000000000000000011110100010101;
assign LUT_4[28495] = 32'b11111111111111111101000000001101;
assign LUT_4[28496] = 32'b00000000000000001011111110101110;
assign LUT_4[28497] = 32'b00000000000000000101001010100110;
assign LUT_4[28498] = 32'b00000000000000001011011001010010;
assign LUT_4[28499] = 32'b00000000000000000100100101001010;
assign LUT_4[28500] = 32'b00000000000000001000111111001010;
assign LUT_4[28501] = 32'b00000000000000000010001011000010;
assign LUT_4[28502] = 32'b00000000000000001000011001101110;
assign LUT_4[28503] = 32'b00000000000000000001100101100110;
assign LUT_4[28504] = 32'b00000000000000000101001011000011;
assign LUT_4[28505] = 32'b11111111111111111110010110111011;
assign LUT_4[28506] = 32'b00000000000000000100100101100111;
assign LUT_4[28507] = 32'b11111111111111111101110001011111;
assign LUT_4[28508] = 32'b00000000000000000010001011011111;
assign LUT_4[28509] = 32'b11111111111111111011010111010111;
assign LUT_4[28510] = 32'b00000000000000000001100110000011;
assign LUT_4[28511] = 32'b11111111111111111010110001111011;
assign LUT_4[28512] = 32'b00000000000000001100101000000111;
assign LUT_4[28513] = 32'b00000000000000000101110011111111;
assign LUT_4[28514] = 32'b00000000000000001100000010101011;
assign LUT_4[28515] = 32'b00000000000000000101001110100011;
assign LUT_4[28516] = 32'b00000000000000001001101000100011;
assign LUT_4[28517] = 32'b00000000000000000010110100011011;
assign LUT_4[28518] = 32'b00000000000000001001000011000111;
assign LUT_4[28519] = 32'b00000000000000000010001110111111;
assign LUT_4[28520] = 32'b00000000000000000101110100011100;
assign LUT_4[28521] = 32'b11111111111111111111000000010100;
assign LUT_4[28522] = 32'b00000000000000000101001111000000;
assign LUT_4[28523] = 32'b11111111111111111110011010111000;
assign LUT_4[28524] = 32'b00000000000000000010110100111000;
assign LUT_4[28525] = 32'b11111111111111111100000000110000;
assign LUT_4[28526] = 32'b00000000000000000010001111011100;
assign LUT_4[28527] = 32'b11111111111111111011011011010100;
assign LUT_4[28528] = 32'b00000000000000001010011001110101;
assign LUT_4[28529] = 32'b00000000000000000011100101101101;
assign LUT_4[28530] = 32'b00000000000000001001110100011001;
assign LUT_4[28531] = 32'b00000000000000000011000000010001;
assign LUT_4[28532] = 32'b00000000000000000111011010010001;
assign LUT_4[28533] = 32'b00000000000000000000100110001001;
assign LUT_4[28534] = 32'b00000000000000000110110100110101;
assign LUT_4[28535] = 32'b00000000000000000000000000101101;
assign LUT_4[28536] = 32'b00000000000000000011100110001010;
assign LUT_4[28537] = 32'b11111111111111111100110010000010;
assign LUT_4[28538] = 32'b00000000000000000011000000101110;
assign LUT_4[28539] = 32'b11111111111111111100001100100110;
assign LUT_4[28540] = 32'b00000000000000000000100110100110;
assign LUT_4[28541] = 32'b11111111111111111001110010011110;
assign LUT_4[28542] = 32'b00000000000000000000000001001010;
assign LUT_4[28543] = 32'b11111111111111111001001101000010;
assign LUT_4[28544] = 32'b00000000000000001111011011110100;
assign LUT_4[28545] = 32'b00000000000000001000100111101100;
assign LUT_4[28546] = 32'b00000000000000001110110110011000;
assign LUT_4[28547] = 32'b00000000000000001000000010010000;
assign LUT_4[28548] = 32'b00000000000000001100011100010000;
assign LUT_4[28549] = 32'b00000000000000000101101000001000;
assign LUT_4[28550] = 32'b00000000000000001011110110110100;
assign LUT_4[28551] = 32'b00000000000000000101000010101100;
assign LUT_4[28552] = 32'b00000000000000001000101000001001;
assign LUT_4[28553] = 32'b00000000000000000001110100000001;
assign LUT_4[28554] = 32'b00000000000000001000000010101101;
assign LUT_4[28555] = 32'b00000000000000000001001110100101;
assign LUT_4[28556] = 32'b00000000000000000101101000100101;
assign LUT_4[28557] = 32'b11111111111111111110110100011101;
assign LUT_4[28558] = 32'b00000000000000000101000011001001;
assign LUT_4[28559] = 32'b11111111111111111110001111000001;
assign LUT_4[28560] = 32'b00000000000000001101001101100010;
assign LUT_4[28561] = 32'b00000000000000000110011001011010;
assign LUT_4[28562] = 32'b00000000000000001100101000000110;
assign LUT_4[28563] = 32'b00000000000000000101110011111110;
assign LUT_4[28564] = 32'b00000000000000001010001101111110;
assign LUT_4[28565] = 32'b00000000000000000011011001110110;
assign LUT_4[28566] = 32'b00000000000000001001101000100010;
assign LUT_4[28567] = 32'b00000000000000000010110100011010;
assign LUT_4[28568] = 32'b00000000000000000110011001110111;
assign LUT_4[28569] = 32'b11111111111111111111100101101111;
assign LUT_4[28570] = 32'b00000000000000000101110100011011;
assign LUT_4[28571] = 32'b11111111111111111111000000010011;
assign LUT_4[28572] = 32'b00000000000000000011011010010011;
assign LUT_4[28573] = 32'b11111111111111111100100110001011;
assign LUT_4[28574] = 32'b00000000000000000010110100110111;
assign LUT_4[28575] = 32'b11111111111111111100000000101111;
assign LUT_4[28576] = 32'b00000000000000001101110110111011;
assign LUT_4[28577] = 32'b00000000000000000111000010110011;
assign LUT_4[28578] = 32'b00000000000000001101010001011111;
assign LUT_4[28579] = 32'b00000000000000000110011101010111;
assign LUT_4[28580] = 32'b00000000000000001010110111010111;
assign LUT_4[28581] = 32'b00000000000000000100000011001111;
assign LUT_4[28582] = 32'b00000000000000001010010001111011;
assign LUT_4[28583] = 32'b00000000000000000011011101110011;
assign LUT_4[28584] = 32'b00000000000000000111000011010000;
assign LUT_4[28585] = 32'b00000000000000000000001111001000;
assign LUT_4[28586] = 32'b00000000000000000110011101110100;
assign LUT_4[28587] = 32'b11111111111111111111101001101100;
assign LUT_4[28588] = 32'b00000000000000000100000011101100;
assign LUT_4[28589] = 32'b11111111111111111101001111100100;
assign LUT_4[28590] = 32'b00000000000000000011011110010000;
assign LUT_4[28591] = 32'b11111111111111111100101010001000;
assign LUT_4[28592] = 32'b00000000000000001011101000101001;
assign LUT_4[28593] = 32'b00000000000000000100110100100001;
assign LUT_4[28594] = 32'b00000000000000001011000011001101;
assign LUT_4[28595] = 32'b00000000000000000100001111000101;
assign LUT_4[28596] = 32'b00000000000000001000101001000101;
assign LUT_4[28597] = 32'b00000000000000000001110100111101;
assign LUT_4[28598] = 32'b00000000000000001000000011101001;
assign LUT_4[28599] = 32'b00000000000000000001001111100001;
assign LUT_4[28600] = 32'b00000000000000000100110100111110;
assign LUT_4[28601] = 32'b11111111111111111110000000110110;
assign LUT_4[28602] = 32'b00000000000000000100001111100010;
assign LUT_4[28603] = 32'b11111111111111111101011011011010;
assign LUT_4[28604] = 32'b00000000000000000001110101011010;
assign LUT_4[28605] = 32'b11111111111111111011000001010010;
assign LUT_4[28606] = 32'b00000000000000000001001111111110;
assign LUT_4[28607] = 32'b11111111111111111010011011110110;
assign LUT_4[28608] = 32'b00000000000000010000110011001000;
assign LUT_4[28609] = 32'b00000000000000001001111111000000;
assign LUT_4[28610] = 32'b00000000000000010000001101101100;
assign LUT_4[28611] = 32'b00000000000000001001011001100100;
assign LUT_4[28612] = 32'b00000000000000001101110011100100;
assign LUT_4[28613] = 32'b00000000000000000110111111011100;
assign LUT_4[28614] = 32'b00000000000000001101001110001000;
assign LUT_4[28615] = 32'b00000000000000000110011010000000;
assign LUT_4[28616] = 32'b00000000000000001001111111011101;
assign LUT_4[28617] = 32'b00000000000000000011001011010101;
assign LUT_4[28618] = 32'b00000000000000001001011010000001;
assign LUT_4[28619] = 32'b00000000000000000010100101111001;
assign LUT_4[28620] = 32'b00000000000000000110111111111001;
assign LUT_4[28621] = 32'b00000000000000000000001011110001;
assign LUT_4[28622] = 32'b00000000000000000110011010011101;
assign LUT_4[28623] = 32'b11111111111111111111100110010101;
assign LUT_4[28624] = 32'b00000000000000001110100100110110;
assign LUT_4[28625] = 32'b00000000000000000111110000101110;
assign LUT_4[28626] = 32'b00000000000000001101111111011010;
assign LUT_4[28627] = 32'b00000000000000000111001011010010;
assign LUT_4[28628] = 32'b00000000000000001011100101010010;
assign LUT_4[28629] = 32'b00000000000000000100110001001010;
assign LUT_4[28630] = 32'b00000000000000001010111111110110;
assign LUT_4[28631] = 32'b00000000000000000100001011101110;
assign LUT_4[28632] = 32'b00000000000000000111110001001011;
assign LUT_4[28633] = 32'b00000000000000000000111101000011;
assign LUT_4[28634] = 32'b00000000000000000111001011101111;
assign LUT_4[28635] = 32'b00000000000000000000010111100111;
assign LUT_4[28636] = 32'b00000000000000000100110001100111;
assign LUT_4[28637] = 32'b11111111111111111101111101011111;
assign LUT_4[28638] = 32'b00000000000000000100001100001011;
assign LUT_4[28639] = 32'b11111111111111111101011000000011;
assign LUT_4[28640] = 32'b00000000000000001111001110001111;
assign LUT_4[28641] = 32'b00000000000000001000011010000111;
assign LUT_4[28642] = 32'b00000000000000001110101000110011;
assign LUT_4[28643] = 32'b00000000000000000111110100101011;
assign LUT_4[28644] = 32'b00000000000000001100001110101011;
assign LUT_4[28645] = 32'b00000000000000000101011010100011;
assign LUT_4[28646] = 32'b00000000000000001011101001001111;
assign LUT_4[28647] = 32'b00000000000000000100110101000111;
assign LUT_4[28648] = 32'b00000000000000001000011010100100;
assign LUT_4[28649] = 32'b00000000000000000001100110011100;
assign LUT_4[28650] = 32'b00000000000000000111110101001000;
assign LUT_4[28651] = 32'b00000000000000000001000001000000;
assign LUT_4[28652] = 32'b00000000000000000101011011000000;
assign LUT_4[28653] = 32'b11111111111111111110100110111000;
assign LUT_4[28654] = 32'b00000000000000000100110101100100;
assign LUT_4[28655] = 32'b11111111111111111110000001011100;
assign LUT_4[28656] = 32'b00000000000000001100111111111101;
assign LUT_4[28657] = 32'b00000000000000000110001011110101;
assign LUT_4[28658] = 32'b00000000000000001100011010100001;
assign LUT_4[28659] = 32'b00000000000000000101100110011001;
assign LUT_4[28660] = 32'b00000000000000001010000000011001;
assign LUT_4[28661] = 32'b00000000000000000011001100010001;
assign LUT_4[28662] = 32'b00000000000000001001011010111101;
assign LUT_4[28663] = 32'b00000000000000000010100110110101;
assign LUT_4[28664] = 32'b00000000000000000110001100010010;
assign LUT_4[28665] = 32'b11111111111111111111011000001010;
assign LUT_4[28666] = 32'b00000000000000000101100110110110;
assign LUT_4[28667] = 32'b11111111111111111110110010101110;
assign LUT_4[28668] = 32'b00000000000000000011001100101110;
assign LUT_4[28669] = 32'b11111111111111111100011000100110;
assign LUT_4[28670] = 32'b00000000000000000010100111010010;
assign LUT_4[28671] = 32'b11111111111111111011110011001010;
assign LUT_4[28672] = 32'b00000000000000000111111100001001;
assign LUT_4[28673] = 32'b00000000000000000001001000000001;
assign LUT_4[28674] = 32'b00000000000000000111010110101101;
assign LUT_4[28675] = 32'b00000000000000000000100010100101;
assign LUT_4[28676] = 32'b00000000000000000100111100100101;
assign LUT_4[28677] = 32'b11111111111111111110001000011101;
assign LUT_4[28678] = 32'b00000000000000000100010111001001;
assign LUT_4[28679] = 32'b11111111111111111101100011000001;
assign LUT_4[28680] = 32'b00000000000000000001001000011110;
assign LUT_4[28681] = 32'b11111111111111111010010100010110;
assign LUT_4[28682] = 32'b00000000000000000000100011000010;
assign LUT_4[28683] = 32'b11111111111111111001101110111010;
assign LUT_4[28684] = 32'b11111111111111111110001000111010;
assign LUT_4[28685] = 32'b11111111111111110111010100110010;
assign LUT_4[28686] = 32'b11111111111111111101100011011110;
assign LUT_4[28687] = 32'b11111111111111110110101111010110;
assign LUT_4[28688] = 32'b00000000000000000101101101110111;
assign LUT_4[28689] = 32'b11111111111111111110111001101111;
assign LUT_4[28690] = 32'b00000000000000000101001000011011;
assign LUT_4[28691] = 32'b11111111111111111110010100010011;
assign LUT_4[28692] = 32'b00000000000000000010101110010011;
assign LUT_4[28693] = 32'b11111111111111111011111010001011;
assign LUT_4[28694] = 32'b00000000000000000010001000110111;
assign LUT_4[28695] = 32'b11111111111111111011010100101111;
assign LUT_4[28696] = 32'b11111111111111111110111010001100;
assign LUT_4[28697] = 32'b11111111111111111000000110000100;
assign LUT_4[28698] = 32'b11111111111111111110010100110000;
assign LUT_4[28699] = 32'b11111111111111110111100000101000;
assign LUT_4[28700] = 32'b11111111111111111011111010101000;
assign LUT_4[28701] = 32'b11111111111111110101000110100000;
assign LUT_4[28702] = 32'b11111111111111111011010101001100;
assign LUT_4[28703] = 32'b11111111111111110100100001000100;
assign LUT_4[28704] = 32'b00000000000000000110010111010000;
assign LUT_4[28705] = 32'b11111111111111111111100011001000;
assign LUT_4[28706] = 32'b00000000000000000101110001110100;
assign LUT_4[28707] = 32'b11111111111111111110111101101100;
assign LUT_4[28708] = 32'b00000000000000000011010111101100;
assign LUT_4[28709] = 32'b11111111111111111100100011100100;
assign LUT_4[28710] = 32'b00000000000000000010110010010000;
assign LUT_4[28711] = 32'b11111111111111111011111110001000;
assign LUT_4[28712] = 32'b11111111111111111111100011100101;
assign LUT_4[28713] = 32'b11111111111111111000101111011101;
assign LUT_4[28714] = 32'b11111111111111111110111110001001;
assign LUT_4[28715] = 32'b11111111111111111000001010000001;
assign LUT_4[28716] = 32'b11111111111111111100100100000001;
assign LUT_4[28717] = 32'b11111111111111110101101111111001;
assign LUT_4[28718] = 32'b11111111111111111011111110100101;
assign LUT_4[28719] = 32'b11111111111111110101001010011101;
assign LUT_4[28720] = 32'b00000000000000000100001000111110;
assign LUT_4[28721] = 32'b11111111111111111101010100110110;
assign LUT_4[28722] = 32'b00000000000000000011100011100010;
assign LUT_4[28723] = 32'b11111111111111111100101111011010;
assign LUT_4[28724] = 32'b00000000000000000001001001011010;
assign LUT_4[28725] = 32'b11111111111111111010010101010010;
assign LUT_4[28726] = 32'b00000000000000000000100011111110;
assign LUT_4[28727] = 32'b11111111111111111001101111110110;
assign LUT_4[28728] = 32'b11111111111111111101010101010011;
assign LUT_4[28729] = 32'b11111111111111110110100001001011;
assign LUT_4[28730] = 32'b11111111111111111100101111110111;
assign LUT_4[28731] = 32'b11111111111111110101111011101111;
assign LUT_4[28732] = 32'b11111111111111111010010101101111;
assign LUT_4[28733] = 32'b11111111111111110011100001100111;
assign LUT_4[28734] = 32'b11111111111111111001110000010011;
assign LUT_4[28735] = 32'b11111111111111110010111100001011;
assign LUT_4[28736] = 32'b00000000000000001001010011011101;
assign LUT_4[28737] = 32'b00000000000000000010011111010101;
assign LUT_4[28738] = 32'b00000000000000001000101110000001;
assign LUT_4[28739] = 32'b00000000000000000001111001111001;
assign LUT_4[28740] = 32'b00000000000000000110010011111001;
assign LUT_4[28741] = 32'b11111111111111111111011111110001;
assign LUT_4[28742] = 32'b00000000000000000101101110011101;
assign LUT_4[28743] = 32'b11111111111111111110111010010101;
assign LUT_4[28744] = 32'b00000000000000000010011111110010;
assign LUT_4[28745] = 32'b11111111111111111011101011101010;
assign LUT_4[28746] = 32'b00000000000000000001111010010110;
assign LUT_4[28747] = 32'b11111111111111111011000110001110;
assign LUT_4[28748] = 32'b11111111111111111111100000001110;
assign LUT_4[28749] = 32'b11111111111111111000101100000110;
assign LUT_4[28750] = 32'b11111111111111111110111010110010;
assign LUT_4[28751] = 32'b11111111111111111000000110101010;
assign LUT_4[28752] = 32'b00000000000000000111000101001011;
assign LUT_4[28753] = 32'b00000000000000000000010001000011;
assign LUT_4[28754] = 32'b00000000000000000110011111101111;
assign LUT_4[28755] = 32'b11111111111111111111101011100111;
assign LUT_4[28756] = 32'b00000000000000000100000101100111;
assign LUT_4[28757] = 32'b11111111111111111101010001011111;
assign LUT_4[28758] = 32'b00000000000000000011100000001011;
assign LUT_4[28759] = 32'b11111111111111111100101100000011;
assign LUT_4[28760] = 32'b00000000000000000000010001100000;
assign LUT_4[28761] = 32'b11111111111111111001011101011000;
assign LUT_4[28762] = 32'b11111111111111111111101100000100;
assign LUT_4[28763] = 32'b11111111111111111000110111111100;
assign LUT_4[28764] = 32'b11111111111111111101010001111100;
assign LUT_4[28765] = 32'b11111111111111110110011101110100;
assign LUT_4[28766] = 32'b11111111111111111100101100100000;
assign LUT_4[28767] = 32'b11111111111111110101111000011000;
assign LUT_4[28768] = 32'b00000000000000000111101110100100;
assign LUT_4[28769] = 32'b00000000000000000000111010011100;
assign LUT_4[28770] = 32'b00000000000000000111001001001000;
assign LUT_4[28771] = 32'b00000000000000000000010101000000;
assign LUT_4[28772] = 32'b00000000000000000100101111000000;
assign LUT_4[28773] = 32'b11111111111111111101111010111000;
assign LUT_4[28774] = 32'b00000000000000000100001001100100;
assign LUT_4[28775] = 32'b11111111111111111101010101011100;
assign LUT_4[28776] = 32'b00000000000000000000111010111001;
assign LUT_4[28777] = 32'b11111111111111111010000110110001;
assign LUT_4[28778] = 32'b00000000000000000000010101011101;
assign LUT_4[28779] = 32'b11111111111111111001100001010101;
assign LUT_4[28780] = 32'b11111111111111111101111011010101;
assign LUT_4[28781] = 32'b11111111111111110111000111001101;
assign LUT_4[28782] = 32'b11111111111111111101010101111001;
assign LUT_4[28783] = 32'b11111111111111110110100001110001;
assign LUT_4[28784] = 32'b00000000000000000101100000010010;
assign LUT_4[28785] = 32'b11111111111111111110101100001010;
assign LUT_4[28786] = 32'b00000000000000000100111010110110;
assign LUT_4[28787] = 32'b11111111111111111110000110101110;
assign LUT_4[28788] = 32'b00000000000000000010100000101110;
assign LUT_4[28789] = 32'b11111111111111111011101100100110;
assign LUT_4[28790] = 32'b00000000000000000001111011010010;
assign LUT_4[28791] = 32'b11111111111111111011000111001010;
assign LUT_4[28792] = 32'b11111111111111111110101100100111;
assign LUT_4[28793] = 32'b11111111111111110111111000011111;
assign LUT_4[28794] = 32'b11111111111111111110000111001011;
assign LUT_4[28795] = 32'b11111111111111110111010011000011;
assign LUT_4[28796] = 32'b11111111111111111011101101000011;
assign LUT_4[28797] = 32'b11111111111111110100111000111011;
assign LUT_4[28798] = 32'b11111111111111111011000111100111;
assign LUT_4[28799] = 32'b11111111111111110100010011011111;
assign LUT_4[28800] = 32'b00000000000000001010100010010001;
assign LUT_4[28801] = 32'b00000000000000000011101110001001;
assign LUT_4[28802] = 32'b00000000000000001001111100110101;
assign LUT_4[28803] = 32'b00000000000000000011001000101101;
assign LUT_4[28804] = 32'b00000000000000000111100010101101;
assign LUT_4[28805] = 32'b00000000000000000000101110100101;
assign LUT_4[28806] = 32'b00000000000000000110111101010001;
assign LUT_4[28807] = 32'b00000000000000000000001001001001;
assign LUT_4[28808] = 32'b00000000000000000011101110100110;
assign LUT_4[28809] = 32'b11111111111111111100111010011110;
assign LUT_4[28810] = 32'b00000000000000000011001001001010;
assign LUT_4[28811] = 32'b11111111111111111100010101000010;
assign LUT_4[28812] = 32'b00000000000000000000101111000010;
assign LUT_4[28813] = 32'b11111111111111111001111010111010;
assign LUT_4[28814] = 32'b00000000000000000000001001100110;
assign LUT_4[28815] = 32'b11111111111111111001010101011110;
assign LUT_4[28816] = 32'b00000000000000001000010011111111;
assign LUT_4[28817] = 32'b00000000000000000001011111110111;
assign LUT_4[28818] = 32'b00000000000000000111101110100011;
assign LUT_4[28819] = 32'b00000000000000000000111010011011;
assign LUT_4[28820] = 32'b00000000000000000101010100011011;
assign LUT_4[28821] = 32'b11111111111111111110100000010011;
assign LUT_4[28822] = 32'b00000000000000000100101110111111;
assign LUT_4[28823] = 32'b11111111111111111101111010110111;
assign LUT_4[28824] = 32'b00000000000000000001100000010100;
assign LUT_4[28825] = 32'b11111111111111111010101100001100;
assign LUT_4[28826] = 32'b00000000000000000000111010111000;
assign LUT_4[28827] = 32'b11111111111111111010000110110000;
assign LUT_4[28828] = 32'b11111111111111111110100000110000;
assign LUT_4[28829] = 32'b11111111111111110111101100101000;
assign LUT_4[28830] = 32'b11111111111111111101111011010100;
assign LUT_4[28831] = 32'b11111111111111110111000111001100;
assign LUT_4[28832] = 32'b00000000000000001000111101011000;
assign LUT_4[28833] = 32'b00000000000000000010001001010000;
assign LUT_4[28834] = 32'b00000000000000001000010111111100;
assign LUT_4[28835] = 32'b00000000000000000001100011110100;
assign LUT_4[28836] = 32'b00000000000000000101111101110100;
assign LUT_4[28837] = 32'b11111111111111111111001001101100;
assign LUT_4[28838] = 32'b00000000000000000101011000011000;
assign LUT_4[28839] = 32'b11111111111111111110100100010000;
assign LUT_4[28840] = 32'b00000000000000000010001001101101;
assign LUT_4[28841] = 32'b11111111111111111011010101100101;
assign LUT_4[28842] = 32'b00000000000000000001100100010001;
assign LUT_4[28843] = 32'b11111111111111111010110000001001;
assign LUT_4[28844] = 32'b11111111111111111111001010001001;
assign LUT_4[28845] = 32'b11111111111111111000010110000001;
assign LUT_4[28846] = 32'b11111111111111111110100100101101;
assign LUT_4[28847] = 32'b11111111111111110111110000100101;
assign LUT_4[28848] = 32'b00000000000000000110101111000110;
assign LUT_4[28849] = 32'b11111111111111111111111010111110;
assign LUT_4[28850] = 32'b00000000000000000110001001101010;
assign LUT_4[28851] = 32'b11111111111111111111010101100010;
assign LUT_4[28852] = 32'b00000000000000000011101111100010;
assign LUT_4[28853] = 32'b11111111111111111100111011011010;
assign LUT_4[28854] = 32'b00000000000000000011001010000110;
assign LUT_4[28855] = 32'b11111111111111111100010101111110;
assign LUT_4[28856] = 32'b11111111111111111111111011011011;
assign LUT_4[28857] = 32'b11111111111111111001000111010011;
assign LUT_4[28858] = 32'b11111111111111111111010101111111;
assign LUT_4[28859] = 32'b11111111111111111000100001110111;
assign LUT_4[28860] = 32'b11111111111111111100111011110111;
assign LUT_4[28861] = 32'b11111111111111110110000111101111;
assign LUT_4[28862] = 32'b11111111111111111100010110011011;
assign LUT_4[28863] = 32'b11111111111111110101100010010011;
assign LUT_4[28864] = 32'b00000000000000001011111001100101;
assign LUT_4[28865] = 32'b00000000000000000101000101011101;
assign LUT_4[28866] = 32'b00000000000000001011010100001001;
assign LUT_4[28867] = 32'b00000000000000000100100000000001;
assign LUT_4[28868] = 32'b00000000000000001000111010000001;
assign LUT_4[28869] = 32'b00000000000000000010000101111001;
assign LUT_4[28870] = 32'b00000000000000001000010100100101;
assign LUT_4[28871] = 32'b00000000000000000001100000011101;
assign LUT_4[28872] = 32'b00000000000000000101000101111010;
assign LUT_4[28873] = 32'b11111111111111111110010001110010;
assign LUT_4[28874] = 32'b00000000000000000100100000011110;
assign LUT_4[28875] = 32'b11111111111111111101101100010110;
assign LUT_4[28876] = 32'b00000000000000000010000110010110;
assign LUT_4[28877] = 32'b11111111111111111011010010001110;
assign LUT_4[28878] = 32'b00000000000000000001100000111010;
assign LUT_4[28879] = 32'b11111111111111111010101100110010;
assign LUT_4[28880] = 32'b00000000000000001001101011010011;
assign LUT_4[28881] = 32'b00000000000000000010110111001011;
assign LUT_4[28882] = 32'b00000000000000001001000101110111;
assign LUT_4[28883] = 32'b00000000000000000010010001101111;
assign LUT_4[28884] = 32'b00000000000000000110101011101111;
assign LUT_4[28885] = 32'b11111111111111111111110111100111;
assign LUT_4[28886] = 32'b00000000000000000110000110010011;
assign LUT_4[28887] = 32'b11111111111111111111010010001011;
assign LUT_4[28888] = 32'b00000000000000000010110111101000;
assign LUT_4[28889] = 32'b11111111111111111100000011100000;
assign LUT_4[28890] = 32'b00000000000000000010010010001100;
assign LUT_4[28891] = 32'b11111111111111111011011110000100;
assign LUT_4[28892] = 32'b11111111111111111111111000000100;
assign LUT_4[28893] = 32'b11111111111111111001000011111100;
assign LUT_4[28894] = 32'b11111111111111111111010010101000;
assign LUT_4[28895] = 32'b11111111111111111000011110100000;
assign LUT_4[28896] = 32'b00000000000000001010010100101100;
assign LUT_4[28897] = 32'b00000000000000000011100000100100;
assign LUT_4[28898] = 32'b00000000000000001001101111010000;
assign LUT_4[28899] = 32'b00000000000000000010111011001000;
assign LUT_4[28900] = 32'b00000000000000000111010101001000;
assign LUT_4[28901] = 32'b00000000000000000000100001000000;
assign LUT_4[28902] = 32'b00000000000000000110101111101100;
assign LUT_4[28903] = 32'b11111111111111111111111011100100;
assign LUT_4[28904] = 32'b00000000000000000011100001000001;
assign LUT_4[28905] = 32'b11111111111111111100101100111001;
assign LUT_4[28906] = 32'b00000000000000000010111011100101;
assign LUT_4[28907] = 32'b11111111111111111100000111011101;
assign LUT_4[28908] = 32'b00000000000000000000100001011101;
assign LUT_4[28909] = 32'b11111111111111111001101101010101;
assign LUT_4[28910] = 32'b11111111111111111111111100000001;
assign LUT_4[28911] = 32'b11111111111111111001000111111001;
assign LUT_4[28912] = 32'b00000000000000001000000110011010;
assign LUT_4[28913] = 32'b00000000000000000001010010010010;
assign LUT_4[28914] = 32'b00000000000000000111100000111110;
assign LUT_4[28915] = 32'b00000000000000000000101100110110;
assign LUT_4[28916] = 32'b00000000000000000101000110110110;
assign LUT_4[28917] = 32'b11111111111111111110010010101110;
assign LUT_4[28918] = 32'b00000000000000000100100001011010;
assign LUT_4[28919] = 32'b11111111111111111101101101010010;
assign LUT_4[28920] = 32'b00000000000000000001010010101111;
assign LUT_4[28921] = 32'b11111111111111111010011110100111;
assign LUT_4[28922] = 32'b00000000000000000000101101010011;
assign LUT_4[28923] = 32'b11111111111111111001111001001011;
assign LUT_4[28924] = 32'b11111111111111111110010011001011;
assign LUT_4[28925] = 32'b11111111111111110111011111000011;
assign LUT_4[28926] = 32'b11111111111111111101101101101111;
assign LUT_4[28927] = 32'b11111111111111110110111001100111;
assign LUT_4[28928] = 32'b00000000000000001100110111101100;
assign LUT_4[28929] = 32'b00000000000000000110000011100100;
assign LUT_4[28930] = 32'b00000000000000001100010010010000;
assign LUT_4[28931] = 32'b00000000000000000101011110001000;
assign LUT_4[28932] = 32'b00000000000000001001111000001000;
assign LUT_4[28933] = 32'b00000000000000000011000100000000;
assign LUT_4[28934] = 32'b00000000000000001001010010101100;
assign LUT_4[28935] = 32'b00000000000000000010011110100100;
assign LUT_4[28936] = 32'b00000000000000000110000100000001;
assign LUT_4[28937] = 32'b11111111111111111111001111111001;
assign LUT_4[28938] = 32'b00000000000000000101011110100101;
assign LUT_4[28939] = 32'b11111111111111111110101010011101;
assign LUT_4[28940] = 32'b00000000000000000011000100011101;
assign LUT_4[28941] = 32'b11111111111111111100010000010101;
assign LUT_4[28942] = 32'b00000000000000000010011111000001;
assign LUT_4[28943] = 32'b11111111111111111011101010111001;
assign LUT_4[28944] = 32'b00000000000000001010101001011010;
assign LUT_4[28945] = 32'b00000000000000000011110101010010;
assign LUT_4[28946] = 32'b00000000000000001010000011111110;
assign LUT_4[28947] = 32'b00000000000000000011001111110110;
assign LUT_4[28948] = 32'b00000000000000000111101001110110;
assign LUT_4[28949] = 32'b00000000000000000000110101101110;
assign LUT_4[28950] = 32'b00000000000000000111000100011010;
assign LUT_4[28951] = 32'b00000000000000000000010000010010;
assign LUT_4[28952] = 32'b00000000000000000011110101101111;
assign LUT_4[28953] = 32'b11111111111111111101000001100111;
assign LUT_4[28954] = 32'b00000000000000000011010000010011;
assign LUT_4[28955] = 32'b11111111111111111100011100001011;
assign LUT_4[28956] = 32'b00000000000000000000110110001011;
assign LUT_4[28957] = 32'b11111111111111111010000010000011;
assign LUT_4[28958] = 32'b00000000000000000000010000101111;
assign LUT_4[28959] = 32'b11111111111111111001011100100111;
assign LUT_4[28960] = 32'b00000000000000001011010010110011;
assign LUT_4[28961] = 32'b00000000000000000100011110101011;
assign LUT_4[28962] = 32'b00000000000000001010101101010111;
assign LUT_4[28963] = 32'b00000000000000000011111001001111;
assign LUT_4[28964] = 32'b00000000000000001000010011001111;
assign LUT_4[28965] = 32'b00000000000000000001011111000111;
assign LUT_4[28966] = 32'b00000000000000000111101101110011;
assign LUT_4[28967] = 32'b00000000000000000000111001101011;
assign LUT_4[28968] = 32'b00000000000000000100011111001000;
assign LUT_4[28969] = 32'b11111111111111111101101011000000;
assign LUT_4[28970] = 32'b00000000000000000011111001101100;
assign LUT_4[28971] = 32'b11111111111111111101000101100100;
assign LUT_4[28972] = 32'b00000000000000000001011111100100;
assign LUT_4[28973] = 32'b11111111111111111010101011011100;
assign LUT_4[28974] = 32'b00000000000000000000111010001000;
assign LUT_4[28975] = 32'b11111111111111111010000110000000;
assign LUT_4[28976] = 32'b00000000000000001001000100100001;
assign LUT_4[28977] = 32'b00000000000000000010010000011001;
assign LUT_4[28978] = 32'b00000000000000001000011111000101;
assign LUT_4[28979] = 32'b00000000000000000001101010111101;
assign LUT_4[28980] = 32'b00000000000000000110000100111101;
assign LUT_4[28981] = 32'b11111111111111111111010000110101;
assign LUT_4[28982] = 32'b00000000000000000101011111100001;
assign LUT_4[28983] = 32'b11111111111111111110101011011001;
assign LUT_4[28984] = 32'b00000000000000000010010000110110;
assign LUT_4[28985] = 32'b11111111111111111011011100101110;
assign LUT_4[28986] = 32'b00000000000000000001101011011010;
assign LUT_4[28987] = 32'b11111111111111111010110111010010;
assign LUT_4[28988] = 32'b11111111111111111111010001010010;
assign LUT_4[28989] = 32'b11111111111111111000011101001010;
assign LUT_4[28990] = 32'b11111111111111111110101011110110;
assign LUT_4[28991] = 32'b11111111111111110111110111101110;
assign LUT_4[28992] = 32'b00000000000000001110001111000000;
assign LUT_4[28993] = 32'b00000000000000000111011010111000;
assign LUT_4[28994] = 32'b00000000000000001101101001100100;
assign LUT_4[28995] = 32'b00000000000000000110110101011100;
assign LUT_4[28996] = 32'b00000000000000001011001111011100;
assign LUT_4[28997] = 32'b00000000000000000100011011010100;
assign LUT_4[28998] = 32'b00000000000000001010101010000000;
assign LUT_4[28999] = 32'b00000000000000000011110101111000;
assign LUT_4[29000] = 32'b00000000000000000111011011010101;
assign LUT_4[29001] = 32'b00000000000000000000100111001101;
assign LUT_4[29002] = 32'b00000000000000000110110101111001;
assign LUT_4[29003] = 32'b00000000000000000000000001110001;
assign LUT_4[29004] = 32'b00000000000000000100011011110001;
assign LUT_4[29005] = 32'b11111111111111111101100111101001;
assign LUT_4[29006] = 32'b00000000000000000011110110010101;
assign LUT_4[29007] = 32'b11111111111111111101000010001101;
assign LUT_4[29008] = 32'b00000000000000001100000000101110;
assign LUT_4[29009] = 32'b00000000000000000101001100100110;
assign LUT_4[29010] = 32'b00000000000000001011011011010010;
assign LUT_4[29011] = 32'b00000000000000000100100111001010;
assign LUT_4[29012] = 32'b00000000000000001001000001001010;
assign LUT_4[29013] = 32'b00000000000000000010001101000010;
assign LUT_4[29014] = 32'b00000000000000001000011011101110;
assign LUT_4[29015] = 32'b00000000000000000001100111100110;
assign LUT_4[29016] = 32'b00000000000000000101001101000011;
assign LUT_4[29017] = 32'b11111111111111111110011000111011;
assign LUT_4[29018] = 32'b00000000000000000100100111100111;
assign LUT_4[29019] = 32'b11111111111111111101110011011111;
assign LUT_4[29020] = 32'b00000000000000000010001101011111;
assign LUT_4[29021] = 32'b11111111111111111011011001010111;
assign LUT_4[29022] = 32'b00000000000000000001101000000011;
assign LUT_4[29023] = 32'b11111111111111111010110011111011;
assign LUT_4[29024] = 32'b00000000000000001100101010000111;
assign LUT_4[29025] = 32'b00000000000000000101110101111111;
assign LUT_4[29026] = 32'b00000000000000001100000100101011;
assign LUT_4[29027] = 32'b00000000000000000101010000100011;
assign LUT_4[29028] = 32'b00000000000000001001101010100011;
assign LUT_4[29029] = 32'b00000000000000000010110110011011;
assign LUT_4[29030] = 32'b00000000000000001001000101000111;
assign LUT_4[29031] = 32'b00000000000000000010010000111111;
assign LUT_4[29032] = 32'b00000000000000000101110110011100;
assign LUT_4[29033] = 32'b11111111111111111111000010010100;
assign LUT_4[29034] = 32'b00000000000000000101010001000000;
assign LUT_4[29035] = 32'b11111111111111111110011100111000;
assign LUT_4[29036] = 32'b00000000000000000010110110111000;
assign LUT_4[29037] = 32'b11111111111111111100000010110000;
assign LUT_4[29038] = 32'b00000000000000000010010001011100;
assign LUT_4[29039] = 32'b11111111111111111011011101010100;
assign LUT_4[29040] = 32'b00000000000000001010011011110101;
assign LUT_4[29041] = 32'b00000000000000000011100111101101;
assign LUT_4[29042] = 32'b00000000000000001001110110011001;
assign LUT_4[29043] = 32'b00000000000000000011000010010001;
assign LUT_4[29044] = 32'b00000000000000000111011100010001;
assign LUT_4[29045] = 32'b00000000000000000000101000001001;
assign LUT_4[29046] = 32'b00000000000000000110110110110101;
assign LUT_4[29047] = 32'b00000000000000000000000010101101;
assign LUT_4[29048] = 32'b00000000000000000011101000001010;
assign LUT_4[29049] = 32'b11111111111111111100110100000010;
assign LUT_4[29050] = 32'b00000000000000000011000010101110;
assign LUT_4[29051] = 32'b11111111111111111100001110100110;
assign LUT_4[29052] = 32'b00000000000000000000101000100110;
assign LUT_4[29053] = 32'b11111111111111111001110100011110;
assign LUT_4[29054] = 32'b00000000000000000000000011001010;
assign LUT_4[29055] = 32'b11111111111111111001001111000010;
assign LUT_4[29056] = 32'b00000000000000001111011101110100;
assign LUT_4[29057] = 32'b00000000000000001000101001101100;
assign LUT_4[29058] = 32'b00000000000000001110111000011000;
assign LUT_4[29059] = 32'b00000000000000001000000100010000;
assign LUT_4[29060] = 32'b00000000000000001100011110010000;
assign LUT_4[29061] = 32'b00000000000000000101101010001000;
assign LUT_4[29062] = 32'b00000000000000001011111000110100;
assign LUT_4[29063] = 32'b00000000000000000101000100101100;
assign LUT_4[29064] = 32'b00000000000000001000101010001001;
assign LUT_4[29065] = 32'b00000000000000000001110110000001;
assign LUT_4[29066] = 32'b00000000000000001000000100101101;
assign LUT_4[29067] = 32'b00000000000000000001010000100101;
assign LUT_4[29068] = 32'b00000000000000000101101010100101;
assign LUT_4[29069] = 32'b11111111111111111110110110011101;
assign LUT_4[29070] = 32'b00000000000000000101000101001001;
assign LUT_4[29071] = 32'b11111111111111111110010001000001;
assign LUT_4[29072] = 32'b00000000000000001101001111100010;
assign LUT_4[29073] = 32'b00000000000000000110011011011010;
assign LUT_4[29074] = 32'b00000000000000001100101010000110;
assign LUT_4[29075] = 32'b00000000000000000101110101111110;
assign LUT_4[29076] = 32'b00000000000000001010001111111110;
assign LUT_4[29077] = 32'b00000000000000000011011011110110;
assign LUT_4[29078] = 32'b00000000000000001001101010100010;
assign LUT_4[29079] = 32'b00000000000000000010110110011010;
assign LUT_4[29080] = 32'b00000000000000000110011011110111;
assign LUT_4[29081] = 32'b11111111111111111111100111101111;
assign LUT_4[29082] = 32'b00000000000000000101110110011011;
assign LUT_4[29083] = 32'b11111111111111111111000010010011;
assign LUT_4[29084] = 32'b00000000000000000011011100010011;
assign LUT_4[29085] = 32'b11111111111111111100101000001011;
assign LUT_4[29086] = 32'b00000000000000000010110110110111;
assign LUT_4[29087] = 32'b11111111111111111100000010101111;
assign LUT_4[29088] = 32'b00000000000000001101111000111011;
assign LUT_4[29089] = 32'b00000000000000000111000100110011;
assign LUT_4[29090] = 32'b00000000000000001101010011011111;
assign LUT_4[29091] = 32'b00000000000000000110011111010111;
assign LUT_4[29092] = 32'b00000000000000001010111001010111;
assign LUT_4[29093] = 32'b00000000000000000100000101001111;
assign LUT_4[29094] = 32'b00000000000000001010010011111011;
assign LUT_4[29095] = 32'b00000000000000000011011111110011;
assign LUT_4[29096] = 32'b00000000000000000111000101010000;
assign LUT_4[29097] = 32'b00000000000000000000010001001000;
assign LUT_4[29098] = 32'b00000000000000000110011111110100;
assign LUT_4[29099] = 32'b11111111111111111111101011101100;
assign LUT_4[29100] = 32'b00000000000000000100000101101100;
assign LUT_4[29101] = 32'b11111111111111111101010001100100;
assign LUT_4[29102] = 32'b00000000000000000011100000010000;
assign LUT_4[29103] = 32'b11111111111111111100101100001000;
assign LUT_4[29104] = 32'b00000000000000001011101010101001;
assign LUT_4[29105] = 32'b00000000000000000100110110100001;
assign LUT_4[29106] = 32'b00000000000000001011000101001101;
assign LUT_4[29107] = 32'b00000000000000000100010001000101;
assign LUT_4[29108] = 32'b00000000000000001000101011000101;
assign LUT_4[29109] = 32'b00000000000000000001110110111101;
assign LUT_4[29110] = 32'b00000000000000001000000101101001;
assign LUT_4[29111] = 32'b00000000000000000001010001100001;
assign LUT_4[29112] = 32'b00000000000000000100110110111110;
assign LUT_4[29113] = 32'b11111111111111111110000010110110;
assign LUT_4[29114] = 32'b00000000000000000100010001100010;
assign LUT_4[29115] = 32'b11111111111111111101011101011010;
assign LUT_4[29116] = 32'b00000000000000000001110111011010;
assign LUT_4[29117] = 32'b11111111111111111011000011010010;
assign LUT_4[29118] = 32'b00000000000000000001010001111110;
assign LUT_4[29119] = 32'b11111111111111111010011101110110;
assign LUT_4[29120] = 32'b00000000000000010000110101001000;
assign LUT_4[29121] = 32'b00000000000000001010000001000000;
assign LUT_4[29122] = 32'b00000000000000010000001111101100;
assign LUT_4[29123] = 32'b00000000000000001001011011100100;
assign LUT_4[29124] = 32'b00000000000000001101110101100100;
assign LUT_4[29125] = 32'b00000000000000000111000001011100;
assign LUT_4[29126] = 32'b00000000000000001101010000001000;
assign LUT_4[29127] = 32'b00000000000000000110011100000000;
assign LUT_4[29128] = 32'b00000000000000001010000001011101;
assign LUT_4[29129] = 32'b00000000000000000011001101010101;
assign LUT_4[29130] = 32'b00000000000000001001011100000001;
assign LUT_4[29131] = 32'b00000000000000000010100111111001;
assign LUT_4[29132] = 32'b00000000000000000111000001111001;
assign LUT_4[29133] = 32'b00000000000000000000001101110001;
assign LUT_4[29134] = 32'b00000000000000000110011100011101;
assign LUT_4[29135] = 32'b11111111111111111111101000010101;
assign LUT_4[29136] = 32'b00000000000000001110100110110110;
assign LUT_4[29137] = 32'b00000000000000000111110010101110;
assign LUT_4[29138] = 32'b00000000000000001110000001011010;
assign LUT_4[29139] = 32'b00000000000000000111001101010010;
assign LUT_4[29140] = 32'b00000000000000001011100111010010;
assign LUT_4[29141] = 32'b00000000000000000100110011001010;
assign LUT_4[29142] = 32'b00000000000000001011000001110110;
assign LUT_4[29143] = 32'b00000000000000000100001101101110;
assign LUT_4[29144] = 32'b00000000000000000111110011001011;
assign LUT_4[29145] = 32'b00000000000000000000111111000011;
assign LUT_4[29146] = 32'b00000000000000000111001101101111;
assign LUT_4[29147] = 32'b00000000000000000000011001100111;
assign LUT_4[29148] = 32'b00000000000000000100110011100111;
assign LUT_4[29149] = 32'b11111111111111111101111111011111;
assign LUT_4[29150] = 32'b00000000000000000100001110001011;
assign LUT_4[29151] = 32'b11111111111111111101011010000011;
assign LUT_4[29152] = 32'b00000000000000001111010000001111;
assign LUT_4[29153] = 32'b00000000000000001000011100000111;
assign LUT_4[29154] = 32'b00000000000000001110101010110011;
assign LUT_4[29155] = 32'b00000000000000000111110110101011;
assign LUT_4[29156] = 32'b00000000000000001100010000101011;
assign LUT_4[29157] = 32'b00000000000000000101011100100011;
assign LUT_4[29158] = 32'b00000000000000001011101011001111;
assign LUT_4[29159] = 32'b00000000000000000100110111000111;
assign LUT_4[29160] = 32'b00000000000000001000011100100100;
assign LUT_4[29161] = 32'b00000000000000000001101000011100;
assign LUT_4[29162] = 32'b00000000000000000111110111001000;
assign LUT_4[29163] = 32'b00000000000000000001000011000000;
assign LUT_4[29164] = 32'b00000000000000000101011101000000;
assign LUT_4[29165] = 32'b11111111111111111110101000111000;
assign LUT_4[29166] = 32'b00000000000000000100110111100100;
assign LUT_4[29167] = 32'b11111111111111111110000011011100;
assign LUT_4[29168] = 32'b00000000000000001101000001111101;
assign LUT_4[29169] = 32'b00000000000000000110001101110101;
assign LUT_4[29170] = 32'b00000000000000001100011100100001;
assign LUT_4[29171] = 32'b00000000000000000101101000011001;
assign LUT_4[29172] = 32'b00000000000000001010000010011001;
assign LUT_4[29173] = 32'b00000000000000000011001110010001;
assign LUT_4[29174] = 32'b00000000000000001001011100111101;
assign LUT_4[29175] = 32'b00000000000000000010101000110101;
assign LUT_4[29176] = 32'b00000000000000000110001110010010;
assign LUT_4[29177] = 32'b11111111111111111111011010001010;
assign LUT_4[29178] = 32'b00000000000000000101101000110110;
assign LUT_4[29179] = 32'b11111111111111111110110100101110;
assign LUT_4[29180] = 32'b00000000000000000011001110101110;
assign LUT_4[29181] = 32'b11111111111111111100011010100110;
assign LUT_4[29182] = 32'b00000000000000000010101001010010;
assign LUT_4[29183] = 32'b11111111111111111011110101001010;
assign LUT_4[29184] = 32'b00000000000000000111000000010001;
assign LUT_4[29185] = 32'b00000000000000000000001100001001;
assign LUT_4[29186] = 32'b00000000000000000110011010110101;
assign LUT_4[29187] = 32'b11111111111111111111100110101101;
assign LUT_4[29188] = 32'b00000000000000000100000000101101;
assign LUT_4[29189] = 32'b11111111111111111101001100100101;
assign LUT_4[29190] = 32'b00000000000000000011011011010001;
assign LUT_4[29191] = 32'b11111111111111111100100111001001;
assign LUT_4[29192] = 32'b00000000000000000000001100100110;
assign LUT_4[29193] = 32'b11111111111111111001011000011110;
assign LUT_4[29194] = 32'b11111111111111111111100111001010;
assign LUT_4[29195] = 32'b11111111111111111000110011000010;
assign LUT_4[29196] = 32'b11111111111111111101001101000010;
assign LUT_4[29197] = 32'b11111111111111110110011000111010;
assign LUT_4[29198] = 32'b11111111111111111100100111100110;
assign LUT_4[29199] = 32'b11111111111111110101110011011110;
assign LUT_4[29200] = 32'b00000000000000000100110001111111;
assign LUT_4[29201] = 32'b11111111111111111101111101110111;
assign LUT_4[29202] = 32'b00000000000000000100001100100011;
assign LUT_4[29203] = 32'b11111111111111111101011000011011;
assign LUT_4[29204] = 32'b00000000000000000001110010011011;
assign LUT_4[29205] = 32'b11111111111111111010111110010011;
assign LUT_4[29206] = 32'b00000000000000000001001100111111;
assign LUT_4[29207] = 32'b11111111111111111010011000110111;
assign LUT_4[29208] = 32'b11111111111111111101111110010100;
assign LUT_4[29209] = 32'b11111111111111110111001010001100;
assign LUT_4[29210] = 32'b11111111111111111101011000111000;
assign LUT_4[29211] = 32'b11111111111111110110100100110000;
assign LUT_4[29212] = 32'b11111111111111111010111110110000;
assign LUT_4[29213] = 32'b11111111111111110100001010101000;
assign LUT_4[29214] = 32'b11111111111111111010011001010100;
assign LUT_4[29215] = 32'b11111111111111110011100101001100;
assign LUT_4[29216] = 32'b00000000000000000101011011011000;
assign LUT_4[29217] = 32'b11111111111111111110100111010000;
assign LUT_4[29218] = 32'b00000000000000000100110101111100;
assign LUT_4[29219] = 32'b11111111111111111110000001110100;
assign LUT_4[29220] = 32'b00000000000000000010011011110100;
assign LUT_4[29221] = 32'b11111111111111111011100111101100;
assign LUT_4[29222] = 32'b00000000000000000001110110011000;
assign LUT_4[29223] = 32'b11111111111111111011000010010000;
assign LUT_4[29224] = 32'b11111111111111111110100111101101;
assign LUT_4[29225] = 32'b11111111111111110111110011100101;
assign LUT_4[29226] = 32'b11111111111111111110000010010001;
assign LUT_4[29227] = 32'b11111111111111110111001110001001;
assign LUT_4[29228] = 32'b11111111111111111011101000001001;
assign LUT_4[29229] = 32'b11111111111111110100110100000001;
assign LUT_4[29230] = 32'b11111111111111111011000010101101;
assign LUT_4[29231] = 32'b11111111111111110100001110100101;
assign LUT_4[29232] = 32'b00000000000000000011001101000110;
assign LUT_4[29233] = 32'b11111111111111111100011000111110;
assign LUT_4[29234] = 32'b00000000000000000010100111101010;
assign LUT_4[29235] = 32'b11111111111111111011110011100010;
assign LUT_4[29236] = 32'b00000000000000000000001101100010;
assign LUT_4[29237] = 32'b11111111111111111001011001011010;
assign LUT_4[29238] = 32'b11111111111111111111101000000110;
assign LUT_4[29239] = 32'b11111111111111111000110011111110;
assign LUT_4[29240] = 32'b11111111111111111100011001011011;
assign LUT_4[29241] = 32'b11111111111111110101100101010011;
assign LUT_4[29242] = 32'b11111111111111111011110011111111;
assign LUT_4[29243] = 32'b11111111111111110100111111110111;
assign LUT_4[29244] = 32'b11111111111111111001011001110111;
assign LUT_4[29245] = 32'b11111111111111110010100101101111;
assign LUT_4[29246] = 32'b11111111111111111000110100011011;
assign LUT_4[29247] = 32'b11111111111111110010000000010011;
assign LUT_4[29248] = 32'b00000000000000001000010111100101;
assign LUT_4[29249] = 32'b00000000000000000001100011011101;
assign LUT_4[29250] = 32'b00000000000000000111110010001001;
assign LUT_4[29251] = 32'b00000000000000000000111110000001;
assign LUT_4[29252] = 32'b00000000000000000101011000000001;
assign LUT_4[29253] = 32'b11111111111111111110100011111001;
assign LUT_4[29254] = 32'b00000000000000000100110010100101;
assign LUT_4[29255] = 32'b11111111111111111101111110011101;
assign LUT_4[29256] = 32'b00000000000000000001100011111010;
assign LUT_4[29257] = 32'b11111111111111111010101111110010;
assign LUT_4[29258] = 32'b00000000000000000000111110011110;
assign LUT_4[29259] = 32'b11111111111111111010001010010110;
assign LUT_4[29260] = 32'b11111111111111111110100100010110;
assign LUT_4[29261] = 32'b11111111111111110111110000001110;
assign LUT_4[29262] = 32'b11111111111111111101111110111010;
assign LUT_4[29263] = 32'b11111111111111110111001010110010;
assign LUT_4[29264] = 32'b00000000000000000110001001010011;
assign LUT_4[29265] = 32'b11111111111111111111010101001011;
assign LUT_4[29266] = 32'b00000000000000000101100011110111;
assign LUT_4[29267] = 32'b11111111111111111110101111101111;
assign LUT_4[29268] = 32'b00000000000000000011001001101111;
assign LUT_4[29269] = 32'b11111111111111111100010101100111;
assign LUT_4[29270] = 32'b00000000000000000010100100010011;
assign LUT_4[29271] = 32'b11111111111111111011110000001011;
assign LUT_4[29272] = 32'b11111111111111111111010101101000;
assign LUT_4[29273] = 32'b11111111111111111000100001100000;
assign LUT_4[29274] = 32'b11111111111111111110110000001100;
assign LUT_4[29275] = 32'b11111111111111110111111100000100;
assign LUT_4[29276] = 32'b11111111111111111100010110000100;
assign LUT_4[29277] = 32'b11111111111111110101100001111100;
assign LUT_4[29278] = 32'b11111111111111111011110000101000;
assign LUT_4[29279] = 32'b11111111111111110100111100100000;
assign LUT_4[29280] = 32'b00000000000000000110110010101100;
assign LUT_4[29281] = 32'b11111111111111111111111110100100;
assign LUT_4[29282] = 32'b00000000000000000110001101010000;
assign LUT_4[29283] = 32'b11111111111111111111011001001000;
assign LUT_4[29284] = 32'b00000000000000000011110011001000;
assign LUT_4[29285] = 32'b11111111111111111100111111000000;
assign LUT_4[29286] = 32'b00000000000000000011001101101100;
assign LUT_4[29287] = 32'b11111111111111111100011001100100;
assign LUT_4[29288] = 32'b11111111111111111111111111000001;
assign LUT_4[29289] = 32'b11111111111111111001001010111001;
assign LUT_4[29290] = 32'b11111111111111111111011001100101;
assign LUT_4[29291] = 32'b11111111111111111000100101011101;
assign LUT_4[29292] = 32'b11111111111111111100111111011101;
assign LUT_4[29293] = 32'b11111111111111110110001011010101;
assign LUT_4[29294] = 32'b11111111111111111100011010000001;
assign LUT_4[29295] = 32'b11111111111111110101100101111001;
assign LUT_4[29296] = 32'b00000000000000000100100100011010;
assign LUT_4[29297] = 32'b11111111111111111101110000010010;
assign LUT_4[29298] = 32'b00000000000000000011111110111110;
assign LUT_4[29299] = 32'b11111111111111111101001010110110;
assign LUT_4[29300] = 32'b00000000000000000001100100110110;
assign LUT_4[29301] = 32'b11111111111111111010110000101110;
assign LUT_4[29302] = 32'b00000000000000000000111111011010;
assign LUT_4[29303] = 32'b11111111111111111010001011010010;
assign LUT_4[29304] = 32'b11111111111111111101110000101111;
assign LUT_4[29305] = 32'b11111111111111110110111100100111;
assign LUT_4[29306] = 32'b11111111111111111101001011010011;
assign LUT_4[29307] = 32'b11111111111111110110010111001011;
assign LUT_4[29308] = 32'b11111111111111111010110001001011;
assign LUT_4[29309] = 32'b11111111111111110011111101000011;
assign LUT_4[29310] = 32'b11111111111111111010001011101111;
assign LUT_4[29311] = 32'b11111111111111110011010111100111;
assign LUT_4[29312] = 32'b00000000000000001001100110011001;
assign LUT_4[29313] = 32'b00000000000000000010110010010001;
assign LUT_4[29314] = 32'b00000000000000001001000000111101;
assign LUT_4[29315] = 32'b00000000000000000010001100110101;
assign LUT_4[29316] = 32'b00000000000000000110100110110101;
assign LUT_4[29317] = 32'b11111111111111111111110010101101;
assign LUT_4[29318] = 32'b00000000000000000110000001011001;
assign LUT_4[29319] = 32'b11111111111111111111001101010001;
assign LUT_4[29320] = 32'b00000000000000000010110010101110;
assign LUT_4[29321] = 32'b11111111111111111011111110100110;
assign LUT_4[29322] = 32'b00000000000000000010001101010010;
assign LUT_4[29323] = 32'b11111111111111111011011001001010;
assign LUT_4[29324] = 32'b11111111111111111111110011001010;
assign LUT_4[29325] = 32'b11111111111111111000111111000010;
assign LUT_4[29326] = 32'b11111111111111111111001101101110;
assign LUT_4[29327] = 32'b11111111111111111000011001100110;
assign LUT_4[29328] = 32'b00000000000000000111011000000111;
assign LUT_4[29329] = 32'b00000000000000000000100011111111;
assign LUT_4[29330] = 32'b00000000000000000110110010101011;
assign LUT_4[29331] = 32'b11111111111111111111111110100011;
assign LUT_4[29332] = 32'b00000000000000000100011000100011;
assign LUT_4[29333] = 32'b11111111111111111101100100011011;
assign LUT_4[29334] = 32'b00000000000000000011110011000111;
assign LUT_4[29335] = 32'b11111111111111111100111110111111;
assign LUT_4[29336] = 32'b00000000000000000000100100011100;
assign LUT_4[29337] = 32'b11111111111111111001110000010100;
assign LUT_4[29338] = 32'b11111111111111111111111111000000;
assign LUT_4[29339] = 32'b11111111111111111001001010111000;
assign LUT_4[29340] = 32'b11111111111111111101100100111000;
assign LUT_4[29341] = 32'b11111111111111110110110000110000;
assign LUT_4[29342] = 32'b11111111111111111100111111011100;
assign LUT_4[29343] = 32'b11111111111111110110001011010100;
assign LUT_4[29344] = 32'b00000000000000001000000001100000;
assign LUT_4[29345] = 32'b00000000000000000001001101011000;
assign LUT_4[29346] = 32'b00000000000000000111011100000100;
assign LUT_4[29347] = 32'b00000000000000000000100111111100;
assign LUT_4[29348] = 32'b00000000000000000101000001111100;
assign LUT_4[29349] = 32'b11111111111111111110001101110100;
assign LUT_4[29350] = 32'b00000000000000000100011100100000;
assign LUT_4[29351] = 32'b11111111111111111101101000011000;
assign LUT_4[29352] = 32'b00000000000000000001001101110101;
assign LUT_4[29353] = 32'b11111111111111111010011001101101;
assign LUT_4[29354] = 32'b00000000000000000000101000011001;
assign LUT_4[29355] = 32'b11111111111111111001110100010001;
assign LUT_4[29356] = 32'b11111111111111111110001110010001;
assign LUT_4[29357] = 32'b11111111111111110111011010001001;
assign LUT_4[29358] = 32'b11111111111111111101101000110101;
assign LUT_4[29359] = 32'b11111111111111110110110100101101;
assign LUT_4[29360] = 32'b00000000000000000101110011001110;
assign LUT_4[29361] = 32'b11111111111111111110111111000110;
assign LUT_4[29362] = 32'b00000000000000000101001101110010;
assign LUT_4[29363] = 32'b11111111111111111110011001101010;
assign LUT_4[29364] = 32'b00000000000000000010110011101010;
assign LUT_4[29365] = 32'b11111111111111111011111111100010;
assign LUT_4[29366] = 32'b00000000000000000010001110001110;
assign LUT_4[29367] = 32'b11111111111111111011011010000110;
assign LUT_4[29368] = 32'b11111111111111111110111111100011;
assign LUT_4[29369] = 32'b11111111111111111000001011011011;
assign LUT_4[29370] = 32'b11111111111111111110011010000111;
assign LUT_4[29371] = 32'b11111111111111110111100101111111;
assign LUT_4[29372] = 32'b11111111111111111011111111111111;
assign LUT_4[29373] = 32'b11111111111111110101001011110111;
assign LUT_4[29374] = 32'b11111111111111111011011010100011;
assign LUT_4[29375] = 32'b11111111111111110100100110011011;
assign LUT_4[29376] = 32'b00000000000000001010111101101101;
assign LUT_4[29377] = 32'b00000000000000000100001001100101;
assign LUT_4[29378] = 32'b00000000000000001010011000010001;
assign LUT_4[29379] = 32'b00000000000000000011100100001001;
assign LUT_4[29380] = 32'b00000000000000000111111110001001;
assign LUT_4[29381] = 32'b00000000000000000001001010000001;
assign LUT_4[29382] = 32'b00000000000000000111011000101101;
assign LUT_4[29383] = 32'b00000000000000000000100100100101;
assign LUT_4[29384] = 32'b00000000000000000100001010000010;
assign LUT_4[29385] = 32'b11111111111111111101010101111010;
assign LUT_4[29386] = 32'b00000000000000000011100100100110;
assign LUT_4[29387] = 32'b11111111111111111100110000011110;
assign LUT_4[29388] = 32'b00000000000000000001001010011110;
assign LUT_4[29389] = 32'b11111111111111111010010110010110;
assign LUT_4[29390] = 32'b00000000000000000000100101000010;
assign LUT_4[29391] = 32'b11111111111111111001110000111010;
assign LUT_4[29392] = 32'b00000000000000001000101111011011;
assign LUT_4[29393] = 32'b00000000000000000001111011010011;
assign LUT_4[29394] = 32'b00000000000000001000001001111111;
assign LUT_4[29395] = 32'b00000000000000000001010101110111;
assign LUT_4[29396] = 32'b00000000000000000101101111110111;
assign LUT_4[29397] = 32'b11111111111111111110111011101111;
assign LUT_4[29398] = 32'b00000000000000000101001010011011;
assign LUT_4[29399] = 32'b11111111111111111110010110010011;
assign LUT_4[29400] = 32'b00000000000000000001111011110000;
assign LUT_4[29401] = 32'b11111111111111111011000111101000;
assign LUT_4[29402] = 32'b00000000000000000001010110010100;
assign LUT_4[29403] = 32'b11111111111111111010100010001100;
assign LUT_4[29404] = 32'b11111111111111111110111100001100;
assign LUT_4[29405] = 32'b11111111111111111000001000000100;
assign LUT_4[29406] = 32'b11111111111111111110010110110000;
assign LUT_4[29407] = 32'b11111111111111110111100010101000;
assign LUT_4[29408] = 32'b00000000000000001001011000110100;
assign LUT_4[29409] = 32'b00000000000000000010100100101100;
assign LUT_4[29410] = 32'b00000000000000001000110011011000;
assign LUT_4[29411] = 32'b00000000000000000001111111010000;
assign LUT_4[29412] = 32'b00000000000000000110011001010000;
assign LUT_4[29413] = 32'b11111111111111111111100101001000;
assign LUT_4[29414] = 32'b00000000000000000101110011110100;
assign LUT_4[29415] = 32'b11111111111111111110111111101100;
assign LUT_4[29416] = 32'b00000000000000000010100101001001;
assign LUT_4[29417] = 32'b11111111111111111011110001000001;
assign LUT_4[29418] = 32'b00000000000000000001111111101101;
assign LUT_4[29419] = 32'b11111111111111111011001011100101;
assign LUT_4[29420] = 32'b11111111111111111111100101100101;
assign LUT_4[29421] = 32'b11111111111111111000110001011101;
assign LUT_4[29422] = 32'b11111111111111111111000000001001;
assign LUT_4[29423] = 32'b11111111111111111000001100000001;
assign LUT_4[29424] = 32'b00000000000000000111001010100010;
assign LUT_4[29425] = 32'b00000000000000000000010110011010;
assign LUT_4[29426] = 32'b00000000000000000110100101000110;
assign LUT_4[29427] = 32'b11111111111111111111110000111110;
assign LUT_4[29428] = 32'b00000000000000000100001010111110;
assign LUT_4[29429] = 32'b11111111111111111101010110110110;
assign LUT_4[29430] = 32'b00000000000000000011100101100010;
assign LUT_4[29431] = 32'b11111111111111111100110001011010;
assign LUT_4[29432] = 32'b00000000000000000000010110110111;
assign LUT_4[29433] = 32'b11111111111111111001100010101111;
assign LUT_4[29434] = 32'b11111111111111111111110001011011;
assign LUT_4[29435] = 32'b11111111111111111000111101010011;
assign LUT_4[29436] = 32'b11111111111111111101010111010011;
assign LUT_4[29437] = 32'b11111111111111110110100011001011;
assign LUT_4[29438] = 32'b11111111111111111100110001110111;
assign LUT_4[29439] = 32'b11111111111111110101111101101111;
assign LUT_4[29440] = 32'b00000000000000001011111011110100;
assign LUT_4[29441] = 32'b00000000000000000101000111101100;
assign LUT_4[29442] = 32'b00000000000000001011010110011000;
assign LUT_4[29443] = 32'b00000000000000000100100010010000;
assign LUT_4[29444] = 32'b00000000000000001000111100010000;
assign LUT_4[29445] = 32'b00000000000000000010001000001000;
assign LUT_4[29446] = 32'b00000000000000001000010110110100;
assign LUT_4[29447] = 32'b00000000000000000001100010101100;
assign LUT_4[29448] = 32'b00000000000000000101001000001001;
assign LUT_4[29449] = 32'b11111111111111111110010100000001;
assign LUT_4[29450] = 32'b00000000000000000100100010101101;
assign LUT_4[29451] = 32'b11111111111111111101101110100101;
assign LUT_4[29452] = 32'b00000000000000000010001000100101;
assign LUT_4[29453] = 32'b11111111111111111011010100011101;
assign LUT_4[29454] = 32'b00000000000000000001100011001001;
assign LUT_4[29455] = 32'b11111111111111111010101111000001;
assign LUT_4[29456] = 32'b00000000000000001001101101100010;
assign LUT_4[29457] = 32'b00000000000000000010111001011010;
assign LUT_4[29458] = 32'b00000000000000001001001000000110;
assign LUT_4[29459] = 32'b00000000000000000010010011111110;
assign LUT_4[29460] = 32'b00000000000000000110101101111110;
assign LUT_4[29461] = 32'b11111111111111111111111001110110;
assign LUT_4[29462] = 32'b00000000000000000110001000100010;
assign LUT_4[29463] = 32'b11111111111111111111010100011010;
assign LUT_4[29464] = 32'b00000000000000000010111001110111;
assign LUT_4[29465] = 32'b11111111111111111100000101101111;
assign LUT_4[29466] = 32'b00000000000000000010010100011011;
assign LUT_4[29467] = 32'b11111111111111111011100000010011;
assign LUT_4[29468] = 32'b11111111111111111111111010010011;
assign LUT_4[29469] = 32'b11111111111111111001000110001011;
assign LUT_4[29470] = 32'b11111111111111111111010100110111;
assign LUT_4[29471] = 32'b11111111111111111000100000101111;
assign LUT_4[29472] = 32'b00000000000000001010010110111011;
assign LUT_4[29473] = 32'b00000000000000000011100010110011;
assign LUT_4[29474] = 32'b00000000000000001001110001011111;
assign LUT_4[29475] = 32'b00000000000000000010111101010111;
assign LUT_4[29476] = 32'b00000000000000000111010111010111;
assign LUT_4[29477] = 32'b00000000000000000000100011001111;
assign LUT_4[29478] = 32'b00000000000000000110110001111011;
assign LUT_4[29479] = 32'b11111111111111111111111101110011;
assign LUT_4[29480] = 32'b00000000000000000011100011010000;
assign LUT_4[29481] = 32'b11111111111111111100101111001000;
assign LUT_4[29482] = 32'b00000000000000000010111101110100;
assign LUT_4[29483] = 32'b11111111111111111100001001101100;
assign LUT_4[29484] = 32'b00000000000000000000100011101100;
assign LUT_4[29485] = 32'b11111111111111111001101111100100;
assign LUT_4[29486] = 32'b11111111111111111111111110010000;
assign LUT_4[29487] = 32'b11111111111111111001001010001000;
assign LUT_4[29488] = 32'b00000000000000001000001000101001;
assign LUT_4[29489] = 32'b00000000000000000001010100100001;
assign LUT_4[29490] = 32'b00000000000000000111100011001101;
assign LUT_4[29491] = 32'b00000000000000000000101111000101;
assign LUT_4[29492] = 32'b00000000000000000101001001000101;
assign LUT_4[29493] = 32'b11111111111111111110010100111101;
assign LUT_4[29494] = 32'b00000000000000000100100011101001;
assign LUT_4[29495] = 32'b11111111111111111101101111100001;
assign LUT_4[29496] = 32'b00000000000000000001010100111110;
assign LUT_4[29497] = 32'b11111111111111111010100000110110;
assign LUT_4[29498] = 32'b00000000000000000000101111100010;
assign LUT_4[29499] = 32'b11111111111111111001111011011010;
assign LUT_4[29500] = 32'b11111111111111111110010101011010;
assign LUT_4[29501] = 32'b11111111111111110111100001010010;
assign LUT_4[29502] = 32'b11111111111111111101101111111110;
assign LUT_4[29503] = 32'b11111111111111110110111011110110;
assign LUT_4[29504] = 32'b00000000000000001101010011001000;
assign LUT_4[29505] = 32'b00000000000000000110011111000000;
assign LUT_4[29506] = 32'b00000000000000001100101101101100;
assign LUT_4[29507] = 32'b00000000000000000101111001100100;
assign LUT_4[29508] = 32'b00000000000000001010010011100100;
assign LUT_4[29509] = 32'b00000000000000000011011111011100;
assign LUT_4[29510] = 32'b00000000000000001001101110001000;
assign LUT_4[29511] = 32'b00000000000000000010111010000000;
assign LUT_4[29512] = 32'b00000000000000000110011111011101;
assign LUT_4[29513] = 32'b11111111111111111111101011010101;
assign LUT_4[29514] = 32'b00000000000000000101111010000001;
assign LUT_4[29515] = 32'b11111111111111111111000101111001;
assign LUT_4[29516] = 32'b00000000000000000011011111111001;
assign LUT_4[29517] = 32'b11111111111111111100101011110001;
assign LUT_4[29518] = 32'b00000000000000000010111010011101;
assign LUT_4[29519] = 32'b11111111111111111100000110010101;
assign LUT_4[29520] = 32'b00000000000000001011000100110110;
assign LUT_4[29521] = 32'b00000000000000000100010000101110;
assign LUT_4[29522] = 32'b00000000000000001010011111011010;
assign LUT_4[29523] = 32'b00000000000000000011101011010010;
assign LUT_4[29524] = 32'b00000000000000001000000101010010;
assign LUT_4[29525] = 32'b00000000000000000001010001001010;
assign LUT_4[29526] = 32'b00000000000000000111011111110110;
assign LUT_4[29527] = 32'b00000000000000000000101011101110;
assign LUT_4[29528] = 32'b00000000000000000100010001001011;
assign LUT_4[29529] = 32'b11111111111111111101011101000011;
assign LUT_4[29530] = 32'b00000000000000000011101011101111;
assign LUT_4[29531] = 32'b11111111111111111100110111100111;
assign LUT_4[29532] = 32'b00000000000000000001010001100111;
assign LUT_4[29533] = 32'b11111111111111111010011101011111;
assign LUT_4[29534] = 32'b00000000000000000000101100001011;
assign LUT_4[29535] = 32'b11111111111111111001111000000011;
assign LUT_4[29536] = 32'b00000000000000001011101110001111;
assign LUT_4[29537] = 32'b00000000000000000100111010000111;
assign LUT_4[29538] = 32'b00000000000000001011001000110011;
assign LUT_4[29539] = 32'b00000000000000000100010100101011;
assign LUT_4[29540] = 32'b00000000000000001000101110101011;
assign LUT_4[29541] = 32'b00000000000000000001111010100011;
assign LUT_4[29542] = 32'b00000000000000001000001001001111;
assign LUT_4[29543] = 32'b00000000000000000001010101000111;
assign LUT_4[29544] = 32'b00000000000000000100111010100100;
assign LUT_4[29545] = 32'b11111111111111111110000110011100;
assign LUT_4[29546] = 32'b00000000000000000100010101001000;
assign LUT_4[29547] = 32'b11111111111111111101100001000000;
assign LUT_4[29548] = 32'b00000000000000000001111011000000;
assign LUT_4[29549] = 32'b11111111111111111011000110111000;
assign LUT_4[29550] = 32'b00000000000000000001010101100100;
assign LUT_4[29551] = 32'b11111111111111111010100001011100;
assign LUT_4[29552] = 32'b00000000000000001001011111111101;
assign LUT_4[29553] = 32'b00000000000000000010101011110101;
assign LUT_4[29554] = 32'b00000000000000001000111010100001;
assign LUT_4[29555] = 32'b00000000000000000010000110011001;
assign LUT_4[29556] = 32'b00000000000000000110100000011001;
assign LUT_4[29557] = 32'b11111111111111111111101100010001;
assign LUT_4[29558] = 32'b00000000000000000101111010111101;
assign LUT_4[29559] = 32'b11111111111111111111000110110101;
assign LUT_4[29560] = 32'b00000000000000000010101100010010;
assign LUT_4[29561] = 32'b11111111111111111011111000001010;
assign LUT_4[29562] = 32'b00000000000000000010000110110110;
assign LUT_4[29563] = 32'b11111111111111111011010010101110;
assign LUT_4[29564] = 32'b11111111111111111111101100101110;
assign LUT_4[29565] = 32'b11111111111111111000111000100110;
assign LUT_4[29566] = 32'b11111111111111111111000111010010;
assign LUT_4[29567] = 32'b11111111111111111000010011001010;
assign LUT_4[29568] = 32'b00000000000000001110100001111100;
assign LUT_4[29569] = 32'b00000000000000000111101101110100;
assign LUT_4[29570] = 32'b00000000000000001101111100100000;
assign LUT_4[29571] = 32'b00000000000000000111001000011000;
assign LUT_4[29572] = 32'b00000000000000001011100010011000;
assign LUT_4[29573] = 32'b00000000000000000100101110010000;
assign LUT_4[29574] = 32'b00000000000000001010111100111100;
assign LUT_4[29575] = 32'b00000000000000000100001000110100;
assign LUT_4[29576] = 32'b00000000000000000111101110010001;
assign LUT_4[29577] = 32'b00000000000000000000111010001001;
assign LUT_4[29578] = 32'b00000000000000000111001000110101;
assign LUT_4[29579] = 32'b00000000000000000000010100101101;
assign LUT_4[29580] = 32'b00000000000000000100101110101101;
assign LUT_4[29581] = 32'b11111111111111111101111010100101;
assign LUT_4[29582] = 32'b00000000000000000100001001010001;
assign LUT_4[29583] = 32'b11111111111111111101010101001001;
assign LUT_4[29584] = 32'b00000000000000001100010011101010;
assign LUT_4[29585] = 32'b00000000000000000101011111100010;
assign LUT_4[29586] = 32'b00000000000000001011101110001110;
assign LUT_4[29587] = 32'b00000000000000000100111010000110;
assign LUT_4[29588] = 32'b00000000000000001001010100000110;
assign LUT_4[29589] = 32'b00000000000000000010011111111110;
assign LUT_4[29590] = 32'b00000000000000001000101110101010;
assign LUT_4[29591] = 32'b00000000000000000001111010100010;
assign LUT_4[29592] = 32'b00000000000000000101011111111111;
assign LUT_4[29593] = 32'b11111111111111111110101011110111;
assign LUT_4[29594] = 32'b00000000000000000100111010100011;
assign LUT_4[29595] = 32'b11111111111111111110000110011011;
assign LUT_4[29596] = 32'b00000000000000000010100000011011;
assign LUT_4[29597] = 32'b11111111111111111011101100010011;
assign LUT_4[29598] = 32'b00000000000000000001111010111111;
assign LUT_4[29599] = 32'b11111111111111111011000110110111;
assign LUT_4[29600] = 32'b00000000000000001100111101000011;
assign LUT_4[29601] = 32'b00000000000000000110001000111011;
assign LUT_4[29602] = 32'b00000000000000001100010111100111;
assign LUT_4[29603] = 32'b00000000000000000101100011011111;
assign LUT_4[29604] = 32'b00000000000000001001111101011111;
assign LUT_4[29605] = 32'b00000000000000000011001001010111;
assign LUT_4[29606] = 32'b00000000000000001001011000000011;
assign LUT_4[29607] = 32'b00000000000000000010100011111011;
assign LUT_4[29608] = 32'b00000000000000000110001001011000;
assign LUT_4[29609] = 32'b11111111111111111111010101010000;
assign LUT_4[29610] = 32'b00000000000000000101100011111100;
assign LUT_4[29611] = 32'b11111111111111111110101111110100;
assign LUT_4[29612] = 32'b00000000000000000011001001110100;
assign LUT_4[29613] = 32'b11111111111111111100010101101100;
assign LUT_4[29614] = 32'b00000000000000000010100100011000;
assign LUT_4[29615] = 32'b11111111111111111011110000010000;
assign LUT_4[29616] = 32'b00000000000000001010101110110001;
assign LUT_4[29617] = 32'b00000000000000000011111010101001;
assign LUT_4[29618] = 32'b00000000000000001010001001010101;
assign LUT_4[29619] = 32'b00000000000000000011010101001101;
assign LUT_4[29620] = 32'b00000000000000000111101111001101;
assign LUT_4[29621] = 32'b00000000000000000000111011000101;
assign LUT_4[29622] = 32'b00000000000000000111001001110001;
assign LUT_4[29623] = 32'b00000000000000000000010101101001;
assign LUT_4[29624] = 32'b00000000000000000011111011000110;
assign LUT_4[29625] = 32'b11111111111111111101000110111110;
assign LUT_4[29626] = 32'b00000000000000000011010101101010;
assign LUT_4[29627] = 32'b11111111111111111100100001100010;
assign LUT_4[29628] = 32'b00000000000000000000111011100010;
assign LUT_4[29629] = 32'b11111111111111111010000111011010;
assign LUT_4[29630] = 32'b00000000000000000000010110000110;
assign LUT_4[29631] = 32'b11111111111111111001100001111110;
assign LUT_4[29632] = 32'b00000000000000001111111001010000;
assign LUT_4[29633] = 32'b00000000000000001001000101001000;
assign LUT_4[29634] = 32'b00000000000000001111010011110100;
assign LUT_4[29635] = 32'b00000000000000001000011111101100;
assign LUT_4[29636] = 32'b00000000000000001100111001101100;
assign LUT_4[29637] = 32'b00000000000000000110000101100100;
assign LUT_4[29638] = 32'b00000000000000001100010100010000;
assign LUT_4[29639] = 32'b00000000000000000101100000001000;
assign LUT_4[29640] = 32'b00000000000000001001000101100101;
assign LUT_4[29641] = 32'b00000000000000000010010001011101;
assign LUT_4[29642] = 32'b00000000000000001000100000001001;
assign LUT_4[29643] = 32'b00000000000000000001101100000001;
assign LUT_4[29644] = 32'b00000000000000000110000110000001;
assign LUT_4[29645] = 32'b11111111111111111111010001111001;
assign LUT_4[29646] = 32'b00000000000000000101100000100101;
assign LUT_4[29647] = 32'b11111111111111111110101100011101;
assign LUT_4[29648] = 32'b00000000000000001101101010111110;
assign LUT_4[29649] = 32'b00000000000000000110110110110110;
assign LUT_4[29650] = 32'b00000000000000001101000101100010;
assign LUT_4[29651] = 32'b00000000000000000110010001011010;
assign LUT_4[29652] = 32'b00000000000000001010101011011010;
assign LUT_4[29653] = 32'b00000000000000000011110111010010;
assign LUT_4[29654] = 32'b00000000000000001010000101111110;
assign LUT_4[29655] = 32'b00000000000000000011010001110110;
assign LUT_4[29656] = 32'b00000000000000000110110111010011;
assign LUT_4[29657] = 32'b00000000000000000000000011001011;
assign LUT_4[29658] = 32'b00000000000000000110010001110111;
assign LUT_4[29659] = 32'b11111111111111111111011101101111;
assign LUT_4[29660] = 32'b00000000000000000011110111101111;
assign LUT_4[29661] = 32'b11111111111111111101000011100111;
assign LUT_4[29662] = 32'b00000000000000000011010010010011;
assign LUT_4[29663] = 32'b11111111111111111100011110001011;
assign LUT_4[29664] = 32'b00000000000000001110010100010111;
assign LUT_4[29665] = 32'b00000000000000000111100000001111;
assign LUT_4[29666] = 32'b00000000000000001101101110111011;
assign LUT_4[29667] = 32'b00000000000000000110111010110011;
assign LUT_4[29668] = 32'b00000000000000001011010100110011;
assign LUT_4[29669] = 32'b00000000000000000100100000101011;
assign LUT_4[29670] = 32'b00000000000000001010101111010111;
assign LUT_4[29671] = 32'b00000000000000000011111011001111;
assign LUT_4[29672] = 32'b00000000000000000111100000101100;
assign LUT_4[29673] = 32'b00000000000000000000101100100100;
assign LUT_4[29674] = 32'b00000000000000000110111011010000;
assign LUT_4[29675] = 32'b00000000000000000000000111001000;
assign LUT_4[29676] = 32'b00000000000000000100100001001000;
assign LUT_4[29677] = 32'b11111111111111111101101101000000;
assign LUT_4[29678] = 32'b00000000000000000011111011101100;
assign LUT_4[29679] = 32'b11111111111111111101000111100100;
assign LUT_4[29680] = 32'b00000000000000001100000110000101;
assign LUT_4[29681] = 32'b00000000000000000101010001111101;
assign LUT_4[29682] = 32'b00000000000000001011100000101001;
assign LUT_4[29683] = 32'b00000000000000000100101100100001;
assign LUT_4[29684] = 32'b00000000000000001001000110100001;
assign LUT_4[29685] = 32'b00000000000000000010010010011001;
assign LUT_4[29686] = 32'b00000000000000001000100001000101;
assign LUT_4[29687] = 32'b00000000000000000001101100111101;
assign LUT_4[29688] = 32'b00000000000000000101010010011010;
assign LUT_4[29689] = 32'b11111111111111111110011110010010;
assign LUT_4[29690] = 32'b00000000000000000100101100111110;
assign LUT_4[29691] = 32'b11111111111111111101111000110110;
assign LUT_4[29692] = 32'b00000000000000000010010010110110;
assign LUT_4[29693] = 32'b11111111111111111011011110101110;
assign LUT_4[29694] = 32'b00000000000000000001101101011010;
assign LUT_4[29695] = 32'b11111111111111111010111001010010;
assign LUT_4[29696] = 32'b00000000000000001001100110101000;
assign LUT_4[29697] = 32'b00000000000000000010110010100000;
assign LUT_4[29698] = 32'b00000000000000001001000001001100;
assign LUT_4[29699] = 32'b00000000000000000010001101000100;
assign LUT_4[29700] = 32'b00000000000000000110100111000100;
assign LUT_4[29701] = 32'b11111111111111111111110010111100;
assign LUT_4[29702] = 32'b00000000000000000110000001101000;
assign LUT_4[29703] = 32'b11111111111111111111001101100000;
assign LUT_4[29704] = 32'b00000000000000000010110010111101;
assign LUT_4[29705] = 32'b11111111111111111011111110110101;
assign LUT_4[29706] = 32'b00000000000000000010001101100001;
assign LUT_4[29707] = 32'b11111111111111111011011001011001;
assign LUT_4[29708] = 32'b11111111111111111111110011011001;
assign LUT_4[29709] = 32'b11111111111111111000111111010001;
assign LUT_4[29710] = 32'b11111111111111111111001101111101;
assign LUT_4[29711] = 32'b11111111111111111000011001110101;
assign LUT_4[29712] = 32'b00000000000000000111011000010110;
assign LUT_4[29713] = 32'b00000000000000000000100100001110;
assign LUT_4[29714] = 32'b00000000000000000110110010111010;
assign LUT_4[29715] = 32'b11111111111111111111111110110010;
assign LUT_4[29716] = 32'b00000000000000000100011000110010;
assign LUT_4[29717] = 32'b11111111111111111101100100101010;
assign LUT_4[29718] = 32'b00000000000000000011110011010110;
assign LUT_4[29719] = 32'b11111111111111111100111111001110;
assign LUT_4[29720] = 32'b00000000000000000000100100101011;
assign LUT_4[29721] = 32'b11111111111111111001110000100011;
assign LUT_4[29722] = 32'b11111111111111111111111111001111;
assign LUT_4[29723] = 32'b11111111111111111001001011000111;
assign LUT_4[29724] = 32'b11111111111111111101100101000111;
assign LUT_4[29725] = 32'b11111111111111110110110000111111;
assign LUT_4[29726] = 32'b11111111111111111100111111101011;
assign LUT_4[29727] = 32'b11111111111111110110001011100011;
assign LUT_4[29728] = 32'b00000000000000001000000001101111;
assign LUT_4[29729] = 32'b00000000000000000001001101100111;
assign LUT_4[29730] = 32'b00000000000000000111011100010011;
assign LUT_4[29731] = 32'b00000000000000000000101000001011;
assign LUT_4[29732] = 32'b00000000000000000101000010001011;
assign LUT_4[29733] = 32'b11111111111111111110001110000011;
assign LUT_4[29734] = 32'b00000000000000000100011100101111;
assign LUT_4[29735] = 32'b11111111111111111101101000100111;
assign LUT_4[29736] = 32'b00000000000000000001001110000100;
assign LUT_4[29737] = 32'b11111111111111111010011001111100;
assign LUT_4[29738] = 32'b00000000000000000000101000101000;
assign LUT_4[29739] = 32'b11111111111111111001110100100000;
assign LUT_4[29740] = 32'b11111111111111111110001110100000;
assign LUT_4[29741] = 32'b11111111111111110111011010011000;
assign LUT_4[29742] = 32'b11111111111111111101101001000100;
assign LUT_4[29743] = 32'b11111111111111110110110100111100;
assign LUT_4[29744] = 32'b00000000000000000101110011011101;
assign LUT_4[29745] = 32'b11111111111111111110111111010101;
assign LUT_4[29746] = 32'b00000000000000000101001110000001;
assign LUT_4[29747] = 32'b11111111111111111110011001111001;
assign LUT_4[29748] = 32'b00000000000000000010110011111001;
assign LUT_4[29749] = 32'b11111111111111111011111111110001;
assign LUT_4[29750] = 32'b00000000000000000010001110011101;
assign LUT_4[29751] = 32'b11111111111111111011011010010101;
assign LUT_4[29752] = 32'b11111111111111111110111111110010;
assign LUT_4[29753] = 32'b11111111111111111000001011101010;
assign LUT_4[29754] = 32'b11111111111111111110011010010110;
assign LUT_4[29755] = 32'b11111111111111110111100110001110;
assign LUT_4[29756] = 32'b11111111111111111100000000001110;
assign LUT_4[29757] = 32'b11111111111111110101001100000110;
assign LUT_4[29758] = 32'b11111111111111111011011010110010;
assign LUT_4[29759] = 32'b11111111111111110100100110101010;
assign LUT_4[29760] = 32'b00000000000000001010111101111100;
assign LUT_4[29761] = 32'b00000000000000000100001001110100;
assign LUT_4[29762] = 32'b00000000000000001010011000100000;
assign LUT_4[29763] = 32'b00000000000000000011100100011000;
assign LUT_4[29764] = 32'b00000000000000000111111110011000;
assign LUT_4[29765] = 32'b00000000000000000001001010010000;
assign LUT_4[29766] = 32'b00000000000000000111011000111100;
assign LUT_4[29767] = 32'b00000000000000000000100100110100;
assign LUT_4[29768] = 32'b00000000000000000100001010010001;
assign LUT_4[29769] = 32'b11111111111111111101010110001001;
assign LUT_4[29770] = 32'b00000000000000000011100100110101;
assign LUT_4[29771] = 32'b11111111111111111100110000101101;
assign LUT_4[29772] = 32'b00000000000000000001001010101101;
assign LUT_4[29773] = 32'b11111111111111111010010110100101;
assign LUT_4[29774] = 32'b00000000000000000000100101010001;
assign LUT_4[29775] = 32'b11111111111111111001110001001001;
assign LUT_4[29776] = 32'b00000000000000001000101111101010;
assign LUT_4[29777] = 32'b00000000000000000001111011100010;
assign LUT_4[29778] = 32'b00000000000000001000001010001110;
assign LUT_4[29779] = 32'b00000000000000000001010110000110;
assign LUT_4[29780] = 32'b00000000000000000101110000000110;
assign LUT_4[29781] = 32'b11111111111111111110111011111110;
assign LUT_4[29782] = 32'b00000000000000000101001010101010;
assign LUT_4[29783] = 32'b11111111111111111110010110100010;
assign LUT_4[29784] = 32'b00000000000000000001111011111111;
assign LUT_4[29785] = 32'b11111111111111111011000111110111;
assign LUT_4[29786] = 32'b00000000000000000001010110100011;
assign LUT_4[29787] = 32'b11111111111111111010100010011011;
assign LUT_4[29788] = 32'b11111111111111111110111100011011;
assign LUT_4[29789] = 32'b11111111111111111000001000010011;
assign LUT_4[29790] = 32'b11111111111111111110010110111111;
assign LUT_4[29791] = 32'b11111111111111110111100010110111;
assign LUT_4[29792] = 32'b00000000000000001001011001000011;
assign LUT_4[29793] = 32'b00000000000000000010100100111011;
assign LUT_4[29794] = 32'b00000000000000001000110011100111;
assign LUT_4[29795] = 32'b00000000000000000001111111011111;
assign LUT_4[29796] = 32'b00000000000000000110011001011111;
assign LUT_4[29797] = 32'b11111111111111111111100101010111;
assign LUT_4[29798] = 32'b00000000000000000101110100000011;
assign LUT_4[29799] = 32'b11111111111111111110111111111011;
assign LUT_4[29800] = 32'b00000000000000000010100101011000;
assign LUT_4[29801] = 32'b11111111111111111011110001010000;
assign LUT_4[29802] = 32'b00000000000000000001111111111100;
assign LUT_4[29803] = 32'b11111111111111111011001011110100;
assign LUT_4[29804] = 32'b11111111111111111111100101110100;
assign LUT_4[29805] = 32'b11111111111111111000110001101100;
assign LUT_4[29806] = 32'b11111111111111111111000000011000;
assign LUT_4[29807] = 32'b11111111111111111000001100010000;
assign LUT_4[29808] = 32'b00000000000000000111001010110001;
assign LUT_4[29809] = 32'b00000000000000000000010110101001;
assign LUT_4[29810] = 32'b00000000000000000110100101010101;
assign LUT_4[29811] = 32'b11111111111111111111110001001101;
assign LUT_4[29812] = 32'b00000000000000000100001011001101;
assign LUT_4[29813] = 32'b11111111111111111101010111000101;
assign LUT_4[29814] = 32'b00000000000000000011100101110001;
assign LUT_4[29815] = 32'b11111111111111111100110001101001;
assign LUT_4[29816] = 32'b00000000000000000000010111000110;
assign LUT_4[29817] = 32'b11111111111111111001100010111110;
assign LUT_4[29818] = 32'b11111111111111111111110001101010;
assign LUT_4[29819] = 32'b11111111111111111000111101100010;
assign LUT_4[29820] = 32'b11111111111111111101010111100010;
assign LUT_4[29821] = 32'b11111111111111110110100011011010;
assign LUT_4[29822] = 32'b11111111111111111100110010000110;
assign LUT_4[29823] = 32'b11111111111111110101111101111110;
assign LUT_4[29824] = 32'b00000000000000001100001100110000;
assign LUT_4[29825] = 32'b00000000000000000101011000101000;
assign LUT_4[29826] = 32'b00000000000000001011100111010100;
assign LUT_4[29827] = 32'b00000000000000000100110011001100;
assign LUT_4[29828] = 32'b00000000000000001001001101001100;
assign LUT_4[29829] = 32'b00000000000000000010011001000100;
assign LUT_4[29830] = 32'b00000000000000001000100111110000;
assign LUT_4[29831] = 32'b00000000000000000001110011101000;
assign LUT_4[29832] = 32'b00000000000000000101011001000101;
assign LUT_4[29833] = 32'b11111111111111111110100100111101;
assign LUT_4[29834] = 32'b00000000000000000100110011101001;
assign LUT_4[29835] = 32'b11111111111111111101111111100001;
assign LUT_4[29836] = 32'b00000000000000000010011001100001;
assign LUT_4[29837] = 32'b11111111111111111011100101011001;
assign LUT_4[29838] = 32'b00000000000000000001110100000101;
assign LUT_4[29839] = 32'b11111111111111111010111111111101;
assign LUT_4[29840] = 32'b00000000000000001001111110011110;
assign LUT_4[29841] = 32'b00000000000000000011001010010110;
assign LUT_4[29842] = 32'b00000000000000001001011001000010;
assign LUT_4[29843] = 32'b00000000000000000010100100111010;
assign LUT_4[29844] = 32'b00000000000000000110111110111010;
assign LUT_4[29845] = 32'b00000000000000000000001010110010;
assign LUT_4[29846] = 32'b00000000000000000110011001011110;
assign LUT_4[29847] = 32'b11111111111111111111100101010110;
assign LUT_4[29848] = 32'b00000000000000000011001010110011;
assign LUT_4[29849] = 32'b11111111111111111100010110101011;
assign LUT_4[29850] = 32'b00000000000000000010100101010111;
assign LUT_4[29851] = 32'b11111111111111111011110001001111;
assign LUT_4[29852] = 32'b00000000000000000000001011001111;
assign LUT_4[29853] = 32'b11111111111111111001010111000111;
assign LUT_4[29854] = 32'b11111111111111111111100101110011;
assign LUT_4[29855] = 32'b11111111111111111000110001101011;
assign LUT_4[29856] = 32'b00000000000000001010100111110111;
assign LUT_4[29857] = 32'b00000000000000000011110011101111;
assign LUT_4[29858] = 32'b00000000000000001010000010011011;
assign LUT_4[29859] = 32'b00000000000000000011001110010011;
assign LUT_4[29860] = 32'b00000000000000000111101000010011;
assign LUT_4[29861] = 32'b00000000000000000000110100001011;
assign LUT_4[29862] = 32'b00000000000000000111000010110111;
assign LUT_4[29863] = 32'b00000000000000000000001110101111;
assign LUT_4[29864] = 32'b00000000000000000011110100001100;
assign LUT_4[29865] = 32'b11111111111111111101000000000100;
assign LUT_4[29866] = 32'b00000000000000000011001110110000;
assign LUT_4[29867] = 32'b11111111111111111100011010101000;
assign LUT_4[29868] = 32'b00000000000000000000110100101000;
assign LUT_4[29869] = 32'b11111111111111111010000000100000;
assign LUT_4[29870] = 32'b00000000000000000000001111001100;
assign LUT_4[29871] = 32'b11111111111111111001011011000100;
assign LUT_4[29872] = 32'b00000000000000001000011001100101;
assign LUT_4[29873] = 32'b00000000000000000001100101011101;
assign LUT_4[29874] = 32'b00000000000000000111110100001001;
assign LUT_4[29875] = 32'b00000000000000000001000000000001;
assign LUT_4[29876] = 32'b00000000000000000101011010000001;
assign LUT_4[29877] = 32'b11111111111111111110100101111001;
assign LUT_4[29878] = 32'b00000000000000000100110100100101;
assign LUT_4[29879] = 32'b11111111111111111110000000011101;
assign LUT_4[29880] = 32'b00000000000000000001100101111010;
assign LUT_4[29881] = 32'b11111111111111111010110001110010;
assign LUT_4[29882] = 32'b00000000000000000001000000011110;
assign LUT_4[29883] = 32'b11111111111111111010001100010110;
assign LUT_4[29884] = 32'b11111111111111111110100110010110;
assign LUT_4[29885] = 32'b11111111111111110111110010001110;
assign LUT_4[29886] = 32'b11111111111111111110000000111010;
assign LUT_4[29887] = 32'b11111111111111110111001100110010;
assign LUT_4[29888] = 32'b00000000000000001101100100000100;
assign LUT_4[29889] = 32'b00000000000000000110101111111100;
assign LUT_4[29890] = 32'b00000000000000001100111110101000;
assign LUT_4[29891] = 32'b00000000000000000110001010100000;
assign LUT_4[29892] = 32'b00000000000000001010100100100000;
assign LUT_4[29893] = 32'b00000000000000000011110000011000;
assign LUT_4[29894] = 32'b00000000000000001001111111000100;
assign LUT_4[29895] = 32'b00000000000000000011001010111100;
assign LUT_4[29896] = 32'b00000000000000000110110000011001;
assign LUT_4[29897] = 32'b11111111111111111111111100010001;
assign LUT_4[29898] = 32'b00000000000000000110001010111101;
assign LUT_4[29899] = 32'b11111111111111111111010110110101;
assign LUT_4[29900] = 32'b00000000000000000011110000110101;
assign LUT_4[29901] = 32'b11111111111111111100111100101101;
assign LUT_4[29902] = 32'b00000000000000000011001011011001;
assign LUT_4[29903] = 32'b11111111111111111100010111010001;
assign LUT_4[29904] = 32'b00000000000000001011010101110010;
assign LUT_4[29905] = 32'b00000000000000000100100001101010;
assign LUT_4[29906] = 32'b00000000000000001010110000010110;
assign LUT_4[29907] = 32'b00000000000000000011111100001110;
assign LUT_4[29908] = 32'b00000000000000001000010110001110;
assign LUT_4[29909] = 32'b00000000000000000001100010000110;
assign LUT_4[29910] = 32'b00000000000000000111110000110010;
assign LUT_4[29911] = 32'b00000000000000000000111100101010;
assign LUT_4[29912] = 32'b00000000000000000100100010000111;
assign LUT_4[29913] = 32'b11111111111111111101101101111111;
assign LUT_4[29914] = 32'b00000000000000000011111100101011;
assign LUT_4[29915] = 32'b11111111111111111101001000100011;
assign LUT_4[29916] = 32'b00000000000000000001100010100011;
assign LUT_4[29917] = 32'b11111111111111111010101110011011;
assign LUT_4[29918] = 32'b00000000000000000000111101000111;
assign LUT_4[29919] = 32'b11111111111111111010001000111111;
assign LUT_4[29920] = 32'b00000000000000001011111111001011;
assign LUT_4[29921] = 32'b00000000000000000101001011000011;
assign LUT_4[29922] = 32'b00000000000000001011011001101111;
assign LUT_4[29923] = 32'b00000000000000000100100101100111;
assign LUT_4[29924] = 32'b00000000000000001000111111100111;
assign LUT_4[29925] = 32'b00000000000000000010001011011111;
assign LUT_4[29926] = 32'b00000000000000001000011010001011;
assign LUT_4[29927] = 32'b00000000000000000001100110000011;
assign LUT_4[29928] = 32'b00000000000000000101001011100000;
assign LUT_4[29929] = 32'b11111111111111111110010111011000;
assign LUT_4[29930] = 32'b00000000000000000100100110000100;
assign LUT_4[29931] = 32'b11111111111111111101110001111100;
assign LUT_4[29932] = 32'b00000000000000000010001011111100;
assign LUT_4[29933] = 32'b11111111111111111011010111110100;
assign LUT_4[29934] = 32'b00000000000000000001100110100000;
assign LUT_4[29935] = 32'b11111111111111111010110010011000;
assign LUT_4[29936] = 32'b00000000000000001001110000111001;
assign LUT_4[29937] = 32'b00000000000000000010111100110001;
assign LUT_4[29938] = 32'b00000000000000001001001011011101;
assign LUT_4[29939] = 32'b00000000000000000010010111010101;
assign LUT_4[29940] = 32'b00000000000000000110110001010101;
assign LUT_4[29941] = 32'b11111111111111111111111101001101;
assign LUT_4[29942] = 32'b00000000000000000110001011111001;
assign LUT_4[29943] = 32'b11111111111111111111010111110001;
assign LUT_4[29944] = 32'b00000000000000000010111101001110;
assign LUT_4[29945] = 32'b11111111111111111100001001000110;
assign LUT_4[29946] = 32'b00000000000000000010010111110010;
assign LUT_4[29947] = 32'b11111111111111111011100011101010;
assign LUT_4[29948] = 32'b11111111111111111111111101101010;
assign LUT_4[29949] = 32'b11111111111111111001001001100010;
assign LUT_4[29950] = 32'b11111111111111111111011000001110;
assign LUT_4[29951] = 32'b11111111111111111000100100000110;
assign LUT_4[29952] = 32'b00000000000000001110100010001011;
assign LUT_4[29953] = 32'b00000000000000000111101110000011;
assign LUT_4[29954] = 32'b00000000000000001101111100101111;
assign LUT_4[29955] = 32'b00000000000000000111001000100111;
assign LUT_4[29956] = 32'b00000000000000001011100010100111;
assign LUT_4[29957] = 32'b00000000000000000100101110011111;
assign LUT_4[29958] = 32'b00000000000000001010111101001011;
assign LUT_4[29959] = 32'b00000000000000000100001001000011;
assign LUT_4[29960] = 32'b00000000000000000111101110100000;
assign LUT_4[29961] = 32'b00000000000000000000111010011000;
assign LUT_4[29962] = 32'b00000000000000000111001001000100;
assign LUT_4[29963] = 32'b00000000000000000000010100111100;
assign LUT_4[29964] = 32'b00000000000000000100101110111100;
assign LUT_4[29965] = 32'b11111111111111111101111010110100;
assign LUT_4[29966] = 32'b00000000000000000100001001100000;
assign LUT_4[29967] = 32'b11111111111111111101010101011000;
assign LUT_4[29968] = 32'b00000000000000001100010011111001;
assign LUT_4[29969] = 32'b00000000000000000101011111110001;
assign LUT_4[29970] = 32'b00000000000000001011101110011101;
assign LUT_4[29971] = 32'b00000000000000000100111010010101;
assign LUT_4[29972] = 32'b00000000000000001001010100010101;
assign LUT_4[29973] = 32'b00000000000000000010100000001101;
assign LUT_4[29974] = 32'b00000000000000001000101110111001;
assign LUT_4[29975] = 32'b00000000000000000001111010110001;
assign LUT_4[29976] = 32'b00000000000000000101100000001110;
assign LUT_4[29977] = 32'b11111111111111111110101100000110;
assign LUT_4[29978] = 32'b00000000000000000100111010110010;
assign LUT_4[29979] = 32'b11111111111111111110000110101010;
assign LUT_4[29980] = 32'b00000000000000000010100000101010;
assign LUT_4[29981] = 32'b11111111111111111011101100100010;
assign LUT_4[29982] = 32'b00000000000000000001111011001110;
assign LUT_4[29983] = 32'b11111111111111111011000111000110;
assign LUT_4[29984] = 32'b00000000000000001100111101010010;
assign LUT_4[29985] = 32'b00000000000000000110001001001010;
assign LUT_4[29986] = 32'b00000000000000001100010111110110;
assign LUT_4[29987] = 32'b00000000000000000101100011101110;
assign LUT_4[29988] = 32'b00000000000000001001111101101110;
assign LUT_4[29989] = 32'b00000000000000000011001001100110;
assign LUT_4[29990] = 32'b00000000000000001001011000010010;
assign LUT_4[29991] = 32'b00000000000000000010100100001010;
assign LUT_4[29992] = 32'b00000000000000000110001001100111;
assign LUT_4[29993] = 32'b11111111111111111111010101011111;
assign LUT_4[29994] = 32'b00000000000000000101100100001011;
assign LUT_4[29995] = 32'b11111111111111111110110000000011;
assign LUT_4[29996] = 32'b00000000000000000011001010000011;
assign LUT_4[29997] = 32'b11111111111111111100010101111011;
assign LUT_4[29998] = 32'b00000000000000000010100100100111;
assign LUT_4[29999] = 32'b11111111111111111011110000011111;
assign LUT_4[30000] = 32'b00000000000000001010101111000000;
assign LUT_4[30001] = 32'b00000000000000000011111010111000;
assign LUT_4[30002] = 32'b00000000000000001010001001100100;
assign LUT_4[30003] = 32'b00000000000000000011010101011100;
assign LUT_4[30004] = 32'b00000000000000000111101111011100;
assign LUT_4[30005] = 32'b00000000000000000000111011010100;
assign LUT_4[30006] = 32'b00000000000000000111001010000000;
assign LUT_4[30007] = 32'b00000000000000000000010101111000;
assign LUT_4[30008] = 32'b00000000000000000011111011010101;
assign LUT_4[30009] = 32'b11111111111111111101000111001101;
assign LUT_4[30010] = 32'b00000000000000000011010101111001;
assign LUT_4[30011] = 32'b11111111111111111100100001110001;
assign LUT_4[30012] = 32'b00000000000000000000111011110001;
assign LUT_4[30013] = 32'b11111111111111111010000111101001;
assign LUT_4[30014] = 32'b00000000000000000000010110010101;
assign LUT_4[30015] = 32'b11111111111111111001100010001101;
assign LUT_4[30016] = 32'b00000000000000001111111001011111;
assign LUT_4[30017] = 32'b00000000000000001001000101010111;
assign LUT_4[30018] = 32'b00000000000000001111010100000011;
assign LUT_4[30019] = 32'b00000000000000001000011111111011;
assign LUT_4[30020] = 32'b00000000000000001100111001111011;
assign LUT_4[30021] = 32'b00000000000000000110000101110011;
assign LUT_4[30022] = 32'b00000000000000001100010100011111;
assign LUT_4[30023] = 32'b00000000000000000101100000010111;
assign LUT_4[30024] = 32'b00000000000000001001000101110100;
assign LUT_4[30025] = 32'b00000000000000000010010001101100;
assign LUT_4[30026] = 32'b00000000000000001000100000011000;
assign LUT_4[30027] = 32'b00000000000000000001101100010000;
assign LUT_4[30028] = 32'b00000000000000000110000110010000;
assign LUT_4[30029] = 32'b11111111111111111111010010001000;
assign LUT_4[30030] = 32'b00000000000000000101100000110100;
assign LUT_4[30031] = 32'b11111111111111111110101100101100;
assign LUT_4[30032] = 32'b00000000000000001101101011001101;
assign LUT_4[30033] = 32'b00000000000000000110110111000101;
assign LUT_4[30034] = 32'b00000000000000001101000101110001;
assign LUT_4[30035] = 32'b00000000000000000110010001101001;
assign LUT_4[30036] = 32'b00000000000000001010101011101001;
assign LUT_4[30037] = 32'b00000000000000000011110111100001;
assign LUT_4[30038] = 32'b00000000000000001010000110001101;
assign LUT_4[30039] = 32'b00000000000000000011010010000101;
assign LUT_4[30040] = 32'b00000000000000000110110111100010;
assign LUT_4[30041] = 32'b00000000000000000000000011011010;
assign LUT_4[30042] = 32'b00000000000000000110010010000110;
assign LUT_4[30043] = 32'b11111111111111111111011101111110;
assign LUT_4[30044] = 32'b00000000000000000011110111111110;
assign LUT_4[30045] = 32'b11111111111111111101000011110110;
assign LUT_4[30046] = 32'b00000000000000000011010010100010;
assign LUT_4[30047] = 32'b11111111111111111100011110011010;
assign LUT_4[30048] = 32'b00000000000000001110010100100110;
assign LUT_4[30049] = 32'b00000000000000000111100000011110;
assign LUT_4[30050] = 32'b00000000000000001101101111001010;
assign LUT_4[30051] = 32'b00000000000000000110111011000010;
assign LUT_4[30052] = 32'b00000000000000001011010101000010;
assign LUT_4[30053] = 32'b00000000000000000100100000111010;
assign LUT_4[30054] = 32'b00000000000000001010101111100110;
assign LUT_4[30055] = 32'b00000000000000000011111011011110;
assign LUT_4[30056] = 32'b00000000000000000111100000111011;
assign LUT_4[30057] = 32'b00000000000000000000101100110011;
assign LUT_4[30058] = 32'b00000000000000000110111011011111;
assign LUT_4[30059] = 32'b00000000000000000000000111010111;
assign LUT_4[30060] = 32'b00000000000000000100100001010111;
assign LUT_4[30061] = 32'b11111111111111111101101101001111;
assign LUT_4[30062] = 32'b00000000000000000011111011111011;
assign LUT_4[30063] = 32'b11111111111111111101000111110011;
assign LUT_4[30064] = 32'b00000000000000001100000110010100;
assign LUT_4[30065] = 32'b00000000000000000101010010001100;
assign LUT_4[30066] = 32'b00000000000000001011100000111000;
assign LUT_4[30067] = 32'b00000000000000000100101100110000;
assign LUT_4[30068] = 32'b00000000000000001001000110110000;
assign LUT_4[30069] = 32'b00000000000000000010010010101000;
assign LUT_4[30070] = 32'b00000000000000001000100001010100;
assign LUT_4[30071] = 32'b00000000000000000001101101001100;
assign LUT_4[30072] = 32'b00000000000000000101010010101001;
assign LUT_4[30073] = 32'b11111111111111111110011110100001;
assign LUT_4[30074] = 32'b00000000000000000100101101001101;
assign LUT_4[30075] = 32'b11111111111111111101111001000101;
assign LUT_4[30076] = 32'b00000000000000000010010011000101;
assign LUT_4[30077] = 32'b11111111111111111011011110111101;
assign LUT_4[30078] = 32'b00000000000000000001101101101001;
assign LUT_4[30079] = 32'b11111111111111111010111001100001;
assign LUT_4[30080] = 32'b00000000000000010001001000010011;
assign LUT_4[30081] = 32'b00000000000000001010010100001011;
assign LUT_4[30082] = 32'b00000000000000010000100010110111;
assign LUT_4[30083] = 32'b00000000000000001001101110101111;
assign LUT_4[30084] = 32'b00000000000000001110001000101111;
assign LUT_4[30085] = 32'b00000000000000000111010100100111;
assign LUT_4[30086] = 32'b00000000000000001101100011010011;
assign LUT_4[30087] = 32'b00000000000000000110101111001011;
assign LUT_4[30088] = 32'b00000000000000001010010100101000;
assign LUT_4[30089] = 32'b00000000000000000011100000100000;
assign LUT_4[30090] = 32'b00000000000000001001101111001100;
assign LUT_4[30091] = 32'b00000000000000000010111011000100;
assign LUT_4[30092] = 32'b00000000000000000111010101000100;
assign LUT_4[30093] = 32'b00000000000000000000100000111100;
assign LUT_4[30094] = 32'b00000000000000000110101111101000;
assign LUT_4[30095] = 32'b11111111111111111111111011100000;
assign LUT_4[30096] = 32'b00000000000000001110111010000001;
assign LUT_4[30097] = 32'b00000000000000001000000101111001;
assign LUT_4[30098] = 32'b00000000000000001110010100100101;
assign LUT_4[30099] = 32'b00000000000000000111100000011101;
assign LUT_4[30100] = 32'b00000000000000001011111010011101;
assign LUT_4[30101] = 32'b00000000000000000101000110010101;
assign LUT_4[30102] = 32'b00000000000000001011010101000001;
assign LUT_4[30103] = 32'b00000000000000000100100000111001;
assign LUT_4[30104] = 32'b00000000000000001000000110010110;
assign LUT_4[30105] = 32'b00000000000000000001010010001110;
assign LUT_4[30106] = 32'b00000000000000000111100000111010;
assign LUT_4[30107] = 32'b00000000000000000000101100110010;
assign LUT_4[30108] = 32'b00000000000000000101000110110010;
assign LUT_4[30109] = 32'b11111111111111111110010010101010;
assign LUT_4[30110] = 32'b00000000000000000100100001010110;
assign LUT_4[30111] = 32'b11111111111111111101101101001110;
assign LUT_4[30112] = 32'b00000000000000001111100011011010;
assign LUT_4[30113] = 32'b00000000000000001000101111010010;
assign LUT_4[30114] = 32'b00000000000000001110111101111110;
assign LUT_4[30115] = 32'b00000000000000001000001001110110;
assign LUT_4[30116] = 32'b00000000000000001100100011110110;
assign LUT_4[30117] = 32'b00000000000000000101101111101110;
assign LUT_4[30118] = 32'b00000000000000001011111110011010;
assign LUT_4[30119] = 32'b00000000000000000101001010010010;
assign LUT_4[30120] = 32'b00000000000000001000101111101111;
assign LUT_4[30121] = 32'b00000000000000000001111011100111;
assign LUT_4[30122] = 32'b00000000000000001000001010010011;
assign LUT_4[30123] = 32'b00000000000000000001010110001011;
assign LUT_4[30124] = 32'b00000000000000000101110000001011;
assign LUT_4[30125] = 32'b11111111111111111110111100000011;
assign LUT_4[30126] = 32'b00000000000000000101001010101111;
assign LUT_4[30127] = 32'b11111111111111111110010110100111;
assign LUT_4[30128] = 32'b00000000000000001101010101001000;
assign LUT_4[30129] = 32'b00000000000000000110100001000000;
assign LUT_4[30130] = 32'b00000000000000001100101111101100;
assign LUT_4[30131] = 32'b00000000000000000101111011100100;
assign LUT_4[30132] = 32'b00000000000000001010010101100100;
assign LUT_4[30133] = 32'b00000000000000000011100001011100;
assign LUT_4[30134] = 32'b00000000000000001001110000001000;
assign LUT_4[30135] = 32'b00000000000000000010111100000000;
assign LUT_4[30136] = 32'b00000000000000000110100001011101;
assign LUT_4[30137] = 32'b11111111111111111111101101010101;
assign LUT_4[30138] = 32'b00000000000000000101111100000001;
assign LUT_4[30139] = 32'b11111111111111111111000111111001;
assign LUT_4[30140] = 32'b00000000000000000011100001111001;
assign LUT_4[30141] = 32'b11111111111111111100101101110001;
assign LUT_4[30142] = 32'b00000000000000000010111100011101;
assign LUT_4[30143] = 32'b11111111111111111100001000010101;
assign LUT_4[30144] = 32'b00000000000000010010011111100111;
assign LUT_4[30145] = 32'b00000000000000001011101011011111;
assign LUT_4[30146] = 32'b00000000000000010001111010001011;
assign LUT_4[30147] = 32'b00000000000000001011000110000011;
assign LUT_4[30148] = 32'b00000000000000001111100000000011;
assign LUT_4[30149] = 32'b00000000000000001000101011111011;
assign LUT_4[30150] = 32'b00000000000000001110111010100111;
assign LUT_4[30151] = 32'b00000000000000001000000110011111;
assign LUT_4[30152] = 32'b00000000000000001011101011111100;
assign LUT_4[30153] = 32'b00000000000000000100110111110100;
assign LUT_4[30154] = 32'b00000000000000001011000110100000;
assign LUT_4[30155] = 32'b00000000000000000100010010011000;
assign LUT_4[30156] = 32'b00000000000000001000101100011000;
assign LUT_4[30157] = 32'b00000000000000000001111000010000;
assign LUT_4[30158] = 32'b00000000000000001000000110111100;
assign LUT_4[30159] = 32'b00000000000000000001010010110100;
assign LUT_4[30160] = 32'b00000000000000010000010001010101;
assign LUT_4[30161] = 32'b00000000000000001001011101001101;
assign LUT_4[30162] = 32'b00000000000000001111101011111001;
assign LUT_4[30163] = 32'b00000000000000001000110111110001;
assign LUT_4[30164] = 32'b00000000000000001101010001110001;
assign LUT_4[30165] = 32'b00000000000000000110011101101001;
assign LUT_4[30166] = 32'b00000000000000001100101100010101;
assign LUT_4[30167] = 32'b00000000000000000101111000001101;
assign LUT_4[30168] = 32'b00000000000000001001011101101010;
assign LUT_4[30169] = 32'b00000000000000000010101001100010;
assign LUT_4[30170] = 32'b00000000000000001000111000001110;
assign LUT_4[30171] = 32'b00000000000000000010000100000110;
assign LUT_4[30172] = 32'b00000000000000000110011110000110;
assign LUT_4[30173] = 32'b11111111111111111111101001111110;
assign LUT_4[30174] = 32'b00000000000000000101111000101010;
assign LUT_4[30175] = 32'b11111111111111111111000100100010;
assign LUT_4[30176] = 32'b00000000000000010000111010101110;
assign LUT_4[30177] = 32'b00000000000000001010000110100110;
assign LUT_4[30178] = 32'b00000000000000010000010101010010;
assign LUT_4[30179] = 32'b00000000000000001001100001001010;
assign LUT_4[30180] = 32'b00000000000000001101111011001010;
assign LUT_4[30181] = 32'b00000000000000000111000111000010;
assign LUT_4[30182] = 32'b00000000000000001101010101101110;
assign LUT_4[30183] = 32'b00000000000000000110100001100110;
assign LUT_4[30184] = 32'b00000000000000001010000111000011;
assign LUT_4[30185] = 32'b00000000000000000011010010111011;
assign LUT_4[30186] = 32'b00000000000000001001100001100111;
assign LUT_4[30187] = 32'b00000000000000000010101101011111;
assign LUT_4[30188] = 32'b00000000000000000111000111011111;
assign LUT_4[30189] = 32'b00000000000000000000010011010111;
assign LUT_4[30190] = 32'b00000000000000000110100010000011;
assign LUT_4[30191] = 32'b11111111111111111111101101111011;
assign LUT_4[30192] = 32'b00000000000000001110101100011100;
assign LUT_4[30193] = 32'b00000000000000000111111000010100;
assign LUT_4[30194] = 32'b00000000000000001110000111000000;
assign LUT_4[30195] = 32'b00000000000000000111010010111000;
assign LUT_4[30196] = 32'b00000000000000001011101100111000;
assign LUT_4[30197] = 32'b00000000000000000100111000110000;
assign LUT_4[30198] = 32'b00000000000000001011000111011100;
assign LUT_4[30199] = 32'b00000000000000000100010011010100;
assign LUT_4[30200] = 32'b00000000000000000111111000110001;
assign LUT_4[30201] = 32'b00000000000000000001000100101001;
assign LUT_4[30202] = 32'b00000000000000000111010011010101;
assign LUT_4[30203] = 32'b00000000000000000000011111001101;
assign LUT_4[30204] = 32'b00000000000000000100111001001101;
assign LUT_4[30205] = 32'b11111111111111111110000101000101;
assign LUT_4[30206] = 32'b00000000000000000100010011110001;
assign LUT_4[30207] = 32'b11111111111111111101011111101001;
assign LUT_4[30208] = 32'b00000000000000001000101010110000;
assign LUT_4[30209] = 32'b00000000000000000001110110101000;
assign LUT_4[30210] = 32'b00000000000000001000000101010100;
assign LUT_4[30211] = 32'b00000000000000000001010001001100;
assign LUT_4[30212] = 32'b00000000000000000101101011001100;
assign LUT_4[30213] = 32'b11111111111111111110110111000100;
assign LUT_4[30214] = 32'b00000000000000000101000101110000;
assign LUT_4[30215] = 32'b11111111111111111110010001101000;
assign LUT_4[30216] = 32'b00000000000000000001110111000101;
assign LUT_4[30217] = 32'b11111111111111111011000010111101;
assign LUT_4[30218] = 32'b00000000000000000001010001101001;
assign LUT_4[30219] = 32'b11111111111111111010011101100001;
assign LUT_4[30220] = 32'b11111111111111111110110111100001;
assign LUT_4[30221] = 32'b11111111111111111000000011011001;
assign LUT_4[30222] = 32'b11111111111111111110010010000101;
assign LUT_4[30223] = 32'b11111111111111110111011101111101;
assign LUT_4[30224] = 32'b00000000000000000110011100011110;
assign LUT_4[30225] = 32'b11111111111111111111101000010110;
assign LUT_4[30226] = 32'b00000000000000000101110111000010;
assign LUT_4[30227] = 32'b11111111111111111111000010111010;
assign LUT_4[30228] = 32'b00000000000000000011011100111010;
assign LUT_4[30229] = 32'b11111111111111111100101000110010;
assign LUT_4[30230] = 32'b00000000000000000010110111011110;
assign LUT_4[30231] = 32'b11111111111111111100000011010110;
assign LUT_4[30232] = 32'b11111111111111111111101000110011;
assign LUT_4[30233] = 32'b11111111111111111000110100101011;
assign LUT_4[30234] = 32'b11111111111111111111000011010111;
assign LUT_4[30235] = 32'b11111111111111111000001111001111;
assign LUT_4[30236] = 32'b11111111111111111100101001001111;
assign LUT_4[30237] = 32'b11111111111111110101110101000111;
assign LUT_4[30238] = 32'b11111111111111111100000011110011;
assign LUT_4[30239] = 32'b11111111111111110101001111101011;
assign LUT_4[30240] = 32'b00000000000000000111000101110111;
assign LUT_4[30241] = 32'b00000000000000000000010001101111;
assign LUT_4[30242] = 32'b00000000000000000110100000011011;
assign LUT_4[30243] = 32'b11111111111111111111101100010011;
assign LUT_4[30244] = 32'b00000000000000000100000110010011;
assign LUT_4[30245] = 32'b11111111111111111101010010001011;
assign LUT_4[30246] = 32'b00000000000000000011100000110111;
assign LUT_4[30247] = 32'b11111111111111111100101100101111;
assign LUT_4[30248] = 32'b00000000000000000000010010001100;
assign LUT_4[30249] = 32'b11111111111111111001011110000100;
assign LUT_4[30250] = 32'b11111111111111111111101100110000;
assign LUT_4[30251] = 32'b11111111111111111000111000101000;
assign LUT_4[30252] = 32'b11111111111111111101010010101000;
assign LUT_4[30253] = 32'b11111111111111110110011110100000;
assign LUT_4[30254] = 32'b11111111111111111100101101001100;
assign LUT_4[30255] = 32'b11111111111111110101111001000100;
assign LUT_4[30256] = 32'b00000000000000000100110111100101;
assign LUT_4[30257] = 32'b11111111111111111110000011011101;
assign LUT_4[30258] = 32'b00000000000000000100010010001001;
assign LUT_4[30259] = 32'b11111111111111111101011110000001;
assign LUT_4[30260] = 32'b00000000000000000001111000000001;
assign LUT_4[30261] = 32'b11111111111111111011000011111001;
assign LUT_4[30262] = 32'b00000000000000000001010010100101;
assign LUT_4[30263] = 32'b11111111111111111010011110011101;
assign LUT_4[30264] = 32'b11111111111111111110000011111010;
assign LUT_4[30265] = 32'b11111111111111110111001111110010;
assign LUT_4[30266] = 32'b11111111111111111101011110011110;
assign LUT_4[30267] = 32'b11111111111111110110101010010110;
assign LUT_4[30268] = 32'b11111111111111111011000100010110;
assign LUT_4[30269] = 32'b11111111111111110100010000001110;
assign LUT_4[30270] = 32'b11111111111111111010011110111010;
assign LUT_4[30271] = 32'b11111111111111110011101010110010;
assign LUT_4[30272] = 32'b00000000000000001010000010000100;
assign LUT_4[30273] = 32'b00000000000000000011001101111100;
assign LUT_4[30274] = 32'b00000000000000001001011100101000;
assign LUT_4[30275] = 32'b00000000000000000010101000100000;
assign LUT_4[30276] = 32'b00000000000000000111000010100000;
assign LUT_4[30277] = 32'b00000000000000000000001110011000;
assign LUT_4[30278] = 32'b00000000000000000110011101000100;
assign LUT_4[30279] = 32'b11111111111111111111101000111100;
assign LUT_4[30280] = 32'b00000000000000000011001110011001;
assign LUT_4[30281] = 32'b11111111111111111100011010010001;
assign LUT_4[30282] = 32'b00000000000000000010101000111101;
assign LUT_4[30283] = 32'b11111111111111111011110100110101;
assign LUT_4[30284] = 32'b00000000000000000000001110110101;
assign LUT_4[30285] = 32'b11111111111111111001011010101101;
assign LUT_4[30286] = 32'b11111111111111111111101001011001;
assign LUT_4[30287] = 32'b11111111111111111000110101010001;
assign LUT_4[30288] = 32'b00000000000000000111110011110010;
assign LUT_4[30289] = 32'b00000000000000000000111111101010;
assign LUT_4[30290] = 32'b00000000000000000111001110010110;
assign LUT_4[30291] = 32'b00000000000000000000011010001110;
assign LUT_4[30292] = 32'b00000000000000000100110100001110;
assign LUT_4[30293] = 32'b11111111111111111110000000000110;
assign LUT_4[30294] = 32'b00000000000000000100001110110010;
assign LUT_4[30295] = 32'b11111111111111111101011010101010;
assign LUT_4[30296] = 32'b00000000000000000001000000000111;
assign LUT_4[30297] = 32'b11111111111111111010001011111111;
assign LUT_4[30298] = 32'b00000000000000000000011010101011;
assign LUT_4[30299] = 32'b11111111111111111001100110100011;
assign LUT_4[30300] = 32'b11111111111111111110000000100011;
assign LUT_4[30301] = 32'b11111111111111110111001100011011;
assign LUT_4[30302] = 32'b11111111111111111101011011000111;
assign LUT_4[30303] = 32'b11111111111111110110100110111111;
assign LUT_4[30304] = 32'b00000000000000001000011101001011;
assign LUT_4[30305] = 32'b00000000000000000001101001000011;
assign LUT_4[30306] = 32'b00000000000000000111110111101111;
assign LUT_4[30307] = 32'b00000000000000000001000011100111;
assign LUT_4[30308] = 32'b00000000000000000101011101100111;
assign LUT_4[30309] = 32'b11111111111111111110101001011111;
assign LUT_4[30310] = 32'b00000000000000000100111000001011;
assign LUT_4[30311] = 32'b11111111111111111110000100000011;
assign LUT_4[30312] = 32'b00000000000000000001101001100000;
assign LUT_4[30313] = 32'b11111111111111111010110101011000;
assign LUT_4[30314] = 32'b00000000000000000001000100000100;
assign LUT_4[30315] = 32'b11111111111111111010001111111100;
assign LUT_4[30316] = 32'b11111111111111111110101001111100;
assign LUT_4[30317] = 32'b11111111111111110111110101110100;
assign LUT_4[30318] = 32'b11111111111111111110000100100000;
assign LUT_4[30319] = 32'b11111111111111110111010000011000;
assign LUT_4[30320] = 32'b00000000000000000110001110111001;
assign LUT_4[30321] = 32'b11111111111111111111011010110001;
assign LUT_4[30322] = 32'b00000000000000000101101001011101;
assign LUT_4[30323] = 32'b11111111111111111110110101010101;
assign LUT_4[30324] = 32'b00000000000000000011001111010101;
assign LUT_4[30325] = 32'b11111111111111111100011011001101;
assign LUT_4[30326] = 32'b00000000000000000010101001111001;
assign LUT_4[30327] = 32'b11111111111111111011110101110001;
assign LUT_4[30328] = 32'b11111111111111111111011011001110;
assign LUT_4[30329] = 32'b11111111111111111000100111000110;
assign LUT_4[30330] = 32'b11111111111111111110110101110010;
assign LUT_4[30331] = 32'b11111111111111111000000001101010;
assign LUT_4[30332] = 32'b11111111111111111100011011101010;
assign LUT_4[30333] = 32'b11111111111111110101100111100010;
assign LUT_4[30334] = 32'b11111111111111111011110110001110;
assign LUT_4[30335] = 32'b11111111111111110101000010000110;
assign LUT_4[30336] = 32'b00000000000000001011010000111000;
assign LUT_4[30337] = 32'b00000000000000000100011100110000;
assign LUT_4[30338] = 32'b00000000000000001010101011011100;
assign LUT_4[30339] = 32'b00000000000000000011110111010100;
assign LUT_4[30340] = 32'b00000000000000001000010001010100;
assign LUT_4[30341] = 32'b00000000000000000001011101001100;
assign LUT_4[30342] = 32'b00000000000000000111101011111000;
assign LUT_4[30343] = 32'b00000000000000000000110111110000;
assign LUT_4[30344] = 32'b00000000000000000100011101001101;
assign LUT_4[30345] = 32'b11111111111111111101101001000101;
assign LUT_4[30346] = 32'b00000000000000000011110111110001;
assign LUT_4[30347] = 32'b11111111111111111101000011101001;
assign LUT_4[30348] = 32'b00000000000000000001011101101001;
assign LUT_4[30349] = 32'b11111111111111111010101001100001;
assign LUT_4[30350] = 32'b00000000000000000000111000001101;
assign LUT_4[30351] = 32'b11111111111111111010000100000101;
assign LUT_4[30352] = 32'b00000000000000001001000010100110;
assign LUT_4[30353] = 32'b00000000000000000010001110011110;
assign LUT_4[30354] = 32'b00000000000000001000011101001010;
assign LUT_4[30355] = 32'b00000000000000000001101001000010;
assign LUT_4[30356] = 32'b00000000000000000110000011000010;
assign LUT_4[30357] = 32'b11111111111111111111001110111010;
assign LUT_4[30358] = 32'b00000000000000000101011101100110;
assign LUT_4[30359] = 32'b11111111111111111110101001011110;
assign LUT_4[30360] = 32'b00000000000000000010001110111011;
assign LUT_4[30361] = 32'b11111111111111111011011010110011;
assign LUT_4[30362] = 32'b00000000000000000001101001011111;
assign LUT_4[30363] = 32'b11111111111111111010110101010111;
assign LUT_4[30364] = 32'b11111111111111111111001111010111;
assign LUT_4[30365] = 32'b11111111111111111000011011001111;
assign LUT_4[30366] = 32'b11111111111111111110101001111011;
assign LUT_4[30367] = 32'b11111111111111110111110101110011;
assign LUT_4[30368] = 32'b00000000000000001001101011111111;
assign LUT_4[30369] = 32'b00000000000000000010110111110111;
assign LUT_4[30370] = 32'b00000000000000001001000110100011;
assign LUT_4[30371] = 32'b00000000000000000010010010011011;
assign LUT_4[30372] = 32'b00000000000000000110101100011011;
assign LUT_4[30373] = 32'b11111111111111111111111000010011;
assign LUT_4[30374] = 32'b00000000000000000110000110111111;
assign LUT_4[30375] = 32'b11111111111111111111010010110111;
assign LUT_4[30376] = 32'b00000000000000000010111000010100;
assign LUT_4[30377] = 32'b11111111111111111100000100001100;
assign LUT_4[30378] = 32'b00000000000000000010010010111000;
assign LUT_4[30379] = 32'b11111111111111111011011110110000;
assign LUT_4[30380] = 32'b11111111111111111111111000110000;
assign LUT_4[30381] = 32'b11111111111111111001000100101000;
assign LUT_4[30382] = 32'b11111111111111111111010011010100;
assign LUT_4[30383] = 32'b11111111111111111000011111001100;
assign LUT_4[30384] = 32'b00000000000000000111011101101101;
assign LUT_4[30385] = 32'b00000000000000000000101001100101;
assign LUT_4[30386] = 32'b00000000000000000110111000010001;
assign LUT_4[30387] = 32'b00000000000000000000000100001001;
assign LUT_4[30388] = 32'b00000000000000000100011110001001;
assign LUT_4[30389] = 32'b11111111111111111101101010000001;
assign LUT_4[30390] = 32'b00000000000000000011111000101101;
assign LUT_4[30391] = 32'b11111111111111111101000100100101;
assign LUT_4[30392] = 32'b00000000000000000000101010000010;
assign LUT_4[30393] = 32'b11111111111111111001110101111010;
assign LUT_4[30394] = 32'b00000000000000000000000100100110;
assign LUT_4[30395] = 32'b11111111111111111001010000011110;
assign LUT_4[30396] = 32'b11111111111111111101101010011110;
assign LUT_4[30397] = 32'b11111111111111110110110110010110;
assign LUT_4[30398] = 32'b11111111111111111101000101000010;
assign LUT_4[30399] = 32'b11111111111111110110010000111010;
assign LUT_4[30400] = 32'b00000000000000001100101000001100;
assign LUT_4[30401] = 32'b00000000000000000101110100000100;
assign LUT_4[30402] = 32'b00000000000000001100000010110000;
assign LUT_4[30403] = 32'b00000000000000000101001110101000;
assign LUT_4[30404] = 32'b00000000000000001001101000101000;
assign LUT_4[30405] = 32'b00000000000000000010110100100000;
assign LUT_4[30406] = 32'b00000000000000001001000011001100;
assign LUT_4[30407] = 32'b00000000000000000010001111000100;
assign LUT_4[30408] = 32'b00000000000000000101110100100001;
assign LUT_4[30409] = 32'b11111111111111111111000000011001;
assign LUT_4[30410] = 32'b00000000000000000101001111000101;
assign LUT_4[30411] = 32'b11111111111111111110011010111101;
assign LUT_4[30412] = 32'b00000000000000000010110100111101;
assign LUT_4[30413] = 32'b11111111111111111100000000110101;
assign LUT_4[30414] = 32'b00000000000000000010001111100001;
assign LUT_4[30415] = 32'b11111111111111111011011011011001;
assign LUT_4[30416] = 32'b00000000000000001010011001111010;
assign LUT_4[30417] = 32'b00000000000000000011100101110010;
assign LUT_4[30418] = 32'b00000000000000001001110100011110;
assign LUT_4[30419] = 32'b00000000000000000011000000010110;
assign LUT_4[30420] = 32'b00000000000000000111011010010110;
assign LUT_4[30421] = 32'b00000000000000000000100110001110;
assign LUT_4[30422] = 32'b00000000000000000110110100111010;
assign LUT_4[30423] = 32'b00000000000000000000000000110010;
assign LUT_4[30424] = 32'b00000000000000000011100110001111;
assign LUT_4[30425] = 32'b11111111111111111100110010000111;
assign LUT_4[30426] = 32'b00000000000000000011000000110011;
assign LUT_4[30427] = 32'b11111111111111111100001100101011;
assign LUT_4[30428] = 32'b00000000000000000000100110101011;
assign LUT_4[30429] = 32'b11111111111111111001110010100011;
assign LUT_4[30430] = 32'b00000000000000000000000001001111;
assign LUT_4[30431] = 32'b11111111111111111001001101000111;
assign LUT_4[30432] = 32'b00000000000000001011000011010011;
assign LUT_4[30433] = 32'b00000000000000000100001111001011;
assign LUT_4[30434] = 32'b00000000000000001010011101110111;
assign LUT_4[30435] = 32'b00000000000000000011101001101111;
assign LUT_4[30436] = 32'b00000000000000001000000011101111;
assign LUT_4[30437] = 32'b00000000000000000001001111100111;
assign LUT_4[30438] = 32'b00000000000000000111011110010011;
assign LUT_4[30439] = 32'b00000000000000000000101010001011;
assign LUT_4[30440] = 32'b00000000000000000100001111101000;
assign LUT_4[30441] = 32'b11111111111111111101011011100000;
assign LUT_4[30442] = 32'b00000000000000000011101010001100;
assign LUT_4[30443] = 32'b11111111111111111100110110000100;
assign LUT_4[30444] = 32'b00000000000000000001010000000100;
assign LUT_4[30445] = 32'b11111111111111111010011011111100;
assign LUT_4[30446] = 32'b00000000000000000000101010101000;
assign LUT_4[30447] = 32'b11111111111111111001110110100000;
assign LUT_4[30448] = 32'b00000000000000001000110101000001;
assign LUT_4[30449] = 32'b00000000000000000010000000111001;
assign LUT_4[30450] = 32'b00000000000000001000001111100101;
assign LUT_4[30451] = 32'b00000000000000000001011011011101;
assign LUT_4[30452] = 32'b00000000000000000101110101011101;
assign LUT_4[30453] = 32'b11111111111111111111000001010101;
assign LUT_4[30454] = 32'b00000000000000000101010000000001;
assign LUT_4[30455] = 32'b11111111111111111110011011111001;
assign LUT_4[30456] = 32'b00000000000000000010000001010110;
assign LUT_4[30457] = 32'b11111111111111111011001101001110;
assign LUT_4[30458] = 32'b00000000000000000001011011111010;
assign LUT_4[30459] = 32'b11111111111111111010100111110010;
assign LUT_4[30460] = 32'b11111111111111111111000001110010;
assign LUT_4[30461] = 32'b11111111111111111000001101101010;
assign LUT_4[30462] = 32'b11111111111111111110011100010110;
assign LUT_4[30463] = 32'b11111111111111110111101000001110;
assign LUT_4[30464] = 32'b00000000000000001101100110010011;
assign LUT_4[30465] = 32'b00000000000000000110110010001011;
assign LUT_4[30466] = 32'b00000000000000001101000000110111;
assign LUT_4[30467] = 32'b00000000000000000110001100101111;
assign LUT_4[30468] = 32'b00000000000000001010100110101111;
assign LUT_4[30469] = 32'b00000000000000000011110010100111;
assign LUT_4[30470] = 32'b00000000000000001010000001010011;
assign LUT_4[30471] = 32'b00000000000000000011001101001011;
assign LUT_4[30472] = 32'b00000000000000000110110010101000;
assign LUT_4[30473] = 32'b11111111111111111111111110100000;
assign LUT_4[30474] = 32'b00000000000000000110001101001100;
assign LUT_4[30475] = 32'b11111111111111111111011001000100;
assign LUT_4[30476] = 32'b00000000000000000011110011000100;
assign LUT_4[30477] = 32'b11111111111111111100111110111100;
assign LUT_4[30478] = 32'b00000000000000000011001101101000;
assign LUT_4[30479] = 32'b11111111111111111100011001100000;
assign LUT_4[30480] = 32'b00000000000000001011011000000001;
assign LUT_4[30481] = 32'b00000000000000000100100011111001;
assign LUT_4[30482] = 32'b00000000000000001010110010100101;
assign LUT_4[30483] = 32'b00000000000000000011111110011101;
assign LUT_4[30484] = 32'b00000000000000001000011000011101;
assign LUT_4[30485] = 32'b00000000000000000001100100010101;
assign LUT_4[30486] = 32'b00000000000000000111110011000001;
assign LUT_4[30487] = 32'b00000000000000000000111110111001;
assign LUT_4[30488] = 32'b00000000000000000100100100010110;
assign LUT_4[30489] = 32'b11111111111111111101110000001110;
assign LUT_4[30490] = 32'b00000000000000000011111110111010;
assign LUT_4[30491] = 32'b11111111111111111101001010110010;
assign LUT_4[30492] = 32'b00000000000000000001100100110010;
assign LUT_4[30493] = 32'b11111111111111111010110000101010;
assign LUT_4[30494] = 32'b00000000000000000000111111010110;
assign LUT_4[30495] = 32'b11111111111111111010001011001110;
assign LUT_4[30496] = 32'b00000000000000001100000001011010;
assign LUT_4[30497] = 32'b00000000000000000101001101010010;
assign LUT_4[30498] = 32'b00000000000000001011011011111110;
assign LUT_4[30499] = 32'b00000000000000000100100111110110;
assign LUT_4[30500] = 32'b00000000000000001001000001110110;
assign LUT_4[30501] = 32'b00000000000000000010001101101110;
assign LUT_4[30502] = 32'b00000000000000001000011100011010;
assign LUT_4[30503] = 32'b00000000000000000001101000010010;
assign LUT_4[30504] = 32'b00000000000000000101001101101111;
assign LUT_4[30505] = 32'b11111111111111111110011001100111;
assign LUT_4[30506] = 32'b00000000000000000100101000010011;
assign LUT_4[30507] = 32'b11111111111111111101110100001011;
assign LUT_4[30508] = 32'b00000000000000000010001110001011;
assign LUT_4[30509] = 32'b11111111111111111011011010000011;
assign LUT_4[30510] = 32'b00000000000000000001101000101111;
assign LUT_4[30511] = 32'b11111111111111111010110100100111;
assign LUT_4[30512] = 32'b00000000000000001001110011001000;
assign LUT_4[30513] = 32'b00000000000000000010111111000000;
assign LUT_4[30514] = 32'b00000000000000001001001101101100;
assign LUT_4[30515] = 32'b00000000000000000010011001100100;
assign LUT_4[30516] = 32'b00000000000000000110110011100100;
assign LUT_4[30517] = 32'b11111111111111111111111111011100;
assign LUT_4[30518] = 32'b00000000000000000110001110001000;
assign LUT_4[30519] = 32'b11111111111111111111011010000000;
assign LUT_4[30520] = 32'b00000000000000000010111111011101;
assign LUT_4[30521] = 32'b11111111111111111100001011010101;
assign LUT_4[30522] = 32'b00000000000000000010011010000001;
assign LUT_4[30523] = 32'b11111111111111111011100101111001;
assign LUT_4[30524] = 32'b11111111111111111111111111111001;
assign LUT_4[30525] = 32'b11111111111111111001001011110001;
assign LUT_4[30526] = 32'b11111111111111111111011010011101;
assign LUT_4[30527] = 32'b11111111111111111000100110010101;
assign LUT_4[30528] = 32'b00000000000000001110111101100111;
assign LUT_4[30529] = 32'b00000000000000001000001001011111;
assign LUT_4[30530] = 32'b00000000000000001110011000001011;
assign LUT_4[30531] = 32'b00000000000000000111100100000011;
assign LUT_4[30532] = 32'b00000000000000001011111110000011;
assign LUT_4[30533] = 32'b00000000000000000101001001111011;
assign LUT_4[30534] = 32'b00000000000000001011011000100111;
assign LUT_4[30535] = 32'b00000000000000000100100100011111;
assign LUT_4[30536] = 32'b00000000000000001000001001111100;
assign LUT_4[30537] = 32'b00000000000000000001010101110100;
assign LUT_4[30538] = 32'b00000000000000000111100100100000;
assign LUT_4[30539] = 32'b00000000000000000000110000011000;
assign LUT_4[30540] = 32'b00000000000000000101001010011000;
assign LUT_4[30541] = 32'b11111111111111111110010110010000;
assign LUT_4[30542] = 32'b00000000000000000100100100111100;
assign LUT_4[30543] = 32'b11111111111111111101110000110100;
assign LUT_4[30544] = 32'b00000000000000001100101111010101;
assign LUT_4[30545] = 32'b00000000000000000101111011001101;
assign LUT_4[30546] = 32'b00000000000000001100001001111001;
assign LUT_4[30547] = 32'b00000000000000000101010101110001;
assign LUT_4[30548] = 32'b00000000000000001001101111110001;
assign LUT_4[30549] = 32'b00000000000000000010111011101001;
assign LUT_4[30550] = 32'b00000000000000001001001010010101;
assign LUT_4[30551] = 32'b00000000000000000010010110001101;
assign LUT_4[30552] = 32'b00000000000000000101111011101010;
assign LUT_4[30553] = 32'b11111111111111111111000111100010;
assign LUT_4[30554] = 32'b00000000000000000101010110001110;
assign LUT_4[30555] = 32'b11111111111111111110100010000110;
assign LUT_4[30556] = 32'b00000000000000000010111100000110;
assign LUT_4[30557] = 32'b11111111111111111100000111111110;
assign LUT_4[30558] = 32'b00000000000000000010010110101010;
assign LUT_4[30559] = 32'b11111111111111111011100010100010;
assign LUT_4[30560] = 32'b00000000000000001101011000101110;
assign LUT_4[30561] = 32'b00000000000000000110100100100110;
assign LUT_4[30562] = 32'b00000000000000001100110011010010;
assign LUT_4[30563] = 32'b00000000000000000101111111001010;
assign LUT_4[30564] = 32'b00000000000000001010011001001010;
assign LUT_4[30565] = 32'b00000000000000000011100101000010;
assign LUT_4[30566] = 32'b00000000000000001001110011101110;
assign LUT_4[30567] = 32'b00000000000000000010111111100110;
assign LUT_4[30568] = 32'b00000000000000000110100101000011;
assign LUT_4[30569] = 32'b11111111111111111111110000111011;
assign LUT_4[30570] = 32'b00000000000000000101111111100111;
assign LUT_4[30571] = 32'b11111111111111111111001011011111;
assign LUT_4[30572] = 32'b00000000000000000011100101011111;
assign LUT_4[30573] = 32'b11111111111111111100110001010111;
assign LUT_4[30574] = 32'b00000000000000000011000000000011;
assign LUT_4[30575] = 32'b11111111111111111100001011111011;
assign LUT_4[30576] = 32'b00000000000000001011001010011100;
assign LUT_4[30577] = 32'b00000000000000000100010110010100;
assign LUT_4[30578] = 32'b00000000000000001010100101000000;
assign LUT_4[30579] = 32'b00000000000000000011110000111000;
assign LUT_4[30580] = 32'b00000000000000001000001010111000;
assign LUT_4[30581] = 32'b00000000000000000001010110110000;
assign LUT_4[30582] = 32'b00000000000000000111100101011100;
assign LUT_4[30583] = 32'b00000000000000000000110001010100;
assign LUT_4[30584] = 32'b00000000000000000100010110110001;
assign LUT_4[30585] = 32'b11111111111111111101100010101001;
assign LUT_4[30586] = 32'b00000000000000000011110001010101;
assign LUT_4[30587] = 32'b11111111111111111100111101001101;
assign LUT_4[30588] = 32'b00000000000000000001010111001101;
assign LUT_4[30589] = 32'b11111111111111111010100011000101;
assign LUT_4[30590] = 32'b00000000000000000000110001110001;
assign LUT_4[30591] = 32'b11111111111111111001111101101001;
assign LUT_4[30592] = 32'b00000000000000010000001100011011;
assign LUT_4[30593] = 32'b00000000000000001001011000010011;
assign LUT_4[30594] = 32'b00000000000000001111100110111111;
assign LUT_4[30595] = 32'b00000000000000001000110010110111;
assign LUT_4[30596] = 32'b00000000000000001101001100110111;
assign LUT_4[30597] = 32'b00000000000000000110011000101111;
assign LUT_4[30598] = 32'b00000000000000001100100111011011;
assign LUT_4[30599] = 32'b00000000000000000101110011010011;
assign LUT_4[30600] = 32'b00000000000000001001011000110000;
assign LUT_4[30601] = 32'b00000000000000000010100100101000;
assign LUT_4[30602] = 32'b00000000000000001000110011010100;
assign LUT_4[30603] = 32'b00000000000000000001111111001100;
assign LUT_4[30604] = 32'b00000000000000000110011001001100;
assign LUT_4[30605] = 32'b11111111111111111111100101000100;
assign LUT_4[30606] = 32'b00000000000000000101110011110000;
assign LUT_4[30607] = 32'b11111111111111111110111111101000;
assign LUT_4[30608] = 32'b00000000000000001101111110001001;
assign LUT_4[30609] = 32'b00000000000000000111001010000001;
assign LUT_4[30610] = 32'b00000000000000001101011000101101;
assign LUT_4[30611] = 32'b00000000000000000110100100100101;
assign LUT_4[30612] = 32'b00000000000000001010111110100101;
assign LUT_4[30613] = 32'b00000000000000000100001010011101;
assign LUT_4[30614] = 32'b00000000000000001010011001001001;
assign LUT_4[30615] = 32'b00000000000000000011100101000001;
assign LUT_4[30616] = 32'b00000000000000000111001010011110;
assign LUT_4[30617] = 32'b00000000000000000000010110010110;
assign LUT_4[30618] = 32'b00000000000000000110100101000010;
assign LUT_4[30619] = 32'b11111111111111111111110000111010;
assign LUT_4[30620] = 32'b00000000000000000100001010111010;
assign LUT_4[30621] = 32'b11111111111111111101010110110010;
assign LUT_4[30622] = 32'b00000000000000000011100101011110;
assign LUT_4[30623] = 32'b11111111111111111100110001010110;
assign LUT_4[30624] = 32'b00000000000000001110100111100010;
assign LUT_4[30625] = 32'b00000000000000000111110011011010;
assign LUT_4[30626] = 32'b00000000000000001110000010000110;
assign LUT_4[30627] = 32'b00000000000000000111001101111110;
assign LUT_4[30628] = 32'b00000000000000001011100111111110;
assign LUT_4[30629] = 32'b00000000000000000100110011110110;
assign LUT_4[30630] = 32'b00000000000000001011000010100010;
assign LUT_4[30631] = 32'b00000000000000000100001110011010;
assign LUT_4[30632] = 32'b00000000000000000111110011110111;
assign LUT_4[30633] = 32'b00000000000000000000111111101111;
assign LUT_4[30634] = 32'b00000000000000000111001110011011;
assign LUT_4[30635] = 32'b00000000000000000000011010010011;
assign LUT_4[30636] = 32'b00000000000000000100110100010011;
assign LUT_4[30637] = 32'b11111111111111111110000000001011;
assign LUT_4[30638] = 32'b00000000000000000100001110110111;
assign LUT_4[30639] = 32'b11111111111111111101011010101111;
assign LUT_4[30640] = 32'b00000000000000001100011001010000;
assign LUT_4[30641] = 32'b00000000000000000101100101001000;
assign LUT_4[30642] = 32'b00000000000000001011110011110100;
assign LUT_4[30643] = 32'b00000000000000000100111111101100;
assign LUT_4[30644] = 32'b00000000000000001001011001101100;
assign LUT_4[30645] = 32'b00000000000000000010100101100100;
assign LUT_4[30646] = 32'b00000000000000001000110100010000;
assign LUT_4[30647] = 32'b00000000000000000010000000001000;
assign LUT_4[30648] = 32'b00000000000000000101100101100101;
assign LUT_4[30649] = 32'b11111111111111111110110001011101;
assign LUT_4[30650] = 32'b00000000000000000101000000001001;
assign LUT_4[30651] = 32'b11111111111111111110001100000001;
assign LUT_4[30652] = 32'b00000000000000000010100110000001;
assign LUT_4[30653] = 32'b11111111111111111011110001111001;
assign LUT_4[30654] = 32'b00000000000000000010000000100101;
assign LUT_4[30655] = 32'b11111111111111111011001100011101;
assign LUT_4[30656] = 32'b00000000000000010001100011101111;
assign LUT_4[30657] = 32'b00000000000000001010101111100111;
assign LUT_4[30658] = 32'b00000000000000010000111110010011;
assign LUT_4[30659] = 32'b00000000000000001010001010001011;
assign LUT_4[30660] = 32'b00000000000000001110100100001011;
assign LUT_4[30661] = 32'b00000000000000000111110000000011;
assign LUT_4[30662] = 32'b00000000000000001101111110101111;
assign LUT_4[30663] = 32'b00000000000000000111001010100111;
assign LUT_4[30664] = 32'b00000000000000001010110000000100;
assign LUT_4[30665] = 32'b00000000000000000011111011111100;
assign LUT_4[30666] = 32'b00000000000000001010001010101000;
assign LUT_4[30667] = 32'b00000000000000000011010110100000;
assign LUT_4[30668] = 32'b00000000000000000111110000100000;
assign LUT_4[30669] = 32'b00000000000000000000111100011000;
assign LUT_4[30670] = 32'b00000000000000000111001011000100;
assign LUT_4[30671] = 32'b00000000000000000000010110111100;
assign LUT_4[30672] = 32'b00000000000000001111010101011101;
assign LUT_4[30673] = 32'b00000000000000001000100001010101;
assign LUT_4[30674] = 32'b00000000000000001110110000000001;
assign LUT_4[30675] = 32'b00000000000000000111111011111001;
assign LUT_4[30676] = 32'b00000000000000001100010101111001;
assign LUT_4[30677] = 32'b00000000000000000101100001110001;
assign LUT_4[30678] = 32'b00000000000000001011110000011101;
assign LUT_4[30679] = 32'b00000000000000000100111100010101;
assign LUT_4[30680] = 32'b00000000000000001000100001110010;
assign LUT_4[30681] = 32'b00000000000000000001101101101010;
assign LUT_4[30682] = 32'b00000000000000000111111100010110;
assign LUT_4[30683] = 32'b00000000000000000001001000001110;
assign LUT_4[30684] = 32'b00000000000000000101100010001110;
assign LUT_4[30685] = 32'b11111111111111111110101110000110;
assign LUT_4[30686] = 32'b00000000000000000100111100110010;
assign LUT_4[30687] = 32'b11111111111111111110001000101010;
assign LUT_4[30688] = 32'b00000000000000001111111110110110;
assign LUT_4[30689] = 32'b00000000000000001001001010101110;
assign LUT_4[30690] = 32'b00000000000000001111011001011010;
assign LUT_4[30691] = 32'b00000000000000001000100101010010;
assign LUT_4[30692] = 32'b00000000000000001100111111010010;
assign LUT_4[30693] = 32'b00000000000000000110001011001010;
assign LUT_4[30694] = 32'b00000000000000001100011001110110;
assign LUT_4[30695] = 32'b00000000000000000101100101101110;
assign LUT_4[30696] = 32'b00000000000000001001001011001011;
assign LUT_4[30697] = 32'b00000000000000000010010111000011;
assign LUT_4[30698] = 32'b00000000000000001000100101101111;
assign LUT_4[30699] = 32'b00000000000000000001110001100111;
assign LUT_4[30700] = 32'b00000000000000000110001011100111;
assign LUT_4[30701] = 32'b11111111111111111111010111011111;
assign LUT_4[30702] = 32'b00000000000000000101100110001011;
assign LUT_4[30703] = 32'b11111111111111111110110010000011;
assign LUT_4[30704] = 32'b00000000000000001101110000100100;
assign LUT_4[30705] = 32'b00000000000000000110111100011100;
assign LUT_4[30706] = 32'b00000000000000001101001011001000;
assign LUT_4[30707] = 32'b00000000000000000110010111000000;
assign LUT_4[30708] = 32'b00000000000000001010110001000000;
assign LUT_4[30709] = 32'b00000000000000000011111100111000;
assign LUT_4[30710] = 32'b00000000000000001010001011100100;
assign LUT_4[30711] = 32'b00000000000000000011010111011100;
assign LUT_4[30712] = 32'b00000000000000000110111100111001;
assign LUT_4[30713] = 32'b00000000000000000000001000110001;
assign LUT_4[30714] = 32'b00000000000000000110010111011101;
assign LUT_4[30715] = 32'b11111111111111111111100011010101;
assign LUT_4[30716] = 32'b00000000000000000011111101010101;
assign LUT_4[30717] = 32'b11111111111111111101001001001101;
assign LUT_4[30718] = 32'b00000000000000000011010111111001;
assign LUT_4[30719] = 32'b11111111111111111100100011110001;
assign LUT_4[30720] = 32'b00000000000000000011011011010011;
assign LUT_4[30721] = 32'b11111111111111111100100111001011;
assign LUT_4[30722] = 32'b00000000000000000010110101110111;
assign LUT_4[30723] = 32'b11111111111111111100000001101111;
assign LUT_4[30724] = 32'b00000000000000000000011011101111;
assign LUT_4[30725] = 32'b11111111111111111001100111100111;
assign LUT_4[30726] = 32'b11111111111111111111110110010011;
assign LUT_4[30727] = 32'b11111111111111111001000010001011;
assign LUT_4[30728] = 32'b11111111111111111100100111101000;
assign LUT_4[30729] = 32'b11111111111111110101110011100000;
assign LUT_4[30730] = 32'b11111111111111111100000010001100;
assign LUT_4[30731] = 32'b11111111111111110101001110000100;
assign LUT_4[30732] = 32'b11111111111111111001101000000100;
assign LUT_4[30733] = 32'b11111111111111110010110011111100;
assign LUT_4[30734] = 32'b11111111111111111001000010101000;
assign LUT_4[30735] = 32'b11111111111111110010001110100000;
assign LUT_4[30736] = 32'b00000000000000000001001101000001;
assign LUT_4[30737] = 32'b11111111111111111010011000111001;
assign LUT_4[30738] = 32'b00000000000000000000100111100101;
assign LUT_4[30739] = 32'b11111111111111111001110011011101;
assign LUT_4[30740] = 32'b11111111111111111110001101011101;
assign LUT_4[30741] = 32'b11111111111111110111011001010101;
assign LUT_4[30742] = 32'b11111111111111111101101000000001;
assign LUT_4[30743] = 32'b11111111111111110110110011111001;
assign LUT_4[30744] = 32'b11111111111111111010011001010110;
assign LUT_4[30745] = 32'b11111111111111110011100101001110;
assign LUT_4[30746] = 32'b11111111111111111001110011111010;
assign LUT_4[30747] = 32'b11111111111111110010111111110010;
assign LUT_4[30748] = 32'b11111111111111110111011001110010;
assign LUT_4[30749] = 32'b11111111111111110000100101101010;
assign LUT_4[30750] = 32'b11111111111111110110110100010110;
assign LUT_4[30751] = 32'b11111111111111110000000000001110;
assign LUT_4[30752] = 32'b00000000000000000001110110011010;
assign LUT_4[30753] = 32'b11111111111111111011000010010010;
assign LUT_4[30754] = 32'b00000000000000000001010000111110;
assign LUT_4[30755] = 32'b11111111111111111010011100110110;
assign LUT_4[30756] = 32'b11111111111111111110110110110110;
assign LUT_4[30757] = 32'b11111111111111111000000010101110;
assign LUT_4[30758] = 32'b11111111111111111110010001011010;
assign LUT_4[30759] = 32'b11111111111111110111011101010010;
assign LUT_4[30760] = 32'b11111111111111111011000010101111;
assign LUT_4[30761] = 32'b11111111111111110100001110100111;
assign LUT_4[30762] = 32'b11111111111111111010011101010011;
assign LUT_4[30763] = 32'b11111111111111110011101001001011;
assign LUT_4[30764] = 32'b11111111111111111000000011001011;
assign LUT_4[30765] = 32'b11111111111111110001001111000011;
assign LUT_4[30766] = 32'b11111111111111110111011101101111;
assign LUT_4[30767] = 32'b11111111111111110000101001100111;
assign LUT_4[30768] = 32'b11111111111111111111101000001000;
assign LUT_4[30769] = 32'b11111111111111111000110100000000;
assign LUT_4[30770] = 32'b11111111111111111111000010101100;
assign LUT_4[30771] = 32'b11111111111111111000001110100100;
assign LUT_4[30772] = 32'b11111111111111111100101000100100;
assign LUT_4[30773] = 32'b11111111111111110101110100011100;
assign LUT_4[30774] = 32'b11111111111111111100000011001000;
assign LUT_4[30775] = 32'b11111111111111110101001111000000;
assign LUT_4[30776] = 32'b11111111111111111000110100011101;
assign LUT_4[30777] = 32'b11111111111111110010000000010101;
assign LUT_4[30778] = 32'b11111111111111111000001111000001;
assign LUT_4[30779] = 32'b11111111111111110001011010111001;
assign LUT_4[30780] = 32'b11111111111111110101110100111001;
assign LUT_4[30781] = 32'b11111111111111101111000000110001;
assign LUT_4[30782] = 32'b11111111111111110101001111011101;
assign LUT_4[30783] = 32'b11111111111111101110011011010101;
assign LUT_4[30784] = 32'b00000000000000000100110010100111;
assign LUT_4[30785] = 32'b11111111111111111101111110011111;
assign LUT_4[30786] = 32'b00000000000000000100001101001011;
assign LUT_4[30787] = 32'b11111111111111111101011001000011;
assign LUT_4[30788] = 32'b00000000000000000001110011000011;
assign LUT_4[30789] = 32'b11111111111111111010111110111011;
assign LUT_4[30790] = 32'b00000000000000000001001101100111;
assign LUT_4[30791] = 32'b11111111111111111010011001011111;
assign LUT_4[30792] = 32'b11111111111111111101111110111100;
assign LUT_4[30793] = 32'b11111111111111110111001010110100;
assign LUT_4[30794] = 32'b11111111111111111101011001100000;
assign LUT_4[30795] = 32'b11111111111111110110100101011000;
assign LUT_4[30796] = 32'b11111111111111111010111111011000;
assign LUT_4[30797] = 32'b11111111111111110100001011010000;
assign LUT_4[30798] = 32'b11111111111111111010011001111100;
assign LUT_4[30799] = 32'b11111111111111110011100101110100;
assign LUT_4[30800] = 32'b00000000000000000010100100010101;
assign LUT_4[30801] = 32'b11111111111111111011110000001101;
assign LUT_4[30802] = 32'b00000000000000000001111110111001;
assign LUT_4[30803] = 32'b11111111111111111011001010110001;
assign LUT_4[30804] = 32'b11111111111111111111100100110001;
assign LUT_4[30805] = 32'b11111111111111111000110000101001;
assign LUT_4[30806] = 32'b11111111111111111110111111010101;
assign LUT_4[30807] = 32'b11111111111111111000001011001101;
assign LUT_4[30808] = 32'b11111111111111111011110000101010;
assign LUT_4[30809] = 32'b11111111111111110100111100100010;
assign LUT_4[30810] = 32'b11111111111111111011001011001110;
assign LUT_4[30811] = 32'b11111111111111110100010111000110;
assign LUT_4[30812] = 32'b11111111111111111000110001000110;
assign LUT_4[30813] = 32'b11111111111111110001111100111110;
assign LUT_4[30814] = 32'b11111111111111111000001011101010;
assign LUT_4[30815] = 32'b11111111111111110001010111100010;
assign LUT_4[30816] = 32'b00000000000000000011001101101110;
assign LUT_4[30817] = 32'b11111111111111111100011001100110;
assign LUT_4[30818] = 32'b00000000000000000010101000010010;
assign LUT_4[30819] = 32'b11111111111111111011110100001010;
assign LUT_4[30820] = 32'b00000000000000000000001110001010;
assign LUT_4[30821] = 32'b11111111111111111001011010000010;
assign LUT_4[30822] = 32'b11111111111111111111101000101110;
assign LUT_4[30823] = 32'b11111111111111111000110100100110;
assign LUT_4[30824] = 32'b11111111111111111100011010000011;
assign LUT_4[30825] = 32'b11111111111111110101100101111011;
assign LUT_4[30826] = 32'b11111111111111111011110100100111;
assign LUT_4[30827] = 32'b11111111111111110101000000011111;
assign LUT_4[30828] = 32'b11111111111111111001011010011111;
assign LUT_4[30829] = 32'b11111111111111110010100110010111;
assign LUT_4[30830] = 32'b11111111111111111000110101000011;
assign LUT_4[30831] = 32'b11111111111111110010000000111011;
assign LUT_4[30832] = 32'b00000000000000000000111111011100;
assign LUT_4[30833] = 32'b11111111111111111010001011010100;
assign LUT_4[30834] = 32'b00000000000000000000011010000000;
assign LUT_4[30835] = 32'b11111111111111111001100101111000;
assign LUT_4[30836] = 32'b11111111111111111101111111111000;
assign LUT_4[30837] = 32'b11111111111111110111001011110000;
assign LUT_4[30838] = 32'b11111111111111111101011010011100;
assign LUT_4[30839] = 32'b11111111111111110110100110010100;
assign LUT_4[30840] = 32'b11111111111111111010001011110001;
assign LUT_4[30841] = 32'b11111111111111110011010111101001;
assign LUT_4[30842] = 32'b11111111111111111001100110010101;
assign LUT_4[30843] = 32'b11111111111111110010110010001101;
assign LUT_4[30844] = 32'b11111111111111110111001100001101;
assign LUT_4[30845] = 32'b11111111111111110000011000000101;
assign LUT_4[30846] = 32'b11111111111111110110100110110001;
assign LUT_4[30847] = 32'b11111111111111101111110010101001;
assign LUT_4[30848] = 32'b00000000000000000110000001011011;
assign LUT_4[30849] = 32'b11111111111111111111001101010011;
assign LUT_4[30850] = 32'b00000000000000000101011011111111;
assign LUT_4[30851] = 32'b11111111111111111110100111110111;
assign LUT_4[30852] = 32'b00000000000000000011000001110111;
assign LUT_4[30853] = 32'b11111111111111111100001101101111;
assign LUT_4[30854] = 32'b00000000000000000010011100011011;
assign LUT_4[30855] = 32'b11111111111111111011101000010011;
assign LUT_4[30856] = 32'b11111111111111111111001101110000;
assign LUT_4[30857] = 32'b11111111111111111000011001101000;
assign LUT_4[30858] = 32'b11111111111111111110101000010100;
assign LUT_4[30859] = 32'b11111111111111110111110100001100;
assign LUT_4[30860] = 32'b11111111111111111100001110001100;
assign LUT_4[30861] = 32'b11111111111111110101011010000100;
assign LUT_4[30862] = 32'b11111111111111111011101000110000;
assign LUT_4[30863] = 32'b11111111111111110100110100101000;
assign LUT_4[30864] = 32'b00000000000000000011110011001001;
assign LUT_4[30865] = 32'b11111111111111111100111111000001;
assign LUT_4[30866] = 32'b00000000000000000011001101101101;
assign LUT_4[30867] = 32'b11111111111111111100011001100101;
assign LUT_4[30868] = 32'b00000000000000000000110011100101;
assign LUT_4[30869] = 32'b11111111111111111001111111011101;
assign LUT_4[30870] = 32'b00000000000000000000001110001001;
assign LUT_4[30871] = 32'b11111111111111111001011010000001;
assign LUT_4[30872] = 32'b11111111111111111100111111011110;
assign LUT_4[30873] = 32'b11111111111111110110001011010110;
assign LUT_4[30874] = 32'b11111111111111111100011010000010;
assign LUT_4[30875] = 32'b11111111111111110101100101111010;
assign LUT_4[30876] = 32'b11111111111111111001111111111010;
assign LUT_4[30877] = 32'b11111111111111110011001011110010;
assign LUT_4[30878] = 32'b11111111111111111001011010011110;
assign LUT_4[30879] = 32'b11111111111111110010100110010110;
assign LUT_4[30880] = 32'b00000000000000000100011100100010;
assign LUT_4[30881] = 32'b11111111111111111101101000011010;
assign LUT_4[30882] = 32'b00000000000000000011110111000110;
assign LUT_4[30883] = 32'b11111111111111111101000010111110;
assign LUT_4[30884] = 32'b00000000000000000001011100111110;
assign LUT_4[30885] = 32'b11111111111111111010101000110110;
assign LUT_4[30886] = 32'b00000000000000000000110111100010;
assign LUT_4[30887] = 32'b11111111111111111010000011011010;
assign LUT_4[30888] = 32'b11111111111111111101101000110111;
assign LUT_4[30889] = 32'b11111111111111110110110100101111;
assign LUT_4[30890] = 32'b11111111111111111101000011011011;
assign LUT_4[30891] = 32'b11111111111111110110001111010011;
assign LUT_4[30892] = 32'b11111111111111111010101001010011;
assign LUT_4[30893] = 32'b11111111111111110011110101001011;
assign LUT_4[30894] = 32'b11111111111111111010000011110111;
assign LUT_4[30895] = 32'b11111111111111110011001111101111;
assign LUT_4[30896] = 32'b00000000000000000010001110010000;
assign LUT_4[30897] = 32'b11111111111111111011011010001000;
assign LUT_4[30898] = 32'b00000000000000000001101000110100;
assign LUT_4[30899] = 32'b11111111111111111010110100101100;
assign LUT_4[30900] = 32'b11111111111111111111001110101100;
assign LUT_4[30901] = 32'b11111111111111111000011010100100;
assign LUT_4[30902] = 32'b11111111111111111110101001010000;
assign LUT_4[30903] = 32'b11111111111111110111110101001000;
assign LUT_4[30904] = 32'b11111111111111111011011010100101;
assign LUT_4[30905] = 32'b11111111111111110100100110011101;
assign LUT_4[30906] = 32'b11111111111111111010110101001001;
assign LUT_4[30907] = 32'b11111111111111110100000001000001;
assign LUT_4[30908] = 32'b11111111111111111000011011000001;
assign LUT_4[30909] = 32'b11111111111111110001100110111001;
assign LUT_4[30910] = 32'b11111111111111110111110101100101;
assign LUT_4[30911] = 32'b11111111111111110001000001011101;
assign LUT_4[30912] = 32'b00000000000000000111011000101111;
assign LUT_4[30913] = 32'b00000000000000000000100100100111;
assign LUT_4[30914] = 32'b00000000000000000110110011010011;
assign LUT_4[30915] = 32'b11111111111111111111111111001011;
assign LUT_4[30916] = 32'b00000000000000000100011001001011;
assign LUT_4[30917] = 32'b11111111111111111101100101000011;
assign LUT_4[30918] = 32'b00000000000000000011110011101111;
assign LUT_4[30919] = 32'b11111111111111111100111111100111;
assign LUT_4[30920] = 32'b00000000000000000000100101000100;
assign LUT_4[30921] = 32'b11111111111111111001110000111100;
assign LUT_4[30922] = 32'b11111111111111111111111111101000;
assign LUT_4[30923] = 32'b11111111111111111001001011100000;
assign LUT_4[30924] = 32'b11111111111111111101100101100000;
assign LUT_4[30925] = 32'b11111111111111110110110001011000;
assign LUT_4[30926] = 32'b11111111111111111101000000000100;
assign LUT_4[30927] = 32'b11111111111111110110001011111100;
assign LUT_4[30928] = 32'b00000000000000000101001010011101;
assign LUT_4[30929] = 32'b11111111111111111110010110010101;
assign LUT_4[30930] = 32'b00000000000000000100100101000001;
assign LUT_4[30931] = 32'b11111111111111111101110000111001;
assign LUT_4[30932] = 32'b00000000000000000010001010111001;
assign LUT_4[30933] = 32'b11111111111111111011010110110001;
assign LUT_4[30934] = 32'b00000000000000000001100101011101;
assign LUT_4[30935] = 32'b11111111111111111010110001010101;
assign LUT_4[30936] = 32'b11111111111111111110010110110010;
assign LUT_4[30937] = 32'b11111111111111110111100010101010;
assign LUT_4[30938] = 32'b11111111111111111101110001010110;
assign LUT_4[30939] = 32'b11111111111111110110111101001110;
assign LUT_4[30940] = 32'b11111111111111111011010111001110;
assign LUT_4[30941] = 32'b11111111111111110100100011000110;
assign LUT_4[30942] = 32'b11111111111111111010110001110010;
assign LUT_4[30943] = 32'b11111111111111110011111101101010;
assign LUT_4[30944] = 32'b00000000000000000101110011110110;
assign LUT_4[30945] = 32'b11111111111111111110111111101110;
assign LUT_4[30946] = 32'b00000000000000000101001110011010;
assign LUT_4[30947] = 32'b11111111111111111110011010010010;
assign LUT_4[30948] = 32'b00000000000000000010110100010010;
assign LUT_4[30949] = 32'b11111111111111111100000000001010;
assign LUT_4[30950] = 32'b00000000000000000010001110110110;
assign LUT_4[30951] = 32'b11111111111111111011011010101110;
assign LUT_4[30952] = 32'b11111111111111111111000000001011;
assign LUT_4[30953] = 32'b11111111111111111000001100000011;
assign LUT_4[30954] = 32'b11111111111111111110011010101111;
assign LUT_4[30955] = 32'b11111111111111110111100110100111;
assign LUT_4[30956] = 32'b11111111111111111100000000100111;
assign LUT_4[30957] = 32'b11111111111111110101001100011111;
assign LUT_4[30958] = 32'b11111111111111111011011011001011;
assign LUT_4[30959] = 32'b11111111111111110100100111000011;
assign LUT_4[30960] = 32'b00000000000000000011100101100100;
assign LUT_4[30961] = 32'b11111111111111111100110001011100;
assign LUT_4[30962] = 32'b00000000000000000011000000001000;
assign LUT_4[30963] = 32'b11111111111111111100001100000000;
assign LUT_4[30964] = 32'b00000000000000000000100110000000;
assign LUT_4[30965] = 32'b11111111111111111001110001111000;
assign LUT_4[30966] = 32'b00000000000000000000000000100100;
assign LUT_4[30967] = 32'b11111111111111111001001100011100;
assign LUT_4[30968] = 32'b11111111111111111100110001111001;
assign LUT_4[30969] = 32'b11111111111111110101111101110001;
assign LUT_4[30970] = 32'b11111111111111111100001100011101;
assign LUT_4[30971] = 32'b11111111111111110101011000010101;
assign LUT_4[30972] = 32'b11111111111111111001110010010101;
assign LUT_4[30973] = 32'b11111111111111110010111110001101;
assign LUT_4[30974] = 32'b11111111111111111001001100111001;
assign LUT_4[30975] = 32'b11111111111111110010011000110001;
assign LUT_4[30976] = 32'b00000000000000001000010110110110;
assign LUT_4[30977] = 32'b00000000000000000001100010101110;
assign LUT_4[30978] = 32'b00000000000000000111110001011010;
assign LUT_4[30979] = 32'b00000000000000000000111101010010;
assign LUT_4[30980] = 32'b00000000000000000101010111010010;
assign LUT_4[30981] = 32'b11111111111111111110100011001010;
assign LUT_4[30982] = 32'b00000000000000000100110001110110;
assign LUT_4[30983] = 32'b11111111111111111101111101101110;
assign LUT_4[30984] = 32'b00000000000000000001100011001011;
assign LUT_4[30985] = 32'b11111111111111111010101111000011;
assign LUT_4[30986] = 32'b00000000000000000000111101101111;
assign LUT_4[30987] = 32'b11111111111111111010001001100111;
assign LUT_4[30988] = 32'b11111111111111111110100011100111;
assign LUT_4[30989] = 32'b11111111111111110111101111011111;
assign LUT_4[30990] = 32'b11111111111111111101111110001011;
assign LUT_4[30991] = 32'b11111111111111110111001010000011;
assign LUT_4[30992] = 32'b00000000000000000110001000100100;
assign LUT_4[30993] = 32'b11111111111111111111010100011100;
assign LUT_4[30994] = 32'b00000000000000000101100011001000;
assign LUT_4[30995] = 32'b11111111111111111110101111000000;
assign LUT_4[30996] = 32'b00000000000000000011001001000000;
assign LUT_4[30997] = 32'b11111111111111111100010100111000;
assign LUT_4[30998] = 32'b00000000000000000010100011100100;
assign LUT_4[30999] = 32'b11111111111111111011101111011100;
assign LUT_4[31000] = 32'b11111111111111111111010100111001;
assign LUT_4[31001] = 32'b11111111111111111000100000110001;
assign LUT_4[31002] = 32'b11111111111111111110101111011101;
assign LUT_4[31003] = 32'b11111111111111110111111011010101;
assign LUT_4[31004] = 32'b11111111111111111100010101010101;
assign LUT_4[31005] = 32'b11111111111111110101100001001101;
assign LUT_4[31006] = 32'b11111111111111111011101111111001;
assign LUT_4[31007] = 32'b11111111111111110100111011110001;
assign LUT_4[31008] = 32'b00000000000000000110110001111101;
assign LUT_4[31009] = 32'b11111111111111111111111101110101;
assign LUT_4[31010] = 32'b00000000000000000110001100100001;
assign LUT_4[31011] = 32'b11111111111111111111011000011001;
assign LUT_4[31012] = 32'b00000000000000000011110010011001;
assign LUT_4[31013] = 32'b11111111111111111100111110010001;
assign LUT_4[31014] = 32'b00000000000000000011001100111101;
assign LUT_4[31015] = 32'b11111111111111111100011000110101;
assign LUT_4[31016] = 32'b11111111111111111111111110010010;
assign LUT_4[31017] = 32'b11111111111111111001001010001010;
assign LUT_4[31018] = 32'b11111111111111111111011000110110;
assign LUT_4[31019] = 32'b11111111111111111000100100101110;
assign LUT_4[31020] = 32'b11111111111111111100111110101110;
assign LUT_4[31021] = 32'b11111111111111110110001010100110;
assign LUT_4[31022] = 32'b11111111111111111100011001010010;
assign LUT_4[31023] = 32'b11111111111111110101100101001010;
assign LUT_4[31024] = 32'b00000000000000000100100011101011;
assign LUT_4[31025] = 32'b11111111111111111101101111100011;
assign LUT_4[31026] = 32'b00000000000000000011111110001111;
assign LUT_4[31027] = 32'b11111111111111111101001010000111;
assign LUT_4[31028] = 32'b00000000000000000001100100000111;
assign LUT_4[31029] = 32'b11111111111111111010101111111111;
assign LUT_4[31030] = 32'b00000000000000000000111110101011;
assign LUT_4[31031] = 32'b11111111111111111010001010100011;
assign LUT_4[31032] = 32'b11111111111111111101110000000000;
assign LUT_4[31033] = 32'b11111111111111110110111011111000;
assign LUT_4[31034] = 32'b11111111111111111101001010100100;
assign LUT_4[31035] = 32'b11111111111111110110010110011100;
assign LUT_4[31036] = 32'b11111111111111111010110000011100;
assign LUT_4[31037] = 32'b11111111111111110011111100010100;
assign LUT_4[31038] = 32'b11111111111111111010001011000000;
assign LUT_4[31039] = 32'b11111111111111110011010110111000;
assign LUT_4[31040] = 32'b00000000000000001001101110001010;
assign LUT_4[31041] = 32'b00000000000000000010111010000010;
assign LUT_4[31042] = 32'b00000000000000001001001000101110;
assign LUT_4[31043] = 32'b00000000000000000010010100100110;
assign LUT_4[31044] = 32'b00000000000000000110101110100110;
assign LUT_4[31045] = 32'b11111111111111111111111010011110;
assign LUT_4[31046] = 32'b00000000000000000110001001001010;
assign LUT_4[31047] = 32'b11111111111111111111010101000010;
assign LUT_4[31048] = 32'b00000000000000000010111010011111;
assign LUT_4[31049] = 32'b11111111111111111100000110010111;
assign LUT_4[31050] = 32'b00000000000000000010010101000011;
assign LUT_4[31051] = 32'b11111111111111111011100000111011;
assign LUT_4[31052] = 32'b11111111111111111111111010111011;
assign LUT_4[31053] = 32'b11111111111111111001000110110011;
assign LUT_4[31054] = 32'b11111111111111111111010101011111;
assign LUT_4[31055] = 32'b11111111111111111000100001010111;
assign LUT_4[31056] = 32'b00000000000000000111011111111000;
assign LUT_4[31057] = 32'b00000000000000000000101011110000;
assign LUT_4[31058] = 32'b00000000000000000110111010011100;
assign LUT_4[31059] = 32'b00000000000000000000000110010100;
assign LUT_4[31060] = 32'b00000000000000000100100000010100;
assign LUT_4[31061] = 32'b11111111111111111101101100001100;
assign LUT_4[31062] = 32'b00000000000000000011111010111000;
assign LUT_4[31063] = 32'b11111111111111111101000110110000;
assign LUT_4[31064] = 32'b00000000000000000000101100001101;
assign LUT_4[31065] = 32'b11111111111111111001111000000101;
assign LUT_4[31066] = 32'b00000000000000000000000110110001;
assign LUT_4[31067] = 32'b11111111111111111001010010101001;
assign LUT_4[31068] = 32'b11111111111111111101101100101001;
assign LUT_4[31069] = 32'b11111111111111110110111000100001;
assign LUT_4[31070] = 32'b11111111111111111101000111001101;
assign LUT_4[31071] = 32'b11111111111111110110010011000101;
assign LUT_4[31072] = 32'b00000000000000001000001001010001;
assign LUT_4[31073] = 32'b00000000000000000001010101001001;
assign LUT_4[31074] = 32'b00000000000000000111100011110101;
assign LUT_4[31075] = 32'b00000000000000000000101111101101;
assign LUT_4[31076] = 32'b00000000000000000101001001101101;
assign LUT_4[31077] = 32'b11111111111111111110010101100101;
assign LUT_4[31078] = 32'b00000000000000000100100100010001;
assign LUT_4[31079] = 32'b11111111111111111101110000001001;
assign LUT_4[31080] = 32'b00000000000000000001010101100110;
assign LUT_4[31081] = 32'b11111111111111111010100001011110;
assign LUT_4[31082] = 32'b00000000000000000000110000001010;
assign LUT_4[31083] = 32'b11111111111111111001111100000010;
assign LUT_4[31084] = 32'b11111111111111111110010110000010;
assign LUT_4[31085] = 32'b11111111111111110111100001111010;
assign LUT_4[31086] = 32'b11111111111111111101110000100110;
assign LUT_4[31087] = 32'b11111111111111110110111100011110;
assign LUT_4[31088] = 32'b00000000000000000101111010111111;
assign LUT_4[31089] = 32'b11111111111111111111000110110111;
assign LUT_4[31090] = 32'b00000000000000000101010101100011;
assign LUT_4[31091] = 32'b11111111111111111110100001011011;
assign LUT_4[31092] = 32'b00000000000000000010111011011011;
assign LUT_4[31093] = 32'b11111111111111111100000111010011;
assign LUT_4[31094] = 32'b00000000000000000010010101111111;
assign LUT_4[31095] = 32'b11111111111111111011100001110111;
assign LUT_4[31096] = 32'b11111111111111111111000111010100;
assign LUT_4[31097] = 32'b11111111111111111000010011001100;
assign LUT_4[31098] = 32'b11111111111111111110100001111000;
assign LUT_4[31099] = 32'b11111111111111110111101101110000;
assign LUT_4[31100] = 32'b11111111111111111100000111110000;
assign LUT_4[31101] = 32'b11111111111111110101010011101000;
assign LUT_4[31102] = 32'b11111111111111111011100010010100;
assign LUT_4[31103] = 32'b11111111111111110100101110001100;
assign LUT_4[31104] = 32'b00000000000000001010111100111110;
assign LUT_4[31105] = 32'b00000000000000000100001000110110;
assign LUT_4[31106] = 32'b00000000000000001010010111100010;
assign LUT_4[31107] = 32'b00000000000000000011100011011010;
assign LUT_4[31108] = 32'b00000000000000000111111101011010;
assign LUT_4[31109] = 32'b00000000000000000001001001010010;
assign LUT_4[31110] = 32'b00000000000000000111010111111110;
assign LUT_4[31111] = 32'b00000000000000000000100011110110;
assign LUT_4[31112] = 32'b00000000000000000100001001010011;
assign LUT_4[31113] = 32'b11111111111111111101010101001011;
assign LUT_4[31114] = 32'b00000000000000000011100011110111;
assign LUT_4[31115] = 32'b11111111111111111100101111101111;
assign LUT_4[31116] = 32'b00000000000000000001001001101111;
assign LUT_4[31117] = 32'b11111111111111111010010101100111;
assign LUT_4[31118] = 32'b00000000000000000000100100010011;
assign LUT_4[31119] = 32'b11111111111111111001110000001011;
assign LUT_4[31120] = 32'b00000000000000001000101110101100;
assign LUT_4[31121] = 32'b00000000000000000001111010100100;
assign LUT_4[31122] = 32'b00000000000000001000001001010000;
assign LUT_4[31123] = 32'b00000000000000000001010101001000;
assign LUT_4[31124] = 32'b00000000000000000101101111001000;
assign LUT_4[31125] = 32'b11111111111111111110111011000000;
assign LUT_4[31126] = 32'b00000000000000000101001001101100;
assign LUT_4[31127] = 32'b11111111111111111110010101100100;
assign LUT_4[31128] = 32'b00000000000000000001111011000001;
assign LUT_4[31129] = 32'b11111111111111111011000110111001;
assign LUT_4[31130] = 32'b00000000000000000001010101100101;
assign LUT_4[31131] = 32'b11111111111111111010100001011101;
assign LUT_4[31132] = 32'b11111111111111111110111011011101;
assign LUT_4[31133] = 32'b11111111111111111000000111010101;
assign LUT_4[31134] = 32'b11111111111111111110010110000001;
assign LUT_4[31135] = 32'b11111111111111110111100001111001;
assign LUT_4[31136] = 32'b00000000000000001001011000000101;
assign LUT_4[31137] = 32'b00000000000000000010100011111101;
assign LUT_4[31138] = 32'b00000000000000001000110010101001;
assign LUT_4[31139] = 32'b00000000000000000001111110100001;
assign LUT_4[31140] = 32'b00000000000000000110011000100001;
assign LUT_4[31141] = 32'b11111111111111111111100100011001;
assign LUT_4[31142] = 32'b00000000000000000101110011000101;
assign LUT_4[31143] = 32'b11111111111111111110111110111101;
assign LUT_4[31144] = 32'b00000000000000000010100100011010;
assign LUT_4[31145] = 32'b11111111111111111011110000010010;
assign LUT_4[31146] = 32'b00000000000000000001111110111110;
assign LUT_4[31147] = 32'b11111111111111111011001010110110;
assign LUT_4[31148] = 32'b11111111111111111111100100110110;
assign LUT_4[31149] = 32'b11111111111111111000110000101110;
assign LUT_4[31150] = 32'b11111111111111111110111111011010;
assign LUT_4[31151] = 32'b11111111111111111000001011010010;
assign LUT_4[31152] = 32'b00000000000000000111001001110011;
assign LUT_4[31153] = 32'b00000000000000000000010101101011;
assign LUT_4[31154] = 32'b00000000000000000110100100010111;
assign LUT_4[31155] = 32'b11111111111111111111110000001111;
assign LUT_4[31156] = 32'b00000000000000000100001010001111;
assign LUT_4[31157] = 32'b11111111111111111101010110000111;
assign LUT_4[31158] = 32'b00000000000000000011100100110011;
assign LUT_4[31159] = 32'b11111111111111111100110000101011;
assign LUT_4[31160] = 32'b00000000000000000000010110001000;
assign LUT_4[31161] = 32'b11111111111111111001100010000000;
assign LUT_4[31162] = 32'b11111111111111111111110000101100;
assign LUT_4[31163] = 32'b11111111111111111000111100100100;
assign LUT_4[31164] = 32'b11111111111111111101010110100100;
assign LUT_4[31165] = 32'b11111111111111110110100010011100;
assign LUT_4[31166] = 32'b11111111111111111100110001001000;
assign LUT_4[31167] = 32'b11111111111111110101111101000000;
assign LUT_4[31168] = 32'b00000000000000001100010100010010;
assign LUT_4[31169] = 32'b00000000000000000101100000001010;
assign LUT_4[31170] = 32'b00000000000000001011101110110110;
assign LUT_4[31171] = 32'b00000000000000000100111010101110;
assign LUT_4[31172] = 32'b00000000000000001001010100101110;
assign LUT_4[31173] = 32'b00000000000000000010100000100110;
assign LUT_4[31174] = 32'b00000000000000001000101111010010;
assign LUT_4[31175] = 32'b00000000000000000001111011001010;
assign LUT_4[31176] = 32'b00000000000000000101100000100111;
assign LUT_4[31177] = 32'b11111111111111111110101100011111;
assign LUT_4[31178] = 32'b00000000000000000100111011001011;
assign LUT_4[31179] = 32'b11111111111111111110000111000011;
assign LUT_4[31180] = 32'b00000000000000000010100001000011;
assign LUT_4[31181] = 32'b11111111111111111011101100111011;
assign LUT_4[31182] = 32'b00000000000000000001111011100111;
assign LUT_4[31183] = 32'b11111111111111111011000111011111;
assign LUT_4[31184] = 32'b00000000000000001010000110000000;
assign LUT_4[31185] = 32'b00000000000000000011010001111000;
assign LUT_4[31186] = 32'b00000000000000001001100000100100;
assign LUT_4[31187] = 32'b00000000000000000010101100011100;
assign LUT_4[31188] = 32'b00000000000000000111000110011100;
assign LUT_4[31189] = 32'b00000000000000000000010010010100;
assign LUT_4[31190] = 32'b00000000000000000110100001000000;
assign LUT_4[31191] = 32'b11111111111111111111101100111000;
assign LUT_4[31192] = 32'b00000000000000000011010010010101;
assign LUT_4[31193] = 32'b11111111111111111100011110001101;
assign LUT_4[31194] = 32'b00000000000000000010101100111001;
assign LUT_4[31195] = 32'b11111111111111111011111000110001;
assign LUT_4[31196] = 32'b00000000000000000000010010110001;
assign LUT_4[31197] = 32'b11111111111111111001011110101001;
assign LUT_4[31198] = 32'b11111111111111111111101101010101;
assign LUT_4[31199] = 32'b11111111111111111000111001001101;
assign LUT_4[31200] = 32'b00000000000000001010101111011001;
assign LUT_4[31201] = 32'b00000000000000000011111011010001;
assign LUT_4[31202] = 32'b00000000000000001010001001111101;
assign LUT_4[31203] = 32'b00000000000000000011010101110101;
assign LUT_4[31204] = 32'b00000000000000000111101111110101;
assign LUT_4[31205] = 32'b00000000000000000000111011101101;
assign LUT_4[31206] = 32'b00000000000000000111001010011001;
assign LUT_4[31207] = 32'b00000000000000000000010110010001;
assign LUT_4[31208] = 32'b00000000000000000011111011101110;
assign LUT_4[31209] = 32'b11111111111111111101000111100110;
assign LUT_4[31210] = 32'b00000000000000000011010110010010;
assign LUT_4[31211] = 32'b11111111111111111100100010001010;
assign LUT_4[31212] = 32'b00000000000000000000111100001010;
assign LUT_4[31213] = 32'b11111111111111111010001000000010;
assign LUT_4[31214] = 32'b00000000000000000000010110101110;
assign LUT_4[31215] = 32'b11111111111111111001100010100110;
assign LUT_4[31216] = 32'b00000000000000001000100001000111;
assign LUT_4[31217] = 32'b00000000000000000001101100111111;
assign LUT_4[31218] = 32'b00000000000000000111111011101011;
assign LUT_4[31219] = 32'b00000000000000000001000111100011;
assign LUT_4[31220] = 32'b00000000000000000101100001100011;
assign LUT_4[31221] = 32'b11111111111111111110101101011011;
assign LUT_4[31222] = 32'b00000000000000000100111100000111;
assign LUT_4[31223] = 32'b11111111111111111110000111111111;
assign LUT_4[31224] = 32'b00000000000000000001101101011100;
assign LUT_4[31225] = 32'b11111111111111111010111001010100;
assign LUT_4[31226] = 32'b00000000000000000001001000000000;
assign LUT_4[31227] = 32'b11111111111111111010010011111000;
assign LUT_4[31228] = 32'b11111111111111111110101101111000;
assign LUT_4[31229] = 32'b11111111111111110111111001110000;
assign LUT_4[31230] = 32'b11111111111111111110001000011100;
assign LUT_4[31231] = 32'b11111111111111110111010100010100;
assign LUT_4[31232] = 32'b00000000000000000010011111011011;
assign LUT_4[31233] = 32'b11111111111111111011101011010011;
assign LUT_4[31234] = 32'b00000000000000000001111001111111;
assign LUT_4[31235] = 32'b11111111111111111011000101110111;
assign LUT_4[31236] = 32'b11111111111111111111011111110111;
assign LUT_4[31237] = 32'b11111111111111111000101011101111;
assign LUT_4[31238] = 32'b11111111111111111110111010011011;
assign LUT_4[31239] = 32'b11111111111111111000000110010011;
assign LUT_4[31240] = 32'b11111111111111111011101011110000;
assign LUT_4[31241] = 32'b11111111111111110100110111101000;
assign LUT_4[31242] = 32'b11111111111111111011000110010100;
assign LUT_4[31243] = 32'b11111111111111110100010010001100;
assign LUT_4[31244] = 32'b11111111111111111000101100001100;
assign LUT_4[31245] = 32'b11111111111111110001111000000100;
assign LUT_4[31246] = 32'b11111111111111111000000110110000;
assign LUT_4[31247] = 32'b11111111111111110001010010101000;
assign LUT_4[31248] = 32'b00000000000000000000010001001001;
assign LUT_4[31249] = 32'b11111111111111111001011101000001;
assign LUT_4[31250] = 32'b11111111111111111111101011101101;
assign LUT_4[31251] = 32'b11111111111111111000110111100101;
assign LUT_4[31252] = 32'b11111111111111111101010001100101;
assign LUT_4[31253] = 32'b11111111111111110110011101011101;
assign LUT_4[31254] = 32'b11111111111111111100101100001001;
assign LUT_4[31255] = 32'b11111111111111110101111000000001;
assign LUT_4[31256] = 32'b11111111111111111001011101011110;
assign LUT_4[31257] = 32'b11111111111111110010101001010110;
assign LUT_4[31258] = 32'b11111111111111111000111000000010;
assign LUT_4[31259] = 32'b11111111111111110010000011111010;
assign LUT_4[31260] = 32'b11111111111111110110011101111010;
assign LUT_4[31261] = 32'b11111111111111101111101001110010;
assign LUT_4[31262] = 32'b11111111111111110101111000011110;
assign LUT_4[31263] = 32'b11111111111111101111000100010110;
assign LUT_4[31264] = 32'b00000000000000000000111010100010;
assign LUT_4[31265] = 32'b11111111111111111010000110011010;
assign LUT_4[31266] = 32'b00000000000000000000010101000110;
assign LUT_4[31267] = 32'b11111111111111111001100000111110;
assign LUT_4[31268] = 32'b11111111111111111101111010111110;
assign LUT_4[31269] = 32'b11111111111111110111000110110110;
assign LUT_4[31270] = 32'b11111111111111111101010101100010;
assign LUT_4[31271] = 32'b11111111111111110110100001011010;
assign LUT_4[31272] = 32'b11111111111111111010000110110111;
assign LUT_4[31273] = 32'b11111111111111110011010010101111;
assign LUT_4[31274] = 32'b11111111111111111001100001011011;
assign LUT_4[31275] = 32'b11111111111111110010101101010011;
assign LUT_4[31276] = 32'b11111111111111110111000111010011;
assign LUT_4[31277] = 32'b11111111111111110000010011001011;
assign LUT_4[31278] = 32'b11111111111111110110100001110111;
assign LUT_4[31279] = 32'b11111111111111101111101101101111;
assign LUT_4[31280] = 32'b11111111111111111110101100010000;
assign LUT_4[31281] = 32'b11111111111111110111111000001000;
assign LUT_4[31282] = 32'b11111111111111111110000110110100;
assign LUT_4[31283] = 32'b11111111111111110111010010101100;
assign LUT_4[31284] = 32'b11111111111111111011101100101100;
assign LUT_4[31285] = 32'b11111111111111110100111000100100;
assign LUT_4[31286] = 32'b11111111111111111011000111010000;
assign LUT_4[31287] = 32'b11111111111111110100010011001000;
assign LUT_4[31288] = 32'b11111111111111110111111000100101;
assign LUT_4[31289] = 32'b11111111111111110001000100011101;
assign LUT_4[31290] = 32'b11111111111111110111010011001001;
assign LUT_4[31291] = 32'b11111111111111110000011111000001;
assign LUT_4[31292] = 32'b11111111111111110100111001000001;
assign LUT_4[31293] = 32'b11111111111111101110000100111001;
assign LUT_4[31294] = 32'b11111111111111110100010011100101;
assign LUT_4[31295] = 32'b11111111111111101101011111011101;
assign LUT_4[31296] = 32'b00000000000000000011110110101111;
assign LUT_4[31297] = 32'b11111111111111111101000010100111;
assign LUT_4[31298] = 32'b00000000000000000011010001010011;
assign LUT_4[31299] = 32'b11111111111111111100011101001011;
assign LUT_4[31300] = 32'b00000000000000000000110111001011;
assign LUT_4[31301] = 32'b11111111111111111010000011000011;
assign LUT_4[31302] = 32'b00000000000000000000010001101111;
assign LUT_4[31303] = 32'b11111111111111111001011101100111;
assign LUT_4[31304] = 32'b11111111111111111101000011000100;
assign LUT_4[31305] = 32'b11111111111111110110001110111100;
assign LUT_4[31306] = 32'b11111111111111111100011101101000;
assign LUT_4[31307] = 32'b11111111111111110101101001100000;
assign LUT_4[31308] = 32'b11111111111111111010000011100000;
assign LUT_4[31309] = 32'b11111111111111110011001111011000;
assign LUT_4[31310] = 32'b11111111111111111001011110000100;
assign LUT_4[31311] = 32'b11111111111111110010101001111100;
assign LUT_4[31312] = 32'b00000000000000000001101000011101;
assign LUT_4[31313] = 32'b11111111111111111010110100010101;
assign LUT_4[31314] = 32'b00000000000000000001000011000001;
assign LUT_4[31315] = 32'b11111111111111111010001110111001;
assign LUT_4[31316] = 32'b11111111111111111110101000111001;
assign LUT_4[31317] = 32'b11111111111111110111110100110001;
assign LUT_4[31318] = 32'b11111111111111111110000011011101;
assign LUT_4[31319] = 32'b11111111111111110111001111010101;
assign LUT_4[31320] = 32'b11111111111111111010110100110010;
assign LUT_4[31321] = 32'b11111111111111110100000000101010;
assign LUT_4[31322] = 32'b11111111111111111010001111010110;
assign LUT_4[31323] = 32'b11111111111111110011011011001110;
assign LUT_4[31324] = 32'b11111111111111110111110101001110;
assign LUT_4[31325] = 32'b11111111111111110001000001000110;
assign LUT_4[31326] = 32'b11111111111111110111001111110010;
assign LUT_4[31327] = 32'b11111111111111110000011011101010;
assign LUT_4[31328] = 32'b00000000000000000010010001110110;
assign LUT_4[31329] = 32'b11111111111111111011011101101110;
assign LUT_4[31330] = 32'b00000000000000000001101100011010;
assign LUT_4[31331] = 32'b11111111111111111010111000010010;
assign LUT_4[31332] = 32'b11111111111111111111010010010010;
assign LUT_4[31333] = 32'b11111111111111111000011110001010;
assign LUT_4[31334] = 32'b11111111111111111110101100110110;
assign LUT_4[31335] = 32'b11111111111111110111111000101110;
assign LUT_4[31336] = 32'b11111111111111111011011110001011;
assign LUT_4[31337] = 32'b11111111111111110100101010000011;
assign LUT_4[31338] = 32'b11111111111111111010111000101111;
assign LUT_4[31339] = 32'b11111111111111110100000100100111;
assign LUT_4[31340] = 32'b11111111111111111000011110100111;
assign LUT_4[31341] = 32'b11111111111111110001101010011111;
assign LUT_4[31342] = 32'b11111111111111110111111001001011;
assign LUT_4[31343] = 32'b11111111111111110001000101000011;
assign LUT_4[31344] = 32'b00000000000000000000000011100100;
assign LUT_4[31345] = 32'b11111111111111111001001111011100;
assign LUT_4[31346] = 32'b11111111111111111111011110001000;
assign LUT_4[31347] = 32'b11111111111111111000101010000000;
assign LUT_4[31348] = 32'b11111111111111111101000100000000;
assign LUT_4[31349] = 32'b11111111111111110110001111111000;
assign LUT_4[31350] = 32'b11111111111111111100011110100100;
assign LUT_4[31351] = 32'b11111111111111110101101010011100;
assign LUT_4[31352] = 32'b11111111111111111001001111111001;
assign LUT_4[31353] = 32'b11111111111111110010011011110001;
assign LUT_4[31354] = 32'b11111111111111111000101010011101;
assign LUT_4[31355] = 32'b11111111111111110001110110010101;
assign LUT_4[31356] = 32'b11111111111111110110010000010101;
assign LUT_4[31357] = 32'b11111111111111101111011100001101;
assign LUT_4[31358] = 32'b11111111111111110101101010111001;
assign LUT_4[31359] = 32'b11111111111111101110110110110001;
assign LUT_4[31360] = 32'b00000000000000000101000101100011;
assign LUT_4[31361] = 32'b11111111111111111110010001011011;
assign LUT_4[31362] = 32'b00000000000000000100100000000111;
assign LUT_4[31363] = 32'b11111111111111111101101011111111;
assign LUT_4[31364] = 32'b00000000000000000010000101111111;
assign LUT_4[31365] = 32'b11111111111111111011010001110111;
assign LUT_4[31366] = 32'b00000000000000000001100000100011;
assign LUT_4[31367] = 32'b11111111111111111010101100011011;
assign LUT_4[31368] = 32'b11111111111111111110010001111000;
assign LUT_4[31369] = 32'b11111111111111110111011101110000;
assign LUT_4[31370] = 32'b11111111111111111101101100011100;
assign LUT_4[31371] = 32'b11111111111111110110111000010100;
assign LUT_4[31372] = 32'b11111111111111111011010010010100;
assign LUT_4[31373] = 32'b11111111111111110100011110001100;
assign LUT_4[31374] = 32'b11111111111111111010101100111000;
assign LUT_4[31375] = 32'b11111111111111110011111000110000;
assign LUT_4[31376] = 32'b00000000000000000010110111010001;
assign LUT_4[31377] = 32'b11111111111111111100000011001001;
assign LUT_4[31378] = 32'b00000000000000000010010001110101;
assign LUT_4[31379] = 32'b11111111111111111011011101101101;
assign LUT_4[31380] = 32'b11111111111111111111110111101101;
assign LUT_4[31381] = 32'b11111111111111111001000011100101;
assign LUT_4[31382] = 32'b11111111111111111111010010010001;
assign LUT_4[31383] = 32'b11111111111111111000011110001001;
assign LUT_4[31384] = 32'b11111111111111111100000011100110;
assign LUT_4[31385] = 32'b11111111111111110101001111011110;
assign LUT_4[31386] = 32'b11111111111111111011011110001010;
assign LUT_4[31387] = 32'b11111111111111110100101010000010;
assign LUT_4[31388] = 32'b11111111111111111001000100000010;
assign LUT_4[31389] = 32'b11111111111111110010001111111010;
assign LUT_4[31390] = 32'b11111111111111111000011110100110;
assign LUT_4[31391] = 32'b11111111111111110001101010011110;
assign LUT_4[31392] = 32'b00000000000000000011100000101010;
assign LUT_4[31393] = 32'b11111111111111111100101100100010;
assign LUT_4[31394] = 32'b00000000000000000010111011001110;
assign LUT_4[31395] = 32'b11111111111111111100000111000110;
assign LUT_4[31396] = 32'b00000000000000000000100001000110;
assign LUT_4[31397] = 32'b11111111111111111001101100111110;
assign LUT_4[31398] = 32'b11111111111111111111111011101010;
assign LUT_4[31399] = 32'b11111111111111111001000111100010;
assign LUT_4[31400] = 32'b11111111111111111100101100111111;
assign LUT_4[31401] = 32'b11111111111111110101111000110111;
assign LUT_4[31402] = 32'b11111111111111111100000111100011;
assign LUT_4[31403] = 32'b11111111111111110101010011011011;
assign LUT_4[31404] = 32'b11111111111111111001101101011011;
assign LUT_4[31405] = 32'b11111111111111110010111001010011;
assign LUT_4[31406] = 32'b11111111111111111001000111111111;
assign LUT_4[31407] = 32'b11111111111111110010010011110111;
assign LUT_4[31408] = 32'b00000000000000000001010010011000;
assign LUT_4[31409] = 32'b11111111111111111010011110010000;
assign LUT_4[31410] = 32'b00000000000000000000101100111100;
assign LUT_4[31411] = 32'b11111111111111111001111000110100;
assign LUT_4[31412] = 32'b11111111111111111110010010110100;
assign LUT_4[31413] = 32'b11111111111111110111011110101100;
assign LUT_4[31414] = 32'b11111111111111111101101101011000;
assign LUT_4[31415] = 32'b11111111111111110110111001010000;
assign LUT_4[31416] = 32'b11111111111111111010011110101101;
assign LUT_4[31417] = 32'b11111111111111110011101010100101;
assign LUT_4[31418] = 32'b11111111111111111001111001010001;
assign LUT_4[31419] = 32'b11111111111111110011000101001001;
assign LUT_4[31420] = 32'b11111111111111110111011111001001;
assign LUT_4[31421] = 32'b11111111111111110000101011000001;
assign LUT_4[31422] = 32'b11111111111111110110111001101101;
assign LUT_4[31423] = 32'b11111111111111110000000101100101;
assign LUT_4[31424] = 32'b00000000000000000110011100110111;
assign LUT_4[31425] = 32'b11111111111111111111101000101111;
assign LUT_4[31426] = 32'b00000000000000000101110111011011;
assign LUT_4[31427] = 32'b11111111111111111111000011010011;
assign LUT_4[31428] = 32'b00000000000000000011011101010011;
assign LUT_4[31429] = 32'b11111111111111111100101001001011;
assign LUT_4[31430] = 32'b00000000000000000010110111110111;
assign LUT_4[31431] = 32'b11111111111111111100000011101111;
assign LUT_4[31432] = 32'b11111111111111111111101001001100;
assign LUT_4[31433] = 32'b11111111111111111000110101000100;
assign LUT_4[31434] = 32'b11111111111111111111000011110000;
assign LUT_4[31435] = 32'b11111111111111111000001111101000;
assign LUT_4[31436] = 32'b11111111111111111100101001101000;
assign LUT_4[31437] = 32'b11111111111111110101110101100000;
assign LUT_4[31438] = 32'b11111111111111111100000100001100;
assign LUT_4[31439] = 32'b11111111111111110101010000000100;
assign LUT_4[31440] = 32'b00000000000000000100001110100101;
assign LUT_4[31441] = 32'b11111111111111111101011010011101;
assign LUT_4[31442] = 32'b00000000000000000011101001001001;
assign LUT_4[31443] = 32'b11111111111111111100110101000001;
assign LUT_4[31444] = 32'b00000000000000000001001111000001;
assign LUT_4[31445] = 32'b11111111111111111010011010111001;
assign LUT_4[31446] = 32'b00000000000000000000101001100101;
assign LUT_4[31447] = 32'b11111111111111111001110101011101;
assign LUT_4[31448] = 32'b11111111111111111101011010111010;
assign LUT_4[31449] = 32'b11111111111111110110100110110010;
assign LUT_4[31450] = 32'b11111111111111111100110101011110;
assign LUT_4[31451] = 32'b11111111111111110110000001010110;
assign LUT_4[31452] = 32'b11111111111111111010011011010110;
assign LUT_4[31453] = 32'b11111111111111110011100111001110;
assign LUT_4[31454] = 32'b11111111111111111001110101111010;
assign LUT_4[31455] = 32'b11111111111111110011000001110010;
assign LUT_4[31456] = 32'b00000000000000000100110111111110;
assign LUT_4[31457] = 32'b11111111111111111110000011110110;
assign LUT_4[31458] = 32'b00000000000000000100010010100010;
assign LUT_4[31459] = 32'b11111111111111111101011110011010;
assign LUT_4[31460] = 32'b00000000000000000001111000011010;
assign LUT_4[31461] = 32'b11111111111111111011000100010010;
assign LUT_4[31462] = 32'b00000000000000000001010010111110;
assign LUT_4[31463] = 32'b11111111111111111010011110110110;
assign LUT_4[31464] = 32'b11111111111111111110000100010011;
assign LUT_4[31465] = 32'b11111111111111110111010000001011;
assign LUT_4[31466] = 32'b11111111111111111101011110110111;
assign LUT_4[31467] = 32'b11111111111111110110101010101111;
assign LUT_4[31468] = 32'b11111111111111111011000100101111;
assign LUT_4[31469] = 32'b11111111111111110100010000100111;
assign LUT_4[31470] = 32'b11111111111111111010011111010011;
assign LUT_4[31471] = 32'b11111111111111110011101011001011;
assign LUT_4[31472] = 32'b00000000000000000010101001101100;
assign LUT_4[31473] = 32'b11111111111111111011110101100100;
assign LUT_4[31474] = 32'b00000000000000000010000100010000;
assign LUT_4[31475] = 32'b11111111111111111011010000001000;
assign LUT_4[31476] = 32'b11111111111111111111101010001000;
assign LUT_4[31477] = 32'b11111111111111111000110110000000;
assign LUT_4[31478] = 32'b11111111111111111111000100101100;
assign LUT_4[31479] = 32'b11111111111111111000010000100100;
assign LUT_4[31480] = 32'b11111111111111111011110110000001;
assign LUT_4[31481] = 32'b11111111111111110101000001111001;
assign LUT_4[31482] = 32'b11111111111111111011010000100101;
assign LUT_4[31483] = 32'b11111111111111110100011100011101;
assign LUT_4[31484] = 32'b11111111111111111000110110011101;
assign LUT_4[31485] = 32'b11111111111111110010000010010101;
assign LUT_4[31486] = 32'b11111111111111111000010001000001;
assign LUT_4[31487] = 32'b11111111111111110001011100111001;
assign LUT_4[31488] = 32'b00000000000000000111011010111110;
assign LUT_4[31489] = 32'b00000000000000000000100110110110;
assign LUT_4[31490] = 32'b00000000000000000110110101100010;
assign LUT_4[31491] = 32'b00000000000000000000000001011010;
assign LUT_4[31492] = 32'b00000000000000000100011011011010;
assign LUT_4[31493] = 32'b11111111111111111101100111010010;
assign LUT_4[31494] = 32'b00000000000000000011110101111110;
assign LUT_4[31495] = 32'b11111111111111111101000001110110;
assign LUT_4[31496] = 32'b00000000000000000000100111010011;
assign LUT_4[31497] = 32'b11111111111111111001110011001011;
assign LUT_4[31498] = 32'b00000000000000000000000001110111;
assign LUT_4[31499] = 32'b11111111111111111001001101101111;
assign LUT_4[31500] = 32'b11111111111111111101100111101111;
assign LUT_4[31501] = 32'b11111111111111110110110011100111;
assign LUT_4[31502] = 32'b11111111111111111101000010010011;
assign LUT_4[31503] = 32'b11111111111111110110001110001011;
assign LUT_4[31504] = 32'b00000000000000000101001100101100;
assign LUT_4[31505] = 32'b11111111111111111110011000100100;
assign LUT_4[31506] = 32'b00000000000000000100100111010000;
assign LUT_4[31507] = 32'b11111111111111111101110011001000;
assign LUT_4[31508] = 32'b00000000000000000010001101001000;
assign LUT_4[31509] = 32'b11111111111111111011011001000000;
assign LUT_4[31510] = 32'b00000000000000000001100111101100;
assign LUT_4[31511] = 32'b11111111111111111010110011100100;
assign LUT_4[31512] = 32'b11111111111111111110011001000001;
assign LUT_4[31513] = 32'b11111111111111110111100100111001;
assign LUT_4[31514] = 32'b11111111111111111101110011100101;
assign LUT_4[31515] = 32'b11111111111111110110111111011101;
assign LUT_4[31516] = 32'b11111111111111111011011001011101;
assign LUT_4[31517] = 32'b11111111111111110100100101010101;
assign LUT_4[31518] = 32'b11111111111111111010110100000001;
assign LUT_4[31519] = 32'b11111111111111110011111111111001;
assign LUT_4[31520] = 32'b00000000000000000101110110000101;
assign LUT_4[31521] = 32'b11111111111111111111000001111101;
assign LUT_4[31522] = 32'b00000000000000000101010000101001;
assign LUT_4[31523] = 32'b11111111111111111110011100100001;
assign LUT_4[31524] = 32'b00000000000000000010110110100001;
assign LUT_4[31525] = 32'b11111111111111111100000010011001;
assign LUT_4[31526] = 32'b00000000000000000010010001000101;
assign LUT_4[31527] = 32'b11111111111111111011011100111101;
assign LUT_4[31528] = 32'b11111111111111111111000010011010;
assign LUT_4[31529] = 32'b11111111111111111000001110010010;
assign LUT_4[31530] = 32'b11111111111111111110011100111110;
assign LUT_4[31531] = 32'b11111111111111110111101000110110;
assign LUT_4[31532] = 32'b11111111111111111100000010110110;
assign LUT_4[31533] = 32'b11111111111111110101001110101110;
assign LUT_4[31534] = 32'b11111111111111111011011101011010;
assign LUT_4[31535] = 32'b11111111111111110100101001010010;
assign LUT_4[31536] = 32'b00000000000000000011100111110011;
assign LUT_4[31537] = 32'b11111111111111111100110011101011;
assign LUT_4[31538] = 32'b00000000000000000011000010010111;
assign LUT_4[31539] = 32'b11111111111111111100001110001111;
assign LUT_4[31540] = 32'b00000000000000000000101000001111;
assign LUT_4[31541] = 32'b11111111111111111001110100000111;
assign LUT_4[31542] = 32'b00000000000000000000000010110011;
assign LUT_4[31543] = 32'b11111111111111111001001110101011;
assign LUT_4[31544] = 32'b11111111111111111100110100001000;
assign LUT_4[31545] = 32'b11111111111111110110000000000000;
assign LUT_4[31546] = 32'b11111111111111111100001110101100;
assign LUT_4[31547] = 32'b11111111111111110101011010100100;
assign LUT_4[31548] = 32'b11111111111111111001110100100100;
assign LUT_4[31549] = 32'b11111111111111110011000000011100;
assign LUT_4[31550] = 32'b11111111111111111001001111001000;
assign LUT_4[31551] = 32'b11111111111111110010011011000000;
assign LUT_4[31552] = 32'b00000000000000001000110010010010;
assign LUT_4[31553] = 32'b00000000000000000001111110001010;
assign LUT_4[31554] = 32'b00000000000000001000001100110110;
assign LUT_4[31555] = 32'b00000000000000000001011000101110;
assign LUT_4[31556] = 32'b00000000000000000101110010101110;
assign LUT_4[31557] = 32'b11111111111111111110111110100110;
assign LUT_4[31558] = 32'b00000000000000000101001101010010;
assign LUT_4[31559] = 32'b11111111111111111110011001001010;
assign LUT_4[31560] = 32'b00000000000000000001111110100111;
assign LUT_4[31561] = 32'b11111111111111111011001010011111;
assign LUT_4[31562] = 32'b00000000000000000001011001001011;
assign LUT_4[31563] = 32'b11111111111111111010100101000011;
assign LUT_4[31564] = 32'b11111111111111111110111111000011;
assign LUT_4[31565] = 32'b11111111111111111000001010111011;
assign LUT_4[31566] = 32'b11111111111111111110011001100111;
assign LUT_4[31567] = 32'b11111111111111110111100101011111;
assign LUT_4[31568] = 32'b00000000000000000110100100000000;
assign LUT_4[31569] = 32'b11111111111111111111101111111000;
assign LUT_4[31570] = 32'b00000000000000000101111110100100;
assign LUT_4[31571] = 32'b11111111111111111111001010011100;
assign LUT_4[31572] = 32'b00000000000000000011100100011100;
assign LUT_4[31573] = 32'b11111111111111111100110000010100;
assign LUT_4[31574] = 32'b00000000000000000010111111000000;
assign LUT_4[31575] = 32'b11111111111111111100001010111000;
assign LUT_4[31576] = 32'b11111111111111111111110000010101;
assign LUT_4[31577] = 32'b11111111111111111000111100001101;
assign LUT_4[31578] = 32'b11111111111111111111001010111001;
assign LUT_4[31579] = 32'b11111111111111111000010110110001;
assign LUT_4[31580] = 32'b11111111111111111100110000110001;
assign LUT_4[31581] = 32'b11111111111111110101111100101001;
assign LUT_4[31582] = 32'b11111111111111111100001011010101;
assign LUT_4[31583] = 32'b11111111111111110101010111001101;
assign LUT_4[31584] = 32'b00000000000000000111001101011001;
assign LUT_4[31585] = 32'b00000000000000000000011001010001;
assign LUT_4[31586] = 32'b00000000000000000110100111111101;
assign LUT_4[31587] = 32'b11111111111111111111110011110101;
assign LUT_4[31588] = 32'b00000000000000000100001101110101;
assign LUT_4[31589] = 32'b11111111111111111101011001101101;
assign LUT_4[31590] = 32'b00000000000000000011101000011001;
assign LUT_4[31591] = 32'b11111111111111111100110100010001;
assign LUT_4[31592] = 32'b00000000000000000000011001101110;
assign LUT_4[31593] = 32'b11111111111111111001100101100110;
assign LUT_4[31594] = 32'b11111111111111111111110100010010;
assign LUT_4[31595] = 32'b11111111111111111001000000001010;
assign LUT_4[31596] = 32'b11111111111111111101011010001010;
assign LUT_4[31597] = 32'b11111111111111110110100110000010;
assign LUT_4[31598] = 32'b11111111111111111100110100101110;
assign LUT_4[31599] = 32'b11111111111111110110000000100110;
assign LUT_4[31600] = 32'b00000000000000000100111111000111;
assign LUT_4[31601] = 32'b11111111111111111110001010111111;
assign LUT_4[31602] = 32'b00000000000000000100011001101011;
assign LUT_4[31603] = 32'b11111111111111111101100101100011;
assign LUT_4[31604] = 32'b00000000000000000001111111100011;
assign LUT_4[31605] = 32'b11111111111111111011001011011011;
assign LUT_4[31606] = 32'b00000000000000000001011010000111;
assign LUT_4[31607] = 32'b11111111111111111010100101111111;
assign LUT_4[31608] = 32'b11111111111111111110001011011100;
assign LUT_4[31609] = 32'b11111111111111110111010111010100;
assign LUT_4[31610] = 32'b11111111111111111101100110000000;
assign LUT_4[31611] = 32'b11111111111111110110110001111000;
assign LUT_4[31612] = 32'b11111111111111111011001011111000;
assign LUT_4[31613] = 32'b11111111111111110100010111110000;
assign LUT_4[31614] = 32'b11111111111111111010100110011100;
assign LUT_4[31615] = 32'b11111111111111110011110010010100;
assign LUT_4[31616] = 32'b00000000000000001010000001000110;
assign LUT_4[31617] = 32'b00000000000000000011001100111110;
assign LUT_4[31618] = 32'b00000000000000001001011011101010;
assign LUT_4[31619] = 32'b00000000000000000010100111100010;
assign LUT_4[31620] = 32'b00000000000000000111000001100010;
assign LUT_4[31621] = 32'b00000000000000000000001101011010;
assign LUT_4[31622] = 32'b00000000000000000110011100000110;
assign LUT_4[31623] = 32'b11111111111111111111100111111110;
assign LUT_4[31624] = 32'b00000000000000000011001101011011;
assign LUT_4[31625] = 32'b11111111111111111100011001010011;
assign LUT_4[31626] = 32'b00000000000000000010100111111111;
assign LUT_4[31627] = 32'b11111111111111111011110011110111;
assign LUT_4[31628] = 32'b00000000000000000000001101110111;
assign LUT_4[31629] = 32'b11111111111111111001011001101111;
assign LUT_4[31630] = 32'b11111111111111111111101000011011;
assign LUT_4[31631] = 32'b11111111111111111000110100010011;
assign LUT_4[31632] = 32'b00000000000000000111110010110100;
assign LUT_4[31633] = 32'b00000000000000000000111110101100;
assign LUT_4[31634] = 32'b00000000000000000111001101011000;
assign LUT_4[31635] = 32'b00000000000000000000011001010000;
assign LUT_4[31636] = 32'b00000000000000000100110011010000;
assign LUT_4[31637] = 32'b11111111111111111101111111001000;
assign LUT_4[31638] = 32'b00000000000000000100001101110100;
assign LUT_4[31639] = 32'b11111111111111111101011001101100;
assign LUT_4[31640] = 32'b00000000000000000000111111001001;
assign LUT_4[31641] = 32'b11111111111111111010001011000001;
assign LUT_4[31642] = 32'b00000000000000000000011001101101;
assign LUT_4[31643] = 32'b11111111111111111001100101100101;
assign LUT_4[31644] = 32'b11111111111111111101111111100101;
assign LUT_4[31645] = 32'b11111111111111110111001011011101;
assign LUT_4[31646] = 32'b11111111111111111101011010001001;
assign LUT_4[31647] = 32'b11111111111111110110100110000001;
assign LUT_4[31648] = 32'b00000000000000001000011100001101;
assign LUT_4[31649] = 32'b00000000000000000001101000000101;
assign LUT_4[31650] = 32'b00000000000000000111110110110001;
assign LUT_4[31651] = 32'b00000000000000000001000010101001;
assign LUT_4[31652] = 32'b00000000000000000101011100101001;
assign LUT_4[31653] = 32'b11111111111111111110101000100001;
assign LUT_4[31654] = 32'b00000000000000000100110111001101;
assign LUT_4[31655] = 32'b11111111111111111110000011000101;
assign LUT_4[31656] = 32'b00000000000000000001101000100010;
assign LUT_4[31657] = 32'b11111111111111111010110100011010;
assign LUT_4[31658] = 32'b00000000000000000001000011000110;
assign LUT_4[31659] = 32'b11111111111111111010001110111110;
assign LUT_4[31660] = 32'b11111111111111111110101000111110;
assign LUT_4[31661] = 32'b11111111111111110111110100110110;
assign LUT_4[31662] = 32'b11111111111111111110000011100010;
assign LUT_4[31663] = 32'b11111111111111110111001111011010;
assign LUT_4[31664] = 32'b00000000000000000110001101111011;
assign LUT_4[31665] = 32'b11111111111111111111011001110011;
assign LUT_4[31666] = 32'b00000000000000000101101000011111;
assign LUT_4[31667] = 32'b11111111111111111110110100010111;
assign LUT_4[31668] = 32'b00000000000000000011001110010111;
assign LUT_4[31669] = 32'b11111111111111111100011010001111;
assign LUT_4[31670] = 32'b00000000000000000010101000111011;
assign LUT_4[31671] = 32'b11111111111111111011110100110011;
assign LUT_4[31672] = 32'b11111111111111111111011010010000;
assign LUT_4[31673] = 32'b11111111111111111000100110001000;
assign LUT_4[31674] = 32'b11111111111111111110110100110100;
assign LUT_4[31675] = 32'b11111111111111111000000000101100;
assign LUT_4[31676] = 32'b11111111111111111100011010101100;
assign LUT_4[31677] = 32'b11111111111111110101100110100100;
assign LUT_4[31678] = 32'b11111111111111111011110101010000;
assign LUT_4[31679] = 32'b11111111111111110101000001001000;
assign LUT_4[31680] = 32'b00000000000000001011011000011010;
assign LUT_4[31681] = 32'b00000000000000000100100100010010;
assign LUT_4[31682] = 32'b00000000000000001010110010111110;
assign LUT_4[31683] = 32'b00000000000000000011111110110110;
assign LUT_4[31684] = 32'b00000000000000001000011000110110;
assign LUT_4[31685] = 32'b00000000000000000001100100101110;
assign LUT_4[31686] = 32'b00000000000000000111110011011010;
assign LUT_4[31687] = 32'b00000000000000000000111111010010;
assign LUT_4[31688] = 32'b00000000000000000100100100101111;
assign LUT_4[31689] = 32'b11111111111111111101110000100111;
assign LUT_4[31690] = 32'b00000000000000000011111111010011;
assign LUT_4[31691] = 32'b11111111111111111101001011001011;
assign LUT_4[31692] = 32'b00000000000000000001100101001011;
assign LUT_4[31693] = 32'b11111111111111111010110001000011;
assign LUT_4[31694] = 32'b00000000000000000000111111101111;
assign LUT_4[31695] = 32'b11111111111111111010001011100111;
assign LUT_4[31696] = 32'b00000000000000001001001010001000;
assign LUT_4[31697] = 32'b00000000000000000010010110000000;
assign LUT_4[31698] = 32'b00000000000000001000100100101100;
assign LUT_4[31699] = 32'b00000000000000000001110000100100;
assign LUT_4[31700] = 32'b00000000000000000110001010100100;
assign LUT_4[31701] = 32'b11111111111111111111010110011100;
assign LUT_4[31702] = 32'b00000000000000000101100101001000;
assign LUT_4[31703] = 32'b11111111111111111110110001000000;
assign LUT_4[31704] = 32'b00000000000000000010010110011101;
assign LUT_4[31705] = 32'b11111111111111111011100010010101;
assign LUT_4[31706] = 32'b00000000000000000001110001000001;
assign LUT_4[31707] = 32'b11111111111111111010111100111001;
assign LUT_4[31708] = 32'b11111111111111111111010110111001;
assign LUT_4[31709] = 32'b11111111111111111000100010110001;
assign LUT_4[31710] = 32'b11111111111111111110110001011101;
assign LUT_4[31711] = 32'b11111111111111110111111101010101;
assign LUT_4[31712] = 32'b00000000000000001001110011100001;
assign LUT_4[31713] = 32'b00000000000000000010111111011001;
assign LUT_4[31714] = 32'b00000000000000001001001110000101;
assign LUT_4[31715] = 32'b00000000000000000010011001111101;
assign LUT_4[31716] = 32'b00000000000000000110110011111101;
assign LUT_4[31717] = 32'b11111111111111111111111111110101;
assign LUT_4[31718] = 32'b00000000000000000110001110100001;
assign LUT_4[31719] = 32'b11111111111111111111011010011001;
assign LUT_4[31720] = 32'b00000000000000000010111111110110;
assign LUT_4[31721] = 32'b11111111111111111100001011101110;
assign LUT_4[31722] = 32'b00000000000000000010011010011010;
assign LUT_4[31723] = 32'b11111111111111111011100110010010;
assign LUT_4[31724] = 32'b00000000000000000000000000010010;
assign LUT_4[31725] = 32'b11111111111111111001001100001010;
assign LUT_4[31726] = 32'b11111111111111111111011010110110;
assign LUT_4[31727] = 32'b11111111111111111000100110101110;
assign LUT_4[31728] = 32'b00000000000000000111100101001111;
assign LUT_4[31729] = 32'b00000000000000000000110001000111;
assign LUT_4[31730] = 32'b00000000000000000110111111110011;
assign LUT_4[31731] = 32'b00000000000000000000001011101011;
assign LUT_4[31732] = 32'b00000000000000000100100101101011;
assign LUT_4[31733] = 32'b11111111111111111101110001100011;
assign LUT_4[31734] = 32'b00000000000000000100000000001111;
assign LUT_4[31735] = 32'b11111111111111111101001100000111;
assign LUT_4[31736] = 32'b00000000000000000000110001100100;
assign LUT_4[31737] = 32'b11111111111111111001111101011100;
assign LUT_4[31738] = 32'b00000000000000000000001100001000;
assign LUT_4[31739] = 32'b11111111111111111001011000000000;
assign LUT_4[31740] = 32'b11111111111111111101110010000000;
assign LUT_4[31741] = 32'b11111111111111110110111101111000;
assign LUT_4[31742] = 32'b11111111111111111101001100100100;
assign LUT_4[31743] = 32'b11111111111111110110011000011100;
assign LUT_4[31744] = 32'b00000000000000000101000101110010;
assign LUT_4[31745] = 32'b11111111111111111110010001101010;
assign LUT_4[31746] = 32'b00000000000000000100100000010110;
assign LUT_4[31747] = 32'b11111111111111111101101100001110;
assign LUT_4[31748] = 32'b00000000000000000010000110001110;
assign LUT_4[31749] = 32'b11111111111111111011010010000110;
assign LUT_4[31750] = 32'b00000000000000000001100000110010;
assign LUT_4[31751] = 32'b11111111111111111010101100101010;
assign LUT_4[31752] = 32'b11111111111111111110010010000111;
assign LUT_4[31753] = 32'b11111111111111110111011101111111;
assign LUT_4[31754] = 32'b11111111111111111101101100101011;
assign LUT_4[31755] = 32'b11111111111111110110111000100011;
assign LUT_4[31756] = 32'b11111111111111111011010010100011;
assign LUT_4[31757] = 32'b11111111111111110100011110011011;
assign LUT_4[31758] = 32'b11111111111111111010101101000111;
assign LUT_4[31759] = 32'b11111111111111110011111000111111;
assign LUT_4[31760] = 32'b00000000000000000010110111100000;
assign LUT_4[31761] = 32'b11111111111111111100000011011000;
assign LUT_4[31762] = 32'b00000000000000000010010010000100;
assign LUT_4[31763] = 32'b11111111111111111011011101111100;
assign LUT_4[31764] = 32'b11111111111111111111110111111100;
assign LUT_4[31765] = 32'b11111111111111111001000011110100;
assign LUT_4[31766] = 32'b11111111111111111111010010100000;
assign LUT_4[31767] = 32'b11111111111111111000011110011000;
assign LUT_4[31768] = 32'b11111111111111111100000011110101;
assign LUT_4[31769] = 32'b11111111111111110101001111101101;
assign LUT_4[31770] = 32'b11111111111111111011011110011001;
assign LUT_4[31771] = 32'b11111111111111110100101010010001;
assign LUT_4[31772] = 32'b11111111111111111001000100010001;
assign LUT_4[31773] = 32'b11111111111111110010010000001001;
assign LUT_4[31774] = 32'b11111111111111111000011110110101;
assign LUT_4[31775] = 32'b11111111111111110001101010101101;
assign LUT_4[31776] = 32'b00000000000000000011100000111001;
assign LUT_4[31777] = 32'b11111111111111111100101100110001;
assign LUT_4[31778] = 32'b00000000000000000010111011011101;
assign LUT_4[31779] = 32'b11111111111111111100000111010101;
assign LUT_4[31780] = 32'b00000000000000000000100001010101;
assign LUT_4[31781] = 32'b11111111111111111001101101001101;
assign LUT_4[31782] = 32'b11111111111111111111111011111001;
assign LUT_4[31783] = 32'b11111111111111111001000111110001;
assign LUT_4[31784] = 32'b11111111111111111100101101001110;
assign LUT_4[31785] = 32'b11111111111111110101111001000110;
assign LUT_4[31786] = 32'b11111111111111111100000111110010;
assign LUT_4[31787] = 32'b11111111111111110101010011101010;
assign LUT_4[31788] = 32'b11111111111111111001101101101010;
assign LUT_4[31789] = 32'b11111111111111110010111001100010;
assign LUT_4[31790] = 32'b11111111111111111001001000001110;
assign LUT_4[31791] = 32'b11111111111111110010010100000110;
assign LUT_4[31792] = 32'b00000000000000000001010010100111;
assign LUT_4[31793] = 32'b11111111111111111010011110011111;
assign LUT_4[31794] = 32'b00000000000000000000101101001011;
assign LUT_4[31795] = 32'b11111111111111111001111001000011;
assign LUT_4[31796] = 32'b11111111111111111110010011000011;
assign LUT_4[31797] = 32'b11111111111111110111011110111011;
assign LUT_4[31798] = 32'b11111111111111111101101101100111;
assign LUT_4[31799] = 32'b11111111111111110110111001011111;
assign LUT_4[31800] = 32'b11111111111111111010011110111100;
assign LUT_4[31801] = 32'b11111111111111110011101010110100;
assign LUT_4[31802] = 32'b11111111111111111001111001100000;
assign LUT_4[31803] = 32'b11111111111111110011000101011000;
assign LUT_4[31804] = 32'b11111111111111110111011111011000;
assign LUT_4[31805] = 32'b11111111111111110000101011010000;
assign LUT_4[31806] = 32'b11111111111111110110111001111100;
assign LUT_4[31807] = 32'b11111111111111110000000101110100;
assign LUT_4[31808] = 32'b00000000000000000110011101000110;
assign LUT_4[31809] = 32'b11111111111111111111101000111110;
assign LUT_4[31810] = 32'b00000000000000000101110111101010;
assign LUT_4[31811] = 32'b11111111111111111111000011100010;
assign LUT_4[31812] = 32'b00000000000000000011011101100010;
assign LUT_4[31813] = 32'b11111111111111111100101001011010;
assign LUT_4[31814] = 32'b00000000000000000010111000000110;
assign LUT_4[31815] = 32'b11111111111111111100000011111110;
assign LUT_4[31816] = 32'b11111111111111111111101001011011;
assign LUT_4[31817] = 32'b11111111111111111000110101010011;
assign LUT_4[31818] = 32'b11111111111111111111000011111111;
assign LUT_4[31819] = 32'b11111111111111111000001111110111;
assign LUT_4[31820] = 32'b11111111111111111100101001110111;
assign LUT_4[31821] = 32'b11111111111111110101110101101111;
assign LUT_4[31822] = 32'b11111111111111111100000100011011;
assign LUT_4[31823] = 32'b11111111111111110101010000010011;
assign LUT_4[31824] = 32'b00000000000000000100001110110100;
assign LUT_4[31825] = 32'b11111111111111111101011010101100;
assign LUT_4[31826] = 32'b00000000000000000011101001011000;
assign LUT_4[31827] = 32'b11111111111111111100110101010000;
assign LUT_4[31828] = 32'b00000000000000000001001111010000;
assign LUT_4[31829] = 32'b11111111111111111010011011001000;
assign LUT_4[31830] = 32'b00000000000000000000101001110100;
assign LUT_4[31831] = 32'b11111111111111111001110101101100;
assign LUT_4[31832] = 32'b11111111111111111101011011001001;
assign LUT_4[31833] = 32'b11111111111111110110100111000001;
assign LUT_4[31834] = 32'b11111111111111111100110101101101;
assign LUT_4[31835] = 32'b11111111111111110110000001100101;
assign LUT_4[31836] = 32'b11111111111111111010011011100101;
assign LUT_4[31837] = 32'b11111111111111110011100111011101;
assign LUT_4[31838] = 32'b11111111111111111001110110001001;
assign LUT_4[31839] = 32'b11111111111111110011000010000001;
assign LUT_4[31840] = 32'b00000000000000000100111000001101;
assign LUT_4[31841] = 32'b11111111111111111110000100000101;
assign LUT_4[31842] = 32'b00000000000000000100010010110001;
assign LUT_4[31843] = 32'b11111111111111111101011110101001;
assign LUT_4[31844] = 32'b00000000000000000001111000101001;
assign LUT_4[31845] = 32'b11111111111111111011000100100001;
assign LUT_4[31846] = 32'b00000000000000000001010011001101;
assign LUT_4[31847] = 32'b11111111111111111010011111000101;
assign LUT_4[31848] = 32'b11111111111111111110000100100010;
assign LUT_4[31849] = 32'b11111111111111110111010000011010;
assign LUT_4[31850] = 32'b11111111111111111101011111000110;
assign LUT_4[31851] = 32'b11111111111111110110101010111110;
assign LUT_4[31852] = 32'b11111111111111111011000100111110;
assign LUT_4[31853] = 32'b11111111111111110100010000110110;
assign LUT_4[31854] = 32'b11111111111111111010011111100010;
assign LUT_4[31855] = 32'b11111111111111110011101011011010;
assign LUT_4[31856] = 32'b00000000000000000010101001111011;
assign LUT_4[31857] = 32'b11111111111111111011110101110011;
assign LUT_4[31858] = 32'b00000000000000000010000100011111;
assign LUT_4[31859] = 32'b11111111111111111011010000010111;
assign LUT_4[31860] = 32'b11111111111111111111101010010111;
assign LUT_4[31861] = 32'b11111111111111111000110110001111;
assign LUT_4[31862] = 32'b11111111111111111111000100111011;
assign LUT_4[31863] = 32'b11111111111111111000010000110011;
assign LUT_4[31864] = 32'b11111111111111111011110110010000;
assign LUT_4[31865] = 32'b11111111111111110101000010001000;
assign LUT_4[31866] = 32'b11111111111111111011010000110100;
assign LUT_4[31867] = 32'b11111111111111110100011100101100;
assign LUT_4[31868] = 32'b11111111111111111000110110101100;
assign LUT_4[31869] = 32'b11111111111111110010000010100100;
assign LUT_4[31870] = 32'b11111111111111111000010001010000;
assign LUT_4[31871] = 32'b11111111111111110001011101001000;
assign LUT_4[31872] = 32'b00000000000000000111101011111010;
assign LUT_4[31873] = 32'b00000000000000000000110111110010;
assign LUT_4[31874] = 32'b00000000000000000111000110011110;
assign LUT_4[31875] = 32'b00000000000000000000010010010110;
assign LUT_4[31876] = 32'b00000000000000000100101100010110;
assign LUT_4[31877] = 32'b11111111111111111101111000001110;
assign LUT_4[31878] = 32'b00000000000000000100000110111010;
assign LUT_4[31879] = 32'b11111111111111111101010010110010;
assign LUT_4[31880] = 32'b00000000000000000000111000001111;
assign LUT_4[31881] = 32'b11111111111111111010000100000111;
assign LUT_4[31882] = 32'b00000000000000000000010010110011;
assign LUT_4[31883] = 32'b11111111111111111001011110101011;
assign LUT_4[31884] = 32'b11111111111111111101111000101011;
assign LUT_4[31885] = 32'b11111111111111110111000100100011;
assign LUT_4[31886] = 32'b11111111111111111101010011001111;
assign LUT_4[31887] = 32'b11111111111111110110011111000111;
assign LUT_4[31888] = 32'b00000000000000000101011101101000;
assign LUT_4[31889] = 32'b11111111111111111110101001100000;
assign LUT_4[31890] = 32'b00000000000000000100111000001100;
assign LUT_4[31891] = 32'b11111111111111111110000100000100;
assign LUT_4[31892] = 32'b00000000000000000010011110000100;
assign LUT_4[31893] = 32'b11111111111111111011101001111100;
assign LUT_4[31894] = 32'b00000000000000000001111000101000;
assign LUT_4[31895] = 32'b11111111111111111011000100100000;
assign LUT_4[31896] = 32'b11111111111111111110101001111101;
assign LUT_4[31897] = 32'b11111111111111110111110101110101;
assign LUT_4[31898] = 32'b11111111111111111110000100100001;
assign LUT_4[31899] = 32'b11111111111111110111010000011001;
assign LUT_4[31900] = 32'b11111111111111111011101010011001;
assign LUT_4[31901] = 32'b11111111111111110100110110010001;
assign LUT_4[31902] = 32'b11111111111111111011000100111101;
assign LUT_4[31903] = 32'b11111111111111110100010000110101;
assign LUT_4[31904] = 32'b00000000000000000110000111000001;
assign LUT_4[31905] = 32'b11111111111111111111010010111001;
assign LUT_4[31906] = 32'b00000000000000000101100001100101;
assign LUT_4[31907] = 32'b11111111111111111110101101011101;
assign LUT_4[31908] = 32'b00000000000000000011000111011101;
assign LUT_4[31909] = 32'b11111111111111111100010011010101;
assign LUT_4[31910] = 32'b00000000000000000010100010000001;
assign LUT_4[31911] = 32'b11111111111111111011101101111001;
assign LUT_4[31912] = 32'b11111111111111111111010011010110;
assign LUT_4[31913] = 32'b11111111111111111000011111001110;
assign LUT_4[31914] = 32'b11111111111111111110101101111010;
assign LUT_4[31915] = 32'b11111111111111110111111001110010;
assign LUT_4[31916] = 32'b11111111111111111100010011110010;
assign LUT_4[31917] = 32'b11111111111111110101011111101010;
assign LUT_4[31918] = 32'b11111111111111111011101110010110;
assign LUT_4[31919] = 32'b11111111111111110100111010001110;
assign LUT_4[31920] = 32'b00000000000000000011111000101111;
assign LUT_4[31921] = 32'b11111111111111111101000100100111;
assign LUT_4[31922] = 32'b00000000000000000011010011010011;
assign LUT_4[31923] = 32'b11111111111111111100011111001011;
assign LUT_4[31924] = 32'b00000000000000000000111001001011;
assign LUT_4[31925] = 32'b11111111111111111010000101000011;
assign LUT_4[31926] = 32'b00000000000000000000010011101111;
assign LUT_4[31927] = 32'b11111111111111111001011111100111;
assign LUT_4[31928] = 32'b11111111111111111101000101000100;
assign LUT_4[31929] = 32'b11111111111111110110010000111100;
assign LUT_4[31930] = 32'b11111111111111111100011111101000;
assign LUT_4[31931] = 32'b11111111111111110101101011100000;
assign LUT_4[31932] = 32'b11111111111111111010000101100000;
assign LUT_4[31933] = 32'b11111111111111110011010001011000;
assign LUT_4[31934] = 32'b11111111111111111001100000000100;
assign LUT_4[31935] = 32'b11111111111111110010101011111100;
assign LUT_4[31936] = 32'b00000000000000001001000011001110;
assign LUT_4[31937] = 32'b00000000000000000010001111000110;
assign LUT_4[31938] = 32'b00000000000000001000011101110010;
assign LUT_4[31939] = 32'b00000000000000000001101001101010;
assign LUT_4[31940] = 32'b00000000000000000110000011101010;
assign LUT_4[31941] = 32'b11111111111111111111001111100010;
assign LUT_4[31942] = 32'b00000000000000000101011110001110;
assign LUT_4[31943] = 32'b11111111111111111110101010000110;
assign LUT_4[31944] = 32'b00000000000000000010001111100011;
assign LUT_4[31945] = 32'b11111111111111111011011011011011;
assign LUT_4[31946] = 32'b00000000000000000001101010000111;
assign LUT_4[31947] = 32'b11111111111111111010110101111111;
assign LUT_4[31948] = 32'b11111111111111111111001111111111;
assign LUT_4[31949] = 32'b11111111111111111000011011110111;
assign LUT_4[31950] = 32'b11111111111111111110101010100011;
assign LUT_4[31951] = 32'b11111111111111110111110110011011;
assign LUT_4[31952] = 32'b00000000000000000110110100111100;
assign LUT_4[31953] = 32'b00000000000000000000000000110100;
assign LUT_4[31954] = 32'b00000000000000000110001111100000;
assign LUT_4[31955] = 32'b11111111111111111111011011011000;
assign LUT_4[31956] = 32'b00000000000000000011110101011000;
assign LUT_4[31957] = 32'b11111111111111111101000001010000;
assign LUT_4[31958] = 32'b00000000000000000011001111111100;
assign LUT_4[31959] = 32'b11111111111111111100011011110100;
assign LUT_4[31960] = 32'b00000000000000000000000001010001;
assign LUT_4[31961] = 32'b11111111111111111001001101001001;
assign LUT_4[31962] = 32'b11111111111111111111011011110101;
assign LUT_4[31963] = 32'b11111111111111111000100111101101;
assign LUT_4[31964] = 32'b11111111111111111101000001101101;
assign LUT_4[31965] = 32'b11111111111111110110001101100101;
assign LUT_4[31966] = 32'b11111111111111111100011100010001;
assign LUT_4[31967] = 32'b11111111111111110101101000001001;
assign LUT_4[31968] = 32'b00000000000000000111011110010101;
assign LUT_4[31969] = 32'b00000000000000000000101010001101;
assign LUT_4[31970] = 32'b00000000000000000110111000111001;
assign LUT_4[31971] = 32'b00000000000000000000000100110001;
assign LUT_4[31972] = 32'b00000000000000000100011110110001;
assign LUT_4[31973] = 32'b11111111111111111101101010101001;
assign LUT_4[31974] = 32'b00000000000000000011111001010101;
assign LUT_4[31975] = 32'b11111111111111111101000101001101;
assign LUT_4[31976] = 32'b00000000000000000000101010101010;
assign LUT_4[31977] = 32'b11111111111111111001110110100010;
assign LUT_4[31978] = 32'b00000000000000000000000101001110;
assign LUT_4[31979] = 32'b11111111111111111001010001000110;
assign LUT_4[31980] = 32'b11111111111111111101101011000110;
assign LUT_4[31981] = 32'b11111111111111110110110110111110;
assign LUT_4[31982] = 32'b11111111111111111101000101101010;
assign LUT_4[31983] = 32'b11111111111111110110010001100010;
assign LUT_4[31984] = 32'b00000000000000000101010000000011;
assign LUT_4[31985] = 32'b11111111111111111110011011111011;
assign LUT_4[31986] = 32'b00000000000000000100101010100111;
assign LUT_4[31987] = 32'b11111111111111111101110110011111;
assign LUT_4[31988] = 32'b00000000000000000010010000011111;
assign LUT_4[31989] = 32'b11111111111111111011011100010111;
assign LUT_4[31990] = 32'b00000000000000000001101011000011;
assign LUT_4[31991] = 32'b11111111111111111010110110111011;
assign LUT_4[31992] = 32'b11111111111111111110011100011000;
assign LUT_4[31993] = 32'b11111111111111110111101000010000;
assign LUT_4[31994] = 32'b11111111111111111101110110111100;
assign LUT_4[31995] = 32'b11111111111111110111000010110100;
assign LUT_4[31996] = 32'b11111111111111111011011100110100;
assign LUT_4[31997] = 32'b11111111111111110100101000101100;
assign LUT_4[31998] = 32'b11111111111111111010110111011000;
assign LUT_4[31999] = 32'b11111111111111110100000011010000;
assign LUT_4[32000] = 32'b00000000000000001010000001010101;
assign LUT_4[32001] = 32'b00000000000000000011001101001101;
assign LUT_4[32002] = 32'b00000000000000001001011011111001;
assign LUT_4[32003] = 32'b00000000000000000010100111110001;
assign LUT_4[32004] = 32'b00000000000000000111000001110001;
assign LUT_4[32005] = 32'b00000000000000000000001101101001;
assign LUT_4[32006] = 32'b00000000000000000110011100010101;
assign LUT_4[32007] = 32'b11111111111111111111101000001101;
assign LUT_4[32008] = 32'b00000000000000000011001101101010;
assign LUT_4[32009] = 32'b11111111111111111100011001100010;
assign LUT_4[32010] = 32'b00000000000000000010101000001110;
assign LUT_4[32011] = 32'b11111111111111111011110100000110;
assign LUT_4[32012] = 32'b00000000000000000000001110000110;
assign LUT_4[32013] = 32'b11111111111111111001011001111110;
assign LUT_4[32014] = 32'b11111111111111111111101000101010;
assign LUT_4[32015] = 32'b11111111111111111000110100100010;
assign LUT_4[32016] = 32'b00000000000000000111110011000011;
assign LUT_4[32017] = 32'b00000000000000000000111110111011;
assign LUT_4[32018] = 32'b00000000000000000111001101100111;
assign LUT_4[32019] = 32'b00000000000000000000011001011111;
assign LUT_4[32020] = 32'b00000000000000000100110011011111;
assign LUT_4[32021] = 32'b11111111111111111101111111010111;
assign LUT_4[32022] = 32'b00000000000000000100001110000011;
assign LUT_4[32023] = 32'b11111111111111111101011001111011;
assign LUT_4[32024] = 32'b00000000000000000000111111011000;
assign LUT_4[32025] = 32'b11111111111111111010001011010000;
assign LUT_4[32026] = 32'b00000000000000000000011001111100;
assign LUT_4[32027] = 32'b11111111111111111001100101110100;
assign LUT_4[32028] = 32'b11111111111111111101111111110100;
assign LUT_4[32029] = 32'b11111111111111110111001011101100;
assign LUT_4[32030] = 32'b11111111111111111101011010011000;
assign LUT_4[32031] = 32'b11111111111111110110100110010000;
assign LUT_4[32032] = 32'b00000000000000001000011100011100;
assign LUT_4[32033] = 32'b00000000000000000001101000010100;
assign LUT_4[32034] = 32'b00000000000000000111110111000000;
assign LUT_4[32035] = 32'b00000000000000000001000010111000;
assign LUT_4[32036] = 32'b00000000000000000101011100111000;
assign LUT_4[32037] = 32'b11111111111111111110101000110000;
assign LUT_4[32038] = 32'b00000000000000000100110111011100;
assign LUT_4[32039] = 32'b11111111111111111110000011010100;
assign LUT_4[32040] = 32'b00000000000000000001101000110001;
assign LUT_4[32041] = 32'b11111111111111111010110100101001;
assign LUT_4[32042] = 32'b00000000000000000001000011010101;
assign LUT_4[32043] = 32'b11111111111111111010001111001101;
assign LUT_4[32044] = 32'b11111111111111111110101001001101;
assign LUT_4[32045] = 32'b11111111111111110111110101000101;
assign LUT_4[32046] = 32'b11111111111111111110000011110001;
assign LUT_4[32047] = 32'b11111111111111110111001111101001;
assign LUT_4[32048] = 32'b00000000000000000110001110001010;
assign LUT_4[32049] = 32'b11111111111111111111011010000010;
assign LUT_4[32050] = 32'b00000000000000000101101000101110;
assign LUT_4[32051] = 32'b11111111111111111110110100100110;
assign LUT_4[32052] = 32'b00000000000000000011001110100110;
assign LUT_4[32053] = 32'b11111111111111111100011010011110;
assign LUT_4[32054] = 32'b00000000000000000010101001001010;
assign LUT_4[32055] = 32'b11111111111111111011110101000010;
assign LUT_4[32056] = 32'b11111111111111111111011010011111;
assign LUT_4[32057] = 32'b11111111111111111000100110010111;
assign LUT_4[32058] = 32'b11111111111111111110110101000011;
assign LUT_4[32059] = 32'b11111111111111111000000000111011;
assign LUT_4[32060] = 32'b11111111111111111100011010111011;
assign LUT_4[32061] = 32'b11111111111111110101100110110011;
assign LUT_4[32062] = 32'b11111111111111111011110101011111;
assign LUT_4[32063] = 32'b11111111111111110101000001010111;
assign LUT_4[32064] = 32'b00000000000000001011011000101001;
assign LUT_4[32065] = 32'b00000000000000000100100100100001;
assign LUT_4[32066] = 32'b00000000000000001010110011001101;
assign LUT_4[32067] = 32'b00000000000000000011111111000101;
assign LUT_4[32068] = 32'b00000000000000001000011001000101;
assign LUT_4[32069] = 32'b00000000000000000001100100111101;
assign LUT_4[32070] = 32'b00000000000000000111110011101001;
assign LUT_4[32071] = 32'b00000000000000000000111111100001;
assign LUT_4[32072] = 32'b00000000000000000100100100111110;
assign LUT_4[32073] = 32'b11111111111111111101110000110110;
assign LUT_4[32074] = 32'b00000000000000000011111111100010;
assign LUT_4[32075] = 32'b11111111111111111101001011011010;
assign LUT_4[32076] = 32'b00000000000000000001100101011010;
assign LUT_4[32077] = 32'b11111111111111111010110001010010;
assign LUT_4[32078] = 32'b00000000000000000000111111111110;
assign LUT_4[32079] = 32'b11111111111111111010001011110110;
assign LUT_4[32080] = 32'b00000000000000001001001010010111;
assign LUT_4[32081] = 32'b00000000000000000010010110001111;
assign LUT_4[32082] = 32'b00000000000000001000100100111011;
assign LUT_4[32083] = 32'b00000000000000000001110000110011;
assign LUT_4[32084] = 32'b00000000000000000110001010110011;
assign LUT_4[32085] = 32'b11111111111111111111010110101011;
assign LUT_4[32086] = 32'b00000000000000000101100101010111;
assign LUT_4[32087] = 32'b11111111111111111110110001001111;
assign LUT_4[32088] = 32'b00000000000000000010010110101100;
assign LUT_4[32089] = 32'b11111111111111111011100010100100;
assign LUT_4[32090] = 32'b00000000000000000001110001010000;
assign LUT_4[32091] = 32'b11111111111111111010111101001000;
assign LUT_4[32092] = 32'b11111111111111111111010111001000;
assign LUT_4[32093] = 32'b11111111111111111000100011000000;
assign LUT_4[32094] = 32'b11111111111111111110110001101100;
assign LUT_4[32095] = 32'b11111111111111110111111101100100;
assign LUT_4[32096] = 32'b00000000000000001001110011110000;
assign LUT_4[32097] = 32'b00000000000000000010111111101000;
assign LUT_4[32098] = 32'b00000000000000001001001110010100;
assign LUT_4[32099] = 32'b00000000000000000010011010001100;
assign LUT_4[32100] = 32'b00000000000000000110110100001100;
assign LUT_4[32101] = 32'b00000000000000000000000000000100;
assign LUT_4[32102] = 32'b00000000000000000110001110110000;
assign LUT_4[32103] = 32'b11111111111111111111011010101000;
assign LUT_4[32104] = 32'b00000000000000000011000000000101;
assign LUT_4[32105] = 32'b11111111111111111100001011111101;
assign LUT_4[32106] = 32'b00000000000000000010011010101001;
assign LUT_4[32107] = 32'b11111111111111111011100110100001;
assign LUT_4[32108] = 32'b00000000000000000000000000100001;
assign LUT_4[32109] = 32'b11111111111111111001001100011001;
assign LUT_4[32110] = 32'b11111111111111111111011011000101;
assign LUT_4[32111] = 32'b11111111111111111000100110111101;
assign LUT_4[32112] = 32'b00000000000000000111100101011110;
assign LUT_4[32113] = 32'b00000000000000000000110001010110;
assign LUT_4[32114] = 32'b00000000000000000111000000000010;
assign LUT_4[32115] = 32'b00000000000000000000001011111010;
assign LUT_4[32116] = 32'b00000000000000000100100101111010;
assign LUT_4[32117] = 32'b11111111111111111101110001110010;
assign LUT_4[32118] = 32'b00000000000000000100000000011110;
assign LUT_4[32119] = 32'b11111111111111111101001100010110;
assign LUT_4[32120] = 32'b00000000000000000000110001110011;
assign LUT_4[32121] = 32'b11111111111111111001111101101011;
assign LUT_4[32122] = 32'b00000000000000000000001100010111;
assign LUT_4[32123] = 32'b11111111111111111001011000001111;
assign LUT_4[32124] = 32'b11111111111111111101110010001111;
assign LUT_4[32125] = 32'b11111111111111110110111110000111;
assign LUT_4[32126] = 32'b11111111111111111101001100110011;
assign LUT_4[32127] = 32'b11111111111111110110011000101011;
assign LUT_4[32128] = 32'b00000000000000001100100111011101;
assign LUT_4[32129] = 32'b00000000000000000101110011010101;
assign LUT_4[32130] = 32'b00000000000000001100000010000001;
assign LUT_4[32131] = 32'b00000000000000000101001101111001;
assign LUT_4[32132] = 32'b00000000000000001001100111111001;
assign LUT_4[32133] = 32'b00000000000000000010110011110001;
assign LUT_4[32134] = 32'b00000000000000001001000010011101;
assign LUT_4[32135] = 32'b00000000000000000010001110010101;
assign LUT_4[32136] = 32'b00000000000000000101110011110010;
assign LUT_4[32137] = 32'b11111111111111111110111111101010;
assign LUT_4[32138] = 32'b00000000000000000101001110010110;
assign LUT_4[32139] = 32'b11111111111111111110011010001110;
assign LUT_4[32140] = 32'b00000000000000000010110100001110;
assign LUT_4[32141] = 32'b11111111111111111100000000000110;
assign LUT_4[32142] = 32'b00000000000000000010001110110010;
assign LUT_4[32143] = 32'b11111111111111111011011010101010;
assign LUT_4[32144] = 32'b00000000000000001010011001001011;
assign LUT_4[32145] = 32'b00000000000000000011100101000011;
assign LUT_4[32146] = 32'b00000000000000001001110011101111;
assign LUT_4[32147] = 32'b00000000000000000010111111100111;
assign LUT_4[32148] = 32'b00000000000000000111011001100111;
assign LUT_4[32149] = 32'b00000000000000000000100101011111;
assign LUT_4[32150] = 32'b00000000000000000110110100001011;
assign LUT_4[32151] = 32'b00000000000000000000000000000011;
assign LUT_4[32152] = 32'b00000000000000000011100101100000;
assign LUT_4[32153] = 32'b11111111111111111100110001011000;
assign LUT_4[32154] = 32'b00000000000000000011000000000100;
assign LUT_4[32155] = 32'b11111111111111111100001011111100;
assign LUT_4[32156] = 32'b00000000000000000000100101111100;
assign LUT_4[32157] = 32'b11111111111111111001110001110100;
assign LUT_4[32158] = 32'b00000000000000000000000000100000;
assign LUT_4[32159] = 32'b11111111111111111001001100011000;
assign LUT_4[32160] = 32'b00000000000000001011000010100100;
assign LUT_4[32161] = 32'b00000000000000000100001110011100;
assign LUT_4[32162] = 32'b00000000000000001010011101001000;
assign LUT_4[32163] = 32'b00000000000000000011101001000000;
assign LUT_4[32164] = 32'b00000000000000001000000011000000;
assign LUT_4[32165] = 32'b00000000000000000001001110111000;
assign LUT_4[32166] = 32'b00000000000000000111011101100100;
assign LUT_4[32167] = 32'b00000000000000000000101001011100;
assign LUT_4[32168] = 32'b00000000000000000100001110111001;
assign LUT_4[32169] = 32'b11111111111111111101011010110001;
assign LUT_4[32170] = 32'b00000000000000000011101001011101;
assign LUT_4[32171] = 32'b11111111111111111100110101010101;
assign LUT_4[32172] = 32'b00000000000000000001001111010101;
assign LUT_4[32173] = 32'b11111111111111111010011011001101;
assign LUT_4[32174] = 32'b00000000000000000000101001111001;
assign LUT_4[32175] = 32'b11111111111111111001110101110001;
assign LUT_4[32176] = 32'b00000000000000001000110100010010;
assign LUT_4[32177] = 32'b00000000000000000010000000001010;
assign LUT_4[32178] = 32'b00000000000000001000001110110110;
assign LUT_4[32179] = 32'b00000000000000000001011010101110;
assign LUT_4[32180] = 32'b00000000000000000101110100101110;
assign LUT_4[32181] = 32'b11111111111111111111000000100110;
assign LUT_4[32182] = 32'b00000000000000000101001111010010;
assign LUT_4[32183] = 32'b11111111111111111110011011001010;
assign LUT_4[32184] = 32'b00000000000000000010000000100111;
assign LUT_4[32185] = 32'b11111111111111111011001100011111;
assign LUT_4[32186] = 32'b00000000000000000001011011001011;
assign LUT_4[32187] = 32'b11111111111111111010100111000011;
assign LUT_4[32188] = 32'b11111111111111111111000001000011;
assign LUT_4[32189] = 32'b11111111111111111000001100111011;
assign LUT_4[32190] = 32'b11111111111111111110011011100111;
assign LUT_4[32191] = 32'b11111111111111110111100111011111;
assign LUT_4[32192] = 32'b00000000000000001101111110110001;
assign LUT_4[32193] = 32'b00000000000000000111001010101001;
assign LUT_4[32194] = 32'b00000000000000001101011001010101;
assign LUT_4[32195] = 32'b00000000000000000110100101001101;
assign LUT_4[32196] = 32'b00000000000000001010111111001101;
assign LUT_4[32197] = 32'b00000000000000000100001011000101;
assign LUT_4[32198] = 32'b00000000000000001010011001110001;
assign LUT_4[32199] = 32'b00000000000000000011100101101001;
assign LUT_4[32200] = 32'b00000000000000000111001011000110;
assign LUT_4[32201] = 32'b00000000000000000000010110111110;
assign LUT_4[32202] = 32'b00000000000000000110100101101010;
assign LUT_4[32203] = 32'b11111111111111111111110001100010;
assign LUT_4[32204] = 32'b00000000000000000100001011100010;
assign LUT_4[32205] = 32'b11111111111111111101010111011010;
assign LUT_4[32206] = 32'b00000000000000000011100110000110;
assign LUT_4[32207] = 32'b11111111111111111100110001111110;
assign LUT_4[32208] = 32'b00000000000000001011110000011111;
assign LUT_4[32209] = 32'b00000000000000000100111100010111;
assign LUT_4[32210] = 32'b00000000000000001011001011000011;
assign LUT_4[32211] = 32'b00000000000000000100010110111011;
assign LUT_4[32212] = 32'b00000000000000001000110000111011;
assign LUT_4[32213] = 32'b00000000000000000001111100110011;
assign LUT_4[32214] = 32'b00000000000000001000001011011111;
assign LUT_4[32215] = 32'b00000000000000000001010111010111;
assign LUT_4[32216] = 32'b00000000000000000100111100110100;
assign LUT_4[32217] = 32'b11111111111111111110001000101100;
assign LUT_4[32218] = 32'b00000000000000000100010111011000;
assign LUT_4[32219] = 32'b11111111111111111101100011010000;
assign LUT_4[32220] = 32'b00000000000000000001111101010000;
assign LUT_4[32221] = 32'b11111111111111111011001001001000;
assign LUT_4[32222] = 32'b00000000000000000001010111110100;
assign LUT_4[32223] = 32'b11111111111111111010100011101100;
assign LUT_4[32224] = 32'b00000000000000001100011001111000;
assign LUT_4[32225] = 32'b00000000000000000101100101110000;
assign LUT_4[32226] = 32'b00000000000000001011110100011100;
assign LUT_4[32227] = 32'b00000000000000000101000000010100;
assign LUT_4[32228] = 32'b00000000000000001001011010010100;
assign LUT_4[32229] = 32'b00000000000000000010100110001100;
assign LUT_4[32230] = 32'b00000000000000001000110100111000;
assign LUT_4[32231] = 32'b00000000000000000010000000110000;
assign LUT_4[32232] = 32'b00000000000000000101100110001101;
assign LUT_4[32233] = 32'b11111111111111111110110010000101;
assign LUT_4[32234] = 32'b00000000000000000101000000110001;
assign LUT_4[32235] = 32'b11111111111111111110001100101001;
assign LUT_4[32236] = 32'b00000000000000000010100110101001;
assign LUT_4[32237] = 32'b11111111111111111011110010100001;
assign LUT_4[32238] = 32'b00000000000000000010000001001101;
assign LUT_4[32239] = 32'b11111111111111111011001101000101;
assign LUT_4[32240] = 32'b00000000000000001010001011100110;
assign LUT_4[32241] = 32'b00000000000000000011010111011110;
assign LUT_4[32242] = 32'b00000000000000001001100110001010;
assign LUT_4[32243] = 32'b00000000000000000010110010000010;
assign LUT_4[32244] = 32'b00000000000000000111001100000010;
assign LUT_4[32245] = 32'b00000000000000000000010111111010;
assign LUT_4[32246] = 32'b00000000000000000110100110100110;
assign LUT_4[32247] = 32'b11111111111111111111110010011110;
assign LUT_4[32248] = 32'b00000000000000000011010111111011;
assign LUT_4[32249] = 32'b11111111111111111100100011110011;
assign LUT_4[32250] = 32'b00000000000000000010110010011111;
assign LUT_4[32251] = 32'b11111111111111111011111110010111;
assign LUT_4[32252] = 32'b00000000000000000000011000010111;
assign LUT_4[32253] = 32'b11111111111111111001100100001111;
assign LUT_4[32254] = 32'b11111111111111111111110010111011;
assign LUT_4[32255] = 32'b11111111111111111000111110110011;
assign LUT_4[32256] = 32'b00000000000000000100001001111010;
assign LUT_4[32257] = 32'b11111111111111111101010101110010;
assign LUT_4[32258] = 32'b00000000000000000011100100011110;
assign LUT_4[32259] = 32'b11111111111111111100110000010110;
assign LUT_4[32260] = 32'b00000000000000000001001010010110;
assign LUT_4[32261] = 32'b11111111111111111010010110001110;
assign LUT_4[32262] = 32'b00000000000000000000100100111010;
assign LUT_4[32263] = 32'b11111111111111111001110000110010;
assign LUT_4[32264] = 32'b11111111111111111101010110001111;
assign LUT_4[32265] = 32'b11111111111111110110100010000111;
assign LUT_4[32266] = 32'b11111111111111111100110000110011;
assign LUT_4[32267] = 32'b11111111111111110101111100101011;
assign LUT_4[32268] = 32'b11111111111111111010010110101011;
assign LUT_4[32269] = 32'b11111111111111110011100010100011;
assign LUT_4[32270] = 32'b11111111111111111001110001001111;
assign LUT_4[32271] = 32'b11111111111111110010111101000111;
assign LUT_4[32272] = 32'b00000000000000000001111011101000;
assign LUT_4[32273] = 32'b11111111111111111011000111100000;
assign LUT_4[32274] = 32'b00000000000000000001010110001100;
assign LUT_4[32275] = 32'b11111111111111111010100010000100;
assign LUT_4[32276] = 32'b11111111111111111110111100000100;
assign LUT_4[32277] = 32'b11111111111111111000000111111100;
assign LUT_4[32278] = 32'b11111111111111111110010110101000;
assign LUT_4[32279] = 32'b11111111111111110111100010100000;
assign LUT_4[32280] = 32'b11111111111111111011000111111101;
assign LUT_4[32281] = 32'b11111111111111110100010011110101;
assign LUT_4[32282] = 32'b11111111111111111010100010100001;
assign LUT_4[32283] = 32'b11111111111111110011101110011001;
assign LUT_4[32284] = 32'b11111111111111111000001000011001;
assign LUT_4[32285] = 32'b11111111111111110001010100010001;
assign LUT_4[32286] = 32'b11111111111111110111100010111101;
assign LUT_4[32287] = 32'b11111111111111110000101110110101;
assign LUT_4[32288] = 32'b00000000000000000010100101000001;
assign LUT_4[32289] = 32'b11111111111111111011110000111001;
assign LUT_4[32290] = 32'b00000000000000000001111111100101;
assign LUT_4[32291] = 32'b11111111111111111011001011011101;
assign LUT_4[32292] = 32'b11111111111111111111100101011101;
assign LUT_4[32293] = 32'b11111111111111111000110001010101;
assign LUT_4[32294] = 32'b11111111111111111111000000000001;
assign LUT_4[32295] = 32'b11111111111111111000001011111001;
assign LUT_4[32296] = 32'b11111111111111111011110001010110;
assign LUT_4[32297] = 32'b11111111111111110100111101001110;
assign LUT_4[32298] = 32'b11111111111111111011001011111010;
assign LUT_4[32299] = 32'b11111111111111110100010111110010;
assign LUT_4[32300] = 32'b11111111111111111000110001110010;
assign LUT_4[32301] = 32'b11111111111111110001111101101010;
assign LUT_4[32302] = 32'b11111111111111111000001100010110;
assign LUT_4[32303] = 32'b11111111111111110001011000001110;
assign LUT_4[32304] = 32'b00000000000000000000010110101111;
assign LUT_4[32305] = 32'b11111111111111111001100010100111;
assign LUT_4[32306] = 32'b11111111111111111111110001010011;
assign LUT_4[32307] = 32'b11111111111111111000111101001011;
assign LUT_4[32308] = 32'b11111111111111111101010111001011;
assign LUT_4[32309] = 32'b11111111111111110110100011000011;
assign LUT_4[32310] = 32'b11111111111111111100110001101111;
assign LUT_4[32311] = 32'b11111111111111110101111101100111;
assign LUT_4[32312] = 32'b11111111111111111001100011000100;
assign LUT_4[32313] = 32'b11111111111111110010101110111100;
assign LUT_4[32314] = 32'b11111111111111111000111101101000;
assign LUT_4[32315] = 32'b11111111111111110010001001100000;
assign LUT_4[32316] = 32'b11111111111111110110100011100000;
assign LUT_4[32317] = 32'b11111111111111101111101111011000;
assign LUT_4[32318] = 32'b11111111111111110101111110000100;
assign LUT_4[32319] = 32'b11111111111111101111001001111100;
assign LUT_4[32320] = 32'b00000000000000000101100001001110;
assign LUT_4[32321] = 32'b11111111111111111110101101000110;
assign LUT_4[32322] = 32'b00000000000000000100111011110010;
assign LUT_4[32323] = 32'b11111111111111111110000111101010;
assign LUT_4[32324] = 32'b00000000000000000010100001101010;
assign LUT_4[32325] = 32'b11111111111111111011101101100010;
assign LUT_4[32326] = 32'b00000000000000000001111100001110;
assign LUT_4[32327] = 32'b11111111111111111011001000000110;
assign LUT_4[32328] = 32'b11111111111111111110101101100011;
assign LUT_4[32329] = 32'b11111111111111110111111001011011;
assign LUT_4[32330] = 32'b11111111111111111110001000000111;
assign LUT_4[32331] = 32'b11111111111111110111010011111111;
assign LUT_4[32332] = 32'b11111111111111111011101101111111;
assign LUT_4[32333] = 32'b11111111111111110100111001110111;
assign LUT_4[32334] = 32'b11111111111111111011001000100011;
assign LUT_4[32335] = 32'b11111111111111110100010100011011;
assign LUT_4[32336] = 32'b00000000000000000011010010111100;
assign LUT_4[32337] = 32'b11111111111111111100011110110100;
assign LUT_4[32338] = 32'b00000000000000000010101101100000;
assign LUT_4[32339] = 32'b11111111111111111011111001011000;
assign LUT_4[32340] = 32'b00000000000000000000010011011000;
assign LUT_4[32341] = 32'b11111111111111111001011111010000;
assign LUT_4[32342] = 32'b11111111111111111111101101111100;
assign LUT_4[32343] = 32'b11111111111111111000111001110100;
assign LUT_4[32344] = 32'b11111111111111111100011111010001;
assign LUT_4[32345] = 32'b11111111111111110101101011001001;
assign LUT_4[32346] = 32'b11111111111111111011111001110101;
assign LUT_4[32347] = 32'b11111111111111110101000101101101;
assign LUT_4[32348] = 32'b11111111111111111001011111101101;
assign LUT_4[32349] = 32'b11111111111111110010101011100101;
assign LUT_4[32350] = 32'b11111111111111111000111010010001;
assign LUT_4[32351] = 32'b11111111111111110010000110001001;
assign LUT_4[32352] = 32'b00000000000000000011111100010101;
assign LUT_4[32353] = 32'b11111111111111111101001000001101;
assign LUT_4[32354] = 32'b00000000000000000011010110111001;
assign LUT_4[32355] = 32'b11111111111111111100100010110001;
assign LUT_4[32356] = 32'b00000000000000000000111100110001;
assign LUT_4[32357] = 32'b11111111111111111010001000101001;
assign LUT_4[32358] = 32'b00000000000000000000010111010101;
assign LUT_4[32359] = 32'b11111111111111111001100011001101;
assign LUT_4[32360] = 32'b11111111111111111101001000101010;
assign LUT_4[32361] = 32'b11111111111111110110010100100010;
assign LUT_4[32362] = 32'b11111111111111111100100011001110;
assign LUT_4[32363] = 32'b11111111111111110101101111000110;
assign LUT_4[32364] = 32'b11111111111111111010001001000110;
assign LUT_4[32365] = 32'b11111111111111110011010100111110;
assign LUT_4[32366] = 32'b11111111111111111001100011101010;
assign LUT_4[32367] = 32'b11111111111111110010101111100010;
assign LUT_4[32368] = 32'b00000000000000000001101110000011;
assign LUT_4[32369] = 32'b11111111111111111010111001111011;
assign LUT_4[32370] = 32'b00000000000000000001001000100111;
assign LUT_4[32371] = 32'b11111111111111111010010100011111;
assign LUT_4[32372] = 32'b11111111111111111110101110011111;
assign LUT_4[32373] = 32'b11111111111111110111111010010111;
assign LUT_4[32374] = 32'b11111111111111111110001001000011;
assign LUT_4[32375] = 32'b11111111111111110111010100111011;
assign LUT_4[32376] = 32'b11111111111111111010111010011000;
assign LUT_4[32377] = 32'b11111111111111110100000110010000;
assign LUT_4[32378] = 32'b11111111111111111010010100111100;
assign LUT_4[32379] = 32'b11111111111111110011100000110100;
assign LUT_4[32380] = 32'b11111111111111110111111010110100;
assign LUT_4[32381] = 32'b11111111111111110001000110101100;
assign LUT_4[32382] = 32'b11111111111111110111010101011000;
assign LUT_4[32383] = 32'b11111111111111110000100001010000;
assign LUT_4[32384] = 32'b00000000000000000110110000000010;
assign LUT_4[32385] = 32'b11111111111111111111111011111010;
assign LUT_4[32386] = 32'b00000000000000000110001010100110;
assign LUT_4[32387] = 32'b11111111111111111111010110011110;
assign LUT_4[32388] = 32'b00000000000000000011110000011110;
assign LUT_4[32389] = 32'b11111111111111111100111100010110;
assign LUT_4[32390] = 32'b00000000000000000011001011000010;
assign LUT_4[32391] = 32'b11111111111111111100010110111010;
assign LUT_4[32392] = 32'b11111111111111111111111100010111;
assign LUT_4[32393] = 32'b11111111111111111001001000001111;
assign LUT_4[32394] = 32'b11111111111111111111010110111011;
assign LUT_4[32395] = 32'b11111111111111111000100010110011;
assign LUT_4[32396] = 32'b11111111111111111100111100110011;
assign LUT_4[32397] = 32'b11111111111111110110001000101011;
assign LUT_4[32398] = 32'b11111111111111111100010111010111;
assign LUT_4[32399] = 32'b11111111111111110101100011001111;
assign LUT_4[32400] = 32'b00000000000000000100100001110000;
assign LUT_4[32401] = 32'b11111111111111111101101101101000;
assign LUT_4[32402] = 32'b00000000000000000011111100010100;
assign LUT_4[32403] = 32'b11111111111111111101001000001100;
assign LUT_4[32404] = 32'b00000000000000000001100010001100;
assign LUT_4[32405] = 32'b11111111111111111010101110000100;
assign LUT_4[32406] = 32'b00000000000000000000111100110000;
assign LUT_4[32407] = 32'b11111111111111111010001000101000;
assign LUT_4[32408] = 32'b11111111111111111101101110000101;
assign LUT_4[32409] = 32'b11111111111111110110111001111101;
assign LUT_4[32410] = 32'b11111111111111111101001000101001;
assign LUT_4[32411] = 32'b11111111111111110110010100100001;
assign LUT_4[32412] = 32'b11111111111111111010101110100001;
assign LUT_4[32413] = 32'b11111111111111110011111010011001;
assign LUT_4[32414] = 32'b11111111111111111010001001000101;
assign LUT_4[32415] = 32'b11111111111111110011010100111101;
assign LUT_4[32416] = 32'b00000000000000000101001011001001;
assign LUT_4[32417] = 32'b11111111111111111110010111000001;
assign LUT_4[32418] = 32'b00000000000000000100100101101101;
assign LUT_4[32419] = 32'b11111111111111111101110001100101;
assign LUT_4[32420] = 32'b00000000000000000010001011100101;
assign LUT_4[32421] = 32'b11111111111111111011010111011101;
assign LUT_4[32422] = 32'b00000000000000000001100110001001;
assign LUT_4[32423] = 32'b11111111111111111010110010000001;
assign LUT_4[32424] = 32'b11111111111111111110010111011110;
assign LUT_4[32425] = 32'b11111111111111110111100011010110;
assign LUT_4[32426] = 32'b11111111111111111101110010000010;
assign LUT_4[32427] = 32'b11111111111111110110111101111010;
assign LUT_4[32428] = 32'b11111111111111111011010111111010;
assign LUT_4[32429] = 32'b11111111111111110100100011110010;
assign LUT_4[32430] = 32'b11111111111111111010110010011110;
assign LUT_4[32431] = 32'b11111111111111110011111110010110;
assign LUT_4[32432] = 32'b00000000000000000010111100110111;
assign LUT_4[32433] = 32'b11111111111111111100001000101111;
assign LUT_4[32434] = 32'b00000000000000000010010111011011;
assign LUT_4[32435] = 32'b11111111111111111011100011010011;
assign LUT_4[32436] = 32'b11111111111111111111111101010011;
assign LUT_4[32437] = 32'b11111111111111111001001001001011;
assign LUT_4[32438] = 32'b11111111111111111111010111110111;
assign LUT_4[32439] = 32'b11111111111111111000100011101111;
assign LUT_4[32440] = 32'b11111111111111111100001001001100;
assign LUT_4[32441] = 32'b11111111111111110101010101000100;
assign LUT_4[32442] = 32'b11111111111111111011100011110000;
assign LUT_4[32443] = 32'b11111111111111110100101111101000;
assign LUT_4[32444] = 32'b11111111111111111001001001101000;
assign LUT_4[32445] = 32'b11111111111111110010010101100000;
assign LUT_4[32446] = 32'b11111111111111111000100100001100;
assign LUT_4[32447] = 32'b11111111111111110001110000000100;
assign LUT_4[32448] = 32'b00000000000000001000000111010110;
assign LUT_4[32449] = 32'b00000000000000000001010011001110;
assign LUT_4[32450] = 32'b00000000000000000111100001111010;
assign LUT_4[32451] = 32'b00000000000000000000101101110010;
assign LUT_4[32452] = 32'b00000000000000000101000111110010;
assign LUT_4[32453] = 32'b11111111111111111110010011101010;
assign LUT_4[32454] = 32'b00000000000000000100100010010110;
assign LUT_4[32455] = 32'b11111111111111111101101110001110;
assign LUT_4[32456] = 32'b00000000000000000001010011101011;
assign LUT_4[32457] = 32'b11111111111111111010011111100011;
assign LUT_4[32458] = 32'b00000000000000000000101110001111;
assign LUT_4[32459] = 32'b11111111111111111001111010000111;
assign LUT_4[32460] = 32'b11111111111111111110010100000111;
assign LUT_4[32461] = 32'b11111111111111110111011111111111;
assign LUT_4[32462] = 32'b11111111111111111101101110101011;
assign LUT_4[32463] = 32'b11111111111111110110111010100011;
assign LUT_4[32464] = 32'b00000000000000000101111001000100;
assign LUT_4[32465] = 32'b11111111111111111111000100111100;
assign LUT_4[32466] = 32'b00000000000000000101010011101000;
assign LUT_4[32467] = 32'b11111111111111111110011111100000;
assign LUT_4[32468] = 32'b00000000000000000010111001100000;
assign LUT_4[32469] = 32'b11111111111111111100000101011000;
assign LUT_4[32470] = 32'b00000000000000000010010100000100;
assign LUT_4[32471] = 32'b11111111111111111011011111111100;
assign LUT_4[32472] = 32'b11111111111111111111000101011001;
assign LUT_4[32473] = 32'b11111111111111111000010001010001;
assign LUT_4[32474] = 32'b11111111111111111110011111111101;
assign LUT_4[32475] = 32'b11111111111111110111101011110101;
assign LUT_4[32476] = 32'b11111111111111111100000101110101;
assign LUT_4[32477] = 32'b11111111111111110101010001101101;
assign LUT_4[32478] = 32'b11111111111111111011100000011001;
assign LUT_4[32479] = 32'b11111111111111110100101100010001;
assign LUT_4[32480] = 32'b00000000000000000110100010011101;
assign LUT_4[32481] = 32'b11111111111111111111101110010101;
assign LUT_4[32482] = 32'b00000000000000000101111101000001;
assign LUT_4[32483] = 32'b11111111111111111111001000111001;
assign LUT_4[32484] = 32'b00000000000000000011100010111001;
assign LUT_4[32485] = 32'b11111111111111111100101110110001;
assign LUT_4[32486] = 32'b00000000000000000010111101011101;
assign LUT_4[32487] = 32'b11111111111111111100001001010101;
assign LUT_4[32488] = 32'b11111111111111111111101110110010;
assign LUT_4[32489] = 32'b11111111111111111000111010101010;
assign LUT_4[32490] = 32'b11111111111111111111001001010110;
assign LUT_4[32491] = 32'b11111111111111111000010101001110;
assign LUT_4[32492] = 32'b11111111111111111100101111001110;
assign LUT_4[32493] = 32'b11111111111111110101111011000110;
assign LUT_4[32494] = 32'b11111111111111111100001001110010;
assign LUT_4[32495] = 32'b11111111111111110101010101101010;
assign LUT_4[32496] = 32'b00000000000000000100010100001011;
assign LUT_4[32497] = 32'b11111111111111111101100000000011;
assign LUT_4[32498] = 32'b00000000000000000011101110101111;
assign LUT_4[32499] = 32'b11111111111111111100111010100111;
assign LUT_4[32500] = 32'b00000000000000000001010100100111;
assign LUT_4[32501] = 32'b11111111111111111010100000011111;
assign LUT_4[32502] = 32'b00000000000000000000101111001011;
assign LUT_4[32503] = 32'b11111111111111111001111011000011;
assign LUT_4[32504] = 32'b11111111111111111101100000100000;
assign LUT_4[32505] = 32'b11111111111111110110101100011000;
assign LUT_4[32506] = 32'b11111111111111111100111011000100;
assign LUT_4[32507] = 32'b11111111111111110110000110111100;
assign LUT_4[32508] = 32'b11111111111111111010100000111100;
assign LUT_4[32509] = 32'b11111111111111110011101100110100;
assign LUT_4[32510] = 32'b11111111111111111001111011100000;
assign LUT_4[32511] = 32'b11111111111111110011000111011000;
assign LUT_4[32512] = 32'b00000000000000001001000101011101;
assign LUT_4[32513] = 32'b00000000000000000010010001010101;
assign LUT_4[32514] = 32'b00000000000000001000100000000001;
assign LUT_4[32515] = 32'b00000000000000000001101011111001;
assign LUT_4[32516] = 32'b00000000000000000110000101111001;
assign LUT_4[32517] = 32'b11111111111111111111010001110001;
assign LUT_4[32518] = 32'b00000000000000000101100000011101;
assign LUT_4[32519] = 32'b11111111111111111110101100010101;
assign LUT_4[32520] = 32'b00000000000000000010010001110010;
assign LUT_4[32521] = 32'b11111111111111111011011101101010;
assign LUT_4[32522] = 32'b00000000000000000001101100010110;
assign LUT_4[32523] = 32'b11111111111111111010111000001110;
assign LUT_4[32524] = 32'b11111111111111111111010010001110;
assign LUT_4[32525] = 32'b11111111111111111000011110000110;
assign LUT_4[32526] = 32'b11111111111111111110101100110010;
assign LUT_4[32527] = 32'b11111111111111110111111000101010;
assign LUT_4[32528] = 32'b00000000000000000110110111001011;
assign LUT_4[32529] = 32'b00000000000000000000000011000011;
assign LUT_4[32530] = 32'b00000000000000000110010001101111;
assign LUT_4[32531] = 32'b11111111111111111111011101100111;
assign LUT_4[32532] = 32'b00000000000000000011110111100111;
assign LUT_4[32533] = 32'b11111111111111111101000011011111;
assign LUT_4[32534] = 32'b00000000000000000011010010001011;
assign LUT_4[32535] = 32'b11111111111111111100011110000011;
assign LUT_4[32536] = 32'b00000000000000000000000011100000;
assign LUT_4[32537] = 32'b11111111111111111001001111011000;
assign LUT_4[32538] = 32'b11111111111111111111011110000100;
assign LUT_4[32539] = 32'b11111111111111111000101001111100;
assign LUT_4[32540] = 32'b11111111111111111101000011111100;
assign LUT_4[32541] = 32'b11111111111111110110001111110100;
assign LUT_4[32542] = 32'b11111111111111111100011110100000;
assign LUT_4[32543] = 32'b11111111111111110101101010011000;
assign LUT_4[32544] = 32'b00000000000000000111100000100100;
assign LUT_4[32545] = 32'b00000000000000000000101100011100;
assign LUT_4[32546] = 32'b00000000000000000110111011001000;
assign LUT_4[32547] = 32'b00000000000000000000000111000000;
assign LUT_4[32548] = 32'b00000000000000000100100001000000;
assign LUT_4[32549] = 32'b11111111111111111101101100111000;
assign LUT_4[32550] = 32'b00000000000000000011111011100100;
assign LUT_4[32551] = 32'b11111111111111111101000111011100;
assign LUT_4[32552] = 32'b00000000000000000000101100111001;
assign LUT_4[32553] = 32'b11111111111111111001111000110001;
assign LUT_4[32554] = 32'b00000000000000000000000111011101;
assign LUT_4[32555] = 32'b11111111111111111001010011010101;
assign LUT_4[32556] = 32'b11111111111111111101101101010101;
assign LUT_4[32557] = 32'b11111111111111110110111001001101;
assign LUT_4[32558] = 32'b11111111111111111101000111111001;
assign LUT_4[32559] = 32'b11111111111111110110010011110001;
assign LUT_4[32560] = 32'b00000000000000000101010010010010;
assign LUT_4[32561] = 32'b11111111111111111110011110001010;
assign LUT_4[32562] = 32'b00000000000000000100101100110110;
assign LUT_4[32563] = 32'b11111111111111111101111000101110;
assign LUT_4[32564] = 32'b00000000000000000010010010101110;
assign LUT_4[32565] = 32'b11111111111111111011011110100110;
assign LUT_4[32566] = 32'b00000000000000000001101101010010;
assign LUT_4[32567] = 32'b11111111111111111010111001001010;
assign LUT_4[32568] = 32'b11111111111111111110011110100111;
assign LUT_4[32569] = 32'b11111111111111110111101010011111;
assign LUT_4[32570] = 32'b11111111111111111101111001001011;
assign LUT_4[32571] = 32'b11111111111111110111000101000011;
assign LUT_4[32572] = 32'b11111111111111111011011111000011;
assign LUT_4[32573] = 32'b11111111111111110100101010111011;
assign LUT_4[32574] = 32'b11111111111111111010111001100111;
assign LUT_4[32575] = 32'b11111111111111110100000101011111;
assign LUT_4[32576] = 32'b00000000000000001010011100110001;
assign LUT_4[32577] = 32'b00000000000000000011101000101001;
assign LUT_4[32578] = 32'b00000000000000001001110111010101;
assign LUT_4[32579] = 32'b00000000000000000011000011001101;
assign LUT_4[32580] = 32'b00000000000000000111011101001101;
assign LUT_4[32581] = 32'b00000000000000000000101001000101;
assign LUT_4[32582] = 32'b00000000000000000110110111110001;
assign LUT_4[32583] = 32'b00000000000000000000000011101001;
assign LUT_4[32584] = 32'b00000000000000000011101001000110;
assign LUT_4[32585] = 32'b11111111111111111100110100111110;
assign LUT_4[32586] = 32'b00000000000000000011000011101010;
assign LUT_4[32587] = 32'b11111111111111111100001111100010;
assign LUT_4[32588] = 32'b00000000000000000000101001100010;
assign LUT_4[32589] = 32'b11111111111111111001110101011010;
assign LUT_4[32590] = 32'b00000000000000000000000100000110;
assign LUT_4[32591] = 32'b11111111111111111001001111111110;
assign LUT_4[32592] = 32'b00000000000000001000001110011111;
assign LUT_4[32593] = 32'b00000000000000000001011010010111;
assign LUT_4[32594] = 32'b00000000000000000111101001000011;
assign LUT_4[32595] = 32'b00000000000000000000110100111011;
assign LUT_4[32596] = 32'b00000000000000000101001110111011;
assign LUT_4[32597] = 32'b11111111111111111110011010110011;
assign LUT_4[32598] = 32'b00000000000000000100101001011111;
assign LUT_4[32599] = 32'b11111111111111111101110101010111;
assign LUT_4[32600] = 32'b00000000000000000001011010110100;
assign LUT_4[32601] = 32'b11111111111111111010100110101100;
assign LUT_4[32602] = 32'b00000000000000000000110101011000;
assign LUT_4[32603] = 32'b11111111111111111010000001010000;
assign LUT_4[32604] = 32'b11111111111111111110011011010000;
assign LUT_4[32605] = 32'b11111111111111110111100111001000;
assign LUT_4[32606] = 32'b11111111111111111101110101110100;
assign LUT_4[32607] = 32'b11111111111111110111000001101100;
assign LUT_4[32608] = 32'b00000000000000001000110111111000;
assign LUT_4[32609] = 32'b00000000000000000010000011110000;
assign LUT_4[32610] = 32'b00000000000000001000010010011100;
assign LUT_4[32611] = 32'b00000000000000000001011110010100;
assign LUT_4[32612] = 32'b00000000000000000101111000010100;
assign LUT_4[32613] = 32'b11111111111111111111000100001100;
assign LUT_4[32614] = 32'b00000000000000000101010010111000;
assign LUT_4[32615] = 32'b11111111111111111110011110110000;
assign LUT_4[32616] = 32'b00000000000000000010000100001101;
assign LUT_4[32617] = 32'b11111111111111111011010000000101;
assign LUT_4[32618] = 32'b00000000000000000001011110110001;
assign LUT_4[32619] = 32'b11111111111111111010101010101001;
assign LUT_4[32620] = 32'b11111111111111111111000100101001;
assign LUT_4[32621] = 32'b11111111111111111000010000100001;
assign LUT_4[32622] = 32'b11111111111111111110011111001101;
assign LUT_4[32623] = 32'b11111111111111110111101011000101;
assign LUT_4[32624] = 32'b00000000000000000110101001100110;
assign LUT_4[32625] = 32'b11111111111111111111110101011110;
assign LUT_4[32626] = 32'b00000000000000000110000100001010;
assign LUT_4[32627] = 32'b11111111111111111111010000000010;
assign LUT_4[32628] = 32'b00000000000000000011101010000010;
assign LUT_4[32629] = 32'b11111111111111111100110101111010;
assign LUT_4[32630] = 32'b00000000000000000011000100100110;
assign LUT_4[32631] = 32'b11111111111111111100010000011110;
assign LUT_4[32632] = 32'b11111111111111111111110101111011;
assign LUT_4[32633] = 32'b11111111111111111001000001110011;
assign LUT_4[32634] = 32'b11111111111111111111010000011111;
assign LUT_4[32635] = 32'b11111111111111111000011100010111;
assign LUT_4[32636] = 32'b11111111111111111100110110010111;
assign LUT_4[32637] = 32'b11111111111111110110000010001111;
assign LUT_4[32638] = 32'b11111111111111111100010000111011;
assign LUT_4[32639] = 32'b11111111111111110101011100110011;
assign LUT_4[32640] = 32'b00000000000000001011101011100101;
assign LUT_4[32641] = 32'b00000000000000000100110111011101;
assign LUT_4[32642] = 32'b00000000000000001011000110001001;
assign LUT_4[32643] = 32'b00000000000000000100010010000001;
assign LUT_4[32644] = 32'b00000000000000001000101100000001;
assign LUT_4[32645] = 32'b00000000000000000001110111111001;
assign LUT_4[32646] = 32'b00000000000000001000000110100101;
assign LUT_4[32647] = 32'b00000000000000000001010010011101;
assign LUT_4[32648] = 32'b00000000000000000100110111111010;
assign LUT_4[32649] = 32'b11111111111111111110000011110010;
assign LUT_4[32650] = 32'b00000000000000000100010010011110;
assign LUT_4[32651] = 32'b11111111111111111101011110010110;
assign LUT_4[32652] = 32'b00000000000000000001111000010110;
assign LUT_4[32653] = 32'b11111111111111111011000100001110;
assign LUT_4[32654] = 32'b00000000000000000001010010111010;
assign LUT_4[32655] = 32'b11111111111111111010011110110010;
assign LUT_4[32656] = 32'b00000000000000001001011101010011;
assign LUT_4[32657] = 32'b00000000000000000010101001001011;
assign LUT_4[32658] = 32'b00000000000000001000110111110111;
assign LUT_4[32659] = 32'b00000000000000000010000011101111;
assign LUT_4[32660] = 32'b00000000000000000110011101101111;
assign LUT_4[32661] = 32'b11111111111111111111101001100111;
assign LUT_4[32662] = 32'b00000000000000000101111000010011;
assign LUT_4[32663] = 32'b11111111111111111111000100001011;
assign LUT_4[32664] = 32'b00000000000000000010101001101000;
assign LUT_4[32665] = 32'b11111111111111111011110101100000;
assign LUT_4[32666] = 32'b00000000000000000010000100001100;
assign LUT_4[32667] = 32'b11111111111111111011010000000100;
assign LUT_4[32668] = 32'b11111111111111111111101010000100;
assign LUT_4[32669] = 32'b11111111111111111000110101111100;
assign LUT_4[32670] = 32'b11111111111111111111000100101000;
assign LUT_4[32671] = 32'b11111111111111111000010000100000;
assign LUT_4[32672] = 32'b00000000000000001010000110101100;
assign LUT_4[32673] = 32'b00000000000000000011010010100100;
assign LUT_4[32674] = 32'b00000000000000001001100001010000;
assign LUT_4[32675] = 32'b00000000000000000010101101001000;
assign LUT_4[32676] = 32'b00000000000000000111000111001000;
assign LUT_4[32677] = 32'b00000000000000000000010011000000;
assign LUT_4[32678] = 32'b00000000000000000110100001101100;
assign LUT_4[32679] = 32'b11111111111111111111101101100100;
assign LUT_4[32680] = 32'b00000000000000000011010011000001;
assign LUT_4[32681] = 32'b11111111111111111100011110111001;
assign LUT_4[32682] = 32'b00000000000000000010101101100101;
assign LUT_4[32683] = 32'b11111111111111111011111001011101;
assign LUT_4[32684] = 32'b00000000000000000000010011011101;
assign LUT_4[32685] = 32'b11111111111111111001011111010101;
assign LUT_4[32686] = 32'b11111111111111111111101110000001;
assign LUT_4[32687] = 32'b11111111111111111000111001111001;
assign LUT_4[32688] = 32'b00000000000000000111111000011010;
assign LUT_4[32689] = 32'b00000000000000000001000100010010;
assign LUT_4[32690] = 32'b00000000000000000111010010111110;
assign LUT_4[32691] = 32'b00000000000000000000011110110110;
assign LUT_4[32692] = 32'b00000000000000000100111000110110;
assign LUT_4[32693] = 32'b11111111111111111110000100101110;
assign LUT_4[32694] = 32'b00000000000000000100010011011010;
assign LUT_4[32695] = 32'b11111111111111111101011111010010;
assign LUT_4[32696] = 32'b00000000000000000001000100101111;
assign LUT_4[32697] = 32'b11111111111111111010010000100111;
assign LUT_4[32698] = 32'b00000000000000000000011111010011;
assign LUT_4[32699] = 32'b11111111111111111001101011001011;
assign LUT_4[32700] = 32'b11111111111111111110000101001011;
assign LUT_4[32701] = 32'b11111111111111110111010001000011;
assign LUT_4[32702] = 32'b11111111111111111101011111101111;
assign LUT_4[32703] = 32'b11111111111111110110101011100111;
assign LUT_4[32704] = 32'b00000000000000001101000010111001;
assign LUT_4[32705] = 32'b00000000000000000110001110110001;
assign LUT_4[32706] = 32'b00000000000000001100011101011101;
assign LUT_4[32707] = 32'b00000000000000000101101001010101;
assign LUT_4[32708] = 32'b00000000000000001010000011010101;
assign LUT_4[32709] = 32'b00000000000000000011001111001101;
assign LUT_4[32710] = 32'b00000000000000001001011101111001;
assign LUT_4[32711] = 32'b00000000000000000010101001110001;
assign LUT_4[32712] = 32'b00000000000000000110001111001110;
assign LUT_4[32713] = 32'b11111111111111111111011011000110;
assign LUT_4[32714] = 32'b00000000000000000101101001110010;
assign LUT_4[32715] = 32'b11111111111111111110110101101010;
assign LUT_4[32716] = 32'b00000000000000000011001111101010;
assign LUT_4[32717] = 32'b11111111111111111100011011100010;
assign LUT_4[32718] = 32'b00000000000000000010101010001110;
assign LUT_4[32719] = 32'b11111111111111111011110110000110;
assign LUT_4[32720] = 32'b00000000000000001010110100100111;
assign LUT_4[32721] = 32'b00000000000000000100000000011111;
assign LUT_4[32722] = 32'b00000000000000001010001111001011;
assign LUT_4[32723] = 32'b00000000000000000011011011000011;
assign LUT_4[32724] = 32'b00000000000000000111110101000011;
assign LUT_4[32725] = 32'b00000000000000000001000000111011;
assign LUT_4[32726] = 32'b00000000000000000111001111100111;
assign LUT_4[32727] = 32'b00000000000000000000011011011111;
assign LUT_4[32728] = 32'b00000000000000000100000000111100;
assign LUT_4[32729] = 32'b11111111111111111101001100110100;
assign LUT_4[32730] = 32'b00000000000000000011011011100000;
assign LUT_4[32731] = 32'b11111111111111111100100111011000;
assign LUT_4[32732] = 32'b00000000000000000001000001011000;
assign LUT_4[32733] = 32'b11111111111111111010001101010000;
assign LUT_4[32734] = 32'b00000000000000000000011011111100;
assign LUT_4[32735] = 32'b11111111111111111001100111110100;
assign LUT_4[32736] = 32'b00000000000000001011011110000000;
assign LUT_4[32737] = 32'b00000000000000000100101001111000;
assign LUT_4[32738] = 32'b00000000000000001010111000100100;
assign LUT_4[32739] = 32'b00000000000000000100000100011100;
assign LUT_4[32740] = 32'b00000000000000001000011110011100;
assign LUT_4[32741] = 32'b00000000000000000001101010010100;
assign LUT_4[32742] = 32'b00000000000000000111111001000000;
assign LUT_4[32743] = 32'b00000000000000000001000100111000;
assign LUT_4[32744] = 32'b00000000000000000100101010010101;
assign LUT_4[32745] = 32'b11111111111111111101110110001101;
assign LUT_4[32746] = 32'b00000000000000000100000100111001;
assign LUT_4[32747] = 32'b11111111111111111101010000110001;
assign LUT_4[32748] = 32'b00000000000000000001101010110001;
assign LUT_4[32749] = 32'b11111111111111111010110110101001;
assign LUT_4[32750] = 32'b00000000000000000001000101010101;
assign LUT_4[32751] = 32'b11111111111111111010010001001101;
assign LUT_4[32752] = 32'b00000000000000001001001111101110;
assign LUT_4[32753] = 32'b00000000000000000010011011100110;
assign LUT_4[32754] = 32'b00000000000000001000101010010010;
assign LUT_4[32755] = 32'b00000000000000000001110110001010;
assign LUT_4[32756] = 32'b00000000000000000110010000001010;
assign LUT_4[32757] = 32'b11111111111111111111011100000010;
assign LUT_4[32758] = 32'b00000000000000000101101010101110;
assign LUT_4[32759] = 32'b11111111111111111110110110100110;
assign LUT_4[32760] = 32'b00000000000000000010011100000011;
assign LUT_4[32761] = 32'b11111111111111111011100111111011;
assign LUT_4[32762] = 32'b00000000000000000001110110100111;
assign LUT_4[32763] = 32'b11111111111111111011000010011111;
assign LUT_4[32764] = 32'b11111111111111111111011100011111;
assign LUT_4[32765] = 32'b11111111111111111000101000010111;
assign LUT_4[32766] = 32'b11111111111111111110110111000011;
assign LUT_4[32767] = 32'b11111111111111111000000010111011;
assign LUT_4[32768] = 32'b00000000000000000111010100010100;
assign LUT_4[32769] = 32'b00000000000000000000100000001100;
assign LUT_4[32770] = 32'b00000000000000000110101110111000;
assign LUT_4[32771] = 32'b11111111111111111111111010110000;
assign LUT_4[32772] = 32'b00000000000000000100010100110000;
assign LUT_4[32773] = 32'b11111111111111111101100000101000;
assign LUT_4[32774] = 32'b00000000000000000011101111010100;
assign LUT_4[32775] = 32'b11111111111111111100111011001100;
assign LUT_4[32776] = 32'b00000000000000000000100000101001;
assign LUT_4[32777] = 32'b11111111111111111001101100100001;
assign LUT_4[32778] = 32'b11111111111111111111111011001101;
assign LUT_4[32779] = 32'b11111111111111111001000111000101;
assign LUT_4[32780] = 32'b11111111111111111101100001000101;
assign LUT_4[32781] = 32'b11111111111111110110101100111101;
assign LUT_4[32782] = 32'b11111111111111111100111011101001;
assign LUT_4[32783] = 32'b11111111111111110110000111100001;
assign LUT_4[32784] = 32'b00000000000000000101000110000010;
assign LUT_4[32785] = 32'b11111111111111111110010001111010;
assign LUT_4[32786] = 32'b00000000000000000100100000100110;
assign LUT_4[32787] = 32'b11111111111111111101101100011110;
assign LUT_4[32788] = 32'b00000000000000000010000110011110;
assign LUT_4[32789] = 32'b11111111111111111011010010010110;
assign LUT_4[32790] = 32'b00000000000000000001100001000010;
assign LUT_4[32791] = 32'b11111111111111111010101100111010;
assign LUT_4[32792] = 32'b11111111111111111110010010010111;
assign LUT_4[32793] = 32'b11111111111111110111011110001111;
assign LUT_4[32794] = 32'b11111111111111111101101100111011;
assign LUT_4[32795] = 32'b11111111111111110110111000110011;
assign LUT_4[32796] = 32'b11111111111111111011010010110011;
assign LUT_4[32797] = 32'b11111111111111110100011110101011;
assign LUT_4[32798] = 32'b11111111111111111010101101010111;
assign LUT_4[32799] = 32'b11111111111111110011111001001111;
assign LUT_4[32800] = 32'b00000000000000000101101111011011;
assign LUT_4[32801] = 32'b11111111111111111110111011010011;
assign LUT_4[32802] = 32'b00000000000000000101001001111111;
assign LUT_4[32803] = 32'b11111111111111111110010101110111;
assign LUT_4[32804] = 32'b00000000000000000010101111110111;
assign LUT_4[32805] = 32'b11111111111111111011111011101111;
assign LUT_4[32806] = 32'b00000000000000000010001010011011;
assign LUT_4[32807] = 32'b11111111111111111011010110010011;
assign LUT_4[32808] = 32'b11111111111111111110111011110000;
assign LUT_4[32809] = 32'b11111111111111111000000111101000;
assign LUT_4[32810] = 32'b11111111111111111110010110010100;
assign LUT_4[32811] = 32'b11111111111111110111100010001100;
assign LUT_4[32812] = 32'b11111111111111111011111100001100;
assign LUT_4[32813] = 32'b11111111111111110101001000000100;
assign LUT_4[32814] = 32'b11111111111111111011010110110000;
assign LUT_4[32815] = 32'b11111111111111110100100010101000;
assign LUT_4[32816] = 32'b00000000000000000011100001001001;
assign LUT_4[32817] = 32'b11111111111111111100101101000001;
assign LUT_4[32818] = 32'b00000000000000000010111011101101;
assign LUT_4[32819] = 32'b11111111111111111100000111100101;
assign LUT_4[32820] = 32'b00000000000000000000100001100101;
assign LUT_4[32821] = 32'b11111111111111111001101101011101;
assign LUT_4[32822] = 32'b11111111111111111111111100001001;
assign LUT_4[32823] = 32'b11111111111111111001001000000001;
assign LUT_4[32824] = 32'b11111111111111111100101101011110;
assign LUT_4[32825] = 32'b11111111111111110101111001010110;
assign LUT_4[32826] = 32'b11111111111111111100001000000010;
assign LUT_4[32827] = 32'b11111111111111110101010011111010;
assign LUT_4[32828] = 32'b11111111111111111001101101111010;
assign LUT_4[32829] = 32'b11111111111111110010111001110010;
assign LUT_4[32830] = 32'b11111111111111111001001000011110;
assign LUT_4[32831] = 32'b11111111111111110010010100010110;
assign LUT_4[32832] = 32'b00000000000000001000101011101000;
assign LUT_4[32833] = 32'b00000000000000000001110111100000;
assign LUT_4[32834] = 32'b00000000000000001000000110001100;
assign LUT_4[32835] = 32'b00000000000000000001010010000100;
assign LUT_4[32836] = 32'b00000000000000000101101100000100;
assign LUT_4[32837] = 32'b11111111111111111110110111111100;
assign LUT_4[32838] = 32'b00000000000000000101000110101000;
assign LUT_4[32839] = 32'b11111111111111111110010010100000;
assign LUT_4[32840] = 32'b00000000000000000001110111111101;
assign LUT_4[32841] = 32'b11111111111111111011000011110101;
assign LUT_4[32842] = 32'b00000000000000000001010010100001;
assign LUT_4[32843] = 32'b11111111111111111010011110011001;
assign LUT_4[32844] = 32'b11111111111111111110111000011001;
assign LUT_4[32845] = 32'b11111111111111111000000100010001;
assign LUT_4[32846] = 32'b11111111111111111110010010111101;
assign LUT_4[32847] = 32'b11111111111111110111011110110101;
assign LUT_4[32848] = 32'b00000000000000000110011101010110;
assign LUT_4[32849] = 32'b11111111111111111111101001001110;
assign LUT_4[32850] = 32'b00000000000000000101110111111010;
assign LUT_4[32851] = 32'b11111111111111111111000011110010;
assign LUT_4[32852] = 32'b00000000000000000011011101110010;
assign LUT_4[32853] = 32'b11111111111111111100101001101010;
assign LUT_4[32854] = 32'b00000000000000000010111000010110;
assign LUT_4[32855] = 32'b11111111111111111100000100001110;
assign LUT_4[32856] = 32'b11111111111111111111101001101011;
assign LUT_4[32857] = 32'b11111111111111111000110101100011;
assign LUT_4[32858] = 32'b11111111111111111111000100001111;
assign LUT_4[32859] = 32'b11111111111111111000010000000111;
assign LUT_4[32860] = 32'b11111111111111111100101010000111;
assign LUT_4[32861] = 32'b11111111111111110101110101111111;
assign LUT_4[32862] = 32'b11111111111111111100000100101011;
assign LUT_4[32863] = 32'b11111111111111110101010000100011;
assign LUT_4[32864] = 32'b00000000000000000111000110101111;
assign LUT_4[32865] = 32'b00000000000000000000010010100111;
assign LUT_4[32866] = 32'b00000000000000000110100001010011;
assign LUT_4[32867] = 32'b11111111111111111111101101001011;
assign LUT_4[32868] = 32'b00000000000000000100000111001011;
assign LUT_4[32869] = 32'b11111111111111111101010011000011;
assign LUT_4[32870] = 32'b00000000000000000011100001101111;
assign LUT_4[32871] = 32'b11111111111111111100101101100111;
assign LUT_4[32872] = 32'b00000000000000000000010011000100;
assign LUT_4[32873] = 32'b11111111111111111001011110111100;
assign LUT_4[32874] = 32'b11111111111111111111101101101000;
assign LUT_4[32875] = 32'b11111111111111111000111001100000;
assign LUT_4[32876] = 32'b11111111111111111101010011100000;
assign LUT_4[32877] = 32'b11111111111111110110011111011000;
assign LUT_4[32878] = 32'b11111111111111111100101110000100;
assign LUT_4[32879] = 32'b11111111111111110101111001111100;
assign LUT_4[32880] = 32'b00000000000000000100111000011101;
assign LUT_4[32881] = 32'b11111111111111111110000100010101;
assign LUT_4[32882] = 32'b00000000000000000100010011000001;
assign LUT_4[32883] = 32'b11111111111111111101011110111001;
assign LUT_4[32884] = 32'b00000000000000000001111000111001;
assign LUT_4[32885] = 32'b11111111111111111011000100110001;
assign LUT_4[32886] = 32'b00000000000000000001010011011101;
assign LUT_4[32887] = 32'b11111111111111111010011111010101;
assign LUT_4[32888] = 32'b11111111111111111110000100110010;
assign LUT_4[32889] = 32'b11111111111111110111010000101010;
assign LUT_4[32890] = 32'b11111111111111111101011111010110;
assign LUT_4[32891] = 32'b11111111111111110110101011001110;
assign LUT_4[32892] = 32'b11111111111111111011000101001110;
assign LUT_4[32893] = 32'b11111111111111110100010001000110;
assign LUT_4[32894] = 32'b11111111111111111010011111110010;
assign LUT_4[32895] = 32'b11111111111111110011101011101010;
assign LUT_4[32896] = 32'b00000000000000001001111010011100;
assign LUT_4[32897] = 32'b00000000000000000011000110010100;
assign LUT_4[32898] = 32'b00000000000000001001010101000000;
assign LUT_4[32899] = 32'b00000000000000000010100000111000;
assign LUT_4[32900] = 32'b00000000000000000110111010111000;
assign LUT_4[32901] = 32'b00000000000000000000000110110000;
assign LUT_4[32902] = 32'b00000000000000000110010101011100;
assign LUT_4[32903] = 32'b11111111111111111111100001010100;
assign LUT_4[32904] = 32'b00000000000000000011000110110001;
assign LUT_4[32905] = 32'b11111111111111111100010010101001;
assign LUT_4[32906] = 32'b00000000000000000010100001010101;
assign LUT_4[32907] = 32'b11111111111111111011101101001101;
assign LUT_4[32908] = 32'b00000000000000000000000111001101;
assign LUT_4[32909] = 32'b11111111111111111001010011000101;
assign LUT_4[32910] = 32'b11111111111111111111100001110001;
assign LUT_4[32911] = 32'b11111111111111111000101101101001;
assign LUT_4[32912] = 32'b00000000000000000111101100001010;
assign LUT_4[32913] = 32'b00000000000000000000111000000010;
assign LUT_4[32914] = 32'b00000000000000000111000110101110;
assign LUT_4[32915] = 32'b00000000000000000000010010100110;
assign LUT_4[32916] = 32'b00000000000000000100101100100110;
assign LUT_4[32917] = 32'b11111111111111111101111000011110;
assign LUT_4[32918] = 32'b00000000000000000100000111001010;
assign LUT_4[32919] = 32'b11111111111111111101010011000010;
assign LUT_4[32920] = 32'b00000000000000000000111000011111;
assign LUT_4[32921] = 32'b11111111111111111010000100010111;
assign LUT_4[32922] = 32'b00000000000000000000010011000011;
assign LUT_4[32923] = 32'b11111111111111111001011110111011;
assign LUT_4[32924] = 32'b11111111111111111101111000111011;
assign LUT_4[32925] = 32'b11111111111111110111000100110011;
assign LUT_4[32926] = 32'b11111111111111111101010011011111;
assign LUT_4[32927] = 32'b11111111111111110110011111010111;
assign LUT_4[32928] = 32'b00000000000000001000010101100011;
assign LUT_4[32929] = 32'b00000000000000000001100001011011;
assign LUT_4[32930] = 32'b00000000000000000111110000000111;
assign LUT_4[32931] = 32'b00000000000000000000111011111111;
assign LUT_4[32932] = 32'b00000000000000000101010101111111;
assign LUT_4[32933] = 32'b11111111111111111110100001110111;
assign LUT_4[32934] = 32'b00000000000000000100110000100011;
assign LUT_4[32935] = 32'b11111111111111111101111100011011;
assign LUT_4[32936] = 32'b00000000000000000001100001111000;
assign LUT_4[32937] = 32'b11111111111111111010101101110000;
assign LUT_4[32938] = 32'b00000000000000000000111100011100;
assign LUT_4[32939] = 32'b11111111111111111010001000010100;
assign LUT_4[32940] = 32'b11111111111111111110100010010100;
assign LUT_4[32941] = 32'b11111111111111110111101110001100;
assign LUT_4[32942] = 32'b11111111111111111101111100111000;
assign LUT_4[32943] = 32'b11111111111111110111001000110000;
assign LUT_4[32944] = 32'b00000000000000000110000111010001;
assign LUT_4[32945] = 32'b11111111111111111111010011001001;
assign LUT_4[32946] = 32'b00000000000000000101100001110101;
assign LUT_4[32947] = 32'b11111111111111111110101101101101;
assign LUT_4[32948] = 32'b00000000000000000011000111101101;
assign LUT_4[32949] = 32'b11111111111111111100010011100101;
assign LUT_4[32950] = 32'b00000000000000000010100010010001;
assign LUT_4[32951] = 32'b11111111111111111011101110001001;
assign LUT_4[32952] = 32'b11111111111111111111010011100110;
assign LUT_4[32953] = 32'b11111111111111111000011111011110;
assign LUT_4[32954] = 32'b11111111111111111110101110001010;
assign LUT_4[32955] = 32'b11111111111111110111111010000010;
assign LUT_4[32956] = 32'b11111111111111111100010100000010;
assign LUT_4[32957] = 32'b11111111111111110101011111111010;
assign LUT_4[32958] = 32'b11111111111111111011101110100110;
assign LUT_4[32959] = 32'b11111111111111110100111010011110;
assign LUT_4[32960] = 32'b00000000000000001011010001110000;
assign LUT_4[32961] = 32'b00000000000000000100011101101000;
assign LUT_4[32962] = 32'b00000000000000001010101100010100;
assign LUT_4[32963] = 32'b00000000000000000011111000001100;
assign LUT_4[32964] = 32'b00000000000000001000010010001100;
assign LUT_4[32965] = 32'b00000000000000000001011110000100;
assign LUT_4[32966] = 32'b00000000000000000111101100110000;
assign LUT_4[32967] = 32'b00000000000000000000111000101000;
assign LUT_4[32968] = 32'b00000000000000000100011110000101;
assign LUT_4[32969] = 32'b11111111111111111101101001111101;
assign LUT_4[32970] = 32'b00000000000000000011111000101001;
assign LUT_4[32971] = 32'b11111111111111111101000100100001;
assign LUT_4[32972] = 32'b00000000000000000001011110100001;
assign LUT_4[32973] = 32'b11111111111111111010101010011001;
assign LUT_4[32974] = 32'b00000000000000000000111001000101;
assign LUT_4[32975] = 32'b11111111111111111010000100111101;
assign LUT_4[32976] = 32'b00000000000000001001000011011110;
assign LUT_4[32977] = 32'b00000000000000000010001111010110;
assign LUT_4[32978] = 32'b00000000000000001000011110000010;
assign LUT_4[32979] = 32'b00000000000000000001101001111010;
assign LUT_4[32980] = 32'b00000000000000000110000011111010;
assign LUT_4[32981] = 32'b11111111111111111111001111110010;
assign LUT_4[32982] = 32'b00000000000000000101011110011110;
assign LUT_4[32983] = 32'b11111111111111111110101010010110;
assign LUT_4[32984] = 32'b00000000000000000010001111110011;
assign LUT_4[32985] = 32'b11111111111111111011011011101011;
assign LUT_4[32986] = 32'b00000000000000000001101010010111;
assign LUT_4[32987] = 32'b11111111111111111010110110001111;
assign LUT_4[32988] = 32'b11111111111111111111010000001111;
assign LUT_4[32989] = 32'b11111111111111111000011100000111;
assign LUT_4[32990] = 32'b11111111111111111110101010110011;
assign LUT_4[32991] = 32'b11111111111111110111110110101011;
assign LUT_4[32992] = 32'b00000000000000001001101100110111;
assign LUT_4[32993] = 32'b00000000000000000010111000101111;
assign LUT_4[32994] = 32'b00000000000000001001000111011011;
assign LUT_4[32995] = 32'b00000000000000000010010011010011;
assign LUT_4[32996] = 32'b00000000000000000110101101010011;
assign LUT_4[32997] = 32'b11111111111111111111111001001011;
assign LUT_4[32998] = 32'b00000000000000000110000111110111;
assign LUT_4[32999] = 32'b11111111111111111111010011101111;
assign LUT_4[33000] = 32'b00000000000000000010111001001100;
assign LUT_4[33001] = 32'b11111111111111111100000101000100;
assign LUT_4[33002] = 32'b00000000000000000010010011110000;
assign LUT_4[33003] = 32'b11111111111111111011011111101000;
assign LUT_4[33004] = 32'b11111111111111111111111001101000;
assign LUT_4[33005] = 32'b11111111111111111001000101100000;
assign LUT_4[33006] = 32'b11111111111111111111010100001100;
assign LUT_4[33007] = 32'b11111111111111111000100000000100;
assign LUT_4[33008] = 32'b00000000000000000111011110100101;
assign LUT_4[33009] = 32'b00000000000000000000101010011101;
assign LUT_4[33010] = 32'b00000000000000000110111001001001;
assign LUT_4[33011] = 32'b00000000000000000000000101000001;
assign LUT_4[33012] = 32'b00000000000000000100011111000001;
assign LUT_4[33013] = 32'b11111111111111111101101010111001;
assign LUT_4[33014] = 32'b00000000000000000011111001100101;
assign LUT_4[33015] = 32'b11111111111111111101000101011101;
assign LUT_4[33016] = 32'b00000000000000000000101010111010;
assign LUT_4[33017] = 32'b11111111111111111001110110110010;
assign LUT_4[33018] = 32'b00000000000000000000000101011110;
assign LUT_4[33019] = 32'b11111111111111111001010001010110;
assign LUT_4[33020] = 32'b11111111111111111101101011010110;
assign LUT_4[33021] = 32'b11111111111111110110110111001110;
assign LUT_4[33022] = 32'b11111111111111111101000101111010;
assign LUT_4[33023] = 32'b11111111111111110110010001110010;
assign LUT_4[33024] = 32'b00000000000000001100001111110111;
assign LUT_4[33025] = 32'b00000000000000000101011011101111;
assign LUT_4[33026] = 32'b00000000000000001011101010011011;
assign LUT_4[33027] = 32'b00000000000000000100110110010011;
assign LUT_4[33028] = 32'b00000000000000001001010000010011;
assign LUT_4[33029] = 32'b00000000000000000010011100001011;
assign LUT_4[33030] = 32'b00000000000000001000101010110111;
assign LUT_4[33031] = 32'b00000000000000000001110110101111;
assign LUT_4[33032] = 32'b00000000000000000101011100001100;
assign LUT_4[33033] = 32'b11111111111111111110101000000100;
assign LUT_4[33034] = 32'b00000000000000000100110110110000;
assign LUT_4[33035] = 32'b11111111111111111110000010101000;
assign LUT_4[33036] = 32'b00000000000000000010011100101000;
assign LUT_4[33037] = 32'b11111111111111111011101000100000;
assign LUT_4[33038] = 32'b00000000000000000001110111001100;
assign LUT_4[33039] = 32'b11111111111111111011000011000100;
assign LUT_4[33040] = 32'b00000000000000001010000001100101;
assign LUT_4[33041] = 32'b00000000000000000011001101011101;
assign LUT_4[33042] = 32'b00000000000000001001011100001001;
assign LUT_4[33043] = 32'b00000000000000000010101000000001;
assign LUT_4[33044] = 32'b00000000000000000111000010000001;
assign LUT_4[33045] = 32'b00000000000000000000001101111001;
assign LUT_4[33046] = 32'b00000000000000000110011100100101;
assign LUT_4[33047] = 32'b11111111111111111111101000011101;
assign LUT_4[33048] = 32'b00000000000000000011001101111010;
assign LUT_4[33049] = 32'b11111111111111111100011001110010;
assign LUT_4[33050] = 32'b00000000000000000010101000011110;
assign LUT_4[33051] = 32'b11111111111111111011110100010110;
assign LUT_4[33052] = 32'b00000000000000000000001110010110;
assign LUT_4[33053] = 32'b11111111111111111001011010001110;
assign LUT_4[33054] = 32'b11111111111111111111101000111010;
assign LUT_4[33055] = 32'b11111111111111111000110100110010;
assign LUT_4[33056] = 32'b00000000000000001010101010111110;
assign LUT_4[33057] = 32'b00000000000000000011110110110110;
assign LUT_4[33058] = 32'b00000000000000001010000101100010;
assign LUT_4[33059] = 32'b00000000000000000011010001011010;
assign LUT_4[33060] = 32'b00000000000000000111101011011010;
assign LUT_4[33061] = 32'b00000000000000000000110111010010;
assign LUT_4[33062] = 32'b00000000000000000111000101111110;
assign LUT_4[33063] = 32'b00000000000000000000010001110110;
assign LUT_4[33064] = 32'b00000000000000000011110111010011;
assign LUT_4[33065] = 32'b11111111111111111101000011001011;
assign LUT_4[33066] = 32'b00000000000000000011010001110111;
assign LUT_4[33067] = 32'b11111111111111111100011101101111;
assign LUT_4[33068] = 32'b00000000000000000000110111101111;
assign LUT_4[33069] = 32'b11111111111111111010000011100111;
assign LUT_4[33070] = 32'b00000000000000000000010010010011;
assign LUT_4[33071] = 32'b11111111111111111001011110001011;
assign LUT_4[33072] = 32'b00000000000000001000011100101100;
assign LUT_4[33073] = 32'b00000000000000000001101000100100;
assign LUT_4[33074] = 32'b00000000000000000111110111010000;
assign LUT_4[33075] = 32'b00000000000000000001000011001000;
assign LUT_4[33076] = 32'b00000000000000000101011101001000;
assign LUT_4[33077] = 32'b11111111111111111110101001000000;
assign LUT_4[33078] = 32'b00000000000000000100110111101100;
assign LUT_4[33079] = 32'b11111111111111111110000011100100;
assign LUT_4[33080] = 32'b00000000000000000001101001000001;
assign LUT_4[33081] = 32'b11111111111111111010110100111001;
assign LUT_4[33082] = 32'b00000000000000000001000011100101;
assign LUT_4[33083] = 32'b11111111111111111010001111011101;
assign LUT_4[33084] = 32'b11111111111111111110101001011101;
assign LUT_4[33085] = 32'b11111111111111110111110101010101;
assign LUT_4[33086] = 32'b11111111111111111110000100000001;
assign LUT_4[33087] = 32'b11111111111111110111001111111001;
assign LUT_4[33088] = 32'b00000000000000001101100111001011;
assign LUT_4[33089] = 32'b00000000000000000110110011000011;
assign LUT_4[33090] = 32'b00000000000000001101000001101111;
assign LUT_4[33091] = 32'b00000000000000000110001101100111;
assign LUT_4[33092] = 32'b00000000000000001010100111100111;
assign LUT_4[33093] = 32'b00000000000000000011110011011111;
assign LUT_4[33094] = 32'b00000000000000001010000010001011;
assign LUT_4[33095] = 32'b00000000000000000011001110000011;
assign LUT_4[33096] = 32'b00000000000000000110110011100000;
assign LUT_4[33097] = 32'b11111111111111111111111111011000;
assign LUT_4[33098] = 32'b00000000000000000110001110000100;
assign LUT_4[33099] = 32'b11111111111111111111011001111100;
assign LUT_4[33100] = 32'b00000000000000000011110011111100;
assign LUT_4[33101] = 32'b11111111111111111100111111110100;
assign LUT_4[33102] = 32'b00000000000000000011001110100000;
assign LUT_4[33103] = 32'b11111111111111111100011010011000;
assign LUT_4[33104] = 32'b00000000000000001011011000111001;
assign LUT_4[33105] = 32'b00000000000000000100100100110001;
assign LUT_4[33106] = 32'b00000000000000001010110011011101;
assign LUT_4[33107] = 32'b00000000000000000011111111010101;
assign LUT_4[33108] = 32'b00000000000000001000011001010101;
assign LUT_4[33109] = 32'b00000000000000000001100101001101;
assign LUT_4[33110] = 32'b00000000000000000111110011111001;
assign LUT_4[33111] = 32'b00000000000000000000111111110001;
assign LUT_4[33112] = 32'b00000000000000000100100101001110;
assign LUT_4[33113] = 32'b11111111111111111101110001000110;
assign LUT_4[33114] = 32'b00000000000000000011111111110010;
assign LUT_4[33115] = 32'b11111111111111111101001011101010;
assign LUT_4[33116] = 32'b00000000000000000001100101101010;
assign LUT_4[33117] = 32'b11111111111111111010110001100010;
assign LUT_4[33118] = 32'b00000000000000000001000000001110;
assign LUT_4[33119] = 32'b11111111111111111010001100000110;
assign LUT_4[33120] = 32'b00000000000000001100000010010010;
assign LUT_4[33121] = 32'b00000000000000000101001110001010;
assign LUT_4[33122] = 32'b00000000000000001011011100110110;
assign LUT_4[33123] = 32'b00000000000000000100101000101110;
assign LUT_4[33124] = 32'b00000000000000001001000010101110;
assign LUT_4[33125] = 32'b00000000000000000010001110100110;
assign LUT_4[33126] = 32'b00000000000000001000011101010010;
assign LUT_4[33127] = 32'b00000000000000000001101001001010;
assign LUT_4[33128] = 32'b00000000000000000101001110100111;
assign LUT_4[33129] = 32'b11111111111111111110011010011111;
assign LUT_4[33130] = 32'b00000000000000000100101001001011;
assign LUT_4[33131] = 32'b11111111111111111101110101000011;
assign LUT_4[33132] = 32'b00000000000000000010001111000011;
assign LUT_4[33133] = 32'b11111111111111111011011010111011;
assign LUT_4[33134] = 32'b00000000000000000001101001100111;
assign LUT_4[33135] = 32'b11111111111111111010110101011111;
assign LUT_4[33136] = 32'b00000000000000001001110100000000;
assign LUT_4[33137] = 32'b00000000000000000010111111111000;
assign LUT_4[33138] = 32'b00000000000000001001001110100100;
assign LUT_4[33139] = 32'b00000000000000000010011010011100;
assign LUT_4[33140] = 32'b00000000000000000110110100011100;
assign LUT_4[33141] = 32'b00000000000000000000000000010100;
assign LUT_4[33142] = 32'b00000000000000000110001111000000;
assign LUT_4[33143] = 32'b11111111111111111111011010111000;
assign LUT_4[33144] = 32'b00000000000000000011000000010101;
assign LUT_4[33145] = 32'b11111111111111111100001100001101;
assign LUT_4[33146] = 32'b00000000000000000010011010111001;
assign LUT_4[33147] = 32'b11111111111111111011100110110001;
assign LUT_4[33148] = 32'b00000000000000000000000000110001;
assign LUT_4[33149] = 32'b11111111111111111001001100101001;
assign LUT_4[33150] = 32'b11111111111111111111011011010101;
assign LUT_4[33151] = 32'b11111111111111111000100111001101;
assign LUT_4[33152] = 32'b00000000000000001110110101111111;
assign LUT_4[33153] = 32'b00000000000000001000000001110111;
assign LUT_4[33154] = 32'b00000000000000001110010000100011;
assign LUT_4[33155] = 32'b00000000000000000111011100011011;
assign LUT_4[33156] = 32'b00000000000000001011110110011011;
assign LUT_4[33157] = 32'b00000000000000000101000010010011;
assign LUT_4[33158] = 32'b00000000000000001011010000111111;
assign LUT_4[33159] = 32'b00000000000000000100011100110111;
assign LUT_4[33160] = 32'b00000000000000001000000010010100;
assign LUT_4[33161] = 32'b00000000000000000001001110001100;
assign LUT_4[33162] = 32'b00000000000000000111011100111000;
assign LUT_4[33163] = 32'b00000000000000000000101000110000;
assign LUT_4[33164] = 32'b00000000000000000101000010110000;
assign LUT_4[33165] = 32'b11111111111111111110001110101000;
assign LUT_4[33166] = 32'b00000000000000000100011101010100;
assign LUT_4[33167] = 32'b11111111111111111101101001001100;
assign LUT_4[33168] = 32'b00000000000000001100100111101101;
assign LUT_4[33169] = 32'b00000000000000000101110011100101;
assign LUT_4[33170] = 32'b00000000000000001100000010010001;
assign LUT_4[33171] = 32'b00000000000000000101001110001001;
assign LUT_4[33172] = 32'b00000000000000001001101000001001;
assign LUT_4[33173] = 32'b00000000000000000010110100000001;
assign LUT_4[33174] = 32'b00000000000000001001000010101101;
assign LUT_4[33175] = 32'b00000000000000000010001110100101;
assign LUT_4[33176] = 32'b00000000000000000101110100000010;
assign LUT_4[33177] = 32'b11111111111111111110111111111010;
assign LUT_4[33178] = 32'b00000000000000000101001110100110;
assign LUT_4[33179] = 32'b11111111111111111110011010011110;
assign LUT_4[33180] = 32'b00000000000000000010110100011110;
assign LUT_4[33181] = 32'b11111111111111111100000000010110;
assign LUT_4[33182] = 32'b00000000000000000010001111000010;
assign LUT_4[33183] = 32'b11111111111111111011011010111010;
assign LUT_4[33184] = 32'b00000000000000001101010001000110;
assign LUT_4[33185] = 32'b00000000000000000110011100111110;
assign LUT_4[33186] = 32'b00000000000000001100101011101010;
assign LUT_4[33187] = 32'b00000000000000000101110111100010;
assign LUT_4[33188] = 32'b00000000000000001010010001100010;
assign LUT_4[33189] = 32'b00000000000000000011011101011010;
assign LUT_4[33190] = 32'b00000000000000001001101100000110;
assign LUT_4[33191] = 32'b00000000000000000010110111111110;
assign LUT_4[33192] = 32'b00000000000000000110011101011011;
assign LUT_4[33193] = 32'b11111111111111111111101001010011;
assign LUT_4[33194] = 32'b00000000000000000101110111111111;
assign LUT_4[33195] = 32'b11111111111111111111000011110111;
assign LUT_4[33196] = 32'b00000000000000000011011101110111;
assign LUT_4[33197] = 32'b11111111111111111100101001101111;
assign LUT_4[33198] = 32'b00000000000000000010111000011011;
assign LUT_4[33199] = 32'b11111111111111111100000100010011;
assign LUT_4[33200] = 32'b00000000000000001011000010110100;
assign LUT_4[33201] = 32'b00000000000000000100001110101100;
assign LUT_4[33202] = 32'b00000000000000001010011101011000;
assign LUT_4[33203] = 32'b00000000000000000011101001010000;
assign LUT_4[33204] = 32'b00000000000000001000000011010000;
assign LUT_4[33205] = 32'b00000000000000000001001111001000;
assign LUT_4[33206] = 32'b00000000000000000111011101110100;
assign LUT_4[33207] = 32'b00000000000000000000101001101100;
assign LUT_4[33208] = 32'b00000000000000000100001111001001;
assign LUT_4[33209] = 32'b11111111111111111101011011000001;
assign LUT_4[33210] = 32'b00000000000000000011101001101101;
assign LUT_4[33211] = 32'b11111111111111111100110101100101;
assign LUT_4[33212] = 32'b00000000000000000001001111100101;
assign LUT_4[33213] = 32'b11111111111111111010011011011101;
assign LUT_4[33214] = 32'b00000000000000000000101010001001;
assign LUT_4[33215] = 32'b11111111111111111001110110000001;
assign LUT_4[33216] = 32'b00000000000000010000001101010011;
assign LUT_4[33217] = 32'b00000000000000001001011001001011;
assign LUT_4[33218] = 32'b00000000000000001111100111110111;
assign LUT_4[33219] = 32'b00000000000000001000110011101111;
assign LUT_4[33220] = 32'b00000000000000001101001101101111;
assign LUT_4[33221] = 32'b00000000000000000110011001100111;
assign LUT_4[33222] = 32'b00000000000000001100101000010011;
assign LUT_4[33223] = 32'b00000000000000000101110100001011;
assign LUT_4[33224] = 32'b00000000000000001001011001101000;
assign LUT_4[33225] = 32'b00000000000000000010100101100000;
assign LUT_4[33226] = 32'b00000000000000001000110100001100;
assign LUT_4[33227] = 32'b00000000000000000010000000000100;
assign LUT_4[33228] = 32'b00000000000000000110011010000100;
assign LUT_4[33229] = 32'b11111111111111111111100101111100;
assign LUT_4[33230] = 32'b00000000000000000101110100101000;
assign LUT_4[33231] = 32'b11111111111111111111000000100000;
assign LUT_4[33232] = 32'b00000000000000001101111111000001;
assign LUT_4[33233] = 32'b00000000000000000111001010111001;
assign LUT_4[33234] = 32'b00000000000000001101011001100101;
assign LUT_4[33235] = 32'b00000000000000000110100101011101;
assign LUT_4[33236] = 32'b00000000000000001010111111011101;
assign LUT_4[33237] = 32'b00000000000000000100001011010101;
assign LUT_4[33238] = 32'b00000000000000001010011010000001;
assign LUT_4[33239] = 32'b00000000000000000011100101111001;
assign LUT_4[33240] = 32'b00000000000000000111001011010110;
assign LUT_4[33241] = 32'b00000000000000000000010111001110;
assign LUT_4[33242] = 32'b00000000000000000110100101111010;
assign LUT_4[33243] = 32'b11111111111111111111110001110010;
assign LUT_4[33244] = 32'b00000000000000000100001011110010;
assign LUT_4[33245] = 32'b11111111111111111101010111101010;
assign LUT_4[33246] = 32'b00000000000000000011100110010110;
assign LUT_4[33247] = 32'b11111111111111111100110010001110;
assign LUT_4[33248] = 32'b00000000000000001110101000011010;
assign LUT_4[33249] = 32'b00000000000000000111110100010010;
assign LUT_4[33250] = 32'b00000000000000001110000010111110;
assign LUT_4[33251] = 32'b00000000000000000111001110110110;
assign LUT_4[33252] = 32'b00000000000000001011101000110110;
assign LUT_4[33253] = 32'b00000000000000000100110100101110;
assign LUT_4[33254] = 32'b00000000000000001011000011011010;
assign LUT_4[33255] = 32'b00000000000000000100001111010010;
assign LUT_4[33256] = 32'b00000000000000000111110100101111;
assign LUT_4[33257] = 32'b00000000000000000001000000100111;
assign LUT_4[33258] = 32'b00000000000000000111001111010011;
assign LUT_4[33259] = 32'b00000000000000000000011011001011;
assign LUT_4[33260] = 32'b00000000000000000100110101001011;
assign LUT_4[33261] = 32'b11111111111111111110000001000011;
assign LUT_4[33262] = 32'b00000000000000000100001111101111;
assign LUT_4[33263] = 32'b11111111111111111101011011100111;
assign LUT_4[33264] = 32'b00000000000000001100011010001000;
assign LUT_4[33265] = 32'b00000000000000000101100110000000;
assign LUT_4[33266] = 32'b00000000000000001011110100101100;
assign LUT_4[33267] = 32'b00000000000000000101000000100100;
assign LUT_4[33268] = 32'b00000000000000001001011010100100;
assign LUT_4[33269] = 32'b00000000000000000010100110011100;
assign LUT_4[33270] = 32'b00000000000000001000110101001000;
assign LUT_4[33271] = 32'b00000000000000000010000001000000;
assign LUT_4[33272] = 32'b00000000000000000101100110011101;
assign LUT_4[33273] = 32'b11111111111111111110110010010101;
assign LUT_4[33274] = 32'b00000000000000000101000001000001;
assign LUT_4[33275] = 32'b11111111111111111110001100111001;
assign LUT_4[33276] = 32'b00000000000000000010100110111001;
assign LUT_4[33277] = 32'b11111111111111111011110010110001;
assign LUT_4[33278] = 32'b00000000000000000010000001011101;
assign LUT_4[33279] = 32'b11111111111111111011001101010101;
assign LUT_4[33280] = 32'b00000000000000000110011000011100;
assign LUT_4[33281] = 32'b11111111111111111111100100010100;
assign LUT_4[33282] = 32'b00000000000000000101110011000000;
assign LUT_4[33283] = 32'b11111111111111111110111110111000;
assign LUT_4[33284] = 32'b00000000000000000011011000111000;
assign LUT_4[33285] = 32'b11111111111111111100100100110000;
assign LUT_4[33286] = 32'b00000000000000000010110011011100;
assign LUT_4[33287] = 32'b11111111111111111011111111010100;
assign LUT_4[33288] = 32'b11111111111111111111100100110001;
assign LUT_4[33289] = 32'b11111111111111111000110000101001;
assign LUT_4[33290] = 32'b11111111111111111110111111010101;
assign LUT_4[33291] = 32'b11111111111111111000001011001101;
assign LUT_4[33292] = 32'b11111111111111111100100101001101;
assign LUT_4[33293] = 32'b11111111111111110101110001000101;
assign LUT_4[33294] = 32'b11111111111111111011111111110001;
assign LUT_4[33295] = 32'b11111111111111110101001011101001;
assign LUT_4[33296] = 32'b00000000000000000100001010001010;
assign LUT_4[33297] = 32'b11111111111111111101010110000010;
assign LUT_4[33298] = 32'b00000000000000000011100100101110;
assign LUT_4[33299] = 32'b11111111111111111100110000100110;
assign LUT_4[33300] = 32'b00000000000000000001001010100110;
assign LUT_4[33301] = 32'b11111111111111111010010110011110;
assign LUT_4[33302] = 32'b00000000000000000000100101001010;
assign LUT_4[33303] = 32'b11111111111111111001110001000010;
assign LUT_4[33304] = 32'b11111111111111111101010110011111;
assign LUT_4[33305] = 32'b11111111111111110110100010010111;
assign LUT_4[33306] = 32'b11111111111111111100110001000011;
assign LUT_4[33307] = 32'b11111111111111110101111100111011;
assign LUT_4[33308] = 32'b11111111111111111010010110111011;
assign LUT_4[33309] = 32'b11111111111111110011100010110011;
assign LUT_4[33310] = 32'b11111111111111111001110001011111;
assign LUT_4[33311] = 32'b11111111111111110010111101010111;
assign LUT_4[33312] = 32'b00000000000000000100110011100011;
assign LUT_4[33313] = 32'b11111111111111111101111111011011;
assign LUT_4[33314] = 32'b00000000000000000100001110000111;
assign LUT_4[33315] = 32'b11111111111111111101011001111111;
assign LUT_4[33316] = 32'b00000000000000000001110011111111;
assign LUT_4[33317] = 32'b11111111111111111010111111110111;
assign LUT_4[33318] = 32'b00000000000000000001001110100011;
assign LUT_4[33319] = 32'b11111111111111111010011010011011;
assign LUT_4[33320] = 32'b11111111111111111101111111111000;
assign LUT_4[33321] = 32'b11111111111111110111001011110000;
assign LUT_4[33322] = 32'b11111111111111111101011010011100;
assign LUT_4[33323] = 32'b11111111111111110110100110010100;
assign LUT_4[33324] = 32'b11111111111111111011000000010100;
assign LUT_4[33325] = 32'b11111111111111110100001100001100;
assign LUT_4[33326] = 32'b11111111111111111010011010111000;
assign LUT_4[33327] = 32'b11111111111111110011100110110000;
assign LUT_4[33328] = 32'b00000000000000000010100101010001;
assign LUT_4[33329] = 32'b11111111111111111011110001001001;
assign LUT_4[33330] = 32'b00000000000000000001111111110101;
assign LUT_4[33331] = 32'b11111111111111111011001011101101;
assign LUT_4[33332] = 32'b11111111111111111111100101101101;
assign LUT_4[33333] = 32'b11111111111111111000110001100101;
assign LUT_4[33334] = 32'b11111111111111111111000000010001;
assign LUT_4[33335] = 32'b11111111111111111000001100001001;
assign LUT_4[33336] = 32'b11111111111111111011110001100110;
assign LUT_4[33337] = 32'b11111111111111110100111101011110;
assign LUT_4[33338] = 32'b11111111111111111011001100001010;
assign LUT_4[33339] = 32'b11111111111111110100011000000010;
assign LUT_4[33340] = 32'b11111111111111111000110010000010;
assign LUT_4[33341] = 32'b11111111111111110001111101111010;
assign LUT_4[33342] = 32'b11111111111111111000001100100110;
assign LUT_4[33343] = 32'b11111111111111110001011000011110;
assign LUT_4[33344] = 32'b00000000000000000111101111110000;
assign LUT_4[33345] = 32'b00000000000000000000111011101000;
assign LUT_4[33346] = 32'b00000000000000000111001010010100;
assign LUT_4[33347] = 32'b00000000000000000000010110001100;
assign LUT_4[33348] = 32'b00000000000000000100110000001100;
assign LUT_4[33349] = 32'b11111111111111111101111100000100;
assign LUT_4[33350] = 32'b00000000000000000100001010110000;
assign LUT_4[33351] = 32'b11111111111111111101010110101000;
assign LUT_4[33352] = 32'b00000000000000000000111100000101;
assign LUT_4[33353] = 32'b11111111111111111010000111111101;
assign LUT_4[33354] = 32'b00000000000000000000010110101001;
assign LUT_4[33355] = 32'b11111111111111111001100010100001;
assign LUT_4[33356] = 32'b11111111111111111101111100100001;
assign LUT_4[33357] = 32'b11111111111111110111001000011001;
assign LUT_4[33358] = 32'b11111111111111111101010111000101;
assign LUT_4[33359] = 32'b11111111111111110110100010111101;
assign LUT_4[33360] = 32'b00000000000000000101100001011110;
assign LUT_4[33361] = 32'b11111111111111111110101101010110;
assign LUT_4[33362] = 32'b00000000000000000100111100000010;
assign LUT_4[33363] = 32'b11111111111111111110000111111010;
assign LUT_4[33364] = 32'b00000000000000000010100001111010;
assign LUT_4[33365] = 32'b11111111111111111011101101110010;
assign LUT_4[33366] = 32'b00000000000000000001111100011110;
assign LUT_4[33367] = 32'b11111111111111111011001000010110;
assign LUT_4[33368] = 32'b11111111111111111110101101110011;
assign LUT_4[33369] = 32'b11111111111111110111111001101011;
assign LUT_4[33370] = 32'b11111111111111111110001000010111;
assign LUT_4[33371] = 32'b11111111111111110111010100001111;
assign LUT_4[33372] = 32'b11111111111111111011101110001111;
assign LUT_4[33373] = 32'b11111111111111110100111010000111;
assign LUT_4[33374] = 32'b11111111111111111011001000110011;
assign LUT_4[33375] = 32'b11111111111111110100010100101011;
assign LUT_4[33376] = 32'b00000000000000000110001010110111;
assign LUT_4[33377] = 32'b11111111111111111111010110101111;
assign LUT_4[33378] = 32'b00000000000000000101100101011011;
assign LUT_4[33379] = 32'b11111111111111111110110001010011;
assign LUT_4[33380] = 32'b00000000000000000011001011010011;
assign LUT_4[33381] = 32'b11111111111111111100010111001011;
assign LUT_4[33382] = 32'b00000000000000000010100101110111;
assign LUT_4[33383] = 32'b11111111111111111011110001101111;
assign LUT_4[33384] = 32'b11111111111111111111010111001100;
assign LUT_4[33385] = 32'b11111111111111111000100011000100;
assign LUT_4[33386] = 32'b11111111111111111110110001110000;
assign LUT_4[33387] = 32'b11111111111111110111111101101000;
assign LUT_4[33388] = 32'b11111111111111111100010111101000;
assign LUT_4[33389] = 32'b11111111111111110101100011100000;
assign LUT_4[33390] = 32'b11111111111111111011110010001100;
assign LUT_4[33391] = 32'b11111111111111110100111110000100;
assign LUT_4[33392] = 32'b00000000000000000011111100100101;
assign LUT_4[33393] = 32'b11111111111111111101001000011101;
assign LUT_4[33394] = 32'b00000000000000000011010111001001;
assign LUT_4[33395] = 32'b11111111111111111100100011000001;
assign LUT_4[33396] = 32'b00000000000000000000111101000001;
assign LUT_4[33397] = 32'b11111111111111111010001000111001;
assign LUT_4[33398] = 32'b00000000000000000000010111100101;
assign LUT_4[33399] = 32'b11111111111111111001100011011101;
assign LUT_4[33400] = 32'b11111111111111111101001000111010;
assign LUT_4[33401] = 32'b11111111111111110110010100110010;
assign LUT_4[33402] = 32'b11111111111111111100100011011110;
assign LUT_4[33403] = 32'b11111111111111110101101111010110;
assign LUT_4[33404] = 32'b11111111111111111010001001010110;
assign LUT_4[33405] = 32'b11111111111111110011010101001110;
assign LUT_4[33406] = 32'b11111111111111111001100011111010;
assign LUT_4[33407] = 32'b11111111111111110010101111110010;
assign LUT_4[33408] = 32'b00000000000000001000111110100100;
assign LUT_4[33409] = 32'b00000000000000000010001010011100;
assign LUT_4[33410] = 32'b00000000000000001000011001001000;
assign LUT_4[33411] = 32'b00000000000000000001100101000000;
assign LUT_4[33412] = 32'b00000000000000000101111111000000;
assign LUT_4[33413] = 32'b11111111111111111111001010111000;
assign LUT_4[33414] = 32'b00000000000000000101011001100100;
assign LUT_4[33415] = 32'b11111111111111111110100101011100;
assign LUT_4[33416] = 32'b00000000000000000010001010111001;
assign LUT_4[33417] = 32'b11111111111111111011010110110001;
assign LUT_4[33418] = 32'b00000000000000000001100101011101;
assign LUT_4[33419] = 32'b11111111111111111010110001010101;
assign LUT_4[33420] = 32'b11111111111111111111001011010101;
assign LUT_4[33421] = 32'b11111111111111111000010111001101;
assign LUT_4[33422] = 32'b11111111111111111110100101111001;
assign LUT_4[33423] = 32'b11111111111111110111110001110001;
assign LUT_4[33424] = 32'b00000000000000000110110000010010;
assign LUT_4[33425] = 32'b11111111111111111111111100001010;
assign LUT_4[33426] = 32'b00000000000000000110001010110110;
assign LUT_4[33427] = 32'b11111111111111111111010110101110;
assign LUT_4[33428] = 32'b00000000000000000011110000101110;
assign LUT_4[33429] = 32'b11111111111111111100111100100110;
assign LUT_4[33430] = 32'b00000000000000000011001011010010;
assign LUT_4[33431] = 32'b11111111111111111100010111001010;
assign LUT_4[33432] = 32'b11111111111111111111111100100111;
assign LUT_4[33433] = 32'b11111111111111111001001000011111;
assign LUT_4[33434] = 32'b11111111111111111111010111001011;
assign LUT_4[33435] = 32'b11111111111111111000100011000011;
assign LUT_4[33436] = 32'b11111111111111111100111101000011;
assign LUT_4[33437] = 32'b11111111111111110110001000111011;
assign LUT_4[33438] = 32'b11111111111111111100010111100111;
assign LUT_4[33439] = 32'b11111111111111110101100011011111;
assign LUT_4[33440] = 32'b00000000000000000111011001101011;
assign LUT_4[33441] = 32'b00000000000000000000100101100011;
assign LUT_4[33442] = 32'b00000000000000000110110100001111;
assign LUT_4[33443] = 32'b00000000000000000000000000000111;
assign LUT_4[33444] = 32'b00000000000000000100011010000111;
assign LUT_4[33445] = 32'b11111111111111111101100101111111;
assign LUT_4[33446] = 32'b00000000000000000011110100101011;
assign LUT_4[33447] = 32'b11111111111111111101000000100011;
assign LUT_4[33448] = 32'b00000000000000000000100110000000;
assign LUT_4[33449] = 32'b11111111111111111001110001111000;
assign LUT_4[33450] = 32'b00000000000000000000000000100100;
assign LUT_4[33451] = 32'b11111111111111111001001100011100;
assign LUT_4[33452] = 32'b11111111111111111101100110011100;
assign LUT_4[33453] = 32'b11111111111111110110110010010100;
assign LUT_4[33454] = 32'b11111111111111111101000001000000;
assign LUT_4[33455] = 32'b11111111111111110110001100111000;
assign LUT_4[33456] = 32'b00000000000000000101001011011001;
assign LUT_4[33457] = 32'b11111111111111111110010111010001;
assign LUT_4[33458] = 32'b00000000000000000100100101111101;
assign LUT_4[33459] = 32'b11111111111111111101110001110101;
assign LUT_4[33460] = 32'b00000000000000000010001011110101;
assign LUT_4[33461] = 32'b11111111111111111011010111101101;
assign LUT_4[33462] = 32'b00000000000000000001100110011001;
assign LUT_4[33463] = 32'b11111111111111111010110010010001;
assign LUT_4[33464] = 32'b11111111111111111110010111101110;
assign LUT_4[33465] = 32'b11111111111111110111100011100110;
assign LUT_4[33466] = 32'b11111111111111111101110010010010;
assign LUT_4[33467] = 32'b11111111111111110110111110001010;
assign LUT_4[33468] = 32'b11111111111111111011011000001010;
assign LUT_4[33469] = 32'b11111111111111110100100100000010;
assign LUT_4[33470] = 32'b11111111111111111010110010101110;
assign LUT_4[33471] = 32'b11111111111111110011111110100110;
assign LUT_4[33472] = 32'b00000000000000001010010101111000;
assign LUT_4[33473] = 32'b00000000000000000011100001110000;
assign LUT_4[33474] = 32'b00000000000000001001110000011100;
assign LUT_4[33475] = 32'b00000000000000000010111100010100;
assign LUT_4[33476] = 32'b00000000000000000111010110010100;
assign LUT_4[33477] = 32'b00000000000000000000100010001100;
assign LUT_4[33478] = 32'b00000000000000000110110000111000;
assign LUT_4[33479] = 32'b11111111111111111111111100110000;
assign LUT_4[33480] = 32'b00000000000000000011100010001101;
assign LUT_4[33481] = 32'b11111111111111111100101110000101;
assign LUT_4[33482] = 32'b00000000000000000010111100110001;
assign LUT_4[33483] = 32'b11111111111111111100001000101001;
assign LUT_4[33484] = 32'b00000000000000000000100010101001;
assign LUT_4[33485] = 32'b11111111111111111001101110100001;
assign LUT_4[33486] = 32'b11111111111111111111111101001101;
assign LUT_4[33487] = 32'b11111111111111111001001001000101;
assign LUT_4[33488] = 32'b00000000000000001000000111100110;
assign LUT_4[33489] = 32'b00000000000000000001010011011110;
assign LUT_4[33490] = 32'b00000000000000000111100010001010;
assign LUT_4[33491] = 32'b00000000000000000000101110000010;
assign LUT_4[33492] = 32'b00000000000000000101001000000010;
assign LUT_4[33493] = 32'b11111111111111111110010011111010;
assign LUT_4[33494] = 32'b00000000000000000100100010100110;
assign LUT_4[33495] = 32'b11111111111111111101101110011110;
assign LUT_4[33496] = 32'b00000000000000000001010011111011;
assign LUT_4[33497] = 32'b11111111111111111010011111110011;
assign LUT_4[33498] = 32'b00000000000000000000101110011111;
assign LUT_4[33499] = 32'b11111111111111111001111010010111;
assign LUT_4[33500] = 32'b11111111111111111110010100010111;
assign LUT_4[33501] = 32'b11111111111111110111100000001111;
assign LUT_4[33502] = 32'b11111111111111111101101110111011;
assign LUT_4[33503] = 32'b11111111111111110110111010110011;
assign LUT_4[33504] = 32'b00000000000000001000110000111111;
assign LUT_4[33505] = 32'b00000000000000000001111100110111;
assign LUT_4[33506] = 32'b00000000000000001000001011100011;
assign LUT_4[33507] = 32'b00000000000000000001010111011011;
assign LUT_4[33508] = 32'b00000000000000000101110001011011;
assign LUT_4[33509] = 32'b11111111111111111110111101010011;
assign LUT_4[33510] = 32'b00000000000000000101001011111111;
assign LUT_4[33511] = 32'b11111111111111111110010111110111;
assign LUT_4[33512] = 32'b00000000000000000001111101010100;
assign LUT_4[33513] = 32'b11111111111111111011001001001100;
assign LUT_4[33514] = 32'b00000000000000000001010111111000;
assign LUT_4[33515] = 32'b11111111111111111010100011110000;
assign LUT_4[33516] = 32'b11111111111111111110111101110000;
assign LUT_4[33517] = 32'b11111111111111111000001001101000;
assign LUT_4[33518] = 32'b11111111111111111110011000010100;
assign LUT_4[33519] = 32'b11111111111111110111100100001100;
assign LUT_4[33520] = 32'b00000000000000000110100010101101;
assign LUT_4[33521] = 32'b11111111111111111111101110100101;
assign LUT_4[33522] = 32'b00000000000000000101111101010001;
assign LUT_4[33523] = 32'b11111111111111111111001001001001;
assign LUT_4[33524] = 32'b00000000000000000011100011001001;
assign LUT_4[33525] = 32'b11111111111111111100101111000001;
assign LUT_4[33526] = 32'b00000000000000000010111101101101;
assign LUT_4[33527] = 32'b11111111111111111100001001100101;
assign LUT_4[33528] = 32'b11111111111111111111101111000010;
assign LUT_4[33529] = 32'b11111111111111111000111010111010;
assign LUT_4[33530] = 32'b11111111111111111111001001100110;
assign LUT_4[33531] = 32'b11111111111111111000010101011110;
assign LUT_4[33532] = 32'b11111111111111111100101111011110;
assign LUT_4[33533] = 32'b11111111111111110101111011010110;
assign LUT_4[33534] = 32'b11111111111111111100001010000010;
assign LUT_4[33535] = 32'b11111111111111110101010101111010;
assign LUT_4[33536] = 32'b00000000000000001011010011111111;
assign LUT_4[33537] = 32'b00000000000000000100011111110111;
assign LUT_4[33538] = 32'b00000000000000001010101110100011;
assign LUT_4[33539] = 32'b00000000000000000011111010011011;
assign LUT_4[33540] = 32'b00000000000000001000010100011011;
assign LUT_4[33541] = 32'b00000000000000000001100000010011;
assign LUT_4[33542] = 32'b00000000000000000111101110111111;
assign LUT_4[33543] = 32'b00000000000000000000111010110111;
assign LUT_4[33544] = 32'b00000000000000000100100000010100;
assign LUT_4[33545] = 32'b11111111111111111101101100001100;
assign LUT_4[33546] = 32'b00000000000000000011111010111000;
assign LUT_4[33547] = 32'b11111111111111111101000110110000;
assign LUT_4[33548] = 32'b00000000000000000001100000110000;
assign LUT_4[33549] = 32'b11111111111111111010101100101000;
assign LUT_4[33550] = 32'b00000000000000000000111011010100;
assign LUT_4[33551] = 32'b11111111111111111010000111001100;
assign LUT_4[33552] = 32'b00000000000000001001000101101101;
assign LUT_4[33553] = 32'b00000000000000000010010001100101;
assign LUT_4[33554] = 32'b00000000000000001000100000010001;
assign LUT_4[33555] = 32'b00000000000000000001101100001001;
assign LUT_4[33556] = 32'b00000000000000000110000110001001;
assign LUT_4[33557] = 32'b11111111111111111111010010000001;
assign LUT_4[33558] = 32'b00000000000000000101100000101101;
assign LUT_4[33559] = 32'b11111111111111111110101100100101;
assign LUT_4[33560] = 32'b00000000000000000010010010000010;
assign LUT_4[33561] = 32'b11111111111111111011011101111010;
assign LUT_4[33562] = 32'b00000000000000000001101100100110;
assign LUT_4[33563] = 32'b11111111111111111010111000011110;
assign LUT_4[33564] = 32'b11111111111111111111010010011110;
assign LUT_4[33565] = 32'b11111111111111111000011110010110;
assign LUT_4[33566] = 32'b11111111111111111110101101000010;
assign LUT_4[33567] = 32'b11111111111111110111111000111010;
assign LUT_4[33568] = 32'b00000000000000001001101111000110;
assign LUT_4[33569] = 32'b00000000000000000010111010111110;
assign LUT_4[33570] = 32'b00000000000000001001001001101010;
assign LUT_4[33571] = 32'b00000000000000000010010101100010;
assign LUT_4[33572] = 32'b00000000000000000110101111100010;
assign LUT_4[33573] = 32'b11111111111111111111111011011010;
assign LUT_4[33574] = 32'b00000000000000000110001010000110;
assign LUT_4[33575] = 32'b11111111111111111111010101111110;
assign LUT_4[33576] = 32'b00000000000000000010111011011011;
assign LUT_4[33577] = 32'b11111111111111111100000111010011;
assign LUT_4[33578] = 32'b00000000000000000010010101111111;
assign LUT_4[33579] = 32'b11111111111111111011100001110111;
assign LUT_4[33580] = 32'b11111111111111111111111011110111;
assign LUT_4[33581] = 32'b11111111111111111001000111101111;
assign LUT_4[33582] = 32'b11111111111111111111010110011011;
assign LUT_4[33583] = 32'b11111111111111111000100010010011;
assign LUT_4[33584] = 32'b00000000000000000111100000110100;
assign LUT_4[33585] = 32'b00000000000000000000101100101100;
assign LUT_4[33586] = 32'b00000000000000000110111011011000;
assign LUT_4[33587] = 32'b00000000000000000000000111010000;
assign LUT_4[33588] = 32'b00000000000000000100100001010000;
assign LUT_4[33589] = 32'b11111111111111111101101101001000;
assign LUT_4[33590] = 32'b00000000000000000011111011110100;
assign LUT_4[33591] = 32'b11111111111111111101000111101100;
assign LUT_4[33592] = 32'b00000000000000000000101101001001;
assign LUT_4[33593] = 32'b11111111111111111001111001000001;
assign LUT_4[33594] = 32'b00000000000000000000000111101101;
assign LUT_4[33595] = 32'b11111111111111111001010011100101;
assign LUT_4[33596] = 32'b11111111111111111101101101100101;
assign LUT_4[33597] = 32'b11111111111111110110111001011101;
assign LUT_4[33598] = 32'b11111111111111111101001000001001;
assign LUT_4[33599] = 32'b11111111111111110110010100000001;
assign LUT_4[33600] = 32'b00000000000000001100101011010011;
assign LUT_4[33601] = 32'b00000000000000000101110111001011;
assign LUT_4[33602] = 32'b00000000000000001100000101110111;
assign LUT_4[33603] = 32'b00000000000000000101010001101111;
assign LUT_4[33604] = 32'b00000000000000001001101011101111;
assign LUT_4[33605] = 32'b00000000000000000010110111100111;
assign LUT_4[33606] = 32'b00000000000000001001000110010011;
assign LUT_4[33607] = 32'b00000000000000000010010010001011;
assign LUT_4[33608] = 32'b00000000000000000101110111101000;
assign LUT_4[33609] = 32'b11111111111111111111000011100000;
assign LUT_4[33610] = 32'b00000000000000000101010010001100;
assign LUT_4[33611] = 32'b11111111111111111110011110000100;
assign LUT_4[33612] = 32'b00000000000000000010111000000100;
assign LUT_4[33613] = 32'b11111111111111111100000011111100;
assign LUT_4[33614] = 32'b00000000000000000010010010101000;
assign LUT_4[33615] = 32'b11111111111111111011011110100000;
assign LUT_4[33616] = 32'b00000000000000001010011101000001;
assign LUT_4[33617] = 32'b00000000000000000011101000111001;
assign LUT_4[33618] = 32'b00000000000000001001110111100101;
assign LUT_4[33619] = 32'b00000000000000000011000011011101;
assign LUT_4[33620] = 32'b00000000000000000111011101011101;
assign LUT_4[33621] = 32'b00000000000000000000101001010101;
assign LUT_4[33622] = 32'b00000000000000000110111000000001;
assign LUT_4[33623] = 32'b00000000000000000000000011111001;
assign LUT_4[33624] = 32'b00000000000000000011101001010110;
assign LUT_4[33625] = 32'b11111111111111111100110101001110;
assign LUT_4[33626] = 32'b00000000000000000011000011111010;
assign LUT_4[33627] = 32'b11111111111111111100001111110010;
assign LUT_4[33628] = 32'b00000000000000000000101001110010;
assign LUT_4[33629] = 32'b11111111111111111001110101101010;
assign LUT_4[33630] = 32'b00000000000000000000000100010110;
assign LUT_4[33631] = 32'b11111111111111111001010000001110;
assign LUT_4[33632] = 32'b00000000000000001011000110011010;
assign LUT_4[33633] = 32'b00000000000000000100010010010010;
assign LUT_4[33634] = 32'b00000000000000001010100000111110;
assign LUT_4[33635] = 32'b00000000000000000011101100110110;
assign LUT_4[33636] = 32'b00000000000000001000000110110110;
assign LUT_4[33637] = 32'b00000000000000000001010010101110;
assign LUT_4[33638] = 32'b00000000000000000111100001011010;
assign LUT_4[33639] = 32'b00000000000000000000101101010010;
assign LUT_4[33640] = 32'b00000000000000000100010010101111;
assign LUT_4[33641] = 32'b11111111111111111101011110100111;
assign LUT_4[33642] = 32'b00000000000000000011101101010011;
assign LUT_4[33643] = 32'b11111111111111111100111001001011;
assign LUT_4[33644] = 32'b00000000000000000001010011001011;
assign LUT_4[33645] = 32'b11111111111111111010011111000011;
assign LUT_4[33646] = 32'b00000000000000000000101101101111;
assign LUT_4[33647] = 32'b11111111111111111001111001100111;
assign LUT_4[33648] = 32'b00000000000000001000111000001000;
assign LUT_4[33649] = 32'b00000000000000000010000100000000;
assign LUT_4[33650] = 32'b00000000000000001000010010101100;
assign LUT_4[33651] = 32'b00000000000000000001011110100100;
assign LUT_4[33652] = 32'b00000000000000000101111000100100;
assign LUT_4[33653] = 32'b11111111111111111111000100011100;
assign LUT_4[33654] = 32'b00000000000000000101010011001000;
assign LUT_4[33655] = 32'b11111111111111111110011111000000;
assign LUT_4[33656] = 32'b00000000000000000010000100011101;
assign LUT_4[33657] = 32'b11111111111111111011010000010101;
assign LUT_4[33658] = 32'b00000000000000000001011111000001;
assign LUT_4[33659] = 32'b11111111111111111010101010111001;
assign LUT_4[33660] = 32'b11111111111111111111000100111001;
assign LUT_4[33661] = 32'b11111111111111111000010000110001;
assign LUT_4[33662] = 32'b11111111111111111110011111011101;
assign LUT_4[33663] = 32'b11111111111111110111101011010101;
assign LUT_4[33664] = 32'b00000000000000001101111010000111;
assign LUT_4[33665] = 32'b00000000000000000111000101111111;
assign LUT_4[33666] = 32'b00000000000000001101010100101011;
assign LUT_4[33667] = 32'b00000000000000000110100000100011;
assign LUT_4[33668] = 32'b00000000000000001010111010100011;
assign LUT_4[33669] = 32'b00000000000000000100000110011011;
assign LUT_4[33670] = 32'b00000000000000001010010101000111;
assign LUT_4[33671] = 32'b00000000000000000011100000111111;
assign LUT_4[33672] = 32'b00000000000000000111000110011100;
assign LUT_4[33673] = 32'b00000000000000000000010010010100;
assign LUT_4[33674] = 32'b00000000000000000110100001000000;
assign LUT_4[33675] = 32'b11111111111111111111101100111000;
assign LUT_4[33676] = 32'b00000000000000000100000110111000;
assign LUT_4[33677] = 32'b11111111111111111101010010110000;
assign LUT_4[33678] = 32'b00000000000000000011100001011100;
assign LUT_4[33679] = 32'b11111111111111111100101101010100;
assign LUT_4[33680] = 32'b00000000000000001011101011110101;
assign LUT_4[33681] = 32'b00000000000000000100110111101101;
assign LUT_4[33682] = 32'b00000000000000001011000110011001;
assign LUT_4[33683] = 32'b00000000000000000100010010010001;
assign LUT_4[33684] = 32'b00000000000000001000101100010001;
assign LUT_4[33685] = 32'b00000000000000000001111000001001;
assign LUT_4[33686] = 32'b00000000000000001000000110110101;
assign LUT_4[33687] = 32'b00000000000000000001010010101101;
assign LUT_4[33688] = 32'b00000000000000000100111000001010;
assign LUT_4[33689] = 32'b11111111111111111110000100000010;
assign LUT_4[33690] = 32'b00000000000000000100010010101110;
assign LUT_4[33691] = 32'b11111111111111111101011110100110;
assign LUT_4[33692] = 32'b00000000000000000001111000100110;
assign LUT_4[33693] = 32'b11111111111111111011000100011110;
assign LUT_4[33694] = 32'b00000000000000000001010011001010;
assign LUT_4[33695] = 32'b11111111111111111010011111000010;
assign LUT_4[33696] = 32'b00000000000000001100010101001110;
assign LUT_4[33697] = 32'b00000000000000000101100001000110;
assign LUT_4[33698] = 32'b00000000000000001011101111110010;
assign LUT_4[33699] = 32'b00000000000000000100111011101010;
assign LUT_4[33700] = 32'b00000000000000001001010101101010;
assign LUT_4[33701] = 32'b00000000000000000010100001100010;
assign LUT_4[33702] = 32'b00000000000000001000110000001110;
assign LUT_4[33703] = 32'b00000000000000000001111100000110;
assign LUT_4[33704] = 32'b00000000000000000101100001100011;
assign LUT_4[33705] = 32'b11111111111111111110101101011011;
assign LUT_4[33706] = 32'b00000000000000000100111100000111;
assign LUT_4[33707] = 32'b11111111111111111110000111111111;
assign LUT_4[33708] = 32'b00000000000000000010100001111111;
assign LUT_4[33709] = 32'b11111111111111111011101101110111;
assign LUT_4[33710] = 32'b00000000000000000001111100100011;
assign LUT_4[33711] = 32'b11111111111111111011001000011011;
assign LUT_4[33712] = 32'b00000000000000001010000110111100;
assign LUT_4[33713] = 32'b00000000000000000011010010110100;
assign LUT_4[33714] = 32'b00000000000000001001100001100000;
assign LUT_4[33715] = 32'b00000000000000000010101101011000;
assign LUT_4[33716] = 32'b00000000000000000111000111011000;
assign LUT_4[33717] = 32'b00000000000000000000010011010000;
assign LUT_4[33718] = 32'b00000000000000000110100001111100;
assign LUT_4[33719] = 32'b11111111111111111111101101110100;
assign LUT_4[33720] = 32'b00000000000000000011010011010001;
assign LUT_4[33721] = 32'b11111111111111111100011111001001;
assign LUT_4[33722] = 32'b00000000000000000010101101110101;
assign LUT_4[33723] = 32'b11111111111111111011111001101101;
assign LUT_4[33724] = 32'b00000000000000000000010011101101;
assign LUT_4[33725] = 32'b11111111111111111001011111100101;
assign LUT_4[33726] = 32'b11111111111111111111101110010001;
assign LUT_4[33727] = 32'b11111111111111111000111010001001;
assign LUT_4[33728] = 32'b00000000000000001111010001011011;
assign LUT_4[33729] = 32'b00000000000000001000011101010011;
assign LUT_4[33730] = 32'b00000000000000001110101011111111;
assign LUT_4[33731] = 32'b00000000000000000111110111110111;
assign LUT_4[33732] = 32'b00000000000000001100010001110111;
assign LUT_4[33733] = 32'b00000000000000000101011101101111;
assign LUT_4[33734] = 32'b00000000000000001011101100011011;
assign LUT_4[33735] = 32'b00000000000000000100111000010011;
assign LUT_4[33736] = 32'b00000000000000001000011101110000;
assign LUT_4[33737] = 32'b00000000000000000001101001101000;
assign LUT_4[33738] = 32'b00000000000000000111111000010100;
assign LUT_4[33739] = 32'b00000000000000000001000100001100;
assign LUT_4[33740] = 32'b00000000000000000101011110001100;
assign LUT_4[33741] = 32'b11111111111111111110101010000100;
assign LUT_4[33742] = 32'b00000000000000000100111000110000;
assign LUT_4[33743] = 32'b11111111111111111110000100101000;
assign LUT_4[33744] = 32'b00000000000000001101000011001001;
assign LUT_4[33745] = 32'b00000000000000000110001111000001;
assign LUT_4[33746] = 32'b00000000000000001100011101101101;
assign LUT_4[33747] = 32'b00000000000000000101101001100101;
assign LUT_4[33748] = 32'b00000000000000001010000011100101;
assign LUT_4[33749] = 32'b00000000000000000011001111011101;
assign LUT_4[33750] = 32'b00000000000000001001011110001001;
assign LUT_4[33751] = 32'b00000000000000000010101010000001;
assign LUT_4[33752] = 32'b00000000000000000110001111011110;
assign LUT_4[33753] = 32'b11111111111111111111011011010110;
assign LUT_4[33754] = 32'b00000000000000000101101010000010;
assign LUT_4[33755] = 32'b11111111111111111110110101111010;
assign LUT_4[33756] = 32'b00000000000000000011001111111010;
assign LUT_4[33757] = 32'b11111111111111111100011011110010;
assign LUT_4[33758] = 32'b00000000000000000010101010011110;
assign LUT_4[33759] = 32'b11111111111111111011110110010110;
assign LUT_4[33760] = 32'b00000000000000001101101100100010;
assign LUT_4[33761] = 32'b00000000000000000110111000011010;
assign LUT_4[33762] = 32'b00000000000000001101000111000110;
assign LUT_4[33763] = 32'b00000000000000000110010010111110;
assign LUT_4[33764] = 32'b00000000000000001010101100111110;
assign LUT_4[33765] = 32'b00000000000000000011111000110110;
assign LUT_4[33766] = 32'b00000000000000001010000111100010;
assign LUT_4[33767] = 32'b00000000000000000011010011011010;
assign LUT_4[33768] = 32'b00000000000000000110111000110111;
assign LUT_4[33769] = 32'b00000000000000000000000100101111;
assign LUT_4[33770] = 32'b00000000000000000110010011011011;
assign LUT_4[33771] = 32'b11111111111111111111011111010011;
assign LUT_4[33772] = 32'b00000000000000000011111001010011;
assign LUT_4[33773] = 32'b11111111111111111101000101001011;
assign LUT_4[33774] = 32'b00000000000000000011010011110111;
assign LUT_4[33775] = 32'b11111111111111111100011111101111;
assign LUT_4[33776] = 32'b00000000000000001011011110010000;
assign LUT_4[33777] = 32'b00000000000000000100101010001000;
assign LUT_4[33778] = 32'b00000000000000001010111000110100;
assign LUT_4[33779] = 32'b00000000000000000100000100101100;
assign LUT_4[33780] = 32'b00000000000000001000011110101100;
assign LUT_4[33781] = 32'b00000000000000000001101010100100;
assign LUT_4[33782] = 32'b00000000000000000111111001010000;
assign LUT_4[33783] = 32'b00000000000000000001000101001000;
assign LUT_4[33784] = 32'b00000000000000000100101010100101;
assign LUT_4[33785] = 32'b11111111111111111101110110011101;
assign LUT_4[33786] = 32'b00000000000000000100000101001001;
assign LUT_4[33787] = 32'b11111111111111111101010001000001;
assign LUT_4[33788] = 32'b00000000000000000001101011000001;
assign LUT_4[33789] = 32'b11111111111111111010110110111001;
assign LUT_4[33790] = 32'b00000000000000000001000101100101;
assign LUT_4[33791] = 32'b11111111111111111010010001011101;
assign LUT_4[33792] = 32'b00000000000000001000111110110011;
assign LUT_4[33793] = 32'b00000000000000000010001010101011;
assign LUT_4[33794] = 32'b00000000000000001000011001010111;
assign LUT_4[33795] = 32'b00000000000000000001100101001111;
assign LUT_4[33796] = 32'b00000000000000000101111111001111;
assign LUT_4[33797] = 32'b11111111111111111111001011000111;
assign LUT_4[33798] = 32'b00000000000000000101011001110011;
assign LUT_4[33799] = 32'b11111111111111111110100101101011;
assign LUT_4[33800] = 32'b00000000000000000010001011001000;
assign LUT_4[33801] = 32'b11111111111111111011010111000000;
assign LUT_4[33802] = 32'b00000000000000000001100101101100;
assign LUT_4[33803] = 32'b11111111111111111010110001100100;
assign LUT_4[33804] = 32'b11111111111111111111001011100100;
assign LUT_4[33805] = 32'b11111111111111111000010111011100;
assign LUT_4[33806] = 32'b11111111111111111110100110001000;
assign LUT_4[33807] = 32'b11111111111111110111110010000000;
assign LUT_4[33808] = 32'b00000000000000000110110000100001;
assign LUT_4[33809] = 32'b11111111111111111111111100011001;
assign LUT_4[33810] = 32'b00000000000000000110001011000101;
assign LUT_4[33811] = 32'b11111111111111111111010110111101;
assign LUT_4[33812] = 32'b00000000000000000011110000111101;
assign LUT_4[33813] = 32'b11111111111111111100111100110101;
assign LUT_4[33814] = 32'b00000000000000000011001011100001;
assign LUT_4[33815] = 32'b11111111111111111100010111011001;
assign LUT_4[33816] = 32'b11111111111111111111111100110110;
assign LUT_4[33817] = 32'b11111111111111111001001000101110;
assign LUT_4[33818] = 32'b11111111111111111111010111011010;
assign LUT_4[33819] = 32'b11111111111111111000100011010010;
assign LUT_4[33820] = 32'b11111111111111111100111101010010;
assign LUT_4[33821] = 32'b11111111111111110110001001001010;
assign LUT_4[33822] = 32'b11111111111111111100010111110110;
assign LUT_4[33823] = 32'b11111111111111110101100011101110;
assign LUT_4[33824] = 32'b00000000000000000111011001111010;
assign LUT_4[33825] = 32'b00000000000000000000100101110010;
assign LUT_4[33826] = 32'b00000000000000000110110100011110;
assign LUT_4[33827] = 32'b00000000000000000000000000010110;
assign LUT_4[33828] = 32'b00000000000000000100011010010110;
assign LUT_4[33829] = 32'b11111111111111111101100110001110;
assign LUT_4[33830] = 32'b00000000000000000011110100111010;
assign LUT_4[33831] = 32'b11111111111111111101000000110010;
assign LUT_4[33832] = 32'b00000000000000000000100110001111;
assign LUT_4[33833] = 32'b11111111111111111001110010000111;
assign LUT_4[33834] = 32'b00000000000000000000000000110011;
assign LUT_4[33835] = 32'b11111111111111111001001100101011;
assign LUT_4[33836] = 32'b11111111111111111101100110101011;
assign LUT_4[33837] = 32'b11111111111111110110110010100011;
assign LUT_4[33838] = 32'b11111111111111111101000001001111;
assign LUT_4[33839] = 32'b11111111111111110110001101000111;
assign LUT_4[33840] = 32'b00000000000000000101001011101000;
assign LUT_4[33841] = 32'b11111111111111111110010111100000;
assign LUT_4[33842] = 32'b00000000000000000100100110001100;
assign LUT_4[33843] = 32'b11111111111111111101110010000100;
assign LUT_4[33844] = 32'b00000000000000000010001100000100;
assign LUT_4[33845] = 32'b11111111111111111011010111111100;
assign LUT_4[33846] = 32'b00000000000000000001100110101000;
assign LUT_4[33847] = 32'b11111111111111111010110010100000;
assign LUT_4[33848] = 32'b11111111111111111110010111111101;
assign LUT_4[33849] = 32'b11111111111111110111100011110101;
assign LUT_4[33850] = 32'b11111111111111111101110010100001;
assign LUT_4[33851] = 32'b11111111111111110110111110011001;
assign LUT_4[33852] = 32'b11111111111111111011011000011001;
assign LUT_4[33853] = 32'b11111111111111110100100100010001;
assign LUT_4[33854] = 32'b11111111111111111010110010111101;
assign LUT_4[33855] = 32'b11111111111111110011111110110101;
assign LUT_4[33856] = 32'b00000000000000001010010110000111;
assign LUT_4[33857] = 32'b00000000000000000011100001111111;
assign LUT_4[33858] = 32'b00000000000000001001110000101011;
assign LUT_4[33859] = 32'b00000000000000000010111100100011;
assign LUT_4[33860] = 32'b00000000000000000111010110100011;
assign LUT_4[33861] = 32'b00000000000000000000100010011011;
assign LUT_4[33862] = 32'b00000000000000000110110001000111;
assign LUT_4[33863] = 32'b11111111111111111111111100111111;
assign LUT_4[33864] = 32'b00000000000000000011100010011100;
assign LUT_4[33865] = 32'b11111111111111111100101110010100;
assign LUT_4[33866] = 32'b00000000000000000010111101000000;
assign LUT_4[33867] = 32'b11111111111111111100001000111000;
assign LUT_4[33868] = 32'b00000000000000000000100010111000;
assign LUT_4[33869] = 32'b11111111111111111001101110110000;
assign LUT_4[33870] = 32'b11111111111111111111111101011100;
assign LUT_4[33871] = 32'b11111111111111111001001001010100;
assign LUT_4[33872] = 32'b00000000000000001000000111110101;
assign LUT_4[33873] = 32'b00000000000000000001010011101101;
assign LUT_4[33874] = 32'b00000000000000000111100010011001;
assign LUT_4[33875] = 32'b00000000000000000000101110010001;
assign LUT_4[33876] = 32'b00000000000000000101001000010001;
assign LUT_4[33877] = 32'b11111111111111111110010100001001;
assign LUT_4[33878] = 32'b00000000000000000100100010110101;
assign LUT_4[33879] = 32'b11111111111111111101101110101101;
assign LUT_4[33880] = 32'b00000000000000000001010100001010;
assign LUT_4[33881] = 32'b11111111111111111010100000000010;
assign LUT_4[33882] = 32'b00000000000000000000101110101110;
assign LUT_4[33883] = 32'b11111111111111111001111010100110;
assign LUT_4[33884] = 32'b11111111111111111110010100100110;
assign LUT_4[33885] = 32'b11111111111111110111100000011110;
assign LUT_4[33886] = 32'b11111111111111111101101111001010;
assign LUT_4[33887] = 32'b11111111111111110110111011000010;
assign LUT_4[33888] = 32'b00000000000000001000110001001110;
assign LUT_4[33889] = 32'b00000000000000000001111101000110;
assign LUT_4[33890] = 32'b00000000000000001000001011110010;
assign LUT_4[33891] = 32'b00000000000000000001010111101010;
assign LUT_4[33892] = 32'b00000000000000000101110001101010;
assign LUT_4[33893] = 32'b11111111111111111110111101100010;
assign LUT_4[33894] = 32'b00000000000000000101001100001110;
assign LUT_4[33895] = 32'b11111111111111111110011000000110;
assign LUT_4[33896] = 32'b00000000000000000001111101100011;
assign LUT_4[33897] = 32'b11111111111111111011001001011011;
assign LUT_4[33898] = 32'b00000000000000000001011000000111;
assign LUT_4[33899] = 32'b11111111111111111010100011111111;
assign LUT_4[33900] = 32'b11111111111111111110111101111111;
assign LUT_4[33901] = 32'b11111111111111111000001001110111;
assign LUT_4[33902] = 32'b11111111111111111110011000100011;
assign LUT_4[33903] = 32'b11111111111111110111100100011011;
assign LUT_4[33904] = 32'b00000000000000000110100010111100;
assign LUT_4[33905] = 32'b11111111111111111111101110110100;
assign LUT_4[33906] = 32'b00000000000000000101111101100000;
assign LUT_4[33907] = 32'b11111111111111111111001001011000;
assign LUT_4[33908] = 32'b00000000000000000011100011011000;
assign LUT_4[33909] = 32'b11111111111111111100101111010000;
assign LUT_4[33910] = 32'b00000000000000000010111101111100;
assign LUT_4[33911] = 32'b11111111111111111100001001110100;
assign LUT_4[33912] = 32'b11111111111111111111101111010001;
assign LUT_4[33913] = 32'b11111111111111111000111011001001;
assign LUT_4[33914] = 32'b11111111111111111111001001110101;
assign LUT_4[33915] = 32'b11111111111111111000010101101101;
assign LUT_4[33916] = 32'b11111111111111111100101111101101;
assign LUT_4[33917] = 32'b11111111111111110101111011100101;
assign LUT_4[33918] = 32'b11111111111111111100001010010001;
assign LUT_4[33919] = 32'b11111111111111110101010110001001;
assign LUT_4[33920] = 32'b00000000000000001011100100111011;
assign LUT_4[33921] = 32'b00000000000000000100110000110011;
assign LUT_4[33922] = 32'b00000000000000001010111111011111;
assign LUT_4[33923] = 32'b00000000000000000100001011010111;
assign LUT_4[33924] = 32'b00000000000000001000100101010111;
assign LUT_4[33925] = 32'b00000000000000000001110001001111;
assign LUT_4[33926] = 32'b00000000000000000111111111111011;
assign LUT_4[33927] = 32'b00000000000000000001001011110011;
assign LUT_4[33928] = 32'b00000000000000000100110001010000;
assign LUT_4[33929] = 32'b11111111111111111101111101001000;
assign LUT_4[33930] = 32'b00000000000000000100001011110100;
assign LUT_4[33931] = 32'b11111111111111111101010111101100;
assign LUT_4[33932] = 32'b00000000000000000001110001101100;
assign LUT_4[33933] = 32'b11111111111111111010111101100100;
assign LUT_4[33934] = 32'b00000000000000000001001100010000;
assign LUT_4[33935] = 32'b11111111111111111010011000001000;
assign LUT_4[33936] = 32'b00000000000000001001010110101001;
assign LUT_4[33937] = 32'b00000000000000000010100010100001;
assign LUT_4[33938] = 32'b00000000000000001000110001001101;
assign LUT_4[33939] = 32'b00000000000000000001111101000101;
assign LUT_4[33940] = 32'b00000000000000000110010111000101;
assign LUT_4[33941] = 32'b11111111111111111111100010111101;
assign LUT_4[33942] = 32'b00000000000000000101110001101001;
assign LUT_4[33943] = 32'b11111111111111111110111101100001;
assign LUT_4[33944] = 32'b00000000000000000010100010111110;
assign LUT_4[33945] = 32'b11111111111111111011101110110110;
assign LUT_4[33946] = 32'b00000000000000000001111101100010;
assign LUT_4[33947] = 32'b11111111111111111011001001011010;
assign LUT_4[33948] = 32'b11111111111111111111100011011010;
assign LUT_4[33949] = 32'b11111111111111111000101111010010;
assign LUT_4[33950] = 32'b11111111111111111110111101111110;
assign LUT_4[33951] = 32'b11111111111111111000001001110110;
assign LUT_4[33952] = 32'b00000000000000001010000000000010;
assign LUT_4[33953] = 32'b00000000000000000011001011111010;
assign LUT_4[33954] = 32'b00000000000000001001011010100110;
assign LUT_4[33955] = 32'b00000000000000000010100110011110;
assign LUT_4[33956] = 32'b00000000000000000111000000011110;
assign LUT_4[33957] = 32'b00000000000000000000001100010110;
assign LUT_4[33958] = 32'b00000000000000000110011011000010;
assign LUT_4[33959] = 32'b11111111111111111111100110111010;
assign LUT_4[33960] = 32'b00000000000000000011001100010111;
assign LUT_4[33961] = 32'b11111111111111111100011000001111;
assign LUT_4[33962] = 32'b00000000000000000010100110111011;
assign LUT_4[33963] = 32'b11111111111111111011110010110011;
assign LUT_4[33964] = 32'b00000000000000000000001100110011;
assign LUT_4[33965] = 32'b11111111111111111001011000101011;
assign LUT_4[33966] = 32'b11111111111111111111100111010111;
assign LUT_4[33967] = 32'b11111111111111111000110011001111;
assign LUT_4[33968] = 32'b00000000000000000111110001110000;
assign LUT_4[33969] = 32'b00000000000000000000111101101000;
assign LUT_4[33970] = 32'b00000000000000000111001100010100;
assign LUT_4[33971] = 32'b00000000000000000000011000001100;
assign LUT_4[33972] = 32'b00000000000000000100110010001100;
assign LUT_4[33973] = 32'b11111111111111111101111110000100;
assign LUT_4[33974] = 32'b00000000000000000100001100110000;
assign LUT_4[33975] = 32'b11111111111111111101011000101000;
assign LUT_4[33976] = 32'b00000000000000000000111110000101;
assign LUT_4[33977] = 32'b11111111111111111010001001111101;
assign LUT_4[33978] = 32'b00000000000000000000011000101001;
assign LUT_4[33979] = 32'b11111111111111111001100100100001;
assign LUT_4[33980] = 32'b11111111111111111101111110100001;
assign LUT_4[33981] = 32'b11111111111111110111001010011001;
assign LUT_4[33982] = 32'b11111111111111111101011001000101;
assign LUT_4[33983] = 32'b11111111111111110110100100111101;
assign LUT_4[33984] = 32'b00000000000000001100111100001111;
assign LUT_4[33985] = 32'b00000000000000000110001000000111;
assign LUT_4[33986] = 32'b00000000000000001100010110110011;
assign LUT_4[33987] = 32'b00000000000000000101100010101011;
assign LUT_4[33988] = 32'b00000000000000001001111100101011;
assign LUT_4[33989] = 32'b00000000000000000011001000100011;
assign LUT_4[33990] = 32'b00000000000000001001010111001111;
assign LUT_4[33991] = 32'b00000000000000000010100011000111;
assign LUT_4[33992] = 32'b00000000000000000110001000100100;
assign LUT_4[33993] = 32'b11111111111111111111010100011100;
assign LUT_4[33994] = 32'b00000000000000000101100011001000;
assign LUT_4[33995] = 32'b11111111111111111110101111000000;
assign LUT_4[33996] = 32'b00000000000000000011001001000000;
assign LUT_4[33997] = 32'b11111111111111111100010100111000;
assign LUT_4[33998] = 32'b00000000000000000010100011100100;
assign LUT_4[33999] = 32'b11111111111111111011101111011100;
assign LUT_4[34000] = 32'b00000000000000001010101101111101;
assign LUT_4[34001] = 32'b00000000000000000011111001110101;
assign LUT_4[34002] = 32'b00000000000000001010001000100001;
assign LUT_4[34003] = 32'b00000000000000000011010100011001;
assign LUT_4[34004] = 32'b00000000000000000111101110011001;
assign LUT_4[34005] = 32'b00000000000000000000111010010001;
assign LUT_4[34006] = 32'b00000000000000000111001000111101;
assign LUT_4[34007] = 32'b00000000000000000000010100110101;
assign LUT_4[34008] = 32'b00000000000000000011111010010010;
assign LUT_4[34009] = 32'b11111111111111111101000110001010;
assign LUT_4[34010] = 32'b00000000000000000011010100110110;
assign LUT_4[34011] = 32'b11111111111111111100100000101110;
assign LUT_4[34012] = 32'b00000000000000000000111010101110;
assign LUT_4[34013] = 32'b11111111111111111010000110100110;
assign LUT_4[34014] = 32'b00000000000000000000010101010010;
assign LUT_4[34015] = 32'b11111111111111111001100001001010;
assign LUT_4[34016] = 32'b00000000000000001011010111010110;
assign LUT_4[34017] = 32'b00000000000000000100100011001110;
assign LUT_4[34018] = 32'b00000000000000001010110001111010;
assign LUT_4[34019] = 32'b00000000000000000011111101110010;
assign LUT_4[34020] = 32'b00000000000000001000010111110010;
assign LUT_4[34021] = 32'b00000000000000000001100011101010;
assign LUT_4[34022] = 32'b00000000000000000111110010010110;
assign LUT_4[34023] = 32'b00000000000000000000111110001110;
assign LUT_4[34024] = 32'b00000000000000000100100011101011;
assign LUT_4[34025] = 32'b11111111111111111101101111100011;
assign LUT_4[34026] = 32'b00000000000000000011111110001111;
assign LUT_4[34027] = 32'b11111111111111111101001010000111;
assign LUT_4[34028] = 32'b00000000000000000001100100000111;
assign LUT_4[34029] = 32'b11111111111111111010101111111111;
assign LUT_4[34030] = 32'b00000000000000000000111110101011;
assign LUT_4[34031] = 32'b11111111111111111010001010100011;
assign LUT_4[34032] = 32'b00000000000000001001001001000100;
assign LUT_4[34033] = 32'b00000000000000000010010100111100;
assign LUT_4[34034] = 32'b00000000000000001000100011101000;
assign LUT_4[34035] = 32'b00000000000000000001101111100000;
assign LUT_4[34036] = 32'b00000000000000000110001001100000;
assign LUT_4[34037] = 32'b11111111111111111111010101011000;
assign LUT_4[34038] = 32'b00000000000000000101100100000100;
assign LUT_4[34039] = 32'b11111111111111111110101111111100;
assign LUT_4[34040] = 32'b00000000000000000010010101011001;
assign LUT_4[34041] = 32'b11111111111111111011100001010001;
assign LUT_4[34042] = 32'b00000000000000000001101111111101;
assign LUT_4[34043] = 32'b11111111111111111010111011110101;
assign LUT_4[34044] = 32'b11111111111111111111010101110101;
assign LUT_4[34045] = 32'b11111111111111111000100001101101;
assign LUT_4[34046] = 32'b11111111111111111110110000011001;
assign LUT_4[34047] = 32'b11111111111111110111111100010001;
assign LUT_4[34048] = 32'b00000000000000001101111010010110;
assign LUT_4[34049] = 32'b00000000000000000111000110001110;
assign LUT_4[34050] = 32'b00000000000000001101010100111010;
assign LUT_4[34051] = 32'b00000000000000000110100000110010;
assign LUT_4[34052] = 32'b00000000000000001010111010110010;
assign LUT_4[34053] = 32'b00000000000000000100000110101010;
assign LUT_4[34054] = 32'b00000000000000001010010101010110;
assign LUT_4[34055] = 32'b00000000000000000011100001001110;
assign LUT_4[34056] = 32'b00000000000000000111000110101011;
assign LUT_4[34057] = 32'b00000000000000000000010010100011;
assign LUT_4[34058] = 32'b00000000000000000110100001001111;
assign LUT_4[34059] = 32'b11111111111111111111101101000111;
assign LUT_4[34060] = 32'b00000000000000000100000111000111;
assign LUT_4[34061] = 32'b11111111111111111101010010111111;
assign LUT_4[34062] = 32'b00000000000000000011100001101011;
assign LUT_4[34063] = 32'b11111111111111111100101101100011;
assign LUT_4[34064] = 32'b00000000000000001011101100000100;
assign LUT_4[34065] = 32'b00000000000000000100110111111100;
assign LUT_4[34066] = 32'b00000000000000001011000110101000;
assign LUT_4[34067] = 32'b00000000000000000100010010100000;
assign LUT_4[34068] = 32'b00000000000000001000101100100000;
assign LUT_4[34069] = 32'b00000000000000000001111000011000;
assign LUT_4[34070] = 32'b00000000000000001000000111000100;
assign LUT_4[34071] = 32'b00000000000000000001010010111100;
assign LUT_4[34072] = 32'b00000000000000000100111000011001;
assign LUT_4[34073] = 32'b11111111111111111110000100010001;
assign LUT_4[34074] = 32'b00000000000000000100010010111101;
assign LUT_4[34075] = 32'b11111111111111111101011110110101;
assign LUT_4[34076] = 32'b00000000000000000001111000110101;
assign LUT_4[34077] = 32'b11111111111111111011000100101101;
assign LUT_4[34078] = 32'b00000000000000000001010011011001;
assign LUT_4[34079] = 32'b11111111111111111010011111010001;
assign LUT_4[34080] = 32'b00000000000000001100010101011101;
assign LUT_4[34081] = 32'b00000000000000000101100001010101;
assign LUT_4[34082] = 32'b00000000000000001011110000000001;
assign LUT_4[34083] = 32'b00000000000000000100111011111001;
assign LUT_4[34084] = 32'b00000000000000001001010101111001;
assign LUT_4[34085] = 32'b00000000000000000010100001110001;
assign LUT_4[34086] = 32'b00000000000000001000110000011101;
assign LUT_4[34087] = 32'b00000000000000000001111100010101;
assign LUT_4[34088] = 32'b00000000000000000101100001110010;
assign LUT_4[34089] = 32'b11111111111111111110101101101010;
assign LUT_4[34090] = 32'b00000000000000000100111100010110;
assign LUT_4[34091] = 32'b11111111111111111110001000001110;
assign LUT_4[34092] = 32'b00000000000000000010100010001110;
assign LUT_4[34093] = 32'b11111111111111111011101110000110;
assign LUT_4[34094] = 32'b00000000000000000001111100110010;
assign LUT_4[34095] = 32'b11111111111111111011001000101010;
assign LUT_4[34096] = 32'b00000000000000001010000111001011;
assign LUT_4[34097] = 32'b00000000000000000011010011000011;
assign LUT_4[34098] = 32'b00000000000000001001100001101111;
assign LUT_4[34099] = 32'b00000000000000000010101101100111;
assign LUT_4[34100] = 32'b00000000000000000111000111100111;
assign LUT_4[34101] = 32'b00000000000000000000010011011111;
assign LUT_4[34102] = 32'b00000000000000000110100010001011;
assign LUT_4[34103] = 32'b11111111111111111111101110000011;
assign LUT_4[34104] = 32'b00000000000000000011010011100000;
assign LUT_4[34105] = 32'b11111111111111111100011111011000;
assign LUT_4[34106] = 32'b00000000000000000010101110000100;
assign LUT_4[34107] = 32'b11111111111111111011111001111100;
assign LUT_4[34108] = 32'b00000000000000000000010011111100;
assign LUT_4[34109] = 32'b11111111111111111001011111110100;
assign LUT_4[34110] = 32'b11111111111111111111101110100000;
assign LUT_4[34111] = 32'b11111111111111111000111010011000;
assign LUT_4[34112] = 32'b00000000000000001111010001101010;
assign LUT_4[34113] = 32'b00000000000000001000011101100010;
assign LUT_4[34114] = 32'b00000000000000001110101100001110;
assign LUT_4[34115] = 32'b00000000000000000111111000000110;
assign LUT_4[34116] = 32'b00000000000000001100010010000110;
assign LUT_4[34117] = 32'b00000000000000000101011101111110;
assign LUT_4[34118] = 32'b00000000000000001011101100101010;
assign LUT_4[34119] = 32'b00000000000000000100111000100010;
assign LUT_4[34120] = 32'b00000000000000001000011101111111;
assign LUT_4[34121] = 32'b00000000000000000001101001110111;
assign LUT_4[34122] = 32'b00000000000000000111111000100011;
assign LUT_4[34123] = 32'b00000000000000000001000100011011;
assign LUT_4[34124] = 32'b00000000000000000101011110011011;
assign LUT_4[34125] = 32'b11111111111111111110101010010011;
assign LUT_4[34126] = 32'b00000000000000000100111000111111;
assign LUT_4[34127] = 32'b11111111111111111110000100110111;
assign LUT_4[34128] = 32'b00000000000000001101000011011000;
assign LUT_4[34129] = 32'b00000000000000000110001111010000;
assign LUT_4[34130] = 32'b00000000000000001100011101111100;
assign LUT_4[34131] = 32'b00000000000000000101101001110100;
assign LUT_4[34132] = 32'b00000000000000001010000011110100;
assign LUT_4[34133] = 32'b00000000000000000011001111101100;
assign LUT_4[34134] = 32'b00000000000000001001011110011000;
assign LUT_4[34135] = 32'b00000000000000000010101010010000;
assign LUT_4[34136] = 32'b00000000000000000110001111101101;
assign LUT_4[34137] = 32'b11111111111111111111011011100101;
assign LUT_4[34138] = 32'b00000000000000000101101010010001;
assign LUT_4[34139] = 32'b11111111111111111110110110001001;
assign LUT_4[34140] = 32'b00000000000000000011010000001001;
assign LUT_4[34141] = 32'b11111111111111111100011100000001;
assign LUT_4[34142] = 32'b00000000000000000010101010101101;
assign LUT_4[34143] = 32'b11111111111111111011110110100101;
assign LUT_4[34144] = 32'b00000000000000001101101100110001;
assign LUT_4[34145] = 32'b00000000000000000110111000101001;
assign LUT_4[34146] = 32'b00000000000000001101000111010101;
assign LUT_4[34147] = 32'b00000000000000000110010011001101;
assign LUT_4[34148] = 32'b00000000000000001010101101001101;
assign LUT_4[34149] = 32'b00000000000000000011111001000101;
assign LUT_4[34150] = 32'b00000000000000001010000111110001;
assign LUT_4[34151] = 32'b00000000000000000011010011101001;
assign LUT_4[34152] = 32'b00000000000000000110111001000110;
assign LUT_4[34153] = 32'b00000000000000000000000100111110;
assign LUT_4[34154] = 32'b00000000000000000110010011101010;
assign LUT_4[34155] = 32'b11111111111111111111011111100010;
assign LUT_4[34156] = 32'b00000000000000000011111001100010;
assign LUT_4[34157] = 32'b11111111111111111101000101011010;
assign LUT_4[34158] = 32'b00000000000000000011010100000110;
assign LUT_4[34159] = 32'b11111111111111111100011111111110;
assign LUT_4[34160] = 32'b00000000000000001011011110011111;
assign LUT_4[34161] = 32'b00000000000000000100101010010111;
assign LUT_4[34162] = 32'b00000000000000001010111001000011;
assign LUT_4[34163] = 32'b00000000000000000100000100111011;
assign LUT_4[34164] = 32'b00000000000000001000011110111011;
assign LUT_4[34165] = 32'b00000000000000000001101010110011;
assign LUT_4[34166] = 32'b00000000000000000111111001011111;
assign LUT_4[34167] = 32'b00000000000000000001000101010111;
assign LUT_4[34168] = 32'b00000000000000000100101010110100;
assign LUT_4[34169] = 32'b11111111111111111101110110101100;
assign LUT_4[34170] = 32'b00000000000000000100000101011000;
assign LUT_4[34171] = 32'b11111111111111111101010001010000;
assign LUT_4[34172] = 32'b00000000000000000001101011010000;
assign LUT_4[34173] = 32'b11111111111111111010110111001000;
assign LUT_4[34174] = 32'b00000000000000000001000101110100;
assign LUT_4[34175] = 32'b11111111111111111010010001101100;
assign LUT_4[34176] = 32'b00000000000000010000100000011110;
assign LUT_4[34177] = 32'b00000000000000001001101100010110;
assign LUT_4[34178] = 32'b00000000000000001111111011000010;
assign LUT_4[34179] = 32'b00000000000000001001000110111010;
assign LUT_4[34180] = 32'b00000000000000001101100000111010;
assign LUT_4[34181] = 32'b00000000000000000110101100110010;
assign LUT_4[34182] = 32'b00000000000000001100111011011110;
assign LUT_4[34183] = 32'b00000000000000000110000111010110;
assign LUT_4[34184] = 32'b00000000000000001001101100110011;
assign LUT_4[34185] = 32'b00000000000000000010111000101011;
assign LUT_4[34186] = 32'b00000000000000001001000111010111;
assign LUT_4[34187] = 32'b00000000000000000010010011001111;
assign LUT_4[34188] = 32'b00000000000000000110101101001111;
assign LUT_4[34189] = 32'b11111111111111111111111001000111;
assign LUT_4[34190] = 32'b00000000000000000110000111110011;
assign LUT_4[34191] = 32'b11111111111111111111010011101011;
assign LUT_4[34192] = 32'b00000000000000001110010010001100;
assign LUT_4[34193] = 32'b00000000000000000111011110000100;
assign LUT_4[34194] = 32'b00000000000000001101101100110000;
assign LUT_4[34195] = 32'b00000000000000000110111000101000;
assign LUT_4[34196] = 32'b00000000000000001011010010101000;
assign LUT_4[34197] = 32'b00000000000000000100011110100000;
assign LUT_4[34198] = 32'b00000000000000001010101101001100;
assign LUT_4[34199] = 32'b00000000000000000011111001000100;
assign LUT_4[34200] = 32'b00000000000000000111011110100001;
assign LUT_4[34201] = 32'b00000000000000000000101010011001;
assign LUT_4[34202] = 32'b00000000000000000110111001000101;
assign LUT_4[34203] = 32'b00000000000000000000000100111101;
assign LUT_4[34204] = 32'b00000000000000000100011110111101;
assign LUT_4[34205] = 32'b11111111111111111101101010110101;
assign LUT_4[34206] = 32'b00000000000000000011111001100001;
assign LUT_4[34207] = 32'b11111111111111111101000101011001;
assign LUT_4[34208] = 32'b00000000000000001110111011100101;
assign LUT_4[34209] = 32'b00000000000000001000000111011101;
assign LUT_4[34210] = 32'b00000000000000001110010110001001;
assign LUT_4[34211] = 32'b00000000000000000111100010000001;
assign LUT_4[34212] = 32'b00000000000000001011111100000001;
assign LUT_4[34213] = 32'b00000000000000000101000111111001;
assign LUT_4[34214] = 32'b00000000000000001011010110100101;
assign LUT_4[34215] = 32'b00000000000000000100100010011101;
assign LUT_4[34216] = 32'b00000000000000001000000111111010;
assign LUT_4[34217] = 32'b00000000000000000001010011110010;
assign LUT_4[34218] = 32'b00000000000000000111100010011110;
assign LUT_4[34219] = 32'b00000000000000000000101110010110;
assign LUT_4[34220] = 32'b00000000000000000101001000010110;
assign LUT_4[34221] = 32'b11111111111111111110010100001110;
assign LUT_4[34222] = 32'b00000000000000000100100010111010;
assign LUT_4[34223] = 32'b11111111111111111101101110110010;
assign LUT_4[34224] = 32'b00000000000000001100101101010011;
assign LUT_4[34225] = 32'b00000000000000000101111001001011;
assign LUT_4[34226] = 32'b00000000000000001100000111110111;
assign LUT_4[34227] = 32'b00000000000000000101010011101111;
assign LUT_4[34228] = 32'b00000000000000001001101101101111;
assign LUT_4[34229] = 32'b00000000000000000010111001100111;
assign LUT_4[34230] = 32'b00000000000000001001001000010011;
assign LUT_4[34231] = 32'b00000000000000000010010100001011;
assign LUT_4[34232] = 32'b00000000000000000101111001101000;
assign LUT_4[34233] = 32'b11111111111111111111000101100000;
assign LUT_4[34234] = 32'b00000000000000000101010100001100;
assign LUT_4[34235] = 32'b11111111111111111110100000000100;
assign LUT_4[34236] = 32'b00000000000000000010111010000100;
assign LUT_4[34237] = 32'b11111111111111111100000101111100;
assign LUT_4[34238] = 32'b00000000000000000010010100101000;
assign LUT_4[34239] = 32'b11111111111111111011100000100000;
assign LUT_4[34240] = 32'b00000000000000010001110111110010;
assign LUT_4[34241] = 32'b00000000000000001011000011101010;
assign LUT_4[34242] = 32'b00000000000000010001010010010110;
assign LUT_4[34243] = 32'b00000000000000001010011110001110;
assign LUT_4[34244] = 32'b00000000000000001110111000001110;
assign LUT_4[34245] = 32'b00000000000000001000000100000110;
assign LUT_4[34246] = 32'b00000000000000001110010010110010;
assign LUT_4[34247] = 32'b00000000000000000111011110101010;
assign LUT_4[34248] = 32'b00000000000000001011000100000111;
assign LUT_4[34249] = 32'b00000000000000000100001111111111;
assign LUT_4[34250] = 32'b00000000000000001010011110101011;
assign LUT_4[34251] = 32'b00000000000000000011101010100011;
assign LUT_4[34252] = 32'b00000000000000001000000100100011;
assign LUT_4[34253] = 32'b00000000000000000001010000011011;
assign LUT_4[34254] = 32'b00000000000000000111011111000111;
assign LUT_4[34255] = 32'b00000000000000000000101010111111;
assign LUT_4[34256] = 32'b00000000000000001111101001100000;
assign LUT_4[34257] = 32'b00000000000000001000110101011000;
assign LUT_4[34258] = 32'b00000000000000001111000100000100;
assign LUT_4[34259] = 32'b00000000000000001000001111111100;
assign LUT_4[34260] = 32'b00000000000000001100101001111100;
assign LUT_4[34261] = 32'b00000000000000000101110101110100;
assign LUT_4[34262] = 32'b00000000000000001100000100100000;
assign LUT_4[34263] = 32'b00000000000000000101010000011000;
assign LUT_4[34264] = 32'b00000000000000001000110101110101;
assign LUT_4[34265] = 32'b00000000000000000010000001101101;
assign LUT_4[34266] = 32'b00000000000000001000010000011001;
assign LUT_4[34267] = 32'b00000000000000000001011100010001;
assign LUT_4[34268] = 32'b00000000000000000101110110010001;
assign LUT_4[34269] = 32'b11111111111111111111000010001001;
assign LUT_4[34270] = 32'b00000000000000000101010000110101;
assign LUT_4[34271] = 32'b11111111111111111110011100101101;
assign LUT_4[34272] = 32'b00000000000000010000010010111001;
assign LUT_4[34273] = 32'b00000000000000001001011110110001;
assign LUT_4[34274] = 32'b00000000000000001111101101011101;
assign LUT_4[34275] = 32'b00000000000000001000111001010101;
assign LUT_4[34276] = 32'b00000000000000001101010011010101;
assign LUT_4[34277] = 32'b00000000000000000110011111001101;
assign LUT_4[34278] = 32'b00000000000000001100101101111001;
assign LUT_4[34279] = 32'b00000000000000000101111001110001;
assign LUT_4[34280] = 32'b00000000000000001001011111001110;
assign LUT_4[34281] = 32'b00000000000000000010101011000110;
assign LUT_4[34282] = 32'b00000000000000001000111001110010;
assign LUT_4[34283] = 32'b00000000000000000010000101101010;
assign LUT_4[34284] = 32'b00000000000000000110011111101010;
assign LUT_4[34285] = 32'b11111111111111111111101011100010;
assign LUT_4[34286] = 32'b00000000000000000101111010001110;
assign LUT_4[34287] = 32'b11111111111111111111000110000110;
assign LUT_4[34288] = 32'b00000000000000001110000100100111;
assign LUT_4[34289] = 32'b00000000000000000111010000011111;
assign LUT_4[34290] = 32'b00000000000000001101011111001011;
assign LUT_4[34291] = 32'b00000000000000000110101011000011;
assign LUT_4[34292] = 32'b00000000000000001011000101000011;
assign LUT_4[34293] = 32'b00000000000000000100010000111011;
assign LUT_4[34294] = 32'b00000000000000001010011111100111;
assign LUT_4[34295] = 32'b00000000000000000011101011011111;
assign LUT_4[34296] = 32'b00000000000000000111010000111100;
assign LUT_4[34297] = 32'b00000000000000000000011100110100;
assign LUT_4[34298] = 32'b00000000000000000110101011100000;
assign LUT_4[34299] = 32'b11111111111111111111110111011000;
assign LUT_4[34300] = 32'b00000000000000000100010001011000;
assign LUT_4[34301] = 32'b11111111111111111101011101010000;
assign LUT_4[34302] = 32'b00000000000000000011101011111100;
assign LUT_4[34303] = 32'b11111111111111111100110111110100;
assign LUT_4[34304] = 32'b00000000000000001000000010111011;
assign LUT_4[34305] = 32'b00000000000000000001001110110011;
assign LUT_4[34306] = 32'b00000000000000000111011101011111;
assign LUT_4[34307] = 32'b00000000000000000000101001010111;
assign LUT_4[34308] = 32'b00000000000000000101000011010111;
assign LUT_4[34309] = 32'b11111111111111111110001111001111;
assign LUT_4[34310] = 32'b00000000000000000100011101111011;
assign LUT_4[34311] = 32'b11111111111111111101101001110011;
assign LUT_4[34312] = 32'b00000000000000000001001111010000;
assign LUT_4[34313] = 32'b11111111111111111010011011001000;
assign LUT_4[34314] = 32'b00000000000000000000101001110100;
assign LUT_4[34315] = 32'b11111111111111111001110101101100;
assign LUT_4[34316] = 32'b11111111111111111110001111101100;
assign LUT_4[34317] = 32'b11111111111111110111011011100100;
assign LUT_4[34318] = 32'b11111111111111111101101010010000;
assign LUT_4[34319] = 32'b11111111111111110110110110001000;
assign LUT_4[34320] = 32'b00000000000000000101110100101001;
assign LUT_4[34321] = 32'b11111111111111111111000000100001;
assign LUT_4[34322] = 32'b00000000000000000101001111001101;
assign LUT_4[34323] = 32'b11111111111111111110011011000101;
assign LUT_4[34324] = 32'b00000000000000000010110101000101;
assign LUT_4[34325] = 32'b11111111111111111100000000111101;
assign LUT_4[34326] = 32'b00000000000000000010001111101001;
assign LUT_4[34327] = 32'b11111111111111111011011011100001;
assign LUT_4[34328] = 32'b11111111111111111111000000111110;
assign LUT_4[34329] = 32'b11111111111111111000001100110110;
assign LUT_4[34330] = 32'b11111111111111111110011011100010;
assign LUT_4[34331] = 32'b11111111111111110111100111011010;
assign LUT_4[34332] = 32'b11111111111111111100000001011010;
assign LUT_4[34333] = 32'b11111111111111110101001101010010;
assign LUT_4[34334] = 32'b11111111111111111011011011111110;
assign LUT_4[34335] = 32'b11111111111111110100100111110110;
assign LUT_4[34336] = 32'b00000000000000000110011110000010;
assign LUT_4[34337] = 32'b11111111111111111111101001111010;
assign LUT_4[34338] = 32'b00000000000000000101111000100110;
assign LUT_4[34339] = 32'b11111111111111111111000100011110;
assign LUT_4[34340] = 32'b00000000000000000011011110011110;
assign LUT_4[34341] = 32'b11111111111111111100101010010110;
assign LUT_4[34342] = 32'b00000000000000000010111001000010;
assign LUT_4[34343] = 32'b11111111111111111100000100111010;
assign LUT_4[34344] = 32'b11111111111111111111101010010111;
assign LUT_4[34345] = 32'b11111111111111111000110110001111;
assign LUT_4[34346] = 32'b11111111111111111111000100111011;
assign LUT_4[34347] = 32'b11111111111111111000010000110011;
assign LUT_4[34348] = 32'b11111111111111111100101010110011;
assign LUT_4[34349] = 32'b11111111111111110101110110101011;
assign LUT_4[34350] = 32'b11111111111111111100000101010111;
assign LUT_4[34351] = 32'b11111111111111110101010001001111;
assign LUT_4[34352] = 32'b00000000000000000100001111110000;
assign LUT_4[34353] = 32'b11111111111111111101011011101000;
assign LUT_4[34354] = 32'b00000000000000000011101010010100;
assign LUT_4[34355] = 32'b11111111111111111100110110001100;
assign LUT_4[34356] = 32'b00000000000000000001010000001100;
assign LUT_4[34357] = 32'b11111111111111111010011100000100;
assign LUT_4[34358] = 32'b00000000000000000000101010110000;
assign LUT_4[34359] = 32'b11111111111111111001110110101000;
assign LUT_4[34360] = 32'b11111111111111111101011100000101;
assign LUT_4[34361] = 32'b11111111111111110110100111111101;
assign LUT_4[34362] = 32'b11111111111111111100110110101001;
assign LUT_4[34363] = 32'b11111111111111110110000010100001;
assign LUT_4[34364] = 32'b11111111111111111010011100100001;
assign LUT_4[34365] = 32'b11111111111111110011101000011001;
assign LUT_4[34366] = 32'b11111111111111111001110111000101;
assign LUT_4[34367] = 32'b11111111111111110011000010111101;
assign LUT_4[34368] = 32'b00000000000000001001011010001111;
assign LUT_4[34369] = 32'b00000000000000000010100110000111;
assign LUT_4[34370] = 32'b00000000000000001000110100110011;
assign LUT_4[34371] = 32'b00000000000000000010000000101011;
assign LUT_4[34372] = 32'b00000000000000000110011010101011;
assign LUT_4[34373] = 32'b11111111111111111111100110100011;
assign LUT_4[34374] = 32'b00000000000000000101110101001111;
assign LUT_4[34375] = 32'b11111111111111111111000001000111;
assign LUT_4[34376] = 32'b00000000000000000010100110100100;
assign LUT_4[34377] = 32'b11111111111111111011110010011100;
assign LUT_4[34378] = 32'b00000000000000000010000001001000;
assign LUT_4[34379] = 32'b11111111111111111011001101000000;
assign LUT_4[34380] = 32'b11111111111111111111100111000000;
assign LUT_4[34381] = 32'b11111111111111111000110010111000;
assign LUT_4[34382] = 32'b11111111111111111111000001100100;
assign LUT_4[34383] = 32'b11111111111111111000001101011100;
assign LUT_4[34384] = 32'b00000000000000000111001011111101;
assign LUT_4[34385] = 32'b00000000000000000000010111110101;
assign LUT_4[34386] = 32'b00000000000000000110100110100001;
assign LUT_4[34387] = 32'b11111111111111111111110010011001;
assign LUT_4[34388] = 32'b00000000000000000100001100011001;
assign LUT_4[34389] = 32'b11111111111111111101011000010001;
assign LUT_4[34390] = 32'b00000000000000000011100110111101;
assign LUT_4[34391] = 32'b11111111111111111100110010110101;
assign LUT_4[34392] = 32'b00000000000000000000011000010010;
assign LUT_4[34393] = 32'b11111111111111111001100100001010;
assign LUT_4[34394] = 32'b11111111111111111111110010110110;
assign LUT_4[34395] = 32'b11111111111111111000111110101110;
assign LUT_4[34396] = 32'b11111111111111111101011000101110;
assign LUT_4[34397] = 32'b11111111111111110110100100100110;
assign LUT_4[34398] = 32'b11111111111111111100110011010010;
assign LUT_4[34399] = 32'b11111111111111110101111111001010;
assign LUT_4[34400] = 32'b00000000000000000111110101010110;
assign LUT_4[34401] = 32'b00000000000000000001000001001110;
assign LUT_4[34402] = 32'b00000000000000000111001111111010;
assign LUT_4[34403] = 32'b00000000000000000000011011110010;
assign LUT_4[34404] = 32'b00000000000000000100110101110010;
assign LUT_4[34405] = 32'b11111111111111111110000001101010;
assign LUT_4[34406] = 32'b00000000000000000100010000010110;
assign LUT_4[34407] = 32'b11111111111111111101011100001110;
assign LUT_4[34408] = 32'b00000000000000000001000001101011;
assign LUT_4[34409] = 32'b11111111111111111010001101100011;
assign LUT_4[34410] = 32'b00000000000000000000011100001111;
assign LUT_4[34411] = 32'b11111111111111111001101000000111;
assign LUT_4[34412] = 32'b11111111111111111110000010000111;
assign LUT_4[34413] = 32'b11111111111111110111001101111111;
assign LUT_4[34414] = 32'b11111111111111111101011100101011;
assign LUT_4[34415] = 32'b11111111111111110110101000100011;
assign LUT_4[34416] = 32'b00000000000000000101100111000100;
assign LUT_4[34417] = 32'b11111111111111111110110010111100;
assign LUT_4[34418] = 32'b00000000000000000101000001101000;
assign LUT_4[34419] = 32'b11111111111111111110001101100000;
assign LUT_4[34420] = 32'b00000000000000000010100111100000;
assign LUT_4[34421] = 32'b11111111111111111011110011011000;
assign LUT_4[34422] = 32'b00000000000000000010000010000100;
assign LUT_4[34423] = 32'b11111111111111111011001101111100;
assign LUT_4[34424] = 32'b11111111111111111110110011011001;
assign LUT_4[34425] = 32'b11111111111111110111111111010001;
assign LUT_4[34426] = 32'b11111111111111111110001101111101;
assign LUT_4[34427] = 32'b11111111111111110111011001110101;
assign LUT_4[34428] = 32'b11111111111111111011110011110101;
assign LUT_4[34429] = 32'b11111111111111110100111111101101;
assign LUT_4[34430] = 32'b11111111111111111011001110011001;
assign LUT_4[34431] = 32'b11111111111111110100011010010001;
assign LUT_4[34432] = 32'b00000000000000001010101001000011;
assign LUT_4[34433] = 32'b00000000000000000011110100111011;
assign LUT_4[34434] = 32'b00000000000000001010000011100111;
assign LUT_4[34435] = 32'b00000000000000000011001111011111;
assign LUT_4[34436] = 32'b00000000000000000111101001011111;
assign LUT_4[34437] = 32'b00000000000000000000110101010111;
assign LUT_4[34438] = 32'b00000000000000000111000100000011;
assign LUT_4[34439] = 32'b00000000000000000000001111111011;
assign LUT_4[34440] = 32'b00000000000000000011110101011000;
assign LUT_4[34441] = 32'b11111111111111111101000001010000;
assign LUT_4[34442] = 32'b00000000000000000011001111111100;
assign LUT_4[34443] = 32'b11111111111111111100011011110100;
assign LUT_4[34444] = 32'b00000000000000000000110101110100;
assign LUT_4[34445] = 32'b11111111111111111010000001101100;
assign LUT_4[34446] = 32'b00000000000000000000010000011000;
assign LUT_4[34447] = 32'b11111111111111111001011100010000;
assign LUT_4[34448] = 32'b00000000000000001000011010110001;
assign LUT_4[34449] = 32'b00000000000000000001100110101001;
assign LUT_4[34450] = 32'b00000000000000000111110101010101;
assign LUT_4[34451] = 32'b00000000000000000001000001001101;
assign LUT_4[34452] = 32'b00000000000000000101011011001101;
assign LUT_4[34453] = 32'b11111111111111111110100111000101;
assign LUT_4[34454] = 32'b00000000000000000100110101110001;
assign LUT_4[34455] = 32'b11111111111111111110000001101001;
assign LUT_4[34456] = 32'b00000000000000000001100111000110;
assign LUT_4[34457] = 32'b11111111111111111010110010111110;
assign LUT_4[34458] = 32'b00000000000000000001000001101010;
assign LUT_4[34459] = 32'b11111111111111111010001101100010;
assign LUT_4[34460] = 32'b11111111111111111110100111100010;
assign LUT_4[34461] = 32'b11111111111111110111110011011010;
assign LUT_4[34462] = 32'b11111111111111111110000010000110;
assign LUT_4[34463] = 32'b11111111111111110111001101111110;
assign LUT_4[34464] = 32'b00000000000000001001000100001010;
assign LUT_4[34465] = 32'b00000000000000000010010000000010;
assign LUT_4[34466] = 32'b00000000000000001000011110101110;
assign LUT_4[34467] = 32'b00000000000000000001101010100110;
assign LUT_4[34468] = 32'b00000000000000000110000100100110;
assign LUT_4[34469] = 32'b11111111111111111111010000011110;
assign LUT_4[34470] = 32'b00000000000000000101011111001010;
assign LUT_4[34471] = 32'b11111111111111111110101011000010;
assign LUT_4[34472] = 32'b00000000000000000010010000011111;
assign LUT_4[34473] = 32'b11111111111111111011011100010111;
assign LUT_4[34474] = 32'b00000000000000000001101011000011;
assign LUT_4[34475] = 32'b11111111111111111010110110111011;
assign LUT_4[34476] = 32'b11111111111111111111010000111011;
assign LUT_4[34477] = 32'b11111111111111111000011100110011;
assign LUT_4[34478] = 32'b11111111111111111110101011011111;
assign LUT_4[34479] = 32'b11111111111111110111110111010111;
assign LUT_4[34480] = 32'b00000000000000000110110101111000;
assign LUT_4[34481] = 32'b00000000000000000000000001110000;
assign LUT_4[34482] = 32'b00000000000000000110010000011100;
assign LUT_4[34483] = 32'b11111111111111111111011100010100;
assign LUT_4[34484] = 32'b00000000000000000011110110010100;
assign LUT_4[34485] = 32'b11111111111111111101000010001100;
assign LUT_4[34486] = 32'b00000000000000000011010000111000;
assign LUT_4[34487] = 32'b11111111111111111100011100110000;
assign LUT_4[34488] = 32'b00000000000000000000000010001101;
assign LUT_4[34489] = 32'b11111111111111111001001110000101;
assign LUT_4[34490] = 32'b11111111111111111111011100110001;
assign LUT_4[34491] = 32'b11111111111111111000101000101001;
assign LUT_4[34492] = 32'b11111111111111111101000010101001;
assign LUT_4[34493] = 32'b11111111111111110110001110100001;
assign LUT_4[34494] = 32'b11111111111111111100011101001101;
assign LUT_4[34495] = 32'b11111111111111110101101001000101;
assign LUT_4[34496] = 32'b00000000000000001100000000010111;
assign LUT_4[34497] = 32'b00000000000000000101001100001111;
assign LUT_4[34498] = 32'b00000000000000001011011010111011;
assign LUT_4[34499] = 32'b00000000000000000100100110110011;
assign LUT_4[34500] = 32'b00000000000000001001000000110011;
assign LUT_4[34501] = 32'b00000000000000000010001100101011;
assign LUT_4[34502] = 32'b00000000000000001000011011010111;
assign LUT_4[34503] = 32'b00000000000000000001100111001111;
assign LUT_4[34504] = 32'b00000000000000000101001100101100;
assign LUT_4[34505] = 32'b11111111111111111110011000100100;
assign LUT_4[34506] = 32'b00000000000000000100100111010000;
assign LUT_4[34507] = 32'b11111111111111111101110011001000;
assign LUT_4[34508] = 32'b00000000000000000010001101001000;
assign LUT_4[34509] = 32'b11111111111111111011011001000000;
assign LUT_4[34510] = 32'b00000000000000000001100111101100;
assign LUT_4[34511] = 32'b11111111111111111010110011100100;
assign LUT_4[34512] = 32'b00000000000000001001110010000101;
assign LUT_4[34513] = 32'b00000000000000000010111101111101;
assign LUT_4[34514] = 32'b00000000000000001001001100101001;
assign LUT_4[34515] = 32'b00000000000000000010011000100001;
assign LUT_4[34516] = 32'b00000000000000000110110010100001;
assign LUT_4[34517] = 32'b11111111111111111111111110011001;
assign LUT_4[34518] = 32'b00000000000000000110001101000101;
assign LUT_4[34519] = 32'b11111111111111111111011000111101;
assign LUT_4[34520] = 32'b00000000000000000010111110011010;
assign LUT_4[34521] = 32'b11111111111111111100001010010010;
assign LUT_4[34522] = 32'b00000000000000000010011000111110;
assign LUT_4[34523] = 32'b11111111111111111011100100110110;
assign LUT_4[34524] = 32'b11111111111111111111111110110110;
assign LUT_4[34525] = 32'b11111111111111111001001010101110;
assign LUT_4[34526] = 32'b11111111111111111111011001011010;
assign LUT_4[34527] = 32'b11111111111111111000100101010010;
assign LUT_4[34528] = 32'b00000000000000001010011011011110;
assign LUT_4[34529] = 32'b00000000000000000011100111010110;
assign LUT_4[34530] = 32'b00000000000000001001110110000010;
assign LUT_4[34531] = 32'b00000000000000000011000001111010;
assign LUT_4[34532] = 32'b00000000000000000111011011111010;
assign LUT_4[34533] = 32'b00000000000000000000100111110010;
assign LUT_4[34534] = 32'b00000000000000000110110110011110;
assign LUT_4[34535] = 32'b00000000000000000000000010010110;
assign LUT_4[34536] = 32'b00000000000000000011100111110011;
assign LUT_4[34537] = 32'b11111111111111111100110011101011;
assign LUT_4[34538] = 32'b00000000000000000011000010010111;
assign LUT_4[34539] = 32'b11111111111111111100001110001111;
assign LUT_4[34540] = 32'b00000000000000000000101000001111;
assign LUT_4[34541] = 32'b11111111111111111001110100000111;
assign LUT_4[34542] = 32'b00000000000000000000000010110011;
assign LUT_4[34543] = 32'b11111111111111111001001110101011;
assign LUT_4[34544] = 32'b00000000000000001000001101001100;
assign LUT_4[34545] = 32'b00000000000000000001011001000100;
assign LUT_4[34546] = 32'b00000000000000000111100111110000;
assign LUT_4[34547] = 32'b00000000000000000000110011101000;
assign LUT_4[34548] = 32'b00000000000000000101001101101000;
assign LUT_4[34549] = 32'b11111111111111111110011001100000;
assign LUT_4[34550] = 32'b00000000000000000100101000001100;
assign LUT_4[34551] = 32'b11111111111111111101110100000100;
assign LUT_4[34552] = 32'b00000000000000000001011001100001;
assign LUT_4[34553] = 32'b11111111111111111010100101011001;
assign LUT_4[34554] = 32'b00000000000000000000110100000101;
assign LUT_4[34555] = 32'b11111111111111111001111111111101;
assign LUT_4[34556] = 32'b11111111111111111110011001111101;
assign LUT_4[34557] = 32'b11111111111111110111100101110101;
assign LUT_4[34558] = 32'b11111111111111111101110100100001;
assign LUT_4[34559] = 32'b11111111111111110111000000011001;
assign LUT_4[34560] = 32'b00000000000000001100111110011110;
assign LUT_4[34561] = 32'b00000000000000000110001010010110;
assign LUT_4[34562] = 32'b00000000000000001100011001000010;
assign LUT_4[34563] = 32'b00000000000000000101100100111010;
assign LUT_4[34564] = 32'b00000000000000001001111110111010;
assign LUT_4[34565] = 32'b00000000000000000011001010110010;
assign LUT_4[34566] = 32'b00000000000000001001011001011110;
assign LUT_4[34567] = 32'b00000000000000000010100101010110;
assign LUT_4[34568] = 32'b00000000000000000110001010110011;
assign LUT_4[34569] = 32'b11111111111111111111010110101011;
assign LUT_4[34570] = 32'b00000000000000000101100101010111;
assign LUT_4[34571] = 32'b11111111111111111110110001001111;
assign LUT_4[34572] = 32'b00000000000000000011001011001111;
assign LUT_4[34573] = 32'b11111111111111111100010111000111;
assign LUT_4[34574] = 32'b00000000000000000010100101110011;
assign LUT_4[34575] = 32'b11111111111111111011110001101011;
assign LUT_4[34576] = 32'b00000000000000001010110000001100;
assign LUT_4[34577] = 32'b00000000000000000011111100000100;
assign LUT_4[34578] = 32'b00000000000000001010001010110000;
assign LUT_4[34579] = 32'b00000000000000000011010110101000;
assign LUT_4[34580] = 32'b00000000000000000111110000101000;
assign LUT_4[34581] = 32'b00000000000000000000111100100000;
assign LUT_4[34582] = 32'b00000000000000000111001011001100;
assign LUT_4[34583] = 32'b00000000000000000000010111000100;
assign LUT_4[34584] = 32'b00000000000000000011111100100001;
assign LUT_4[34585] = 32'b11111111111111111101001000011001;
assign LUT_4[34586] = 32'b00000000000000000011010111000101;
assign LUT_4[34587] = 32'b11111111111111111100100010111101;
assign LUT_4[34588] = 32'b00000000000000000000111100111101;
assign LUT_4[34589] = 32'b11111111111111111010001000110101;
assign LUT_4[34590] = 32'b00000000000000000000010111100001;
assign LUT_4[34591] = 32'b11111111111111111001100011011001;
assign LUT_4[34592] = 32'b00000000000000001011011001100101;
assign LUT_4[34593] = 32'b00000000000000000100100101011101;
assign LUT_4[34594] = 32'b00000000000000001010110100001001;
assign LUT_4[34595] = 32'b00000000000000000100000000000001;
assign LUT_4[34596] = 32'b00000000000000001000011010000001;
assign LUT_4[34597] = 32'b00000000000000000001100101111001;
assign LUT_4[34598] = 32'b00000000000000000111110100100101;
assign LUT_4[34599] = 32'b00000000000000000001000000011101;
assign LUT_4[34600] = 32'b00000000000000000100100101111010;
assign LUT_4[34601] = 32'b11111111111111111101110001110010;
assign LUT_4[34602] = 32'b00000000000000000100000000011110;
assign LUT_4[34603] = 32'b11111111111111111101001100010110;
assign LUT_4[34604] = 32'b00000000000000000001100110010110;
assign LUT_4[34605] = 32'b11111111111111111010110010001110;
assign LUT_4[34606] = 32'b00000000000000000001000000111010;
assign LUT_4[34607] = 32'b11111111111111111010001100110010;
assign LUT_4[34608] = 32'b00000000000000001001001011010011;
assign LUT_4[34609] = 32'b00000000000000000010010111001011;
assign LUT_4[34610] = 32'b00000000000000001000100101110111;
assign LUT_4[34611] = 32'b00000000000000000001110001101111;
assign LUT_4[34612] = 32'b00000000000000000110001011101111;
assign LUT_4[34613] = 32'b11111111111111111111010111100111;
assign LUT_4[34614] = 32'b00000000000000000101100110010011;
assign LUT_4[34615] = 32'b11111111111111111110110010001011;
assign LUT_4[34616] = 32'b00000000000000000010010111101000;
assign LUT_4[34617] = 32'b11111111111111111011100011100000;
assign LUT_4[34618] = 32'b00000000000000000001110010001100;
assign LUT_4[34619] = 32'b11111111111111111010111110000100;
assign LUT_4[34620] = 32'b11111111111111111111011000000100;
assign LUT_4[34621] = 32'b11111111111111111000100011111100;
assign LUT_4[34622] = 32'b11111111111111111110110010101000;
assign LUT_4[34623] = 32'b11111111111111110111111110100000;
assign LUT_4[34624] = 32'b00000000000000001110010101110010;
assign LUT_4[34625] = 32'b00000000000000000111100001101010;
assign LUT_4[34626] = 32'b00000000000000001101110000010110;
assign LUT_4[34627] = 32'b00000000000000000110111100001110;
assign LUT_4[34628] = 32'b00000000000000001011010110001110;
assign LUT_4[34629] = 32'b00000000000000000100100010000110;
assign LUT_4[34630] = 32'b00000000000000001010110000110010;
assign LUT_4[34631] = 32'b00000000000000000011111100101010;
assign LUT_4[34632] = 32'b00000000000000000111100010000111;
assign LUT_4[34633] = 32'b00000000000000000000101101111111;
assign LUT_4[34634] = 32'b00000000000000000110111100101011;
assign LUT_4[34635] = 32'b00000000000000000000001000100011;
assign LUT_4[34636] = 32'b00000000000000000100100010100011;
assign LUT_4[34637] = 32'b11111111111111111101101110011011;
assign LUT_4[34638] = 32'b00000000000000000011111101000111;
assign LUT_4[34639] = 32'b11111111111111111101001000111111;
assign LUT_4[34640] = 32'b00000000000000001100000111100000;
assign LUT_4[34641] = 32'b00000000000000000101010011011000;
assign LUT_4[34642] = 32'b00000000000000001011100010000100;
assign LUT_4[34643] = 32'b00000000000000000100101101111100;
assign LUT_4[34644] = 32'b00000000000000001001000111111100;
assign LUT_4[34645] = 32'b00000000000000000010010011110100;
assign LUT_4[34646] = 32'b00000000000000001000100010100000;
assign LUT_4[34647] = 32'b00000000000000000001101110011000;
assign LUT_4[34648] = 32'b00000000000000000101010011110101;
assign LUT_4[34649] = 32'b11111111111111111110011111101101;
assign LUT_4[34650] = 32'b00000000000000000100101110011001;
assign LUT_4[34651] = 32'b11111111111111111101111010010001;
assign LUT_4[34652] = 32'b00000000000000000010010100010001;
assign LUT_4[34653] = 32'b11111111111111111011100000001001;
assign LUT_4[34654] = 32'b00000000000000000001101110110101;
assign LUT_4[34655] = 32'b11111111111111111010111010101101;
assign LUT_4[34656] = 32'b00000000000000001100110000111001;
assign LUT_4[34657] = 32'b00000000000000000101111100110001;
assign LUT_4[34658] = 32'b00000000000000001100001011011101;
assign LUT_4[34659] = 32'b00000000000000000101010111010101;
assign LUT_4[34660] = 32'b00000000000000001001110001010101;
assign LUT_4[34661] = 32'b00000000000000000010111101001101;
assign LUT_4[34662] = 32'b00000000000000001001001011111001;
assign LUT_4[34663] = 32'b00000000000000000010010111110001;
assign LUT_4[34664] = 32'b00000000000000000101111101001110;
assign LUT_4[34665] = 32'b11111111111111111111001001000110;
assign LUT_4[34666] = 32'b00000000000000000101010111110010;
assign LUT_4[34667] = 32'b11111111111111111110100011101010;
assign LUT_4[34668] = 32'b00000000000000000010111101101010;
assign LUT_4[34669] = 32'b11111111111111111100001001100010;
assign LUT_4[34670] = 32'b00000000000000000010011000001110;
assign LUT_4[34671] = 32'b11111111111111111011100100000110;
assign LUT_4[34672] = 32'b00000000000000001010100010100111;
assign LUT_4[34673] = 32'b00000000000000000011101110011111;
assign LUT_4[34674] = 32'b00000000000000001001111101001011;
assign LUT_4[34675] = 32'b00000000000000000011001001000011;
assign LUT_4[34676] = 32'b00000000000000000111100011000011;
assign LUT_4[34677] = 32'b00000000000000000000101110111011;
assign LUT_4[34678] = 32'b00000000000000000110111101100111;
assign LUT_4[34679] = 32'b00000000000000000000001001011111;
assign LUT_4[34680] = 32'b00000000000000000011101110111100;
assign LUT_4[34681] = 32'b11111111111111111100111010110100;
assign LUT_4[34682] = 32'b00000000000000000011001001100000;
assign LUT_4[34683] = 32'b11111111111111111100010101011000;
assign LUT_4[34684] = 32'b00000000000000000000101111011000;
assign LUT_4[34685] = 32'b11111111111111111001111011010000;
assign LUT_4[34686] = 32'b00000000000000000000001001111100;
assign LUT_4[34687] = 32'b11111111111111111001010101110100;
assign LUT_4[34688] = 32'b00000000000000001111100100100110;
assign LUT_4[34689] = 32'b00000000000000001000110000011110;
assign LUT_4[34690] = 32'b00000000000000001110111111001010;
assign LUT_4[34691] = 32'b00000000000000001000001011000010;
assign LUT_4[34692] = 32'b00000000000000001100100101000010;
assign LUT_4[34693] = 32'b00000000000000000101110000111010;
assign LUT_4[34694] = 32'b00000000000000001011111111100110;
assign LUT_4[34695] = 32'b00000000000000000101001011011110;
assign LUT_4[34696] = 32'b00000000000000001000110000111011;
assign LUT_4[34697] = 32'b00000000000000000001111100110011;
assign LUT_4[34698] = 32'b00000000000000001000001011011111;
assign LUT_4[34699] = 32'b00000000000000000001010111010111;
assign LUT_4[34700] = 32'b00000000000000000101110001010111;
assign LUT_4[34701] = 32'b11111111111111111110111101001111;
assign LUT_4[34702] = 32'b00000000000000000101001011111011;
assign LUT_4[34703] = 32'b11111111111111111110010111110011;
assign LUT_4[34704] = 32'b00000000000000001101010110010100;
assign LUT_4[34705] = 32'b00000000000000000110100010001100;
assign LUT_4[34706] = 32'b00000000000000001100110000111000;
assign LUT_4[34707] = 32'b00000000000000000101111100110000;
assign LUT_4[34708] = 32'b00000000000000001010010110110000;
assign LUT_4[34709] = 32'b00000000000000000011100010101000;
assign LUT_4[34710] = 32'b00000000000000001001110001010100;
assign LUT_4[34711] = 32'b00000000000000000010111101001100;
assign LUT_4[34712] = 32'b00000000000000000110100010101001;
assign LUT_4[34713] = 32'b11111111111111111111101110100001;
assign LUT_4[34714] = 32'b00000000000000000101111101001101;
assign LUT_4[34715] = 32'b11111111111111111111001001000101;
assign LUT_4[34716] = 32'b00000000000000000011100011000101;
assign LUT_4[34717] = 32'b11111111111111111100101110111101;
assign LUT_4[34718] = 32'b00000000000000000010111101101001;
assign LUT_4[34719] = 32'b11111111111111111100001001100001;
assign LUT_4[34720] = 32'b00000000000000001101111111101101;
assign LUT_4[34721] = 32'b00000000000000000111001011100101;
assign LUT_4[34722] = 32'b00000000000000001101011010010001;
assign LUT_4[34723] = 32'b00000000000000000110100110001001;
assign LUT_4[34724] = 32'b00000000000000001011000000001001;
assign LUT_4[34725] = 32'b00000000000000000100001100000001;
assign LUT_4[34726] = 32'b00000000000000001010011010101101;
assign LUT_4[34727] = 32'b00000000000000000011100110100101;
assign LUT_4[34728] = 32'b00000000000000000111001100000010;
assign LUT_4[34729] = 32'b00000000000000000000010111111010;
assign LUT_4[34730] = 32'b00000000000000000110100110100110;
assign LUT_4[34731] = 32'b11111111111111111111110010011110;
assign LUT_4[34732] = 32'b00000000000000000100001100011110;
assign LUT_4[34733] = 32'b11111111111111111101011000010110;
assign LUT_4[34734] = 32'b00000000000000000011100111000010;
assign LUT_4[34735] = 32'b11111111111111111100110010111010;
assign LUT_4[34736] = 32'b00000000000000001011110001011011;
assign LUT_4[34737] = 32'b00000000000000000100111101010011;
assign LUT_4[34738] = 32'b00000000000000001011001011111111;
assign LUT_4[34739] = 32'b00000000000000000100010111110111;
assign LUT_4[34740] = 32'b00000000000000001000110001110111;
assign LUT_4[34741] = 32'b00000000000000000001111101101111;
assign LUT_4[34742] = 32'b00000000000000001000001100011011;
assign LUT_4[34743] = 32'b00000000000000000001011000010011;
assign LUT_4[34744] = 32'b00000000000000000100111101110000;
assign LUT_4[34745] = 32'b11111111111111111110001001101000;
assign LUT_4[34746] = 32'b00000000000000000100011000010100;
assign LUT_4[34747] = 32'b11111111111111111101100100001100;
assign LUT_4[34748] = 32'b00000000000000000001111110001100;
assign LUT_4[34749] = 32'b11111111111111111011001010000100;
assign LUT_4[34750] = 32'b00000000000000000001011000110000;
assign LUT_4[34751] = 32'b11111111111111111010100100101000;
assign LUT_4[34752] = 32'b00000000000000010000111011111010;
assign LUT_4[34753] = 32'b00000000000000001010000111110010;
assign LUT_4[34754] = 32'b00000000000000010000010110011110;
assign LUT_4[34755] = 32'b00000000000000001001100010010110;
assign LUT_4[34756] = 32'b00000000000000001101111100010110;
assign LUT_4[34757] = 32'b00000000000000000111001000001110;
assign LUT_4[34758] = 32'b00000000000000001101010110111010;
assign LUT_4[34759] = 32'b00000000000000000110100010110010;
assign LUT_4[34760] = 32'b00000000000000001010001000001111;
assign LUT_4[34761] = 32'b00000000000000000011010100000111;
assign LUT_4[34762] = 32'b00000000000000001001100010110011;
assign LUT_4[34763] = 32'b00000000000000000010101110101011;
assign LUT_4[34764] = 32'b00000000000000000111001000101011;
assign LUT_4[34765] = 32'b00000000000000000000010100100011;
assign LUT_4[34766] = 32'b00000000000000000110100011001111;
assign LUT_4[34767] = 32'b11111111111111111111101111000111;
assign LUT_4[34768] = 32'b00000000000000001110101101101000;
assign LUT_4[34769] = 32'b00000000000000000111111001100000;
assign LUT_4[34770] = 32'b00000000000000001110001000001100;
assign LUT_4[34771] = 32'b00000000000000000111010100000100;
assign LUT_4[34772] = 32'b00000000000000001011101110000100;
assign LUT_4[34773] = 32'b00000000000000000100111001111100;
assign LUT_4[34774] = 32'b00000000000000001011001000101000;
assign LUT_4[34775] = 32'b00000000000000000100010100100000;
assign LUT_4[34776] = 32'b00000000000000000111111001111101;
assign LUT_4[34777] = 32'b00000000000000000001000101110101;
assign LUT_4[34778] = 32'b00000000000000000111010100100001;
assign LUT_4[34779] = 32'b00000000000000000000100000011001;
assign LUT_4[34780] = 32'b00000000000000000100111010011001;
assign LUT_4[34781] = 32'b11111111111111111110000110010001;
assign LUT_4[34782] = 32'b00000000000000000100010100111101;
assign LUT_4[34783] = 32'b11111111111111111101100000110101;
assign LUT_4[34784] = 32'b00000000000000001111010111000001;
assign LUT_4[34785] = 32'b00000000000000001000100010111001;
assign LUT_4[34786] = 32'b00000000000000001110110001100101;
assign LUT_4[34787] = 32'b00000000000000000111111101011101;
assign LUT_4[34788] = 32'b00000000000000001100010111011101;
assign LUT_4[34789] = 32'b00000000000000000101100011010101;
assign LUT_4[34790] = 32'b00000000000000001011110010000001;
assign LUT_4[34791] = 32'b00000000000000000100111101111001;
assign LUT_4[34792] = 32'b00000000000000001000100011010110;
assign LUT_4[34793] = 32'b00000000000000000001101111001110;
assign LUT_4[34794] = 32'b00000000000000000111111101111010;
assign LUT_4[34795] = 32'b00000000000000000001001001110010;
assign LUT_4[34796] = 32'b00000000000000000101100011110010;
assign LUT_4[34797] = 32'b11111111111111111110101111101010;
assign LUT_4[34798] = 32'b00000000000000000100111110010110;
assign LUT_4[34799] = 32'b11111111111111111110001010001110;
assign LUT_4[34800] = 32'b00000000000000001101001000101111;
assign LUT_4[34801] = 32'b00000000000000000110010100100111;
assign LUT_4[34802] = 32'b00000000000000001100100011010011;
assign LUT_4[34803] = 32'b00000000000000000101101111001011;
assign LUT_4[34804] = 32'b00000000000000001010001001001011;
assign LUT_4[34805] = 32'b00000000000000000011010101000011;
assign LUT_4[34806] = 32'b00000000000000001001100011101111;
assign LUT_4[34807] = 32'b00000000000000000010101111100111;
assign LUT_4[34808] = 32'b00000000000000000110010101000100;
assign LUT_4[34809] = 32'b11111111111111111111100000111100;
assign LUT_4[34810] = 32'b00000000000000000101101111101000;
assign LUT_4[34811] = 32'b11111111111111111110111011100000;
assign LUT_4[34812] = 32'b00000000000000000011010101100000;
assign LUT_4[34813] = 32'b11111111111111111100100001011000;
assign LUT_4[34814] = 32'b00000000000000000010110000000100;
assign LUT_4[34815] = 32'b11111111111111111011111011111100;
assign LUT_4[34816] = 32'b00000000000000000010110011011110;
assign LUT_4[34817] = 32'b11111111111111111011111111010110;
assign LUT_4[34818] = 32'b00000000000000000010001110000010;
assign LUT_4[34819] = 32'b11111111111111111011011001111010;
assign LUT_4[34820] = 32'b11111111111111111111110011111010;
assign LUT_4[34821] = 32'b11111111111111111000111111110010;
assign LUT_4[34822] = 32'b11111111111111111111001110011110;
assign LUT_4[34823] = 32'b11111111111111111000011010010110;
assign LUT_4[34824] = 32'b11111111111111111011111111110011;
assign LUT_4[34825] = 32'b11111111111111110101001011101011;
assign LUT_4[34826] = 32'b11111111111111111011011010010111;
assign LUT_4[34827] = 32'b11111111111111110100100110001111;
assign LUT_4[34828] = 32'b11111111111111111001000000001111;
assign LUT_4[34829] = 32'b11111111111111110010001100000111;
assign LUT_4[34830] = 32'b11111111111111111000011010110011;
assign LUT_4[34831] = 32'b11111111111111110001100110101011;
assign LUT_4[34832] = 32'b00000000000000000000100101001100;
assign LUT_4[34833] = 32'b11111111111111111001110001000100;
assign LUT_4[34834] = 32'b11111111111111111111111111110000;
assign LUT_4[34835] = 32'b11111111111111111001001011101000;
assign LUT_4[34836] = 32'b11111111111111111101100101101000;
assign LUT_4[34837] = 32'b11111111111111110110110001100000;
assign LUT_4[34838] = 32'b11111111111111111101000000001100;
assign LUT_4[34839] = 32'b11111111111111110110001100000100;
assign LUT_4[34840] = 32'b11111111111111111001110001100001;
assign LUT_4[34841] = 32'b11111111111111110010111101011001;
assign LUT_4[34842] = 32'b11111111111111111001001100000101;
assign LUT_4[34843] = 32'b11111111111111110010010111111101;
assign LUT_4[34844] = 32'b11111111111111110110110001111101;
assign LUT_4[34845] = 32'b11111111111111101111111101110101;
assign LUT_4[34846] = 32'b11111111111111110110001100100001;
assign LUT_4[34847] = 32'b11111111111111101111011000011001;
assign LUT_4[34848] = 32'b00000000000000000001001110100101;
assign LUT_4[34849] = 32'b11111111111111111010011010011101;
assign LUT_4[34850] = 32'b00000000000000000000101001001001;
assign LUT_4[34851] = 32'b11111111111111111001110101000001;
assign LUT_4[34852] = 32'b11111111111111111110001111000001;
assign LUT_4[34853] = 32'b11111111111111110111011010111001;
assign LUT_4[34854] = 32'b11111111111111111101101001100101;
assign LUT_4[34855] = 32'b11111111111111110110110101011101;
assign LUT_4[34856] = 32'b11111111111111111010011010111010;
assign LUT_4[34857] = 32'b11111111111111110011100110110010;
assign LUT_4[34858] = 32'b11111111111111111001110101011110;
assign LUT_4[34859] = 32'b11111111111111110011000001010110;
assign LUT_4[34860] = 32'b11111111111111110111011011010110;
assign LUT_4[34861] = 32'b11111111111111110000100111001110;
assign LUT_4[34862] = 32'b11111111111111110110110101111010;
assign LUT_4[34863] = 32'b11111111111111110000000001110010;
assign LUT_4[34864] = 32'b11111111111111111111000000010011;
assign LUT_4[34865] = 32'b11111111111111111000001100001011;
assign LUT_4[34866] = 32'b11111111111111111110011010110111;
assign LUT_4[34867] = 32'b11111111111111110111100110101111;
assign LUT_4[34868] = 32'b11111111111111111100000000101111;
assign LUT_4[34869] = 32'b11111111111111110101001100100111;
assign LUT_4[34870] = 32'b11111111111111111011011011010011;
assign LUT_4[34871] = 32'b11111111111111110100100111001011;
assign LUT_4[34872] = 32'b11111111111111111000001100101000;
assign LUT_4[34873] = 32'b11111111111111110001011000100000;
assign LUT_4[34874] = 32'b11111111111111110111100111001100;
assign LUT_4[34875] = 32'b11111111111111110000110011000100;
assign LUT_4[34876] = 32'b11111111111111110101001101000100;
assign LUT_4[34877] = 32'b11111111111111101110011000111100;
assign LUT_4[34878] = 32'b11111111111111110100100111101000;
assign LUT_4[34879] = 32'b11111111111111101101110011100000;
assign LUT_4[34880] = 32'b00000000000000000100001010110010;
assign LUT_4[34881] = 32'b11111111111111111101010110101010;
assign LUT_4[34882] = 32'b00000000000000000011100101010110;
assign LUT_4[34883] = 32'b11111111111111111100110001001110;
assign LUT_4[34884] = 32'b00000000000000000001001011001110;
assign LUT_4[34885] = 32'b11111111111111111010010111000110;
assign LUT_4[34886] = 32'b00000000000000000000100101110010;
assign LUT_4[34887] = 32'b11111111111111111001110001101010;
assign LUT_4[34888] = 32'b11111111111111111101010111000111;
assign LUT_4[34889] = 32'b11111111111111110110100010111111;
assign LUT_4[34890] = 32'b11111111111111111100110001101011;
assign LUT_4[34891] = 32'b11111111111111110101111101100011;
assign LUT_4[34892] = 32'b11111111111111111010010111100011;
assign LUT_4[34893] = 32'b11111111111111110011100011011011;
assign LUT_4[34894] = 32'b11111111111111111001110010000111;
assign LUT_4[34895] = 32'b11111111111111110010111101111111;
assign LUT_4[34896] = 32'b00000000000000000001111100100000;
assign LUT_4[34897] = 32'b11111111111111111011001000011000;
assign LUT_4[34898] = 32'b00000000000000000001010111000100;
assign LUT_4[34899] = 32'b11111111111111111010100010111100;
assign LUT_4[34900] = 32'b11111111111111111110111100111100;
assign LUT_4[34901] = 32'b11111111111111111000001000110100;
assign LUT_4[34902] = 32'b11111111111111111110010111100000;
assign LUT_4[34903] = 32'b11111111111111110111100011011000;
assign LUT_4[34904] = 32'b11111111111111111011001000110101;
assign LUT_4[34905] = 32'b11111111111111110100010100101101;
assign LUT_4[34906] = 32'b11111111111111111010100011011001;
assign LUT_4[34907] = 32'b11111111111111110011101111010001;
assign LUT_4[34908] = 32'b11111111111111111000001001010001;
assign LUT_4[34909] = 32'b11111111111111110001010101001001;
assign LUT_4[34910] = 32'b11111111111111110111100011110101;
assign LUT_4[34911] = 32'b11111111111111110000101111101101;
assign LUT_4[34912] = 32'b00000000000000000010100101111001;
assign LUT_4[34913] = 32'b11111111111111111011110001110001;
assign LUT_4[34914] = 32'b00000000000000000010000000011101;
assign LUT_4[34915] = 32'b11111111111111111011001100010101;
assign LUT_4[34916] = 32'b11111111111111111111100110010101;
assign LUT_4[34917] = 32'b11111111111111111000110010001101;
assign LUT_4[34918] = 32'b11111111111111111111000000111001;
assign LUT_4[34919] = 32'b11111111111111111000001100110001;
assign LUT_4[34920] = 32'b11111111111111111011110010001110;
assign LUT_4[34921] = 32'b11111111111111110100111110000110;
assign LUT_4[34922] = 32'b11111111111111111011001100110010;
assign LUT_4[34923] = 32'b11111111111111110100011000101010;
assign LUT_4[34924] = 32'b11111111111111111000110010101010;
assign LUT_4[34925] = 32'b11111111111111110001111110100010;
assign LUT_4[34926] = 32'b11111111111111111000001101001110;
assign LUT_4[34927] = 32'b11111111111111110001011001000110;
assign LUT_4[34928] = 32'b00000000000000000000010111100111;
assign LUT_4[34929] = 32'b11111111111111111001100011011111;
assign LUT_4[34930] = 32'b11111111111111111111110010001011;
assign LUT_4[34931] = 32'b11111111111111111000111110000011;
assign LUT_4[34932] = 32'b11111111111111111101011000000011;
assign LUT_4[34933] = 32'b11111111111111110110100011111011;
assign LUT_4[34934] = 32'b11111111111111111100110010100111;
assign LUT_4[34935] = 32'b11111111111111110101111110011111;
assign LUT_4[34936] = 32'b11111111111111111001100011111100;
assign LUT_4[34937] = 32'b11111111111111110010101111110100;
assign LUT_4[34938] = 32'b11111111111111111000111110100000;
assign LUT_4[34939] = 32'b11111111111111110010001010011000;
assign LUT_4[34940] = 32'b11111111111111110110100100011000;
assign LUT_4[34941] = 32'b11111111111111101111110000010000;
assign LUT_4[34942] = 32'b11111111111111110101111110111100;
assign LUT_4[34943] = 32'b11111111111111101111001010110100;
assign LUT_4[34944] = 32'b00000000000000000101011001100110;
assign LUT_4[34945] = 32'b11111111111111111110100101011110;
assign LUT_4[34946] = 32'b00000000000000000100110100001010;
assign LUT_4[34947] = 32'b11111111111111111110000000000010;
assign LUT_4[34948] = 32'b00000000000000000010011010000010;
assign LUT_4[34949] = 32'b11111111111111111011100101111010;
assign LUT_4[34950] = 32'b00000000000000000001110100100110;
assign LUT_4[34951] = 32'b11111111111111111011000000011110;
assign LUT_4[34952] = 32'b11111111111111111110100101111011;
assign LUT_4[34953] = 32'b11111111111111110111110001110011;
assign LUT_4[34954] = 32'b11111111111111111110000000011111;
assign LUT_4[34955] = 32'b11111111111111110111001100010111;
assign LUT_4[34956] = 32'b11111111111111111011100110010111;
assign LUT_4[34957] = 32'b11111111111111110100110010001111;
assign LUT_4[34958] = 32'b11111111111111111011000000111011;
assign LUT_4[34959] = 32'b11111111111111110100001100110011;
assign LUT_4[34960] = 32'b00000000000000000011001011010100;
assign LUT_4[34961] = 32'b11111111111111111100010111001100;
assign LUT_4[34962] = 32'b00000000000000000010100101111000;
assign LUT_4[34963] = 32'b11111111111111111011110001110000;
assign LUT_4[34964] = 32'b00000000000000000000001011110000;
assign LUT_4[34965] = 32'b11111111111111111001010111101000;
assign LUT_4[34966] = 32'b11111111111111111111100110010100;
assign LUT_4[34967] = 32'b11111111111111111000110010001100;
assign LUT_4[34968] = 32'b11111111111111111100010111101001;
assign LUT_4[34969] = 32'b11111111111111110101100011100001;
assign LUT_4[34970] = 32'b11111111111111111011110010001101;
assign LUT_4[34971] = 32'b11111111111111110100111110000101;
assign LUT_4[34972] = 32'b11111111111111111001011000000101;
assign LUT_4[34973] = 32'b11111111111111110010100011111101;
assign LUT_4[34974] = 32'b11111111111111111000110010101001;
assign LUT_4[34975] = 32'b11111111111111110001111110100001;
assign LUT_4[34976] = 32'b00000000000000000011110100101101;
assign LUT_4[34977] = 32'b11111111111111111101000000100101;
assign LUT_4[34978] = 32'b00000000000000000011001111010001;
assign LUT_4[34979] = 32'b11111111111111111100011011001001;
assign LUT_4[34980] = 32'b00000000000000000000110101001001;
assign LUT_4[34981] = 32'b11111111111111111010000001000001;
assign LUT_4[34982] = 32'b00000000000000000000001111101101;
assign LUT_4[34983] = 32'b11111111111111111001011011100101;
assign LUT_4[34984] = 32'b11111111111111111101000001000010;
assign LUT_4[34985] = 32'b11111111111111110110001100111010;
assign LUT_4[34986] = 32'b11111111111111111100011011100110;
assign LUT_4[34987] = 32'b11111111111111110101100111011110;
assign LUT_4[34988] = 32'b11111111111111111010000001011110;
assign LUT_4[34989] = 32'b11111111111111110011001101010110;
assign LUT_4[34990] = 32'b11111111111111111001011100000010;
assign LUT_4[34991] = 32'b11111111111111110010100111111010;
assign LUT_4[34992] = 32'b00000000000000000001100110011011;
assign LUT_4[34993] = 32'b11111111111111111010110010010011;
assign LUT_4[34994] = 32'b00000000000000000001000000111111;
assign LUT_4[34995] = 32'b11111111111111111010001100110111;
assign LUT_4[34996] = 32'b11111111111111111110100110110111;
assign LUT_4[34997] = 32'b11111111111111110111110010101111;
assign LUT_4[34998] = 32'b11111111111111111110000001011011;
assign LUT_4[34999] = 32'b11111111111111110111001101010011;
assign LUT_4[35000] = 32'b11111111111111111010110010110000;
assign LUT_4[35001] = 32'b11111111111111110011111110101000;
assign LUT_4[35002] = 32'b11111111111111111010001101010100;
assign LUT_4[35003] = 32'b11111111111111110011011001001100;
assign LUT_4[35004] = 32'b11111111111111110111110011001100;
assign LUT_4[35005] = 32'b11111111111111110000111111000100;
assign LUT_4[35006] = 32'b11111111111111110111001101110000;
assign LUT_4[35007] = 32'b11111111111111110000011001101000;
assign LUT_4[35008] = 32'b00000000000000000110110000111010;
assign LUT_4[35009] = 32'b11111111111111111111111100110010;
assign LUT_4[35010] = 32'b00000000000000000110001011011110;
assign LUT_4[35011] = 32'b11111111111111111111010111010110;
assign LUT_4[35012] = 32'b00000000000000000011110001010110;
assign LUT_4[35013] = 32'b11111111111111111100111101001110;
assign LUT_4[35014] = 32'b00000000000000000011001011111010;
assign LUT_4[35015] = 32'b11111111111111111100010111110010;
assign LUT_4[35016] = 32'b11111111111111111111111101001111;
assign LUT_4[35017] = 32'b11111111111111111001001001000111;
assign LUT_4[35018] = 32'b11111111111111111111010111110011;
assign LUT_4[35019] = 32'b11111111111111111000100011101011;
assign LUT_4[35020] = 32'b11111111111111111100111101101011;
assign LUT_4[35021] = 32'b11111111111111110110001001100011;
assign LUT_4[35022] = 32'b11111111111111111100011000001111;
assign LUT_4[35023] = 32'b11111111111111110101100100000111;
assign LUT_4[35024] = 32'b00000000000000000100100010101000;
assign LUT_4[35025] = 32'b11111111111111111101101110100000;
assign LUT_4[35026] = 32'b00000000000000000011111101001100;
assign LUT_4[35027] = 32'b11111111111111111101001001000100;
assign LUT_4[35028] = 32'b00000000000000000001100011000100;
assign LUT_4[35029] = 32'b11111111111111111010101110111100;
assign LUT_4[35030] = 32'b00000000000000000000111101101000;
assign LUT_4[35031] = 32'b11111111111111111010001001100000;
assign LUT_4[35032] = 32'b11111111111111111101101110111101;
assign LUT_4[35033] = 32'b11111111111111110110111010110101;
assign LUT_4[35034] = 32'b11111111111111111101001001100001;
assign LUT_4[35035] = 32'b11111111111111110110010101011001;
assign LUT_4[35036] = 32'b11111111111111111010101111011001;
assign LUT_4[35037] = 32'b11111111111111110011111011010001;
assign LUT_4[35038] = 32'b11111111111111111010001001111101;
assign LUT_4[35039] = 32'b11111111111111110011010101110101;
assign LUT_4[35040] = 32'b00000000000000000101001100000001;
assign LUT_4[35041] = 32'b11111111111111111110010111111001;
assign LUT_4[35042] = 32'b00000000000000000100100110100101;
assign LUT_4[35043] = 32'b11111111111111111101110010011101;
assign LUT_4[35044] = 32'b00000000000000000010001100011101;
assign LUT_4[35045] = 32'b11111111111111111011011000010101;
assign LUT_4[35046] = 32'b00000000000000000001100111000001;
assign LUT_4[35047] = 32'b11111111111111111010110010111001;
assign LUT_4[35048] = 32'b11111111111111111110011000010110;
assign LUT_4[35049] = 32'b11111111111111110111100100001110;
assign LUT_4[35050] = 32'b11111111111111111101110010111010;
assign LUT_4[35051] = 32'b11111111111111110110111110110010;
assign LUT_4[35052] = 32'b11111111111111111011011000110010;
assign LUT_4[35053] = 32'b11111111111111110100100100101010;
assign LUT_4[35054] = 32'b11111111111111111010110011010110;
assign LUT_4[35055] = 32'b11111111111111110011111111001110;
assign LUT_4[35056] = 32'b00000000000000000010111101101111;
assign LUT_4[35057] = 32'b11111111111111111100001001100111;
assign LUT_4[35058] = 32'b00000000000000000010011000010011;
assign LUT_4[35059] = 32'b11111111111111111011100100001011;
assign LUT_4[35060] = 32'b11111111111111111111111110001011;
assign LUT_4[35061] = 32'b11111111111111111001001010000011;
assign LUT_4[35062] = 32'b11111111111111111111011000101111;
assign LUT_4[35063] = 32'b11111111111111111000100100100111;
assign LUT_4[35064] = 32'b11111111111111111100001010000100;
assign LUT_4[35065] = 32'b11111111111111110101010101111100;
assign LUT_4[35066] = 32'b11111111111111111011100100101000;
assign LUT_4[35067] = 32'b11111111111111110100110000100000;
assign LUT_4[35068] = 32'b11111111111111111001001010100000;
assign LUT_4[35069] = 32'b11111111111111110010010110011000;
assign LUT_4[35070] = 32'b11111111111111111000100101000100;
assign LUT_4[35071] = 32'b11111111111111110001110000111100;
assign LUT_4[35072] = 32'b00000000000000000111101111000001;
assign LUT_4[35073] = 32'b00000000000000000000111010111001;
assign LUT_4[35074] = 32'b00000000000000000111001001100101;
assign LUT_4[35075] = 32'b00000000000000000000010101011101;
assign LUT_4[35076] = 32'b00000000000000000100101111011101;
assign LUT_4[35077] = 32'b11111111111111111101111011010101;
assign LUT_4[35078] = 32'b00000000000000000100001010000001;
assign LUT_4[35079] = 32'b11111111111111111101010101111001;
assign LUT_4[35080] = 32'b00000000000000000000111011010110;
assign LUT_4[35081] = 32'b11111111111111111010000111001110;
assign LUT_4[35082] = 32'b00000000000000000000010101111010;
assign LUT_4[35083] = 32'b11111111111111111001100001110010;
assign LUT_4[35084] = 32'b11111111111111111101111011110010;
assign LUT_4[35085] = 32'b11111111111111110111000111101010;
assign LUT_4[35086] = 32'b11111111111111111101010110010110;
assign LUT_4[35087] = 32'b11111111111111110110100010001110;
assign LUT_4[35088] = 32'b00000000000000000101100000101111;
assign LUT_4[35089] = 32'b11111111111111111110101100100111;
assign LUT_4[35090] = 32'b00000000000000000100111011010011;
assign LUT_4[35091] = 32'b11111111111111111110000111001011;
assign LUT_4[35092] = 32'b00000000000000000010100001001011;
assign LUT_4[35093] = 32'b11111111111111111011101101000011;
assign LUT_4[35094] = 32'b00000000000000000001111011101111;
assign LUT_4[35095] = 32'b11111111111111111011000111100111;
assign LUT_4[35096] = 32'b11111111111111111110101101000100;
assign LUT_4[35097] = 32'b11111111111111110111111000111100;
assign LUT_4[35098] = 32'b11111111111111111110000111101000;
assign LUT_4[35099] = 32'b11111111111111110111010011100000;
assign LUT_4[35100] = 32'b11111111111111111011101101100000;
assign LUT_4[35101] = 32'b11111111111111110100111001011000;
assign LUT_4[35102] = 32'b11111111111111111011001000000100;
assign LUT_4[35103] = 32'b11111111111111110100010011111100;
assign LUT_4[35104] = 32'b00000000000000000110001010001000;
assign LUT_4[35105] = 32'b11111111111111111111010110000000;
assign LUT_4[35106] = 32'b00000000000000000101100100101100;
assign LUT_4[35107] = 32'b11111111111111111110110000100100;
assign LUT_4[35108] = 32'b00000000000000000011001010100100;
assign LUT_4[35109] = 32'b11111111111111111100010110011100;
assign LUT_4[35110] = 32'b00000000000000000010100101001000;
assign LUT_4[35111] = 32'b11111111111111111011110001000000;
assign LUT_4[35112] = 32'b11111111111111111111010110011101;
assign LUT_4[35113] = 32'b11111111111111111000100010010101;
assign LUT_4[35114] = 32'b11111111111111111110110001000001;
assign LUT_4[35115] = 32'b11111111111111110111111100111001;
assign LUT_4[35116] = 32'b11111111111111111100010110111001;
assign LUT_4[35117] = 32'b11111111111111110101100010110001;
assign LUT_4[35118] = 32'b11111111111111111011110001011101;
assign LUT_4[35119] = 32'b11111111111111110100111101010101;
assign LUT_4[35120] = 32'b00000000000000000011111011110110;
assign LUT_4[35121] = 32'b11111111111111111101000111101110;
assign LUT_4[35122] = 32'b00000000000000000011010110011010;
assign LUT_4[35123] = 32'b11111111111111111100100010010010;
assign LUT_4[35124] = 32'b00000000000000000000111100010010;
assign LUT_4[35125] = 32'b11111111111111111010001000001010;
assign LUT_4[35126] = 32'b00000000000000000000010110110110;
assign LUT_4[35127] = 32'b11111111111111111001100010101110;
assign LUT_4[35128] = 32'b11111111111111111101001000001011;
assign LUT_4[35129] = 32'b11111111111111110110010100000011;
assign LUT_4[35130] = 32'b11111111111111111100100010101111;
assign LUT_4[35131] = 32'b11111111111111110101101110100111;
assign LUT_4[35132] = 32'b11111111111111111010001000100111;
assign LUT_4[35133] = 32'b11111111111111110011010100011111;
assign LUT_4[35134] = 32'b11111111111111111001100011001011;
assign LUT_4[35135] = 32'b11111111111111110010101111000011;
assign LUT_4[35136] = 32'b00000000000000001001000110010101;
assign LUT_4[35137] = 32'b00000000000000000010010010001101;
assign LUT_4[35138] = 32'b00000000000000001000100000111001;
assign LUT_4[35139] = 32'b00000000000000000001101100110001;
assign LUT_4[35140] = 32'b00000000000000000110000110110001;
assign LUT_4[35141] = 32'b11111111111111111111010010101001;
assign LUT_4[35142] = 32'b00000000000000000101100001010101;
assign LUT_4[35143] = 32'b11111111111111111110101101001101;
assign LUT_4[35144] = 32'b00000000000000000010010010101010;
assign LUT_4[35145] = 32'b11111111111111111011011110100010;
assign LUT_4[35146] = 32'b00000000000000000001101101001110;
assign LUT_4[35147] = 32'b11111111111111111010111001000110;
assign LUT_4[35148] = 32'b11111111111111111111010011000110;
assign LUT_4[35149] = 32'b11111111111111111000011110111110;
assign LUT_4[35150] = 32'b11111111111111111110101101101010;
assign LUT_4[35151] = 32'b11111111111111110111111001100010;
assign LUT_4[35152] = 32'b00000000000000000110111000000011;
assign LUT_4[35153] = 32'b00000000000000000000000011111011;
assign LUT_4[35154] = 32'b00000000000000000110010010100111;
assign LUT_4[35155] = 32'b11111111111111111111011110011111;
assign LUT_4[35156] = 32'b00000000000000000011111000011111;
assign LUT_4[35157] = 32'b11111111111111111101000100010111;
assign LUT_4[35158] = 32'b00000000000000000011010011000011;
assign LUT_4[35159] = 32'b11111111111111111100011110111011;
assign LUT_4[35160] = 32'b00000000000000000000000100011000;
assign LUT_4[35161] = 32'b11111111111111111001010000010000;
assign LUT_4[35162] = 32'b11111111111111111111011110111100;
assign LUT_4[35163] = 32'b11111111111111111000101010110100;
assign LUT_4[35164] = 32'b11111111111111111101000100110100;
assign LUT_4[35165] = 32'b11111111111111110110010000101100;
assign LUT_4[35166] = 32'b11111111111111111100011111011000;
assign LUT_4[35167] = 32'b11111111111111110101101011010000;
assign LUT_4[35168] = 32'b00000000000000000111100001011100;
assign LUT_4[35169] = 32'b00000000000000000000101101010100;
assign LUT_4[35170] = 32'b00000000000000000110111100000000;
assign LUT_4[35171] = 32'b00000000000000000000000111111000;
assign LUT_4[35172] = 32'b00000000000000000100100001111000;
assign LUT_4[35173] = 32'b11111111111111111101101101110000;
assign LUT_4[35174] = 32'b00000000000000000011111100011100;
assign LUT_4[35175] = 32'b11111111111111111101001000010100;
assign LUT_4[35176] = 32'b00000000000000000000101101110001;
assign LUT_4[35177] = 32'b11111111111111111001111001101001;
assign LUT_4[35178] = 32'b00000000000000000000001000010101;
assign LUT_4[35179] = 32'b11111111111111111001010100001101;
assign LUT_4[35180] = 32'b11111111111111111101101110001101;
assign LUT_4[35181] = 32'b11111111111111110110111010000101;
assign LUT_4[35182] = 32'b11111111111111111101001000110001;
assign LUT_4[35183] = 32'b11111111111111110110010100101001;
assign LUT_4[35184] = 32'b00000000000000000101010011001010;
assign LUT_4[35185] = 32'b11111111111111111110011111000010;
assign LUT_4[35186] = 32'b00000000000000000100101101101110;
assign LUT_4[35187] = 32'b11111111111111111101111001100110;
assign LUT_4[35188] = 32'b00000000000000000010010011100110;
assign LUT_4[35189] = 32'b11111111111111111011011111011110;
assign LUT_4[35190] = 32'b00000000000000000001101110001010;
assign LUT_4[35191] = 32'b11111111111111111010111010000010;
assign LUT_4[35192] = 32'b11111111111111111110011111011111;
assign LUT_4[35193] = 32'b11111111111111110111101011010111;
assign LUT_4[35194] = 32'b11111111111111111101111010000011;
assign LUT_4[35195] = 32'b11111111111111110111000101111011;
assign LUT_4[35196] = 32'b11111111111111111011011111111011;
assign LUT_4[35197] = 32'b11111111111111110100101011110011;
assign LUT_4[35198] = 32'b11111111111111111010111010011111;
assign LUT_4[35199] = 32'b11111111111111110100000110010111;
assign LUT_4[35200] = 32'b00000000000000001010010101001001;
assign LUT_4[35201] = 32'b00000000000000000011100001000001;
assign LUT_4[35202] = 32'b00000000000000001001101111101101;
assign LUT_4[35203] = 32'b00000000000000000010111011100101;
assign LUT_4[35204] = 32'b00000000000000000111010101100101;
assign LUT_4[35205] = 32'b00000000000000000000100001011101;
assign LUT_4[35206] = 32'b00000000000000000110110000001001;
assign LUT_4[35207] = 32'b11111111111111111111111100000001;
assign LUT_4[35208] = 32'b00000000000000000011100001011110;
assign LUT_4[35209] = 32'b11111111111111111100101101010110;
assign LUT_4[35210] = 32'b00000000000000000010111100000010;
assign LUT_4[35211] = 32'b11111111111111111100000111111010;
assign LUT_4[35212] = 32'b00000000000000000000100001111010;
assign LUT_4[35213] = 32'b11111111111111111001101101110010;
assign LUT_4[35214] = 32'b11111111111111111111111100011110;
assign LUT_4[35215] = 32'b11111111111111111001001000010110;
assign LUT_4[35216] = 32'b00000000000000001000000110110111;
assign LUT_4[35217] = 32'b00000000000000000001010010101111;
assign LUT_4[35218] = 32'b00000000000000000111100001011011;
assign LUT_4[35219] = 32'b00000000000000000000101101010011;
assign LUT_4[35220] = 32'b00000000000000000101000111010011;
assign LUT_4[35221] = 32'b11111111111111111110010011001011;
assign LUT_4[35222] = 32'b00000000000000000100100001110111;
assign LUT_4[35223] = 32'b11111111111111111101101101101111;
assign LUT_4[35224] = 32'b00000000000000000001010011001100;
assign LUT_4[35225] = 32'b11111111111111111010011111000100;
assign LUT_4[35226] = 32'b00000000000000000000101101110000;
assign LUT_4[35227] = 32'b11111111111111111001111001101000;
assign LUT_4[35228] = 32'b11111111111111111110010011101000;
assign LUT_4[35229] = 32'b11111111111111110111011111100000;
assign LUT_4[35230] = 32'b11111111111111111101101110001100;
assign LUT_4[35231] = 32'b11111111111111110110111010000100;
assign LUT_4[35232] = 32'b00000000000000001000110000010000;
assign LUT_4[35233] = 32'b00000000000000000001111100001000;
assign LUT_4[35234] = 32'b00000000000000001000001010110100;
assign LUT_4[35235] = 32'b00000000000000000001010110101100;
assign LUT_4[35236] = 32'b00000000000000000101110000101100;
assign LUT_4[35237] = 32'b11111111111111111110111100100100;
assign LUT_4[35238] = 32'b00000000000000000101001011010000;
assign LUT_4[35239] = 32'b11111111111111111110010111001000;
assign LUT_4[35240] = 32'b00000000000000000001111100100101;
assign LUT_4[35241] = 32'b11111111111111111011001000011101;
assign LUT_4[35242] = 32'b00000000000000000001010111001001;
assign LUT_4[35243] = 32'b11111111111111111010100011000001;
assign LUT_4[35244] = 32'b11111111111111111110111101000001;
assign LUT_4[35245] = 32'b11111111111111111000001000111001;
assign LUT_4[35246] = 32'b11111111111111111110010111100101;
assign LUT_4[35247] = 32'b11111111111111110111100011011101;
assign LUT_4[35248] = 32'b00000000000000000110100001111110;
assign LUT_4[35249] = 32'b11111111111111111111101101110110;
assign LUT_4[35250] = 32'b00000000000000000101111100100010;
assign LUT_4[35251] = 32'b11111111111111111111001000011010;
assign LUT_4[35252] = 32'b00000000000000000011100010011010;
assign LUT_4[35253] = 32'b11111111111111111100101110010010;
assign LUT_4[35254] = 32'b00000000000000000010111100111110;
assign LUT_4[35255] = 32'b11111111111111111100001000110110;
assign LUT_4[35256] = 32'b11111111111111111111101110010011;
assign LUT_4[35257] = 32'b11111111111111111000111010001011;
assign LUT_4[35258] = 32'b11111111111111111111001000110111;
assign LUT_4[35259] = 32'b11111111111111111000010100101111;
assign LUT_4[35260] = 32'b11111111111111111100101110101111;
assign LUT_4[35261] = 32'b11111111111111110101111010100111;
assign LUT_4[35262] = 32'b11111111111111111100001001010011;
assign LUT_4[35263] = 32'b11111111111111110101010101001011;
assign LUT_4[35264] = 32'b00000000000000001011101100011101;
assign LUT_4[35265] = 32'b00000000000000000100111000010101;
assign LUT_4[35266] = 32'b00000000000000001011000111000001;
assign LUT_4[35267] = 32'b00000000000000000100010010111001;
assign LUT_4[35268] = 32'b00000000000000001000101100111001;
assign LUT_4[35269] = 32'b00000000000000000001111000110001;
assign LUT_4[35270] = 32'b00000000000000001000000111011101;
assign LUT_4[35271] = 32'b00000000000000000001010011010101;
assign LUT_4[35272] = 32'b00000000000000000100111000110010;
assign LUT_4[35273] = 32'b11111111111111111110000100101010;
assign LUT_4[35274] = 32'b00000000000000000100010011010110;
assign LUT_4[35275] = 32'b11111111111111111101011111001110;
assign LUT_4[35276] = 32'b00000000000000000001111001001110;
assign LUT_4[35277] = 32'b11111111111111111011000101000110;
assign LUT_4[35278] = 32'b00000000000000000001010011110010;
assign LUT_4[35279] = 32'b11111111111111111010011111101010;
assign LUT_4[35280] = 32'b00000000000000001001011110001011;
assign LUT_4[35281] = 32'b00000000000000000010101010000011;
assign LUT_4[35282] = 32'b00000000000000001000111000101111;
assign LUT_4[35283] = 32'b00000000000000000010000100100111;
assign LUT_4[35284] = 32'b00000000000000000110011110100111;
assign LUT_4[35285] = 32'b11111111111111111111101010011111;
assign LUT_4[35286] = 32'b00000000000000000101111001001011;
assign LUT_4[35287] = 32'b11111111111111111111000101000011;
assign LUT_4[35288] = 32'b00000000000000000010101010100000;
assign LUT_4[35289] = 32'b11111111111111111011110110011000;
assign LUT_4[35290] = 32'b00000000000000000010000101000100;
assign LUT_4[35291] = 32'b11111111111111111011010000111100;
assign LUT_4[35292] = 32'b11111111111111111111101010111100;
assign LUT_4[35293] = 32'b11111111111111111000110110110100;
assign LUT_4[35294] = 32'b11111111111111111111000101100000;
assign LUT_4[35295] = 32'b11111111111111111000010001011000;
assign LUT_4[35296] = 32'b00000000000000001010000111100100;
assign LUT_4[35297] = 32'b00000000000000000011010011011100;
assign LUT_4[35298] = 32'b00000000000000001001100010001000;
assign LUT_4[35299] = 32'b00000000000000000010101110000000;
assign LUT_4[35300] = 32'b00000000000000000111001000000000;
assign LUT_4[35301] = 32'b00000000000000000000010011111000;
assign LUT_4[35302] = 32'b00000000000000000110100010100100;
assign LUT_4[35303] = 32'b11111111111111111111101110011100;
assign LUT_4[35304] = 32'b00000000000000000011010011111001;
assign LUT_4[35305] = 32'b11111111111111111100011111110001;
assign LUT_4[35306] = 32'b00000000000000000010101110011101;
assign LUT_4[35307] = 32'b11111111111111111011111010010101;
assign LUT_4[35308] = 32'b00000000000000000000010100010101;
assign LUT_4[35309] = 32'b11111111111111111001100000001101;
assign LUT_4[35310] = 32'b11111111111111111111101110111001;
assign LUT_4[35311] = 32'b11111111111111111000111010110001;
assign LUT_4[35312] = 32'b00000000000000000111111001010010;
assign LUT_4[35313] = 32'b00000000000000000001000101001010;
assign LUT_4[35314] = 32'b00000000000000000111010011110110;
assign LUT_4[35315] = 32'b00000000000000000000011111101110;
assign LUT_4[35316] = 32'b00000000000000000100111001101110;
assign LUT_4[35317] = 32'b11111111111111111110000101100110;
assign LUT_4[35318] = 32'b00000000000000000100010100010010;
assign LUT_4[35319] = 32'b11111111111111111101100000001010;
assign LUT_4[35320] = 32'b00000000000000000001000101100111;
assign LUT_4[35321] = 32'b11111111111111111010010001011111;
assign LUT_4[35322] = 32'b00000000000000000000100000001011;
assign LUT_4[35323] = 32'b11111111111111111001101100000011;
assign LUT_4[35324] = 32'b11111111111111111110000110000011;
assign LUT_4[35325] = 32'b11111111111111110111010001111011;
assign LUT_4[35326] = 32'b11111111111111111101100000100111;
assign LUT_4[35327] = 32'b11111111111111110110101100011111;
assign LUT_4[35328] = 32'b00000000000000000001110111100110;
assign LUT_4[35329] = 32'b11111111111111111011000011011110;
assign LUT_4[35330] = 32'b00000000000000000001010010001010;
assign LUT_4[35331] = 32'b11111111111111111010011110000010;
assign LUT_4[35332] = 32'b11111111111111111110111000000010;
assign LUT_4[35333] = 32'b11111111111111111000000011111010;
assign LUT_4[35334] = 32'b11111111111111111110010010100110;
assign LUT_4[35335] = 32'b11111111111111110111011110011110;
assign LUT_4[35336] = 32'b11111111111111111011000011111011;
assign LUT_4[35337] = 32'b11111111111111110100001111110011;
assign LUT_4[35338] = 32'b11111111111111111010011110011111;
assign LUT_4[35339] = 32'b11111111111111110011101010010111;
assign LUT_4[35340] = 32'b11111111111111111000000100010111;
assign LUT_4[35341] = 32'b11111111111111110001010000001111;
assign LUT_4[35342] = 32'b11111111111111110111011110111011;
assign LUT_4[35343] = 32'b11111111111111110000101010110011;
assign LUT_4[35344] = 32'b11111111111111111111101001010100;
assign LUT_4[35345] = 32'b11111111111111111000110101001100;
assign LUT_4[35346] = 32'b11111111111111111111000011111000;
assign LUT_4[35347] = 32'b11111111111111111000001111110000;
assign LUT_4[35348] = 32'b11111111111111111100101001110000;
assign LUT_4[35349] = 32'b11111111111111110101110101101000;
assign LUT_4[35350] = 32'b11111111111111111100000100010100;
assign LUT_4[35351] = 32'b11111111111111110101010000001100;
assign LUT_4[35352] = 32'b11111111111111111000110101101001;
assign LUT_4[35353] = 32'b11111111111111110010000001100001;
assign LUT_4[35354] = 32'b11111111111111111000010000001101;
assign LUT_4[35355] = 32'b11111111111111110001011100000101;
assign LUT_4[35356] = 32'b11111111111111110101110110000101;
assign LUT_4[35357] = 32'b11111111111111101111000001111101;
assign LUT_4[35358] = 32'b11111111111111110101010000101001;
assign LUT_4[35359] = 32'b11111111111111101110011100100001;
assign LUT_4[35360] = 32'b00000000000000000000010010101101;
assign LUT_4[35361] = 32'b11111111111111111001011110100101;
assign LUT_4[35362] = 32'b11111111111111111111101101010001;
assign LUT_4[35363] = 32'b11111111111111111000111001001001;
assign LUT_4[35364] = 32'b11111111111111111101010011001001;
assign LUT_4[35365] = 32'b11111111111111110110011111000001;
assign LUT_4[35366] = 32'b11111111111111111100101101101101;
assign LUT_4[35367] = 32'b11111111111111110101111001100101;
assign LUT_4[35368] = 32'b11111111111111111001011111000010;
assign LUT_4[35369] = 32'b11111111111111110010101010111010;
assign LUT_4[35370] = 32'b11111111111111111000111001100110;
assign LUT_4[35371] = 32'b11111111111111110010000101011110;
assign LUT_4[35372] = 32'b11111111111111110110011111011110;
assign LUT_4[35373] = 32'b11111111111111101111101011010110;
assign LUT_4[35374] = 32'b11111111111111110101111010000010;
assign LUT_4[35375] = 32'b11111111111111101111000101111010;
assign LUT_4[35376] = 32'b11111111111111111110000100011011;
assign LUT_4[35377] = 32'b11111111111111110111010000010011;
assign LUT_4[35378] = 32'b11111111111111111101011110111111;
assign LUT_4[35379] = 32'b11111111111111110110101010110111;
assign LUT_4[35380] = 32'b11111111111111111011000100110111;
assign LUT_4[35381] = 32'b11111111111111110100010000101111;
assign LUT_4[35382] = 32'b11111111111111111010011111011011;
assign LUT_4[35383] = 32'b11111111111111110011101011010011;
assign LUT_4[35384] = 32'b11111111111111110111010000110000;
assign LUT_4[35385] = 32'b11111111111111110000011100101000;
assign LUT_4[35386] = 32'b11111111111111110110101011010100;
assign LUT_4[35387] = 32'b11111111111111101111110111001100;
assign LUT_4[35388] = 32'b11111111111111110100010001001100;
assign LUT_4[35389] = 32'b11111111111111101101011101000100;
assign LUT_4[35390] = 32'b11111111111111110011101011110000;
assign LUT_4[35391] = 32'b11111111111111101100110111101000;
assign LUT_4[35392] = 32'b00000000000000000011001110111010;
assign LUT_4[35393] = 32'b11111111111111111100011010110010;
assign LUT_4[35394] = 32'b00000000000000000010101001011110;
assign LUT_4[35395] = 32'b11111111111111111011110101010110;
assign LUT_4[35396] = 32'b00000000000000000000001111010110;
assign LUT_4[35397] = 32'b11111111111111111001011011001110;
assign LUT_4[35398] = 32'b11111111111111111111101001111010;
assign LUT_4[35399] = 32'b11111111111111111000110101110010;
assign LUT_4[35400] = 32'b11111111111111111100011011001111;
assign LUT_4[35401] = 32'b11111111111111110101100111000111;
assign LUT_4[35402] = 32'b11111111111111111011110101110011;
assign LUT_4[35403] = 32'b11111111111111110101000001101011;
assign LUT_4[35404] = 32'b11111111111111111001011011101011;
assign LUT_4[35405] = 32'b11111111111111110010100111100011;
assign LUT_4[35406] = 32'b11111111111111111000110110001111;
assign LUT_4[35407] = 32'b11111111111111110010000010000111;
assign LUT_4[35408] = 32'b00000000000000000001000000101000;
assign LUT_4[35409] = 32'b11111111111111111010001100100000;
assign LUT_4[35410] = 32'b00000000000000000000011011001100;
assign LUT_4[35411] = 32'b11111111111111111001100111000100;
assign LUT_4[35412] = 32'b11111111111111111110000001000100;
assign LUT_4[35413] = 32'b11111111111111110111001100111100;
assign LUT_4[35414] = 32'b11111111111111111101011011101000;
assign LUT_4[35415] = 32'b11111111111111110110100111100000;
assign LUT_4[35416] = 32'b11111111111111111010001100111101;
assign LUT_4[35417] = 32'b11111111111111110011011000110101;
assign LUT_4[35418] = 32'b11111111111111111001100111100001;
assign LUT_4[35419] = 32'b11111111111111110010110011011001;
assign LUT_4[35420] = 32'b11111111111111110111001101011001;
assign LUT_4[35421] = 32'b11111111111111110000011001010001;
assign LUT_4[35422] = 32'b11111111111111110110100111111101;
assign LUT_4[35423] = 32'b11111111111111101111110011110101;
assign LUT_4[35424] = 32'b00000000000000000001101010000001;
assign LUT_4[35425] = 32'b11111111111111111010110101111001;
assign LUT_4[35426] = 32'b00000000000000000001000100100101;
assign LUT_4[35427] = 32'b11111111111111111010010000011101;
assign LUT_4[35428] = 32'b11111111111111111110101010011101;
assign LUT_4[35429] = 32'b11111111111111110111110110010101;
assign LUT_4[35430] = 32'b11111111111111111110000101000001;
assign LUT_4[35431] = 32'b11111111111111110111010000111001;
assign LUT_4[35432] = 32'b11111111111111111010110110010110;
assign LUT_4[35433] = 32'b11111111111111110100000010001110;
assign LUT_4[35434] = 32'b11111111111111111010010000111010;
assign LUT_4[35435] = 32'b11111111111111110011011100110010;
assign LUT_4[35436] = 32'b11111111111111110111110110110010;
assign LUT_4[35437] = 32'b11111111111111110001000010101010;
assign LUT_4[35438] = 32'b11111111111111110111010001010110;
assign LUT_4[35439] = 32'b11111111111111110000011101001110;
assign LUT_4[35440] = 32'b11111111111111111111011011101111;
assign LUT_4[35441] = 32'b11111111111111111000100111100111;
assign LUT_4[35442] = 32'b11111111111111111110110110010011;
assign LUT_4[35443] = 32'b11111111111111111000000010001011;
assign LUT_4[35444] = 32'b11111111111111111100011100001011;
assign LUT_4[35445] = 32'b11111111111111110101101000000011;
assign LUT_4[35446] = 32'b11111111111111111011110110101111;
assign LUT_4[35447] = 32'b11111111111111110101000010100111;
assign LUT_4[35448] = 32'b11111111111111111000101000000100;
assign LUT_4[35449] = 32'b11111111111111110001110011111100;
assign LUT_4[35450] = 32'b11111111111111111000000010101000;
assign LUT_4[35451] = 32'b11111111111111110001001110100000;
assign LUT_4[35452] = 32'b11111111111111110101101000100000;
assign LUT_4[35453] = 32'b11111111111111101110110100011000;
assign LUT_4[35454] = 32'b11111111111111110101000011000100;
assign LUT_4[35455] = 32'b11111111111111101110001110111100;
assign LUT_4[35456] = 32'b00000000000000000100011101101110;
assign LUT_4[35457] = 32'b11111111111111111101101001100110;
assign LUT_4[35458] = 32'b00000000000000000011111000010010;
assign LUT_4[35459] = 32'b11111111111111111101000100001010;
assign LUT_4[35460] = 32'b00000000000000000001011110001010;
assign LUT_4[35461] = 32'b11111111111111111010101010000010;
assign LUT_4[35462] = 32'b00000000000000000000111000101110;
assign LUT_4[35463] = 32'b11111111111111111010000100100110;
assign LUT_4[35464] = 32'b11111111111111111101101010000011;
assign LUT_4[35465] = 32'b11111111111111110110110101111011;
assign LUT_4[35466] = 32'b11111111111111111101000100100111;
assign LUT_4[35467] = 32'b11111111111111110110010000011111;
assign LUT_4[35468] = 32'b11111111111111111010101010011111;
assign LUT_4[35469] = 32'b11111111111111110011110110010111;
assign LUT_4[35470] = 32'b11111111111111111010000101000011;
assign LUT_4[35471] = 32'b11111111111111110011010000111011;
assign LUT_4[35472] = 32'b00000000000000000010001111011100;
assign LUT_4[35473] = 32'b11111111111111111011011011010100;
assign LUT_4[35474] = 32'b00000000000000000001101010000000;
assign LUT_4[35475] = 32'b11111111111111111010110101111000;
assign LUT_4[35476] = 32'b11111111111111111111001111111000;
assign LUT_4[35477] = 32'b11111111111111111000011011110000;
assign LUT_4[35478] = 32'b11111111111111111110101010011100;
assign LUT_4[35479] = 32'b11111111111111110111110110010100;
assign LUT_4[35480] = 32'b11111111111111111011011011110001;
assign LUT_4[35481] = 32'b11111111111111110100100111101001;
assign LUT_4[35482] = 32'b11111111111111111010110110010101;
assign LUT_4[35483] = 32'b11111111111111110100000010001101;
assign LUT_4[35484] = 32'b11111111111111111000011100001101;
assign LUT_4[35485] = 32'b11111111111111110001101000000101;
assign LUT_4[35486] = 32'b11111111111111110111110110110001;
assign LUT_4[35487] = 32'b11111111111111110001000010101001;
assign LUT_4[35488] = 32'b00000000000000000010111000110101;
assign LUT_4[35489] = 32'b11111111111111111100000100101101;
assign LUT_4[35490] = 32'b00000000000000000010010011011001;
assign LUT_4[35491] = 32'b11111111111111111011011111010001;
assign LUT_4[35492] = 32'b11111111111111111111111001010001;
assign LUT_4[35493] = 32'b11111111111111111001000101001001;
assign LUT_4[35494] = 32'b11111111111111111111010011110101;
assign LUT_4[35495] = 32'b11111111111111111000011111101101;
assign LUT_4[35496] = 32'b11111111111111111100000101001010;
assign LUT_4[35497] = 32'b11111111111111110101010001000010;
assign LUT_4[35498] = 32'b11111111111111111011011111101110;
assign LUT_4[35499] = 32'b11111111111111110100101011100110;
assign LUT_4[35500] = 32'b11111111111111111001000101100110;
assign LUT_4[35501] = 32'b11111111111111110010010001011110;
assign LUT_4[35502] = 32'b11111111111111111000100000001010;
assign LUT_4[35503] = 32'b11111111111111110001101100000010;
assign LUT_4[35504] = 32'b00000000000000000000101010100011;
assign LUT_4[35505] = 32'b11111111111111111001110110011011;
assign LUT_4[35506] = 32'b00000000000000000000000101000111;
assign LUT_4[35507] = 32'b11111111111111111001010000111111;
assign LUT_4[35508] = 32'b11111111111111111101101010111111;
assign LUT_4[35509] = 32'b11111111111111110110110110110111;
assign LUT_4[35510] = 32'b11111111111111111101000101100011;
assign LUT_4[35511] = 32'b11111111111111110110010001011011;
assign LUT_4[35512] = 32'b11111111111111111001110110111000;
assign LUT_4[35513] = 32'b11111111111111110011000010110000;
assign LUT_4[35514] = 32'b11111111111111111001010001011100;
assign LUT_4[35515] = 32'b11111111111111110010011101010100;
assign LUT_4[35516] = 32'b11111111111111110110110111010100;
assign LUT_4[35517] = 32'b11111111111111110000000011001100;
assign LUT_4[35518] = 32'b11111111111111110110010001111000;
assign LUT_4[35519] = 32'b11111111111111101111011101110000;
assign LUT_4[35520] = 32'b00000000000000000101110101000010;
assign LUT_4[35521] = 32'b11111111111111111111000000111010;
assign LUT_4[35522] = 32'b00000000000000000101001111100110;
assign LUT_4[35523] = 32'b11111111111111111110011011011110;
assign LUT_4[35524] = 32'b00000000000000000010110101011110;
assign LUT_4[35525] = 32'b11111111111111111100000001010110;
assign LUT_4[35526] = 32'b00000000000000000010010000000010;
assign LUT_4[35527] = 32'b11111111111111111011011011111010;
assign LUT_4[35528] = 32'b11111111111111111111000001010111;
assign LUT_4[35529] = 32'b11111111111111111000001101001111;
assign LUT_4[35530] = 32'b11111111111111111110011011111011;
assign LUT_4[35531] = 32'b11111111111111110111100111110011;
assign LUT_4[35532] = 32'b11111111111111111100000001110011;
assign LUT_4[35533] = 32'b11111111111111110101001101101011;
assign LUT_4[35534] = 32'b11111111111111111011011100010111;
assign LUT_4[35535] = 32'b11111111111111110100101000001111;
assign LUT_4[35536] = 32'b00000000000000000011100110110000;
assign LUT_4[35537] = 32'b11111111111111111100110010101000;
assign LUT_4[35538] = 32'b00000000000000000011000001010100;
assign LUT_4[35539] = 32'b11111111111111111100001101001100;
assign LUT_4[35540] = 32'b00000000000000000000100111001100;
assign LUT_4[35541] = 32'b11111111111111111001110011000100;
assign LUT_4[35542] = 32'b00000000000000000000000001110000;
assign LUT_4[35543] = 32'b11111111111111111001001101101000;
assign LUT_4[35544] = 32'b11111111111111111100110011000101;
assign LUT_4[35545] = 32'b11111111111111110101111110111101;
assign LUT_4[35546] = 32'b11111111111111111100001101101001;
assign LUT_4[35547] = 32'b11111111111111110101011001100001;
assign LUT_4[35548] = 32'b11111111111111111001110011100001;
assign LUT_4[35549] = 32'b11111111111111110010111111011001;
assign LUT_4[35550] = 32'b11111111111111111001001110000101;
assign LUT_4[35551] = 32'b11111111111111110010011001111101;
assign LUT_4[35552] = 32'b00000000000000000100010000001001;
assign LUT_4[35553] = 32'b11111111111111111101011100000001;
assign LUT_4[35554] = 32'b00000000000000000011101010101101;
assign LUT_4[35555] = 32'b11111111111111111100110110100101;
assign LUT_4[35556] = 32'b00000000000000000001010000100101;
assign LUT_4[35557] = 32'b11111111111111111010011100011101;
assign LUT_4[35558] = 32'b00000000000000000000101011001001;
assign LUT_4[35559] = 32'b11111111111111111001110111000001;
assign LUT_4[35560] = 32'b11111111111111111101011100011110;
assign LUT_4[35561] = 32'b11111111111111110110101000010110;
assign LUT_4[35562] = 32'b11111111111111111100110111000010;
assign LUT_4[35563] = 32'b11111111111111110110000010111010;
assign LUT_4[35564] = 32'b11111111111111111010011100111010;
assign LUT_4[35565] = 32'b11111111111111110011101000110010;
assign LUT_4[35566] = 32'b11111111111111111001110111011110;
assign LUT_4[35567] = 32'b11111111111111110011000011010110;
assign LUT_4[35568] = 32'b00000000000000000010000001110111;
assign LUT_4[35569] = 32'b11111111111111111011001101101111;
assign LUT_4[35570] = 32'b00000000000000000001011100011011;
assign LUT_4[35571] = 32'b11111111111111111010101000010011;
assign LUT_4[35572] = 32'b11111111111111111111000010010011;
assign LUT_4[35573] = 32'b11111111111111111000001110001011;
assign LUT_4[35574] = 32'b11111111111111111110011100110111;
assign LUT_4[35575] = 32'b11111111111111110111101000101111;
assign LUT_4[35576] = 32'b11111111111111111011001110001100;
assign LUT_4[35577] = 32'b11111111111111110100011010000100;
assign LUT_4[35578] = 32'b11111111111111111010101000110000;
assign LUT_4[35579] = 32'b11111111111111110011110100101000;
assign LUT_4[35580] = 32'b11111111111111111000001110101000;
assign LUT_4[35581] = 32'b11111111111111110001011010100000;
assign LUT_4[35582] = 32'b11111111111111110111101001001100;
assign LUT_4[35583] = 32'b11111111111111110000110101000100;
assign LUT_4[35584] = 32'b00000000000000000110110011001001;
assign LUT_4[35585] = 32'b11111111111111111111111111000001;
assign LUT_4[35586] = 32'b00000000000000000110001101101101;
assign LUT_4[35587] = 32'b11111111111111111111011001100101;
assign LUT_4[35588] = 32'b00000000000000000011110011100101;
assign LUT_4[35589] = 32'b11111111111111111100111111011101;
assign LUT_4[35590] = 32'b00000000000000000011001110001001;
assign LUT_4[35591] = 32'b11111111111111111100011010000001;
assign LUT_4[35592] = 32'b11111111111111111111111111011110;
assign LUT_4[35593] = 32'b11111111111111111001001011010110;
assign LUT_4[35594] = 32'b11111111111111111111011010000010;
assign LUT_4[35595] = 32'b11111111111111111000100101111010;
assign LUT_4[35596] = 32'b11111111111111111100111111111010;
assign LUT_4[35597] = 32'b11111111111111110110001011110010;
assign LUT_4[35598] = 32'b11111111111111111100011010011110;
assign LUT_4[35599] = 32'b11111111111111110101100110010110;
assign LUT_4[35600] = 32'b00000000000000000100100100110111;
assign LUT_4[35601] = 32'b11111111111111111101110000101111;
assign LUT_4[35602] = 32'b00000000000000000011111111011011;
assign LUT_4[35603] = 32'b11111111111111111101001011010011;
assign LUT_4[35604] = 32'b00000000000000000001100101010011;
assign LUT_4[35605] = 32'b11111111111111111010110001001011;
assign LUT_4[35606] = 32'b00000000000000000000111111110111;
assign LUT_4[35607] = 32'b11111111111111111010001011101111;
assign LUT_4[35608] = 32'b11111111111111111101110001001100;
assign LUT_4[35609] = 32'b11111111111111110110111101000100;
assign LUT_4[35610] = 32'b11111111111111111101001011110000;
assign LUT_4[35611] = 32'b11111111111111110110010111101000;
assign LUT_4[35612] = 32'b11111111111111111010110001101000;
assign LUT_4[35613] = 32'b11111111111111110011111101100000;
assign LUT_4[35614] = 32'b11111111111111111010001100001100;
assign LUT_4[35615] = 32'b11111111111111110011011000000100;
assign LUT_4[35616] = 32'b00000000000000000101001110010000;
assign LUT_4[35617] = 32'b11111111111111111110011010001000;
assign LUT_4[35618] = 32'b00000000000000000100101000110100;
assign LUT_4[35619] = 32'b11111111111111111101110100101100;
assign LUT_4[35620] = 32'b00000000000000000010001110101100;
assign LUT_4[35621] = 32'b11111111111111111011011010100100;
assign LUT_4[35622] = 32'b00000000000000000001101001010000;
assign LUT_4[35623] = 32'b11111111111111111010110101001000;
assign LUT_4[35624] = 32'b11111111111111111110011010100101;
assign LUT_4[35625] = 32'b11111111111111110111100110011101;
assign LUT_4[35626] = 32'b11111111111111111101110101001001;
assign LUT_4[35627] = 32'b11111111111111110111000001000001;
assign LUT_4[35628] = 32'b11111111111111111011011011000001;
assign LUT_4[35629] = 32'b11111111111111110100100110111001;
assign LUT_4[35630] = 32'b11111111111111111010110101100101;
assign LUT_4[35631] = 32'b11111111111111110100000001011101;
assign LUT_4[35632] = 32'b00000000000000000010111111111110;
assign LUT_4[35633] = 32'b11111111111111111100001011110110;
assign LUT_4[35634] = 32'b00000000000000000010011010100010;
assign LUT_4[35635] = 32'b11111111111111111011100110011010;
assign LUT_4[35636] = 32'b00000000000000000000000000011010;
assign LUT_4[35637] = 32'b11111111111111111001001100010010;
assign LUT_4[35638] = 32'b11111111111111111111011010111110;
assign LUT_4[35639] = 32'b11111111111111111000100110110110;
assign LUT_4[35640] = 32'b11111111111111111100001100010011;
assign LUT_4[35641] = 32'b11111111111111110101011000001011;
assign LUT_4[35642] = 32'b11111111111111111011100110110111;
assign LUT_4[35643] = 32'b11111111111111110100110010101111;
assign LUT_4[35644] = 32'b11111111111111111001001100101111;
assign LUT_4[35645] = 32'b11111111111111110010011000100111;
assign LUT_4[35646] = 32'b11111111111111111000100111010011;
assign LUT_4[35647] = 32'b11111111111111110001110011001011;
assign LUT_4[35648] = 32'b00000000000000001000001010011101;
assign LUT_4[35649] = 32'b00000000000000000001010110010101;
assign LUT_4[35650] = 32'b00000000000000000111100101000001;
assign LUT_4[35651] = 32'b00000000000000000000110000111001;
assign LUT_4[35652] = 32'b00000000000000000101001010111001;
assign LUT_4[35653] = 32'b11111111111111111110010110110001;
assign LUT_4[35654] = 32'b00000000000000000100100101011101;
assign LUT_4[35655] = 32'b11111111111111111101110001010101;
assign LUT_4[35656] = 32'b00000000000000000001010110110010;
assign LUT_4[35657] = 32'b11111111111111111010100010101010;
assign LUT_4[35658] = 32'b00000000000000000000110001010110;
assign LUT_4[35659] = 32'b11111111111111111001111101001110;
assign LUT_4[35660] = 32'b11111111111111111110010111001110;
assign LUT_4[35661] = 32'b11111111111111110111100011000110;
assign LUT_4[35662] = 32'b11111111111111111101110001110010;
assign LUT_4[35663] = 32'b11111111111111110110111101101010;
assign LUT_4[35664] = 32'b00000000000000000101111100001011;
assign LUT_4[35665] = 32'b11111111111111111111001000000011;
assign LUT_4[35666] = 32'b00000000000000000101010110101111;
assign LUT_4[35667] = 32'b11111111111111111110100010100111;
assign LUT_4[35668] = 32'b00000000000000000010111100100111;
assign LUT_4[35669] = 32'b11111111111111111100001000011111;
assign LUT_4[35670] = 32'b00000000000000000010010111001011;
assign LUT_4[35671] = 32'b11111111111111111011100011000011;
assign LUT_4[35672] = 32'b11111111111111111111001000100000;
assign LUT_4[35673] = 32'b11111111111111111000010100011000;
assign LUT_4[35674] = 32'b11111111111111111110100011000100;
assign LUT_4[35675] = 32'b11111111111111110111101110111100;
assign LUT_4[35676] = 32'b11111111111111111100001000111100;
assign LUT_4[35677] = 32'b11111111111111110101010100110100;
assign LUT_4[35678] = 32'b11111111111111111011100011100000;
assign LUT_4[35679] = 32'b11111111111111110100101111011000;
assign LUT_4[35680] = 32'b00000000000000000110100101100100;
assign LUT_4[35681] = 32'b11111111111111111111110001011100;
assign LUT_4[35682] = 32'b00000000000000000110000000001000;
assign LUT_4[35683] = 32'b11111111111111111111001100000000;
assign LUT_4[35684] = 32'b00000000000000000011100110000000;
assign LUT_4[35685] = 32'b11111111111111111100110001111000;
assign LUT_4[35686] = 32'b00000000000000000011000000100100;
assign LUT_4[35687] = 32'b11111111111111111100001100011100;
assign LUT_4[35688] = 32'b11111111111111111111110001111001;
assign LUT_4[35689] = 32'b11111111111111111000111101110001;
assign LUT_4[35690] = 32'b11111111111111111111001100011101;
assign LUT_4[35691] = 32'b11111111111111111000011000010101;
assign LUT_4[35692] = 32'b11111111111111111100110010010101;
assign LUT_4[35693] = 32'b11111111111111110101111110001101;
assign LUT_4[35694] = 32'b11111111111111111100001100111001;
assign LUT_4[35695] = 32'b11111111111111110101011000110001;
assign LUT_4[35696] = 32'b00000000000000000100010111010010;
assign LUT_4[35697] = 32'b11111111111111111101100011001010;
assign LUT_4[35698] = 32'b00000000000000000011110001110110;
assign LUT_4[35699] = 32'b11111111111111111100111101101110;
assign LUT_4[35700] = 32'b00000000000000000001010111101110;
assign LUT_4[35701] = 32'b11111111111111111010100011100110;
assign LUT_4[35702] = 32'b00000000000000000000110010010010;
assign LUT_4[35703] = 32'b11111111111111111001111110001010;
assign LUT_4[35704] = 32'b11111111111111111101100011100111;
assign LUT_4[35705] = 32'b11111111111111110110101111011111;
assign LUT_4[35706] = 32'b11111111111111111100111110001011;
assign LUT_4[35707] = 32'b11111111111111110110001010000011;
assign LUT_4[35708] = 32'b11111111111111111010100100000011;
assign LUT_4[35709] = 32'b11111111111111110011101111111011;
assign LUT_4[35710] = 32'b11111111111111111001111110100111;
assign LUT_4[35711] = 32'b11111111111111110011001010011111;
assign LUT_4[35712] = 32'b00000000000000001001011001010001;
assign LUT_4[35713] = 32'b00000000000000000010100101001001;
assign LUT_4[35714] = 32'b00000000000000001000110011110101;
assign LUT_4[35715] = 32'b00000000000000000001111111101101;
assign LUT_4[35716] = 32'b00000000000000000110011001101101;
assign LUT_4[35717] = 32'b11111111111111111111100101100101;
assign LUT_4[35718] = 32'b00000000000000000101110100010001;
assign LUT_4[35719] = 32'b11111111111111111111000000001001;
assign LUT_4[35720] = 32'b00000000000000000010100101100110;
assign LUT_4[35721] = 32'b11111111111111111011110001011110;
assign LUT_4[35722] = 32'b00000000000000000010000000001010;
assign LUT_4[35723] = 32'b11111111111111111011001100000010;
assign LUT_4[35724] = 32'b11111111111111111111100110000010;
assign LUT_4[35725] = 32'b11111111111111111000110001111010;
assign LUT_4[35726] = 32'b11111111111111111111000000100110;
assign LUT_4[35727] = 32'b11111111111111111000001100011110;
assign LUT_4[35728] = 32'b00000000000000000111001010111111;
assign LUT_4[35729] = 32'b00000000000000000000010110110111;
assign LUT_4[35730] = 32'b00000000000000000110100101100011;
assign LUT_4[35731] = 32'b11111111111111111111110001011011;
assign LUT_4[35732] = 32'b00000000000000000100001011011011;
assign LUT_4[35733] = 32'b11111111111111111101010111010011;
assign LUT_4[35734] = 32'b00000000000000000011100101111111;
assign LUT_4[35735] = 32'b11111111111111111100110001110111;
assign LUT_4[35736] = 32'b00000000000000000000010111010100;
assign LUT_4[35737] = 32'b11111111111111111001100011001100;
assign LUT_4[35738] = 32'b11111111111111111111110001111000;
assign LUT_4[35739] = 32'b11111111111111111000111101110000;
assign LUT_4[35740] = 32'b11111111111111111101010111110000;
assign LUT_4[35741] = 32'b11111111111111110110100011101000;
assign LUT_4[35742] = 32'b11111111111111111100110010010100;
assign LUT_4[35743] = 32'b11111111111111110101111110001100;
assign LUT_4[35744] = 32'b00000000000000000111110100011000;
assign LUT_4[35745] = 32'b00000000000000000001000000010000;
assign LUT_4[35746] = 32'b00000000000000000111001110111100;
assign LUT_4[35747] = 32'b00000000000000000000011010110100;
assign LUT_4[35748] = 32'b00000000000000000100110100110100;
assign LUT_4[35749] = 32'b11111111111111111110000000101100;
assign LUT_4[35750] = 32'b00000000000000000100001111011000;
assign LUT_4[35751] = 32'b11111111111111111101011011010000;
assign LUT_4[35752] = 32'b00000000000000000001000000101101;
assign LUT_4[35753] = 32'b11111111111111111010001100100101;
assign LUT_4[35754] = 32'b00000000000000000000011011010001;
assign LUT_4[35755] = 32'b11111111111111111001100111001001;
assign LUT_4[35756] = 32'b11111111111111111110000001001001;
assign LUT_4[35757] = 32'b11111111111111110111001101000001;
assign LUT_4[35758] = 32'b11111111111111111101011011101101;
assign LUT_4[35759] = 32'b11111111111111110110100111100101;
assign LUT_4[35760] = 32'b00000000000000000101100110000110;
assign LUT_4[35761] = 32'b11111111111111111110110001111110;
assign LUT_4[35762] = 32'b00000000000000000101000000101010;
assign LUT_4[35763] = 32'b11111111111111111110001100100010;
assign LUT_4[35764] = 32'b00000000000000000010100110100010;
assign LUT_4[35765] = 32'b11111111111111111011110010011010;
assign LUT_4[35766] = 32'b00000000000000000010000001000110;
assign LUT_4[35767] = 32'b11111111111111111011001100111110;
assign LUT_4[35768] = 32'b11111111111111111110110010011011;
assign LUT_4[35769] = 32'b11111111111111110111111110010011;
assign LUT_4[35770] = 32'b11111111111111111110001100111111;
assign LUT_4[35771] = 32'b11111111111111110111011000110111;
assign LUT_4[35772] = 32'b11111111111111111011110010110111;
assign LUT_4[35773] = 32'b11111111111111110100111110101111;
assign LUT_4[35774] = 32'b11111111111111111011001101011011;
assign LUT_4[35775] = 32'b11111111111111110100011001010011;
assign LUT_4[35776] = 32'b00000000000000001010110000100101;
assign LUT_4[35777] = 32'b00000000000000000011111100011101;
assign LUT_4[35778] = 32'b00000000000000001010001011001001;
assign LUT_4[35779] = 32'b00000000000000000011010111000001;
assign LUT_4[35780] = 32'b00000000000000000111110001000001;
assign LUT_4[35781] = 32'b00000000000000000000111100111001;
assign LUT_4[35782] = 32'b00000000000000000111001011100101;
assign LUT_4[35783] = 32'b00000000000000000000010111011101;
assign LUT_4[35784] = 32'b00000000000000000011111100111010;
assign LUT_4[35785] = 32'b11111111111111111101001000110010;
assign LUT_4[35786] = 32'b00000000000000000011010111011110;
assign LUT_4[35787] = 32'b11111111111111111100100011010110;
assign LUT_4[35788] = 32'b00000000000000000000111101010110;
assign LUT_4[35789] = 32'b11111111111111111010001001001110;
assign LUT_4[35790] = 32'b00000000000000000000010111111010;
assign LUT_4[35791] = 32'b11111111111111111001100011110010;
assign LUT_4[35792] = 32'b00000000000000001000100010010011;
assign LUT_4[35793] = 32'b00000000000000000001101110001011;
assign LUT_4[35794] = 32'b00000000000000000111111100110111;
assign LUT_4[35795] = 32'b00000000000000000001001000101111;
assign LUT_4[35796] = 32'b00000000000000000101100010101111;
assign LUT_4[35797] = 32'b11111111111111111110101110100111;
assign LUT_4[35798] = 32'b00000000000000000100111101010011;
assign LUT_4[35799] = 32'b11111111111111111110001001001011;
assign LUT_4[35800] = 32'b00000000000000000001101110101000;
assign LUT_4[35801] = 32'b11111111111111111010111010100000;
assign LUT_4[35802] = 32'b00000000000000000001001001001100;
assign LUT_4[35803] = 32'b11111111111111111010010101000100;
assign LUT_4[35804] = 32'b11111111111111111110101111000100;
assign LUT_4[35805] = 32'b11111111111111110111111010111100;
assign LUT_4[35806] = 32'b11111111111111111110001001101000;
assign LUT_4[35807] = 32'b11111111111111110111010101100000;
assign LUT_4[35808] = 32'b00000000000000001001001011101100;
assign LUT_4[35809] = 32'b00000000000000000010010111100100;
assign LUT_4[35810] = 32'b00000000000000001000100110010000;
assign LUT_4[35811] = 32'b00000000000000000001110010001000;
assign LUT_4[35812] = 32'b00000000000000000110001100001000;
assign LUT_4[35813] = 32'b11111111111111111111011000000000;
assign LUT_4[35814] = 32'b00000000000000000101100110101100;
assign LUT_4[35815] = 32'b11111111111111111110110010100100;
assign LUT_4[35816] = 32'b00000000000000000010011000000001;
assign LUT_4[35817] = 32'b11111111111111111011100011111001;
assign LUT_4[35818] = 32'b00000000000000000001110010100101;
assign LUT_4[35819] = 32'b11111111111111111010111110011101;
assign LUT_4[35820] = 32'b11111111111111111111011000011101;
assign LUT_4[35821] = 32'b11111111111111111000100100010101;
assign LUT_4[35822] = 32'b11111111111111111110110011000001;
assign LUT_4[35823] = 32'b11111111111111110111111110111001;
assign LUT_4[35824] = 32'b00000000000000000110111101011010;
assign LUT_4[35825] = 32'b00000000000000000000001001010010;
assign LUT_4[35826] = 32'b00000000000000000110010111111110;
assign LUT_4[35827] = 32'b11111111111111111111100011110110;
assign LUT_4[35828] = 32'b00000000000000000011111101110110;
assign LUT_4[35829] = 32'b11111111111111111101001001101110;
assign LUT_4[35830] = 32'b00000000000000000011011000011010;
assign LUT_4[35831] = 32'b11111111111111111100100100010010;
assign LUT_4[35832] = 32'b00000000000000000000001001101111;
assign LUT_4[35833] = 32'b11111111111111111001010101100111;
assign LUT_4[35834] = 32'b11111111111111111111100100010011;
assign LUT_4[35835] = 32'b11111111111111111000110000001011;
assign LUT_4[35836] = 32'b11111111111111111101001010001011;
assign LUT_4[35837] = 32'b11111111111111110110010110000011;
assign LUT_4[35838] = 32'b11111111111111111100100100101111;
assign LUT_4[35839] = 32'b11111111111111110101110000100111;
assign LUT_4[35840] = 32'b00000000000000000100011101111101;
assign LUT_4[35841] = 32'b11111111111111111101101001110101;
assign LUT_4[35842] = 32'b00000000000000000011111000100001;
assign LUT_4[35843] = 32'b11111111111111111101000100011001;
assign LUT_4[35844] = 32'b00000000000000000001011110011001;
assign LUT_4[35845] = 32'b11111111111111111010101010010001;
assign LUT_4[35846] = 32'b00000000000000000000111000111101;
assign LUT_4[35847] = 32'b11111111111111111010000100110101;
assign LUT_4[35848] = 32'b11111111111111111101101010010010;
assign LUT_4[35849] = 32'b11111111111111110110110110001010;
assign LUT_4[35850] = 32'b11111111111111111101000100110110;
assign LUT_4[35851] = 32'b11111111111111110110010000101110;
assign LUT_4[35852] = 32'b11111111111111111010101010101110;
assign LUT_4[35853] = 32'b11111111111111110011110110100110;
assign LUT_4[35854] = 32'b11111111111111111010000101010010;
assign LUT_4[35855] = 32'b11111111111111110011010001001010;
assign LUT_4[35856] = 32'b00000000000000000010001111101011;
assign LUT_4[35857] = 32'b11111111111111111011011011100011;
assign LUT_4[35858] = 32'b00000000000000000001101010001111;
assign LUT_4[35859] = 32'b11111111111111111010110110000111;
assign LUT_4[35860] = 32'b11111111111111111111010000000111;
assign LUT_4[35861] = 32'b11111111111111111000011011111111;
assign LUT_4[35862] = 32'b11111111111111111110101010101011;
assign LUT_4[35863] = 32'b11111111111111110111110110100011;
assign LUT_4[35864] = 32'b11111111111111111011011100000000;
assign LUT_4[35865] = 32'b11111111111111110100100111111000;
assign LUT_4[35866] = 32'b11111111111111111010110110100100;
assign LUT_4[35867] = 32'b11111111111111110100000010011100;
assign LUT_4[35868] = 32'b11111111111111111000011100011100;
assign LUT_4[35869] = 32'b11111111111111110001101000010100;
assign LUT_4[35870] = 32'b11111111111111110111110111000000;
assign LUT_4[35871] = 32'b11111111111111110001000010111000;
assign LUT_4[35872] = 32'b00000000000000000010111001000100;
assign LUT_4[35873] = 32'b11111111111111111100000100111100;
assign LUT_4[35874] = 32'b00000000000000000010010011101000;
assign LUT_4[35875] = 32'b11111111111111111011011111100000;
assign LUT_4[35876] = 32'b11111111111111111111111001100000;
assign LUT_4[35877] = 32'b11111111111111111001000101011000;
assign LUT_4[35878] = 32'b11111111111111111111010100000100;
assign LUT_4[35879] = 32'b11111111111111111000011111111100;
assign LUT_4[35880] = 32'b11111111111111111100000101011001;
assign LUT_4[35881] = 32'b11111111111111110101010001010001;
assign LUT_4[35882] = 32'b11111111111111111011011111111101;
assign LUT_4[35883] = 32'b11111111111111110100101011110101;
assign LUT_4[35884] = 32'b11111111111111111001000101110101;
assign LUT_4[35885] = 32'b11111111111111110010010001101101;
assign LUT_4[35886] = 32'b11111111111111111000100000011001;
assign LUT_4[35887] = 32'b11111111111111110001101100010001;
assign LUT_4[35888] = 32'b00000000000000000000101010110010;
assign LUT_4[35889] = 32'b11111111111111111001110110101010;
assign LUT_4[35890] = 32'b00000000000000000000000101010110;
assign LUT_4[35891] = 32'b11111111111111111001010001001110;
assign LUT_4[35892] = 32'b11111111111111111101101011001110;
assign LUT_4[35893] = 32'b11111111111111110110110111000110;
assign LUT_4[35894] = 32'b11111111111111111101000101110010;
assign LUT_4[35895] = 32'b11111111111111110110010001101010;
assign LUT_4[35896] = 32'b11111111111111111001110111000111;
assign LUT_4[35897] = 32'b11111111111111110011000010111111;
assign LUT_4[35898] = 32'b11111111111111111001010001101011;
assign LUT_4[35899] = 32'b11111111111111110010011101100011;
assign LUT_4[35900] = 32'b11111111111111110110110111100011;
assign LUT_4[35901] = 32'b11111111111111110000000011011011;
assign LUT_4[35902] = 32'b11111111111111110110010010000111;
assign LUT_4[35903] = 32'b11111111111111101111011101111111;
assign LUT_4[35904] = 32'b00000000000000000101110101010001;
assign LUT_4[35905] = 32'b11111111111111111111000001001001;
assign LUT_4[35906] = 32'b00000000000000000101001111110101;
assign LUT_4[35907] = 32'b11111111111111111110011011101101;
assign LUT_4[35908] = 32'b00000000000000000010110101101101;
assign LUT_4[35909] = 32'b11111111111111111100000001100101;
assign LUT_4[35910] = 32'b00000000000000000010010000010001;
assign LUT_4[35911] = 32'b11111111111111111011011100001001;
assign LUT_4[35912] = 32'b11111111111111111111000001100110;
assign LUT_4[35913] = 32'b11111111111111111000001101011110;
assign LUT_4[35914] = 32'b11111111111111111110011100001010;
assign LUT_4[35915] = 32'b11111111111111110111101000000010;
assign LUT_4[35916] = 32'b11111111111111111100000010000010;
assign LUT_4[35917] = 32'b11111111111111110101001101111010;
assign LUT_4[35918] = 32'b11111111111111111011011100100110;
assign LUT_4[35919] = 32'b11111111111111110100101000011110;
assign LUT_4[35920] = 32'b00000000000000000011100110111111;
assign LUT_4[35921] = 32'b11111111111111111100110010110111;
assign LUT_4[35922] = 32'b00000000000000000011000001100011;
assign LUT_4[35923] = 32'b11111111111111111100001101011011;
assign LUT_4[35924] = 32'b00000000000000000000100111011011;
assign LUT_4[35925] = 32'b11111111111111111001110011010011;
assign LUT_4[35926] = 32'b00000000000000000000000001111111;
assign LUT_4[35927] = 32'b11111111111111111001001101110111;
assign LUT_4[35928] = 32'b11111111111111111100110011010100;
assign LUT_4[35929] = 32'b11111111111111110101111111001100;
assign LUT_4[35930] = 32'b11111111111111111100001101111000;
assign LUT_4[35931] = 32'b11111111111111110101011001110000;
assign LUT_4[35932] = 32'b11111111111111111001110011110000;
assign LUT_4[35933] = 32'b11111111111111110010111111101000;
assign LUT_4[35934] = 32'b11111111111111111001001110010100;
assign LUT_4[35935] = 32'b11111111111111110010011010001100;
assign LUT_4[35936] = 32'b00000000000000000100010000011000;
assign LUT_4[35937] = 32'b11111111111111111101011100010000;
assign LUT_4[35938] = 32'b00000000000000000011101010111100;
assign LUT_4[35939] = 32'b11111111111111111100110110110100;
assign LUT_4[35940] = 32'b00000000000000000001010000110100;
assign LUT_4[35941] = 32'b11111111111111111010011100101100;
assign LUT_4[35942] = 32'b00000000000000000000101011011000;
assign LUT_4[35943] = 32'b11111111111111111001110111010000;
assign LUT_4[35944] = 32'b11111111111111111101011100101101;
assign LUT_4[35945] = 32'b11111111111111110110101000100101;
assign LUT_4[35946] = 32'b11111111111111111100110111010001;
assign LUT_4[35947] = 32'b11111111111111110110000011001001;
assign LUT_4[35948] = 32'b11111111111111111010011101001001;
assign LUT_4[35949] = 32'b11111111111111110011101001000001;
assign LUT_4[35950] = 32'b11111111111111111001110111101101;
assign LUT_4[35951] = 32'b11111111111111110011000011100101;
assign LUT_4[35952] = 32'b00000000000000000010000010000110;
assign LUT_4[35953] = 32'b11111111111111111011001101111110;
assign LUT_4[35954] = 32'b00000000000000000001011100101010;
assign LUT_4[35955] = 32'b11111111111111111010101000100010;
assign LUT_4[35956] = 32'b11111111111111111111000010100010;
assign LUT_4[35957] = 32'b11111111111111111000001110011010;
assign LUT_4[35958] = 32'b11111111111111111110011101000110;
assign LUT_4[35959] = 32'b11111111111111110111101000111110;
assign LUT_4[35960] = 32'b11111111111111111011001110011011;
assign LUT_4[35961] = 32'b11111111111111110100011010010011;
assign LUT_4[35962] = 32'b11111111111111111010101000111111;
assign LUT_4[35963] = 32'b11111111111111110011110100110111;
assign LUT_4[35964] = 32'b11111111111111111000001110110111;
assign LUT_4[35965] = 32'b11111111111111110001011010101111;
assign LUT_4[35966] = 32'b11111111111111110111101001011011;
assign LUT_4[35967] = 32'b11111111111111110000110101010011;
assign LUT_4[35968] = 32'b00000000000000000111000100000101;
assign LUT_4[35969] = 32'b00000000000000000000001111111101;
assign LUT_4[35970] = 32'b00000000000000000110011110101001;
assign LUT_4[35971] = 32'b11111111111111111111101010100001;
assign LUT_4[35972] = 32'b00000000000000000100000100100001;
assign LUT_4[35973] = 32'b11111111111111111101010000011001;
assign LUT_4[35974] = 32'b00000000000000000011011111000101;
assign LUT_4[35975] = 32'b11111111111111111100101010111101;
assign LUT_4[35976] = 32'b00000000000000000000010000011010;
assign LUT_4[35977] = 32'b11111111111111111001011100010010;
assign LUT_4[35978] = 32'b11111111111111111111101010111110;
assign LUT_4[35979] = 32'b11111111111111111000110110110110;
assign LUT_4[35980] = 32'b11111111111111111101010000110110;
assign LUT_4[35981] = 32'b11111111111111110110011100101110;
assign LUT_4[35982] = 32'b11111111111111111100101011011010;
assign LUT_4[35983] = 32'b11111111111111110101110111010010;
assign LUT_4[35984] = 32'b00000000000000000100110101110011;
assign LUT_4[35985] = 32'b11111111111111111110000001101011;
assign LUT_4[35986] = 32'b00000000000000000100010000010111;
assign LUT_4[35987] = 32'b11111111111111111101011100001111;
assign LUT_4[35988] = 32'b00000000000000000001110110001111;
assign LUT_4[35989] = 32'b11111111111111111011000010000111;
assign LUT_4[35990] = 32'b00000000000000000001010000110011;
assign LUT_4[35991] = 32'b11111111111111111010011100101011;
assign LUT_4[35992] = 32'b11111111111111111110000010001000;
assign LUT_4[35993] = 32'b11111111111111110111001110000000;
assign LUT_4[35994] = 32'b11111111111111111101011100101100;
assign LUT_4[35995] = 32'b11111111111111110110101000100100;
assign LUT_4[35996] = 32'b11111111111111111011000010100100;
assign LUT_4[35997] = 32'b11111111111111110100001110011100;
assign LUT_4[35998] = 32'b11111111111111111010011101001000;
assign LUT_4[35999] = 32'b11111111111111110011101001000000;
assign LUT_4[36000] = 32'b00000000000000000101011111001100;
assign LUT_4[36001] = 32'b11111111111111111110101011000100;
assign LUT_4[36002] = 32'b00000000000000000100111001110000;
assign LUT_4[36003] = 32'b11111111111111111110000101101000;
assign LUT_4[36004] = 32'b00000000000000000010011111101000;
assign LUT_4[36005] = 32'b11111111111111111011101011100000;
assign LUT_4[36006] = 32'b00000000000000000001111010001100;
assign LUT_4[36007] = 32'b11111111111111111011000110000100;
assign LUT_4[36008] = 32'b11111111111111111110101011100001;
assign LUT_4[36009] = 32'b11111111111111110111110111011001;
assign LUT_4[36010] = 32'b11111111111111111110000110000101;
assign LUT_4[36011] = 32'b11111111111111110111010001111101;
assign LUT_4[36012] = 32'b11111111111111111011101011111101;
assign LUT_4[36013] = 32'b11111111111111110100110111110101;
assign LUT_4[36014] = 32'b11111111111111111011000110100001;
assign LUT_4[36015] = 32'b11111111111111110100010010011001;
assign LUT_4[36016] = 32'b00000000000000000011010000111010;
assign LUT_4[36017] = 32'b11111111111111111100011100110010;
assign LUT_4[36018] = 32'b00000000000000000010101011011110;
assign LUT_4[36019] = 32'b11111111111111111011110111010110;
assign LUT_4[36020] = 32'b00000000000000000000010001010110;
assign LUT_4[36021] = 32'b11111111111111111001011101001110;
assign LUT_4[36022] = 32'b11111111111111111111101011111010;
assign LUT_4[36023] = 32'b11111111111111111000110111110010;
assign LUT_4[36024] = 32'b11111111111111111100011101001111;
assign LUT_4[36025] = 32'b11111111111111110101101001000111;
assign LUT_4[36026] = 32'b11111111111111111011110111110011;
assign LUT_4[36027] = 32'b11111111111111110101000011101011;
assign LUT_4[36028] = 32'b11111111111111111001011101101011;
assign LUT_4[36029] = 32'b11111111111111110010101001100011;
assign LUT_4[36030] = 32'b11111111111111111000111000001111;
assign LUT_4[36031] = 32'b11111111111111110010000100000111;
assign LUT_4[36032] = 32'b00000000000000001000011011011001;
assign LUT_4[36033] = 32'b00000000000000000001100111010001;
assign LUT_4[36034] = 32'b00000000000000000111110101111101;
assign LUT_4[36035] = 32'b00000000000000000001000001110101;
assign LUT_4[36036] = 32'b00000000000000000101011011110101;
assign LUT_4[36037] = 32'b11111111111111111110100111101101;
assign LUT_4[36038] = 32'b00000000000000000100110110011001;
assign LUT_4[36039] = 32'b11111111111111111110000010010001;
assign LUT_4[36040] = 32'b00000000000000000001100111101110;
assign LUT_4[36041] = 32'b11111111111111111010110011100110;
assign LUT_4[36042] = 32'b00000000000000000001000010010010;
assign LUT_4[36043] = 32'b11111111111111111010001110001010;
assign LUT_4[36044] = 32'b11111111111111111110101000001010;
assign LUT_4[36045] = 32'b11111111111111110111110100000010;
assign LUT_4[36046] = 32'b11111111111111111110000010101110;
assign LUT_4[36047] = 32'b11111111111111110111001110100110;
assign LUT_4[36048] = 32'b00000000000000000110001101000111;
assign LUT_4[36049] = 32'b11111111111111111111011000111111;
assign LUT_4[36050] = 32'b00000000000000000101100111101011;
assign LUT_4[36051] = 32'b11111111111111111110110011100011;
assign LUT_4[36052] = 32'b00000000000000000011001101100011;
assign LUT_4[36053] = 32'b11111111111111111100011001011011;
assign LUT_4[36054] = 32'b00000000000000000010101000000111;
assign LUT_4[36055] = 32'b11111111111111111011110011111111;
assign LUT_4[36056] = 32'b11111111111111111111011001011100;
assign LUT_4[36057] = 32'b11111111111111111000100101010100;
assign LUT_4[36058] = 32'b11111111111111111110110100000000;
assign LUT_4[36059] = 32'b11111111111111110111111111111000;
assign LUT_4[36060] = 32'b11111111111111111100011001111000;
assign LUT_4[36061] = 32'b11111111111111110101100101110000;
assign LUT_4[36062] = 32'b11111111111111111011110100011100;
assign LUT_4[36063] = 32'b11111111111111110101000000010100;
assign LUT_4[36064] = 32'b00000000000000000110110110100000;
assign LUT_4[36065] = 32'b00000000000000000000000010011000;
assign LUT_4[36066] = 32'b00000000000000000110010001000100;
assign LUT_4[36067] = 32'b11111111111111111111011100111100;
assign LUT_4[36068] = 32'b00000000000000000011110110111100;
assign LUT_4[36069] = 32'b11111111111111111101000010110100;
assign LUT_4[36070] = 32'b00000000000000000011010001100000;
assign LUT_4[36071] = 32'b11111111111111111100011101011000;
assign LUT_4[36072] = 32'b00000000000000000000000010110101;
assign LUT_4[36073] = 32'b11111111111111111001001110101101;
assign LUT_4[36074] = 32'b11111111111111111111011101011001;
assign LUT_4[36075] = 32'b11111111111111111000101001010001;
assign LUT_4[36076] = 32'b11111111111111111101000011010001;
assign LUT_4[36077] = 32'b11111111111111110110001111001001;
assign LUT_4[36078] = 32'b11111111111111111100011101110101;
assign LUT_4[36079] = 32'b11111111111111110101101001101101;
assign LUT_4[36080] = 32'b00000000000000000100101000001110;
assign LUT_4[36081] = 32'b11111111111111111101110100000110;
assign LUT_4[36082] = 32'b00000000000000000100000010110010;
assign LUT_4[36083] = 32'b11111111111111111101001110101010;
assign LUT_4[36084] = 32'b00000000000000000001101000101010;
assign LUT_4[36085] = 32'b11111111111111111010110100100010;
assign LUT_4[36086] = 32'b00000000000000000001000011001110;
assign LUT_4[36087] = 32'b11111111111111111010001111000110;
assign LUT_4[36088] = 32'b11111111111111111101110100100011;
assign LUT_4[36089] = 32'b11111111111111110111000000011011;
assign LUT_4[36090] = 32'b11111111111111111101001111000111;
assign LUT_4[36091] = 32'b11111111111111110110011010111111;
assign LUT_4[36092] = 32'b11111111111111111010110100111111;
assign LUT_4[36093] = 32'b11111111111111110100000000110111;
assign LUT_4[36094] = 32'b11111111111111111010001111100011;
assign LUT_4[36095] = 32'b11111111111111110011011011011011;
assign LUT_4[36096] = 32'b00000000000000001001011001100000;
assign LUT_4[36097] = 32'b00000000000000000010100101011000;
assign LUT_4[36098] = 32'b00000000000000001000110100000100;
assign LUT_4[36099] = 32'b00000000000000000001111111111100;
assign LUT_4[36100] = 32'b00000000000000000110011001111100;
assign LUT_4[36101] = 32'b11111111111111111111100101110100;
assign LUT_4[36102] = 32'b00000000000000000101110100100000;
assign LUT_4[36103] = 32'b11111111111111111111000000011000;
assign LUT_4[36104] = 32'b00000000000000000010100101110101;
assign LUT_4[36105] = 32'b11111111111111111011110001101101;
assign LUT_4[36106] = 32'b00000000000000000010000000011001;
assign LUT_4[36107] = 32'b11111111111111111011001100010001;
assign LUT_4[36108] = 32'b11111111111111111111100110010001;
assign LUT_4[36109] = 32'b11111111111111111000110010001001;
assign LUT_4[36110] = 32'b11111111111111111111000000110101;
assign LUT_4[36111] = 32'b11111111111111111000001100101101;
assign LUT_4[36112] = 32'b00000000000000000111001011001110;
assign LUT_4[36113] = 32'b00000000000000000000010111000110;
assign LUT_4[36114] = 32'b00000000000000000110100101110010;
assign LUT_4[36115] = 32'b11111111111111111111110001101010;
assign LUT_4[36116] = 32'b00000000000000000100001011101010;
assign LUT_4[36117] = 32'b11111111111111111101010111100010;
assign LUT_4[36118] = 32'b00000000000000000011100110001110;
assign LUT_4[36119] = 32'b11111111111111111100110010000110;
assign LUT_4[36120] = 32'b00000000000000000000010111100011;
assign LUT_4[36121] = 32'b11111111111111111001100011011011;
assign LUT_4[36122] = 32'b11111111111111111111110010000111;
assign LUT_4[36123] = 32'b11111111111111111000111101111111;
assign LUT_4[36124] = 32'b11111111111111111101010111111111;
assign LUT_4[36125] = 32'b11111111111111110110100011110111;
assign LUT_4[36126] = 32'b11111111111111111100110010100011;
assign LUT_4[36127] = 32'b11111111111111110101111110011011;
assign LUT_4[36128] = 32'b00000000000000000111110100100111;
assign LUT_4[36129] = 32'b00000000000000000001000000011111;
assign LUT_4[36130] = 32'b00000000000000000111001111001011;
assign LUT_4[36131] = 32'b00000000000000000000011011000011;
assign LUT_4[36132] = 32'b00000000000000000100110101000011;
assign LUT_4[36133] = 32'b11111111111111111110000000111011;
assign LUT_4[36134] = 32'b00000000000000000100001111100111;
assign LUT_4[36135] = 32'b11111111111111111101011011011111;
assign LUT_4[36136] = 32'b00000000000000000001000000111100;
assign LUT_4[36137] = 32'b11111111111111111010001100110100;
assign LUT_4[36138] = 32'b00000000000000000000011011100000;
assign LUT_4[36139] = 32'b11111111111111111001100111011000;
assign LUT_4[36140] = 32'b11111111111111111110000001011000;
assign LUT_4[36141] = 32'b11111111111111110111001101010000;
assign LUT_4[36142] = 32'b11111111111111111101011011111100;
assign LUT_4[36143] = 32'b11111111111111110110100111110100;
assign LUT_4[36144] = 32'b00000000000000000101100110010101;
assign LUT_4[36145] = 32'b11111111111111111110110010001101;
assign LUT_4[36146] = 32'b00000000000000000101000000111001;
assign LUT_4[36147] = 32'b11111111111111111110001100110001;
assign LUT_4[36148] = 32'b00000000000000000010100110110001;
assign LUT_4[36149] = 32'b11111111111111111011110010101001;
assign LUT_4[36150] = 32'b00000000000000000010000001010101;
assign LUT_4[36151] = 32'b11111111111111111011001101001101;
assign LUT_4[36152] = 32'b11111111111111111110110010101010;
assign LUT_4[36153] = 32'b11111111111111110111111110100010;
assign LUT_4[36154] = 32'b11111111111111111110001101001110;
assign LUT_4[36155] = 32'b11111111111111110111011001000110;
assign LUT_4[36156] = 32'b11111111111111111011110011000110;
assign LUT_4[36157] = 32'b11111111111111110100111110111110;
assign LUT_4[36158] = 32'b11111111111111111011001101101010;
assign LUT_4[36159] = 32'b11111111111111110100011001100010;
assign LUT_4[36160] = 32'b00000000000000001010110000110100;
assign LUT_4[36161] = 32'b00000000000000000011111100101100;
assign LUT_4[36162] = 32'b00000000000000001010001011011000;
assign LUT_4[36163] = 32'b00000000000000000011010111010000;
assign LUT_4[36164] = 32'b00000000000000000111110001010000;
assign LUT_4[36165] = 32'b00000000000000000000111101001000;
assign LUT_4[36166] = 32'b00000000000000000111001011110100;
assign LUT_4[36167] = 32'b00000000000000000000010111101100;
assign LUT_4[36168] = 32'b00000000000000000011111101001001;
assign LUT_4[36169] = 32'b11111111111111111101001001000001;
assign LUT_4[36170] = 32'b00000000000000000011010111101101;
assign LUT_4[36171] = 32'b11111111111111111100100011100101;
assign LUT_4[36172] = 32'b00000000000000000000111101100101;
assign LUT_4[36173] = 32'b11111111111111111010001001011101;
assign LUT_4[36174] = 32'b00000000000000000000011000001001;
assign LUT_4[36175] = 32'b11111111111111111001100100000001;
assign LUT_4[36176] = 32'b00000000000000001000100010100010;
assign LUT_4[36177] = 32'b00000000000000000001101110011010;
assign LUT_4[36178] = 32'b00000000000000000111111101000110;
assign LUT_4[36179] = 32'b00000000000000000001001000111110;
assign LUT_4[36180] = 32'b00000000000000000101100010111110;
assign LUT_4[36181] = 32'b11111111111111111110101110110110;
assign LUT_4[36182] = 32'b00000000000000000100111101100010;
assign LUT_4[36183] = 32'b11111111111111111110001001011010;
assign LUT_4[36184] = 32'b00000000000000000001101110110111;
assign LUT_4[36185] = 32'b11111111111111111010111010101111;
assign LUT_4[36186] = 32'b00000000000000000001001001011011;
assign LUT_4[36187] = 32'b11111111111111111010010101010011;
assign LUT_4[36188] = 32'b11111111111111111110101111010011;
assign LUT_4[36189] = 32'b11111111111111110111111011001011;
assign LUT_4[36190] = 32'b11111111111111111110001001110111;
assign LUT_4[36191] = 32'b11111111111111110111010101101111;
assign LUT_4[36192] = 32'b00000000000000001001001011111011;
assign LUT_4[36193] = 32'b00000000000000000010010111110011;
assign LUT_4[36194] = 32'b00000000000000001000100110011111;
assign LUT_4[36195] = 32'b00000000000000000001110010010111;
assign LUT_4[36196] = 32'b00000000000000000110001100010111;
assign LUT_4[36197] = 32'b11111111111111111111011000001111;
assign LUT_4[36198] = 32'b00000000000000000101100110111011;
assign LUT_4[36199] = 32'b11111111111111111110110010110011;
assign LUT_4[36200] = 32'b00000000000000000010011000010000;
assign LUT_4[36201] = 32'b11111111111111111011100100001000;
assign LUT_4[36202] = 32'b00000000000000000001110010110100;
assign LUT_4[36203] = 32'b11111111111111111010111110101100;
assign LUT_4[36204] = 32'b11111111111111111111011000101100;
assign LUT_4[36205] = 32'b11111111111111111000100100100100;
assign LUT_4[36206] = 32'b11111111111111111110110011010000;
assign LUT_4[36207] = 32'b11111111111111110111111111001000;
assign LUT_4[36208] = 32'b00000000000000000110111101101001;
assign LUT_4[36209] = 32'b00000000000000000000001001100001;
assign LUT_4[36210] = 32'b00000000000000000110011000001101;
assign LUT_4[36211] = 32'b11111111111111111111100100000101;
assign LUT_4[36212] = 32'b00000000000000000011111110000101;
assign LUT_4[36213] = 32'b11111111111111111101001001111101;
assign LUT_4[36214] = 32'b00000000000000000011011000101001;
assign LUT_4[36215] = 32'b11111111111111111100100100100001;
assign LUT_4[36216] = 32'b00000000000000000000001001111110;
assign LUT_4[36217] = 32'b11111111111111111001010101110110;
assign LUT_4[36218] = 32'b11111111111111111111100100100010;
assign LUT_4[36219] = 32'b11111111111111111000110000011010;
assign LUT_4[36220] = 32'b11111111111111111101001010011010;
assign LUT_4[36221] = 32'b11111111111111110110010110010010;
assign LUT_4[36222] = 32'b11111111111111111100100100111110;
assign LUT_4[36223] = 32'b11111111111111110101110000110110;
assign LUT_4[36224] = 32'b00000000000000001011111111101000;
assign LUT_4[36225] = 32'b00000000000000000101001011100000;
assign LUT_4[36226] = 32'b00000000000000001011011010001100;
assign LUT_4[36227] = 32'b00000000000000000100100110000100;
assign LUT_4[36228] = 32'b00000000000000001001000000000100;
assign LUT_4[36229] = 32'b00000000000000000010001011111100;
assign LUT_4[36230] = 32'b00000000000000001000011010101000;
assign LUT_4[36231] = 32'b00000000000000000001100110100000;
assign LUT_4[36232] = 32'b00000000000000000101001011111101;
assign LUT_4[36233] = 32'b11111111111111111110010111110101;
assign LUT_4[36234] = 32'b00000000000000000100100110100001;
assign LUT_4[36235] = 32'b11111111111111111101110010011001;
assign LUT_4[36236] = 32'b00000000000000000010001100011001;
assign LUT_4[36237] = 32'b11111111111111111011011000010001;
assign LUT_4[36238] = 32'b00000000000000000001100110111101;
assign LUT_4[36239] = 32'b11111111111111111010110010110101;
assign LUT_4[36240] = 32'b00000000000000001001110001010110;
assign LUT_4[36241] = 32'b00000000000000000010111101001110;
assign LUT_4[36242] = 32'b00000000000000001001001011111010;
assign LUT_4[36243] = 32'b00000000000000000010010111110010;
assign LUT_4[36244] = 32'b00000000000000000110110001110010;
assign LUT_4[36245] = 32'b11111111111111111111111101101010;
assign LUT_4[36246] = 32'b00000000000000000110001100010110;
assign LUT_4[36247] = 32'b11111111111111111111011000001110;
assign LUT_4[36248] = 32'b00000000000000000010111101101011;
assign LUT_4[36249] = 32'b11111111111111111100001001100011;
assign LUT_4[36250] = 32'b00000000000000000010011000001111;
assign LUT_4[36251] = 32'b11111111111111111011100100000111;
assign LUT_4[36252] = 32'b11111111111111111111111110000111;
assign LUT_4[36253] = 32'b11111111111111111001001001111111;
assign LUT_4[36254] = 32'b11111111111111111111011000101011;
assign LUT_4[36255] = 32'b11111111111111111000100100100011;
assign LUT_4[36256] = 32'b00000000000000001010011010101111;
assign LUT_4[36257] = 32'b00000000000000000011100110100111;
assign LUT_4[36258] = 32'b00000000000000001001110101010011;
assign LUT_4[36259] = 32'b00000000000000000011000001001011;
assign LUT_4[36260] = 32'b00000000000000000111011011001011;
assign LUT_4[36261] = 32'b00000000000000000000100111000011;
assign LUT_4[36262] = 32'b00000000000000000110110101101111;
assign LUT_4[36263] = 32'b00000000000000000000000001100111;
assign LUT_4[36264] = 32'b00000000000000000011100111000100;
assign LUT_4[36265] = 32'b11111111111111111100110010111100;
assign LUT_4[36266] = 32'b00000000000000000011000001101000;
assign LUT_4[36267] = 32'b11111111111111111100001101100000;
assign LUT_4[36268] = 32'b00000000000000000000100111100000;
assign LUT_4[36269] = 32'b11111111111111111001110011011000;
assign LUT_4[36270] = 32'b00000000000000000000000010000100;
assign LUT_4[36271] = 32'b11111111111111111001001101111100;
assign LUT_4[36272] = 32'b00000000000000001000001100011101;
assign LUT_4[36273] = 32'b00000000000000000001011000010101;
assign LUT_4[36274] = 32'b00000000000000000111100111000001;
assign LUT_4[36275] = 32'b00000000000000000000110010111001;
assign LUT_4[36276] = 32'b00000000000000000101001100111001;
assign LUT_4[36277] = 32'b11111111111111111110011000110001;
assign LUT_4[36278] = 32'b00000000000000000100100111011101;
assign LUT_4[36279] = 32'b11111111111111111101110011010101;
assign LUT_4[36280] = 32'b00000000000000000001011000110010;
assign LUT_4[36281] = 32'b11111111111111111010100100101010;
assign LUT_4[36282] = 32'b00000000000000000000110011010110;
assign LUT_4[36283] = 32'b11111111111111111001111111001110;
assign LUT_4[36284] = 32'b11111111111111111110011001001110;
assign LUT_4[36285] = 32'b11111111111111110111100101000110;
assign LUT_4[36286] = 32'b11111111111111111101110011110010;
assign LUT_4[36287] = 32'b11111111111111110110111111101010;
assign LUT_4[36288] = 32'b00000000000000001101010110111100;
assign LUT_4[36289] = 32'b00000000000000000110100010110100;
assign LUT_4[36290] = 32'b00000000000000001100110001100000;
assign LUT_4[36291] = 32'b00000000000000000101111101011000;
assign LUT_4[36292] = 32'b00000000000000001010010111011000;
assign LUT_4[36293] = 32'b00000000000000000011100011010000;
assign LUT_4[36294] = 32'b00000000000000001001110001111100;
assign LUT_4[36295] = 32'b00000000000000000010111101110100;
assign LUT_4[36296] = 32'b00000000000000000110100011010001;
assign LUT_4[36297] = 32'b11111111111111111111101111001001;
assign LUT_4[36298] = 32'b00000000000000000101111101110101;
assign LUT_4[36299] = 32'b11111111111111111111001001101101;
assign LUT_4[36300] = 32'b00000000000000000011100011101101;
assign LUT_4[36301] = 32'b11111111111111111100101111100101;
assign LUT_4[36302] = 32'b00000000000000000010111110010001;
assign LUT_4[36303] = 32'b11111111111111111100001010001001;
assign LUT_4[36304] = 32'b00000000000000001011001000101010;
assign LUT_4[36305] = 32'b00000000000000000100010100100010;
assign LUT_4[36306] = 32'b00000000000000001010100011001110;
assign LUT_4[36307] = 32'b00000000000000000011101111000110;
assign LUT_4[36308] = 32'b00000000000000001000001001000110;
assign LUT_4[36309] = 32'b00000000000000000001010100111110;
assign LUT_4[36310] = 32'b00000000000000000111100011101010;
assign LUT_4[36311] = 32'b00000000000000000000101111100010;
assign LUT_4[36312] = 32'b00000000000000000100010100111111;
assign LUT_4[36313] = 32'b11111111111111111101100000110111;
assign LUT_4[36314] = 32'b00000000000000000011101111100011;
assign LUT_4[36315] = 32'b11111111111111111100111011011011;
assign LUT_4[36316] = 32'b00000000000000000001010101011011;
assign LUT_4[36317] = 32'b11111111111111111010100001010011;
assign LUT_4[36318] = 32'b00000000000000000000101111111111;
assign LUT_4[36319] = 32'b11111111111111111001111011110111;
assign LUT_4[36320] = 32'b00000000000000001011110010000011;
assign LUT_4[36321] = 32'b00000000000000000100111101111011;
assign LUT_4[36322] = 32'b00000000000000001011001100100111;
assign LUT_4[36323] = 32'b00000000000000000100011000011111;
assign LUT_4[36324] = 32'b00000000000000001000110010011111;
assign LUT_4[36325] = 32'b00000000000000000001111110010111;
assign LUT_4[36326] = 32'b00000000000000001000001101000011;
assign LUT_4[36327] = 32'b00000000000000000001011000111011;
assign LUT_4[36328] = 32'b00000000000000000100111110011000;
assign LUT_4[36329] = 32'b11111111111111111110001010010000;
assign LUT_4[36330] = 32'b00000000000000000100011000111100;
assign LUT_4[36331] = 32'b11111111111111111101100100110100;
assign LUT_4[36332] = 32'b00000000000000000001111110110100;
assign LUT_4[36333] = 32'b11111111111111111011001010101100;
assign LUT_4[36334] = 32'b00000000000000000001011001011000;
assign LUT_4[36335] = 32'b11111111111111111010100101010000;
assign LUT_4[36336] = 32'b00000000000000001001100011110001;
assign LUT_4[36337] = 32'b00000000000000000010101111101001;
assign LUT_4[36338] = 32'b00000000000000001000111110010101;
assign LUT_4[36339] = 32'b00000000000000000010001010001101;
assign LUT_4[36340] = 32'b00000000000000000110100100001101;
assign LUT_4[36341] = 32'b11111111111111111111110000000101;
assign LUT_4[36342] = 32'b00000000000000000101111110110001;
assign LUT_4[36343] = 32'b11111111111111111111001010101001;
assign LUT_4[36344] = 32'b00000000000000000010110000000110;
assign LUT_4[36345] = 32'b11111111111111111011111011111110;
assign LUT_4[36346] = 32'b00000000000000000010001010101010;
assign LUT_4[36347] = 32'b11111111111111111011010110100010;
assign LUT_4[36348] = 32'b11111111111111111111110000100010;
assign LUT_4[36349] = 32'b11111111111111111000111100011010;
assign LUT_4[36350] = 32'b11111111111111111111001011000110;
assign LUT_4[36351] = 32'b11111111111111111000010110111110;
assign LUT_4[36352] = 32'b00000000000000000011100010000101;
assign LUT_4[36353] = 32'b11111111111111111100101101111101;
assign LUT_4[36354] = 32'b00000000000000000010111100101001;
assign LUT_4[36355] = 32'b11111111111111111100001000100001;
assign LUT_4[36356] = 32'b00000000000000000000100010100001;
assign LUT_4[36357] = 32'b11111111111111111001101110011001;
assign LUT_4[36358] = 32'b11111111111111111111111101000101;
assign LUT_4[36359] = 32'b11111111111111111001001000111101;
assign LUT_4[36360] = 32'b11111111111111111100101110011010;
assign LUT_4[36361] = 32'b11111111111111110101111010010010;
assign LUT_4[36362] = 32'b11111111111111111100001000111110;
assign LUT_4[36363] = 32'b11111111111111110101010100110110;
assign LUT_4[36364] = 32'b11111111111111111001101110110110;
assign LUT_4[36365] = 32'b11111111111111110010111010101110;
assign LUT_4[36366] = 32'b11111111111111111001001001011010;
assign LUT_4[36367] = 32'b11111111111111110010010101010010;
assign LUT_4[36368] = 32'b00000000000000000001010011110011;
assign LUT_4[36369] = 32'b11111111111111111010011111101011;
assign LUT_4[36370] = 32'b00000000000000000000101110010111;
assign LUT_4[36371] = 32'b11111111111111111001111010001111;
assign LUT_4[36372] = 32'b11111111111111111110010100001111;
assign LUT_4[36373] = 32'b11111111111111110111100000000111;
assign LUT_4[36374] = 32'b11111111111111111101101110110011;
assign LUT_4[36375] = 32'b11111111111111110110111010101011;
assign LUT_4[36376] = 32'b11111111111111111010100000001000;
assign LUT_4[36377] = 32'b11111111111111110011101100000000;
assign LUT_4[36378] = 32'b11111111111111111001111010101100;
assign LUT_4[36379] = 32'b11111111111111110011000110100100;
assign LUT_4[36380] = 32'b11111111111111110111100000100100;
assign LUT_4[36381] = 32'b11111111111111110000101100011100;
assign LUT_4[36382] = 32'b11111111111111110110111011001000;
assign LUT_4[36383] = 32'b11111111111111110000000111000000;
assign LUT_4[36384] = 32'b00000000000000000001111101001100;
assign LUT_4[36385] = 32'b11111111111111111011001001000100;
assign LUT_4[36386] = 32'b00000000000000000001010111110000;
assign LUT_4[36387] = 32'b11111111111111111010100011101000;
assign LUT_4[36388] = 32'b11111111111111111110111101101000;
assign LUT_4[36389] = 32'b11111111111111111000001001100000;
assign LUT_4[36390] = 32'b11111111111111111110011000001100;
assign LUT_4[36391] = 32'b11111111111111110111100100000100;
assign LUT_4[36392] = 32'b11111111111111111011001001100001;
assign LUT_4[36393] = 32'b11111111111111110100010101011001;
assign LUT_4[36394] = 32'b11111111111111111010100100000101;
assign LUT_4[36395] = 32'b11111111111111110011101111111101;
assign LUT_4[36396] = 32'b11111111111111111000001001111101;
assign LUT_4[36397] = 32'b11111111111111110001010101110101;
assign LUT_4[36398] = 32'b11111111111111110111100100100001;
assign LUT_4[36399] = 32'b11111111111111110000110000011001;
assign LUT_4[36400] = 32'b11111111111111111111101110111010;
assign LUT_4[36401] = 32'b11111111111111111000111010110010;
assign LUT_4[36402] = 32'b11111111111111111111001001011110;
assign LUT_4[36403] = 32'b11111111111111111000010101010110;
assign LUT_4[36404] = 32'b11111111111111111100101111010110;
assign LUT_4[36405] = 32'b11111111111111110101111011001110;
assign LUT_4[36406] = 32'b11111111111111111100001001111010;
assign LUT_4[36407] = 32'b11111111111111110101010101110010;
assign LUT_4[36408] = 32'b11111111111111111000111011001111;
assign LUT_4[36409] = 32'b11111111111111110010000111000111;
assign LUT_4[36410] = 32'b11111111111111111000010101110011;
assign LUT_4[36411] = 32'b11111111111111110001100001101011;
assign LUT_4[36412] = 32'b11111111111111110101111011101011;
assign LUT_4[36413] = 32'b11111111111111101111000111100011;
assign LUT_4[36414] = 32'b11111111111111110101010110001111;
assign LUT_4[36415] = 32'b11111111111111101110100010000111;
assign LUT_4[36416] = 32'b00000000000000000100111001011001;
assign LUT_4[36417] = 32'b11111111111111111110000101010001;
assign LUT_4[36418] = 32'b00000000000000000100010011111101;
assign LUT_4[36419] = 32'b11111111111111111101011111110101;
assign LUT_4[36420] = 32'b00000000000000000001111001110101;
assign LUT_4[36421] = 32'b11111111111111111011000101101101;
assign LUT_4[36422] = 32'b00000000000000000001010100011001;
assign LUT_4[36423] = 32'b11111111111111111010100000010001;
assign LUT_4[36424] = 32'b11111111111111111110000101101110;
assign LUT_4[36425] = 32'b11111111111111110111010001100110;
assign LUT_4[36426] = 32'b11111111111111111101100000010010;
assign LUT_4[36427] = 32'b11111111111111110110101100001010;
assign LUT_4[36428] = 32'b11111111111111111011000110001010;
assign LUT_4[36429] = 32'b11111111111111110100010010000010;
assign LUT_4[36430] = 32'b11111111111111111010100000101110;
assign LUT_4[36431] = 32'b11111111111111110011101100100110;
assign LUT_4[36432] = 32'b00000000000000000010101011000111;
assign LUT_4[36433] = 32'b11111111111111111011110110111111;
assign LUT_4[36434] = 32'b00000000000000000010000101101011;
assign LUT_4[36435] = 32'b11111111111111111011010001100011;
assign LUT_4[36436] = 32'b11111111111111111111101011100011;
assign LUT_4[36437] = 32'b11111111111111111000110111011011;
assign LUT_4[36438] = 32'b11111111111111111111000110000111;
assign LUT_4[36439] = 32'b11111111111111111000010001111111;
assign LUT_4[36440] = 32'b11111111111111111011110111011100;
assign LUT_4[36441] = 32'b11111111111111110101000011010100;
assign LUT_4[36442] = 32'b11111111111111111011010010000000;
assign LUT_4[36443] = 32'b11111111111111110100011101111000;
assign LUT_4[36444] = 32'b11111111111111111000110111111000;
assign LUT_4[36445] = 32'b11111111111111110010000011110000;
assign LUT_4[36446] = 32'b11111111111111111000010010011100;
assign LUT_4[36447] = 32'b11111111111111110001011110010100;
assign LUT_4[36448] = 32'b00000000000000000011010100100000;
assign LUT_4[36449] = 32'b11111111111111111100100000011000;
assign LUT_4[36450] = 32'b00000000000000000010101111000100;
assign LUT_4[36451] = 32'b11111111111111111011111010111100;
assign LUT_4[36452] = 32'b00000000000000000000010100111100;
assign LUT_4[36453] = 32'b11111111111111111001100000110100;
assign LUT_4[36454] = 32'b11111111111111111111101111100000;
assign LUT_4[36455] = 32'b11111111111111111000111011011000;
assign LUT_4[36456] = 32'b11111111111111111100100000110101;
assign LUT_4[36457] = 32'b11111111111111110101101100101101;
assign LUT_4[36458] = 32'b11111111111111111011111011011001;
assign LUT_4[36459] = 32'b11111111111111110101000111010001;
assign LUT_4[36460] = 32'b11111111111111111001100001010001;
assign LUT_4[36461] = 32'b11111111111111110010101101001001;
assign LUT_4[36462] = 32'b11111111111111111000111011110101;
assign LUT_4[36463] = 32'b11111111111111110010000111101101;
assign LUT_4[36464] = 32'b00000000000000000001000110001110;
assign LUT_4[36465] = 32'b11111111111111111010010010000110;
assign LUT_4[36466] = 32'b00000000000000000000100000110010;
assign LUT_4[36467] = 32'b11111111111111111001101100101010;
assign LUT_4[36468] = 32'b11111111111111111110000110101010;
assign LUT_4[36469] = 32'b11111111111111110111010010100010;
assign LUT_4[36470] = 32'b11111111111111111101100001001110;
assign LUT_4[36471] = 32'b11111111111111110110101101000110;
assign LUT_4[36472] = 32'b11111111111111111010010010100011;
assign LUT_4[36473] = 32'b11111111111111110011011110011011;
assign LUT_4[36474] = 32'b11111111111111111001101101000111;
assign LUT_4[36475] = 32'b11111111111111110010111000111111;
assign LUT_4[36476] = 32'b11111111111111110111010010111111;
assign LUT_4[36477] = 32'b11111111111111110000011110110111;
assign LUT_4[36478] = 32'b11111111111111110110101101100011;
assign LUT_4[36479] = 32'b11111111111111101111111001011011;
assign LUT_4[36480] = 32'b00000000000000000110001000001101;
assign LUT_4[36481] = 32'b11111111111111111111010100000101;
assign LUT_4[36482] = 32'b00000000000000000101100010110001;
assign LUT_4[36483] = 32'b11111111111111111110101110101001;
assign LUT_4[36484] = 32'b00000000000000000011001000101001;
assign LUT_4[36485] = 32'b11111111111111111100010100100001;
assign LUT_4[36486] = 32'b00000000000000000010100011001101;
assign LUT_4[36487] = 32'b11111111111111111011101111000101;
assign LUT_4[36488] = 32'b11111111111111111111010100100010;
assign LUT_4[36489] = 32'b11111111111111111000100000011010;
assign LUT_4[36490] = 32'b11111111111111111110101111000110;
assign LUT_4[36491] = 32'b11111111111111110111111010111110;
assign LUT_4[36492] = 32'b11111111111111111100010100111110;
assign LUT_4[36493] = 32'b11111111111111110101100000110110;
assign LUT_4[36494] = 32'b11111111111111111011101111100010;
assign LUT_4[36495] = 32'b11111111111111110100111011011010;
assign LUT_4[36496] = 32'b00000000000000000011111001111011;
assign LUT_4[36497] = 32'b11111111111111111101000101110011;
assign LUT_4[36498] = 32'b00000000000000000011010100011111;
assign LUT_4[36499] = 32'b11111111111111111100100000010111;
assign LUT_4[36500] = 32'b00000000000000000000111010010111;
assign LUT_4[36501] = 32'b11111111111111111010000110001111;
assign LUT_4[36502] = 32'b00000000000000000000010100111011;
assign LUT_4[36503] = 32'b11111111111111111001100000110011;
assign LUT_4[36504] = 32'b11111111111111111101000110010000;
assign LUT_4[36505] = 32'b11111111111111110110010010001000;
assign LUT_4[36506] = 32'b11111111111111111100100000110100;
assign LUT_4[36507] = 32'b11111111111111110101101100101100;
assign LUT_4[36508] = 32'b11111111111111111010000110101100;
assign LUT_4[36509] = 32'b11111111111111110011010010100100;
assign LUT_4[36510] = 32'b11111111111111111001100001010000;
assign LUT_4[36511] = 32'b11111111111111110010101101001000;
assign LUT_4[36512] = 32'b00000000000000000100100011010100;
assign LUT_4[36513] = 32'b11111111111111111101101111001100;
assign LUT_4[36514] = 32'b00000000000000000011111101111000;
assign LUT_4[36515] = 32'b11111111111111111101001001110000;
assign LUT_4[36516] = 32'b00000000000000000001100011110000;
assign LUT_4[36517] = 32'b11111111111111111010101111101000;
assign LUT_4[36518] = 32'b00000000000000000000111110010100;
assign LUT_4[36519] = 32'b11111111111111111010001010001100;
assign LUT_4[36520] = 32'b11111111111111111101101111101001;
assign LUT_4[36521] = 32'b11111111111111110110111011100001;
assign LUT_4[36522] = 32'b11111111111111111101001010001101;
assign LUT_4[36523] = 32'b11111111111111110110010110000101;
assign LUT_4[36524] = 32'b11111111111111111010110000000101;
assign LUT_4[36525] = 32'b11111111111111110011111011111101;
assign LUT_4[36526] = 32'b11111111111111111010001010101001;
assign LUT_4[36527] = 32'b11111111111111110011010110100001;
assign LUT_4[36528] = 32'b00000000000000000010010101000010;
assign LUT_4[36529] = 32'b11111111111111111011100000111010;
assign LUT_4[36530] = 32'b00000000000000000001101111100110;
assign LUT_4[36531] = 32'b11111111111111111010111011011110;
assign LUT_4[36532] = 32'b11111111111111111111010101011110;
assign LUT_4[36533] = 32'b11111111111111111000100001010110;
assign LUT_4[36534] = 32'b11111111111111111110110000000010;
assign LUT_4[36535] = 32'b11111111111111110111111011111010;
assign LUT_4[36536] = 32'b11111111111111111011100001010111;
assign LUT_4[36537] = 32'b11111111111111110100101101001111;
assign LUT_4[36538] = 32'b11111111111111111010111011111011;
assign LUT_4[36539] = 32'b11111111111111110100000111110011;
assign LUT_4[36540] = 32'b11111111111111111000100001110011;
assign LUT_4[36541] = 32'b11111111111111110001101101101011;
assign LUT_4[36542] = 32'b11111111111111110111111100010111;
assign LUT_4[36543] = 32'b11111111111111110001001000001111;
assign LUT_4[36544] = 32'b00000000000000000111011111100001;
assign LUT_4[36545] = 32'b00000000000000000000101011011001;
assign LUT_4[36546] = 32'b00000000000000000110111010000101;
assign LUT_4[36547] = 32'b00000000000000000000000101111101;
assign LUT_4[36548] = 32'b00000000000000000100011111111101;
assign LUT_4[36549] = 32'b11111111111111111101101011110101;
assign LUT_4[36550] = 32'b00000000000000000011111010100001;
assign LUT_4[36551] = 32'b11111111111111111101000110011001;
assign LUT_4[36552] = 32'b00000000000000000000101011110110;
assign LUT_4[36553] = 32'b11111111111111111001110111101110;
assign LUT_4[36554] = 32'b00000000000000000000000110011010;
assign LUT_4[36555] = 32'b11111111111111111001010010010010;
assign LUT_4[36556] = 32'b11111111111111111101101100010010;
assign LUT_4[36557] = 32'b11111111111111110110111000001010;
assign LUT_4[36558] = 32'b11111111111111111101000110110110;
assign LUT_4[36559] = 32'b11111111111111110110010010101110;
assign LUT_4[36560] = 32'b00000000000000000101010001001111;
assign LUT_4[36561] = 32'b11111111111111111110011101000111;
assign LUT_4[36562] = 32'b00000000000000000100101011110011;
assign LUT_4[36563] = 32'b11111111111111111101110111101011;
assign LUT_4[36564] = 32'b00000000000000000010010001101011;
assign LUT_4[36565] = 32'b11111111111111111011011101100011;
assign LUT_4[36566] = 32'b00000000000000000001101100001111;
assign LUT_4[36567] = 32'b11111111111111111010111000000111;
assign LUT_4[36568] = 32'b11111111111111111110011101100100;
assign LUT_4[36569] = 32'b11111111111111110111101001011100;
assign LUT_4[36570] = 32'b11111111111111111101111000001000;
assign LUT_4[36571] = 32'b11111111111111110111000100000000;
assign LUT_4[36572] = 32'b11111111111111111011011110000000;
assign LUT_4[36573] = 32'b11111111111111110100101001111000;
assign LUT_4[36574] = 32'b11111111111111111010111000100100;
assign LUT_4[36575] = 32'b11111111111111110100000100011100;
assign LUT_4[36576] = 32'b00000000000000000101111010101000;
assign LUT_4[36577] = 32'b11111111111111111111000110100000;
assign LUT_4[36578] = 32'b00000000000000000101010101001100;
assign LUT_4[36579] = 32'b11111111111111111110100001000100;
assign LUT_4[36580] = 32'b00000000000000000010111011000100;
assign LUT_4[36581] = 32'b11111111111111111100000110111100;
assign LUT_4[36582] = 32'b00000000000000000010010101101000;
assign LUT_4[36583] = 32'b11111111111111111011100001100000;
assign LUT_4[36584] = 32'b11111111111111111111000110111101;
assign LUT_4[36585] = 32'b11111111111111111000010010110101;
assign LUT_4[36586] = 32'b11111111111111111110100001100001;
assign LUT_4[36587] = 32'b11111111111111110111101101011001;
assign LUT_4[36588] = 32'b11111111111111111100000111011001;
assign LUT_4[36589] = 32'b11111111111111110101010011010001;
assign LUT_4[36590] = 32'b11111111111111111011100001111101;
assign LUT_4[36591] = 32'b11111111111111110100101101110101;
assign LUT_4[36592] = 32'b00000000000000000011101100010110;
assign LUT_4[36593] = 32'b11111111111111111100111000001110;
assign LUT_4[36594] = 32'b00000000000000000011000110111010;
assign LUT_4[36595] = 32'b11111111111111111100010010110010;
assign LUT_4[36596] = 32'b00000000000000000000101100110010;
assign LUT_4[36597] = 32'b11111111111111111001111000101010;
assign LUT_4[36598] = 32'b00000000000000000000000111010110;
assign LUT_4[36599] = 32'b11111111111111111001010011001110;
assign LUT_4[36600] = 32'b11111111111111111100111000101011;
assign LUT_4[36601] = 32'b11111111111111110110000100100011;
assign LUT_4[36602] = 32'b11111111111111111100010011001111;
assign LUT_4[36603] = 32'b11111111111111110101011111000111;
assign LUT_4[36604] = 32'b11111111111111111001111001000111;
assign LUT_4[36605] = 32'b11111111111111110011000100111111;
assign LUT_4[36606] = 32'b11111111111111111001010011101011;
assign LUT_4[36607] = 32'b11111111111111110010011111100011;
assign LUT_4[36608] = 32'b00000000000000001000011101101000;
assign LUT_4[36609] = 32'b00000000000000000001101001100000;
assign LUT_4[36610] = 32'b00000000000000000111111000001100;
assign LUT_4[36611] = 32'b00000000000000000001000100000100;
assign LUT_4[36612] = 32'b00000000000000000101011110000100;
assign LUT_4[36613] = 32'b11111111111111111110101001111100;
assign LUT_4[36614] = 32'b00000000000000000100111000101000;
assign LUT_4[36615] = 32'b11111111111111111110000100100000;
assign LUT_4[36616] = 32'b00000000000000000001101001111101;
assign LUT_4[36617] = 32'b11111111111111111010110101110101;
assign LUT_4[36618] = 32'b00000000000000000001000100100001;
assign LUT_4[36619] = 32'b11111111111111111010010000011001;
assign LUT_4[36620] = 32'b11111111111111111110101010011001;
assign LUT_4[36621] = 32'b11111111111111110111110110010001;
assign LUT_4[36622] = 32'b11111111111111111110000100111101;
assign LUT_4[36623] = 32'b11111111111111110111010000110101;
assign LUT_4[36624] = 32'b00000000000000000110001111010110;
assign LUT_4[36625] = 32'b11111111111111111111011011001110;
assign LUT_4[36626] = 32'b00000000000000000101101001111010;
assign LUT_4[36627] = 32'b11111111111111111110110101110010;
assign LUT_4[36628] = 32'b00000000000000000011001111110010;
assign LUT_4[36629] = 32'b11111111111111111100011011101010;
assign LUT_4[36630] = 32'b00000000000000000010101010010110;
assign LUT_4[36631] = 32'b11111111111111111011110110001110;
assign LUT_4[36632] = 32'b11111111111111111111011011101011;
assign LUT_4[36633] = 32'b11111111111111111000100111100011;
assign LUT_4[36634] = 32'b11111111111111111110110110001111;
assign LUT_4[36635] = 32'b11111111111111111000000010000111;
assign LUT_4[36636] = 32'b11111111111111111100011100000111;
assign LUT_4[36637] = 32'b11111111111111110101100111111111;
assign LUT_4[36638] = 32'b11111111111111111011110110101011;
assign LUT_4[36639] = 32'b11111111111111110101000010100011;
assign LUT_4[36640] = 32'b00000000000000000110111000101111;
assign LUT_4[36641] = 32'b00000000000000000000000100100111;
assign LUT_4[36642] = 32'b00000000000000000110010011010011;
assign LUT_4[36643] = 32'b11111111111111111111011111001011;
assign LUT_4[36644] = 32'b00000000000000000011111001001011;
assign LUT_4[36645] = 32'b11111111111111111101000101000011;
assign LUT_4[36646] = 32'b00000000000000000011010011101111;
assign LUT_4[36647] = 32'b11111111111111111100011111100111;
assign LUT_4[36648] = 32'b00000000000000000000000101000100;
assign LUT_4[36649] = 32'b11111111111111111001010000111100;
assign LUT_4[36650] = 32'b11111111111111111111011111101000;
assign LUT_4[36651] = 32'b11111111111111111000101011100000;
assign LUT_4[36652] = 32'b11111111111111111101000101100000;
assign LUT_4[36653] = 32'b11111111111111110110010001011000;
assign LUT_4[36654] = 32'b11111111111111111100100000000100;
assign LUT_4[36655] = 32'b11111111111111110101101011111100;
assign LUT_4[36656] = 32'b00000000000000000100101010011101;
assign LUT_4[36657] = 32'b11111111111111111101110110010101;
assign LUT_4[36658] = 32'b00000000000000000100000101000001;
assign LUT_4[36659] = 32'b11111111111111111101010000111001;
assign LUT_4[36660] = 32'b00000000000000000001101010111001;
assign LUT_4[36661] = 32'b11111111111111111010110110110001;
assign LUT_4[36662] = 32'b00000000000000000001000101011101;
assign LUT_4[36663] = 32'b11111111111111111010010001010101;
assign LUT_4[36664] = 32'b11111111111111111101110110110010;
assign LUT_4[36665] = 32'b11111111111111110111000010101010;
assign LUT_4[36666] = 32'b11111111111111111101010001010110;
assign LUT_4[36667] = 32'b11111111111111110110011101001110;
assign LUT_4[36668] = 32'b11111111111111111010110111001110;
assign LUT_4[36669] = 32'b11111111111111110100000011000110;
assign LUT_4[36670] = 32'b11111111111111111010010001110010;
assign LUT_4[36671] = 32'b11111111111111110011011101101010;
assign LUT_4[36672] = 32'b00000000000000001001110100111100;
assign LUT_4[36673] = 32'b00000000000000000011000000110100;
assign LUT_4[36674] = 32'b00000000000000001001001111100000;
assign LUT_4[36675] = 32'b00000000000000000010011011011000;
assign LUT_4[36676] = 32'b00000000000000000110110101011000;
assign LUT_4[36677] = 32'b00000000000000000000000001010000;
assign LUT_4[36678] = 32'b00000000000000000110001111111100;
assign LUT_4[36679] = 32'b11111111111111111111011011110100;
assign LUT_4[36680] = 32'b00000000000000000011000001010001;
assign LUT_4[36681] = 32'b11111111111111111100001101001001;
assign LUT_4[36682] = 32'b00000000000000000010011011110101;
assign LUT_4[36683] = 32'b11111111111111111011100111101101;
assign LUT_4[36684] = 32'b00000000000000000000000001101101;
assign LUT_4[36685] = 32'b11111111111111111001001101100101;
assign LUT_4[36686] = 32'b11111111111111111111011100010001;
assign LUT_4[36687] = 32'b11111111111111111000101000001001;
assign LUT_4[36688] = 32'b00000000000000000111100110101010;
assign LUT_4[36689] = 32'b00000000000000000000110010100010;
assign LUT_4[36690] = 32'b00000000000000000111000001001110;
assign LUT_4[36691] = 32'b00000000000000000000001101000110;
assign LUT_4[36692] = 32'b00000000000000000100100111000110;
assign LUT_4[36693] = 32'b11111111111111111101110010111110;
assign LUT_4[36694] = 32'b00000000000000000100000001101010;
assign LUT_4[36695] = 32'b11111111111111111101001101100010;
assign LUT_4[36696] = 32'b00000000000000000000110010111111;
assign LUT_4[36697] = 32'b11111111111111111001111110110111;
assign LUT_4[36698] = 32'b00000000000000000000001101100011;
assign LUT_4[36699] = 32'b11111111111111111001011001011011;
assign LUT_4[36700] = 32'b11111111111111111101110011011011;
assign LUT_4[36701] = 32'b11111111111111110110111111010011;
assign LUT_4[36702] = 32'b11111111111111111101001101111111;
assign LUT_4[36703] = 32'b11111111111111110110011001110111;
assign LUT_4[36704] = 32'b00000000000000001000010000000011;
assign LUT_4[36705] = 32'b00000000000000000001011011111011;
assign LUT_4[36706] = 32'b00000000000000000111101010100111;
assign LUT_4[36707] = 32'b00000000000000000000110110011111;
assign LUT_4[36708] = 32'b00000000000000000101010000011111;
assign LUT_4[36709] = 32'b11111111111111111110011100010111;
assign LUT_4[36710] = 32'b00000000000000000100101011000011;
assign LUT_4[36711] = 32'b11111111111111111101110110111011;
assign LUT_4[36712] = 32'b00000000000000000001011100011000;
assign LUT_4[36713] = 32'b11111111111111111010101000010000;
assign LUT_4[36714] = 32'b00000000000000000000110110111100;
assign LUT_4[36715] = 32'b11111111111111111010000010110100;
assign LUT_4[36716] = 32'b11111111111111111110011100110100;
assign LUT_4[36717] = 32'b11111111111111110111101000101100;
assign LUT_4[36718] = 32'b11111111111111111101110111011000;
assign LUT_4[36719] = 32'b11111111111111110111000011010000;
assign LUT_4[36720] = 32'b00000000000000000110000001110001;
assign LUT_4[36721] = 32'b11111111111111111111001101101001;
assign LUT_4[36722] = 32'b00000000000000000101011100010101;
assign LUT_4[36723] = 32'b11111111111111111110101000001101;
assign LUT_4[36724] = 32'b00000000000000000011000010001101;
assign LUT_4[36725] = 32'b11111111111111111100001110000101;
assign LUT_4[36726] = 32'b00000000000000000010011100110001;
assign LUT_4[36727] = 32'b11111111111111111011101000101001;
assign LUT_4[36728] = 32'b11111111111111111111001110000110;
assign LUT_4[36729] = 32'b11111111111111111000011001111110;
assign LUT_4[36730] = 32'b11111111111111111110101000101010;
assign LUT_4[36731] = 32'b11111111111111110111110100100010;
assign LUT_4[36732] = 32'b11111111111111111100001110100010;
assign LUT_4[36733] = 32'b11111111111111110101011010011010;
assign LUT_4[36734] = 32'b11111111111111111011101001000110;
assign LUT_4[36735] = 32'b11111111111111110100110100111110;
assign LUT_4[36736] = 32'b00000000000000001011000011110000;
assign LUT_4[36737] = 32'b00000000000000000100001111101000;
assign LUT_4[36738] = 32'b00000000000000001010011110010100;
assign LUT_4[36739] = 32'b00000000000000000011101010001100;
assign LUT_4[36740] = 32'b00000000000000001000000100001100;
assign LUT_4[36741] = 32'b00000000000000000001010000000100;
assign LUT_4[36742] = 32'b00000000000000000111011110110000;
assign LUT_4[36743] = 32'b00000000000000000000101010101000;
assign LUT_4[36744] = 32'b00000000000000000100010000000101;
assign LUT_4[36745] = 32'b11111111111111111101011011111101;
assign LUT_4[36746] = 32'b00000000000000000011101010101001;
assign LUT_4[36747] = 32'b11111111111111111100110110100001;
assign LUT_4[36748] = 32'b00000000000000000001010000100001;
assign LUT_4[36749] = 32'b11111111111111111010011100011001;
assign LUT_4[36750] = 32'b00000000000000000000101011000101;
assign LUT_4[36751] = 32'b11111111111111111001110110111101;
assign LUT_4[36752] = 32'b00000000000000001000110101011110;
assign LUT_4[36753] = 32'b00000000000000000010000001010110;
assign LUT_4[36754] = 32'b00000000000000001000010000000010;
assign LUT_4[36755] = 32'b00000000000000000001011011111010;
assign LUT_4[36756] = 32'b00000000000000000101110101111010;
assign LUT_4[36757] = 32'b11111111111111111111000001110010;
assign LUT_4[36758] = 32'b00000000000000000101010000011110;
assign LUT_4[36759] = 32'b11111111111111111110011100010110;
assign LUT_4[36760] = 32'b00000000000000000010000001110011;
assign LUT_4[36761] = 32'b11111111111111111011001101101011;
assign LUT_4[36762] = 32'b00000000000000000001011100010111;
assign LUT_4[36763] = 32'b11111111111111111010101000001111;
assign LUT_4[36764] = 32'b11111111111111111111000010001111;
assign LUT_4[36765] = 32'b11111111111111111000001110000111;
assign LUT_4[36766] = 32'b11111111111111111110011100110011;
assign LUT_4[36767] = 32'b11111111111111110111101000101011;
assign LUT_4[36768] = 32'b00000000000000001001011110110111;
assign LUT_4[36769] = 32'b00000000000000000010101010101111;
assign LUT_4[36770] = 32'b00000000000000001000111001011011;
assign LUT_4[36771] = 32'b00000000000000000010000101010011;
assign LUT_4[36772] = 32'b00000000000000000110011111010011;
assign LUT_4[36773] = 32'b11111111111111111111101011001011;
assign LUT_4[36774] = 32'b00000000000000000101111001110111;
assign LUT_4[36775] = 32'b11111111111111111111000101101111;
assign LUT_4[36776] = 32'b00000000000000000010101011001100;
assign LUT_4[36777] = 32'b11111111111111111011110111000100;
assign LUT_4[36778] = 32'b00000000000000000010000101110000;
assign LUT_4[36779] = 32'b11111111111111111011010001101000;
assign LUT_4[36780] = 32'b11111111111111111111101011101000;
assign LUT_4[36781] = 32'b11111111111111111000110111100000;
assign LUT_4[36782] = 32'b11111111111111111111000110001100;
assign LUT_4[36783] = 32'b11111111111111111000010010000100;
assign LUT_4[36784] = 32'b00000000000000000111010000100101;
assign LUT_4[36785] = 32'b00000000000000000000011100011101;
assign LUT_4[36786] = 32'b00000000000000000110101011001001;
assign LUT_4[36787] = 32'b11111111111111111111110111000001;
assign LUT_4[36788] = 32'b00000000000000000100010001000001;
assign LUT_4[36789] = 32'b11111111111111111101011100111001;
assign LUT_4[36790] = 32'b00000000000000000011101011100101;
assign LUT_4[36791] = 32'b11111111111111111100110111011101;
assign LUT_4[36792] = 32'b00000000000000000000011100111010;
assign LUT_4[36793] = 32'b11111111111111111001101000110010;
assign LUT_4[36794] = 32'b11111111111111111111110111011110;
assign LUT_4[36795] = 32'b11111111111111111001000011010110;
assign LUT_4[36796] = 32'b11111111111111111101011101010110;
assign LUT_4[36797] = 32'b11111111111111110110101001001110;
assign LUT_4[36798] = 32'b11111111111111111100110111111010;
assign LUT_4[36799] = 32'b11111111111111110110000011110010;
assign LUT_4[36800] = 32'b00000000000000001100011011000100;
assign LUT_4[36801] = 32'b00000000000000000101100110111100;
assign LUT_4[36802] = 32'b00000000000000001011110101101000;
assign LUT_4[36803] = 32'b00000000000000000101000001100000;
assign LUT_4[36804] = 32'b00000000000000001001011011100000;
assign LUT_4[36805] = 32'b00000000000000000010100111011000;
assign LUT_4[36806] = 32'b00000000000000001000110110000100;
assign LUT_4[36807] = 32'b00000000000000000010000001111100;
assign LUT_4[36808] = 32'b00000000000000000101100111011001;
assign LUT_4[36809] = 32'b11111111111111111110110011010001;
assign LUT_4[36810] = 32'b00000000000000000101000001111101;
assign LUT_4[36811] = 32'b11111111111111111110001101110101;
assign LUT_4[36812] = 32'b00000000000000000010100111110101;
assign LUT_4[36813] = 32'b11111111111111111011110011101101;
assign LUT_4[36814] = 32'b00000000000000000010000010011001;
assign LUT_4[36815] = 32'b11111111111111111011001110010001;
assign LUT_4[36816] = 32'b00000000000000001010001100110010;
assign LUT_4[36817] = 32'b00000000000000000011011000101010;
assign LUT_4[36818] = 32'b00000000000000001001100111010110;
assign LUT_4[36819] = 32'b00000000000000000010110011001110;
assign LUT_4[36820] = 32'b00000000000000000111001101001110;
assign LUT_4[36821] = 32'b00000000000000000000011001000110;
assign LUT_4[36822] = 32'b00000000000000000110100111110010;
assign LUT_4[36823] = 32'b11111111111111111111110011101010;
assign LUT_4[36824] = 32'b00000000000000000011011001000111;
assign LUT_4[36825] = 32'b11111111111111111100100100111111;
assign LUT_4[36826] = 32'b00000000000000000010110011101011;
assign LUT_4[36827] = 32'b11111111111111111011111111100011;
assign LUT_4[36828] = 32'b00000000000000000000011001100011;
assign LUT_4[36829] = 32'b11111111111111111001100101011011;
assign LUT_4[36830] = 32'b11111111111111111111110100000111;
assign LUT_4[36831] = 32'b11111111111111111000111111111111;
assign LUT_4[36832] = 32'b00000000000000001010110110001011;
assign LUT_4[36833] = 32'b00000000000000000100000010000011;
assign LUT_4[36834] = 32'b00000000000000001010010000101111;
assign LUT_4[36835] = 32'b00000000000000000011011100100111;
assign LUT_4[36836] = 32'b00000000000000000111110110100111;
assign LUT_4[36837] = 32'b00000000000000000001000010011111;
assign LUT_4[36838] = 32'b00000000000000000111010001001011;
assign LUT_4[36839] = 32'b00000000000000000000011101000011;
assign LUT_4[36840] = 32'b00000000000000000100000010100000;
assign LUT_4[36841] = 32'b11111111111111111101001110011000;
assign LUT_4[36842] = 32'b00000000000000000011011101000100;
assign LUT_4[36843] = 32'b11111111111111111100101000111100;
assign LUT_4[36844] = 32'b00000000000000000001000010111100;
assign LUT_4[36845] = 32'b11111111111111111010001110110100;
assign LUT_4[36846] = 32'b00000000000000000000011101100000;
assign LUT_4[36847] = 32'b11111111111111111001101001011000;
assign LUT_4[36848] = 32'b00000000000000001000100111111001;
assign LUT_4[36849] = 32'b00000000000000000001110011110001;
assign LUT_4[36850] = 32'b00000000000000001000000010011101;
assign LUT_4[36851] = 32'b00000000000000000001001110010101;
assign LUT_4[36852] = 32'b00000000000000000101101000010101;
assign LUT_4[36853] = 32'b11111111111111111110110100001101;
assign LUT_4[36854] = 32'b00000000000000000101000010111001;
assign LUT_4[36855] = 32'b11111111111111111110001110110001;
assign LUT_4[36856] = 32'b00000000000000000001110100001110;
assign LUT_4[36857] = 32'b11111111111111111011000000000110;
assign LUT_4[36858] = 32'b00000000000000000001001110110010;
assign LUT_4[36859] = 32'b11111111111111111010011010101010;
assign LUT_4[36860] = 32'b11111111111111111110110100101010;
assign LUT_4[36861] = 32'b11111111111111111000000000100010;
assign LUT_4[36862] = 32'b11111111111111111110001111001110;
assign LUT_4[36863] = 32'b11111111111111110111011011000110;
assign LUT_4[36864] = 32'b00000000000000000011100100000101;
assign LUT_4[36865] = 32'b11111111111111111100101111111101;
assign LUT_4[36866] = 32'b00000000000000000010111110101001;
assign LUT_4[36867] = 32'b11111111111111111100001010100001;
assign LUT_4[36868] = 32'b00000000000000000000100100100001;
assign LUT_4[36869] = 32'b11111111111111111001110000011001;
assign LUT_4[36870] = 32'b11111111111111111111111111000101;
assign LUT_4[36871] = 32'b11111111111111111001001010111101;
assign LUT_4[36872] = 32'b11111111111111111100110000011010;
assign LUT_4[36873] = 32'b11111111111111110101111100010010;
assign LUT_4[36874] = 32'b11111111111111111100001010111110;
assign LUT_4[36875] = 32'b11111111111111110101010110110110;
assign LUT_4[36876] = 32'b11111111111111111001110000110110;
assign LUT_4[36877] = 32'b11111111111111110010111100101110;
assign LUT_4[36878] = 32'b11111111111111111001001011011010;
assign LUT_4[36879] = 32'b11111111111111110010010111010010;
assign LUT_4[36880] = 32'b00000000000000000001010101110011;
assign LUT_4[36881] = 32'b11111111111111111010100001101011;
assign LUT_4[36882] = 32'b00000000000000000000110000010111;
assign LUT_4[36883] = 32'b11111111111111111001111100001111;
assign LUT_4[36884] = 32'b11111111111111111110010110001111;
assign LUT_4[36885] = 32'b11111111111111110111100010000111;
assign LUT_4[36886] = 32'b11111111111111111101110000110011;
assign LUT_4[36887] = 32'b11111111111111110110111100101011;
assign LUT_4[36888] = 32'b11111111111111111010100010001000;
assign LUT_4[36889] = 32'b11111111111111110011101110000000;
assign LUT_4[36890] = 32'b11111111111111111001111100101100;
assign LUT_4[36891] = 32'b11111111111111110011001000100100;
assign LUT_4[36892] = 32'b11111111111111110111100010100100;
assign LUT_4[36893] = 32'b11111111111111110000101110011100;
assign LUT_4[36894] = 32'b11111111111111110110111101001000;
assign LUT_4[36895] = 32'b11111111111111110000001001000000;
assign LUT_4[36896] = 32'b00000000000000000001111111001100;
assign LUT_4[36897] = 32'b11111111111111111011001011000100;
assign LUT_4[36898] = 32'b00000000000000000001011001110000;
assign LUT_4[36899] = 32'b11111111111111111010100101101000;
assign LUT_4[36900] = 32'b11111111111111111110111111101000;
assign LUT_4[36901] = 32'b11111111111111111000001011100000;
assign LUT_4[36902] = 32'b11111111111111111110011010001100;
assign LUT_4[36903] = 32'b11111111111111110111100110000100;
assign LUT_4[36904] = 32'b11111111111111111011001011100001;
assign LUT_4[36905] = 32'b11111111111111110100010111011001;
assign LUT_4[36906] = 32'b11111111111111111010100110000101;
assign LUT_4[36907] = 32'b11111111111111110011110001111101;
assign LUT_4[36908] = 32'b11111111111111111000001011111101;
assign LUT_4[36909] = 32'b11111111111111110001010111110101;
assign LUT_4[36910] = 32'b11111111111111110111100110100001;
assign LUT_4[36911] = 32'b11111111111111110000110010011001;
assign LUT_4[36912] = 32'b11111111111111111111110000111010;
assign LUT_4[36913] = 32'b11111111111111111000111100110010;
assign LUT_4[36914] = 32'b11111111111111111111001011011110;
assign LUT_4[36915] = 32'b11111111111111111000010111010110;
assign LUT_4[36916] = 32'b11111111111111111100110001010110;
assign LUT_4[36917] = 32'b11111111111111110101111101001110;
assign LUT_4[36918] = 32'b11111111111111111100001011111010;
assign LUT_4[36919] = 32'b11111111111111110101010111110010;
assign LUT_4[36920] = 32'b11111111111111111000111101001111;
assign LUT_4[36921] = 32'b11111111111111110010001001000111;
assign LUT_4[36922] = 32'b11111111111111111000010111110011;
assign LUT_4[36923] = 32'b11111111111111110001100011101011;
assign LUT_4[36924] = 32'b11111111111111110101111101101011;
assign LUT_4[36925] = 32'b11111111111111101111001001100011;
assign LUT_4[36926] = 32'b11111111111111110101011000001111;
assign LUT_4[36927] = 32'b11111111111111101110100100000111;
assign LUT_4[36928] = 32'b00000000000000000100111011011001;
assign LUT_4[36929] = 32'b11111111111111111110000111010001;
assign LUT_4[36930] = 32'b00000000000000000100010101111101;
assign LUT_4[36931] = 32'b11111111111111111101100001110101;
assign LUT_4[36932] = 32'b00000000000000000001111011110101;
assign LUT_4[36933] = 32'b11111111111111111011000111101101;
assign LUT_4[36934] = 32'b00000000000000000001010110011001;
assign LUT_4[36935] = 32'b11111111111111111010100010010001;
assign LUT_4[36936] = 32'b11111111111111111110000111101110;
assign LUT_4[36937] = 32'b11111111111111110111010011100110;
assign LUT_4[36938] = 32'b11111111111111111101100010010010;
assign LUT_4[36939] = 32'b11111111111111110110101110001010;
assign LUT_4[36940] = 32'b11111111111111111011001000001010;
assign LUT_4[36941] = 32'b11111111111111110100010100000010;
assign LUT_4[36942] = 32'b11111111111111111010100010101110;
assign LUT_4[36943] = 32'b11111111111111110011101110100110;
assign LUT_4[36944] = 32'b00000000000000000010101101000111;
assign LUT_4[36945] = 32'b11111111111111111011111000111111;
assign LUT_4[36946] = 32'b00000000000000000010000111101011;
assign LUT_4[36947] = 32'b11111111111111111011010011100011;
assign LUT_4[36948] = 32'b11111111111111111111101101100011;
assign LUT_4[36949] = 32'b11111111111111111000111001011011;
assign LUT_4[36950] = 32'b11111111111111111111001000000111;
assign LUT_4[36951] = 32'b11111111111111111000010011111111;
assign LUT_4[36952] = 32'b11111111111111111011111001011100;
assign LUT_4[36953] = 32'b11111111111111110101000101010100;
assign LUT_4[36954] = 32'b11111111111111111011010100000000;
assign LUT_4[36955] = 32'b11111111111111110100011111111000;
assign LUT_4[36956] = 32'b11111111111111111000111001111000;
assign LUT_4[36957] = 32'b11111111111111110010000101110000;
assign LUT_4[36958] = 32'b11111111111111111000010100011100;
assign LUT_4[36959] = 32'b11111111111111110001100000010100;
assign LUT_4[36960] = 32'b00000000000000000011010110100000;
assign LUT_4[36961] = 32'b11111111111111111100100010011000;
assign LUT_4[36962] = 32'b00000000000000000010110001000100;
assign LUT_4[36963] = 32'b11111111111111111011111100111100;
assign LUT_4[36964] = 32'b00000000000000000000010110111100;
assign LUT_4[36965] = 32'b11111111111111111001100010110100;
assign LUT_4[36966] = 32'b11111111111111111111110001100000;
assign LUT_4[36967] = 32'b11111111111111111000111101011000;
assign LUT_4[36968] = 32'b11111111111111111100100010110101;
assign LUT_4[36969] = 32'b11111111111111110101101110101101;
assign LUT_4[36970] = 32'b11111111111111111011111101011001;
assign LUT_4[36971] = 32'b11111111111111110101001001010001;
assign LUT_4[36972] = 32'b11111111111111111001100011010001;
assign LUT_4[36973] = 32'b11111111111111110010101111001001;
assign LUT_4[36974] = 32'b11111111111111111000111101110101;
assign LUT_4[36975] = 32'b11111111111111110010001001101101;
assign LUT_4[36976] = 32'b00000000000000000001001000001110;
assign LUT_4[36977] = 32'b11111111111111111010010100000110;
assign LUT_4[36978] = 32'b00000000000000000000100010110010;
assign LUT_4[36979] = 32'b11111111111111111001101110101010;
assign LUT_4[36980] = 32'b11111111111111111110001000101010;
assign LUT_4[36981] = 32'b11111111111111110111010100100010;
assign LUT_4[36982] = 32'b11111111111111111101100011001110;
assign LUT_4[36983] = 32'b11111111111111110110101111000110;
assign LUT_4[36984] = 32'b11111111111111111010010100100011;
assign LUT_4[36985] = 32'b11111111111111110011100000011011;
assign LUT_4[36986] = 32'b11111111111111111001101111000111;
assign LUT_4[36987] = 32'b11111111111111110010111010111111;
assign LUT_4[36988] = 32'b11111111111111110111010100111111;
assign LUT_4[36989] = 32'b11111111111111110000100000110111;
assign LUT_4[36990] = 32'b11111111111111110110101111100011;
assign LUT_4[36991] = 32'b11111111111111101111111011011011;
assign LUT_4[36992] = 32'b00000000000000000110001010001101;
assign LUT_4[36993] = 32'b11111111111111111111010110000101;
assign LUT_4[36994] = 32'b00000000000000000101100100110001;
assign LUT_4[36995] = 32'b11111111111111111110110000101001;
assign LUT_4[36996] = 32'b00000000000000000011001010101001;
assign LUT_4[36997] = 32'b11111111111111111100010110100001;
assign LUT_4[36998] = 32'b00000000000000000010100101001101;
assign LUT_4[36999] = 32'b11111111111111111011110001000101;
assign LUT_4[37000] = 32'b11111111111111111111010110100010;
assign LUT_4[37001] = 32'b11111111111111111000100010011010;
assign LUT_4[37002] = 32'b11111111111111111110110001000110;
assign LUT_4[37003] = 32'b11111111111111110111111100111110;
assign LUT_4[37004] = 32'b11111111111111111100010110111110;
assign LUT_4[37005] = 32'b11111111111111110101100010110110;
assign LUT_4[37006] = 32'b11111111111111111011110001100010;
assign LUT_4[37007] = 32'b11111111111111110100111101011010;
assign LUT_4[37008] = 32'b00000000000000000011111011111011;
assign LUT_4[37009] = 32'b11111111111111111101000111110011;
assign LUT_4[37010] = 32'b00000000000000000011010110011111;
assign LUT_4[37011] = 32'b11111111111111111100100010010111;
assign LUT_4[37012] = 32'b00000000000000000000111100010111;
assign LUT_4[37013] = 32'b11111111111111111010001000001111;
assign LUT_4[37014] = 32'b00000000000000000000010110111011;
assign LUT_4[37015] = 32'b11111111111111111001100010110011;
assign LUT_4[37016] = 32'b11111111111111111101001000010000;
assign LUT_4[37017] = 32'b11111111111111110110010100001000;
assign LUT_4[37018] = 32'b11111111111111111100100010110100;
assign LUT_4[37019] = 32'b11111111111111110101101110101100;
assign LUT_4[37020] = 32'b11111111111111111010001000101100;
assign LUT_4[37021] = 32'b11111111111111110011010100100100;
assign LUT_4[37022] = 32'b11111111111111111001100011010000;
assign LUT_4[37023] = 32'b11111111111111110010101111001000;
assign LUT_4[37024] = 32'b00000000000000000100100101010100;
assign LUT_4[37025] = 32'b11111111111111111101110001001100;
assign LUT_4[37026] = 32'b00000000000000000011111111111000;
assign LUT_4[37027] = 32'b11111111111111111101001011110000;
assign LUT_4[37028] = 32'b00000000000000000001100101110000;
assign LUT_4[37029] = 32'b11111111111111111010110001101000;
assign LUT_4[37030] = 32'b00000000000000000001000000010100;
assign LUT_4[37031] = 32'b11111111111111111010001100001100;
assign LUT_4[37032] = 32'b11111111111111111101110001101001;
assign LUT_4[37033] = 32'b11111111111111110110111101100001;
assign LUT_4[37034] = 32'b11111111111111111101001100001101;
assign LUT_4[37035] = 32'b11111111111111110110011000000101;
assign LUT_4[37036] = 32'b11111111111111111010110010000101;
assign LUT_4[37037] = 32'b11111111111111110011111101111101;
assign LUT_4[37038] = 32'b11111111111111111010001100101001;
assign LUT_4[37039] = 32'b11111111111111110011011000100001;
assign LUT_4[37040] = 32'b00000000000000000010010111000010;
assign LUT_4[37041] = 32'b11111111111111111011100010111010;
assign LUT_4[37042] = 32'b00000000000000000001110001100110;
assign LUT_4[37043] = 32'b11111111111111111010111101011110;
assign LUT_4[37044] = 32'b11111111111111111111010111011110;
assign LUT_4[37045] = 32'b11111111111111111000100011010110;
assign LUT_4[37046] = 32'b11111111111111111110110010000010;
assign LUT_4[37047] = 32'b11111111111111110111111101111010;
assign LUT_4[37048] = 32'b11111111111111111011100011010111;
assign LUT_4[37049] = 32'b11111111111111110100101111001111;
assign LUT_4[37050] = 32'b11111111111111111010111101111011;
assign LUT_4[37051] = 32'b11111111111111110100001001110011;
assign LUT_4[37052] = 32'b11111111111111111000100011110011;
assign LUT_4[37053] = 32'b11111111111111110001101111101011;
assign LUT_4[37054] = 32'b11111111111111110111111110010111;
assign LUT_4[37055] = 32'b11111111111111110001001010001111;
assign LUT_4[37056] = 32'b00000000000000000111100001100001;
assign LUT_4[37057] = 32'b00000000000000000000101101011001;
assign LUT_4[37058] = 32'b00000000000000000110111100000101;
assign LUT_4[37059] = 32'b00000000000000000000000111111101;
assign LUT_4[37060] = 32'b00000000000000000100100001111101;
assign LUT_4[37061] = 32'b11111111111111111101101101110101;
assign LUT_4[37062] = 32'b00000000000000000011111100100001;
assign LUT_4[37063] = 32'b11111111111111111101001000011001;
assign LUT_4[37064] = 32'b00000000000000000000101101110110;
assign LUT_4[37065] = 32'b11111111111111111001111001101110;
assign LUT_4[37066] = 32'b00000000000000000000001000011010;
assign LUT_4[37067] = 32'b11111111111111111001010100010010;
assign LUT_4[37068] = 32'b11111111111111111101101110010010;
assign LUT_4[37069] = 32'b11111111111111110110111010001010;
assign LUT_4[37070] = 32'b11111111111111111101001000110110;
assign LUT_4[37071] = 32'b11111111111111110110010100101110;
assign LUT_4[37072] = 32'b00000000000000000101010011001111;
assign LUT_4[37073] = 32'b11111111111111111110011111000111;
assign LUT_4[37074] = 32'b00000000000000000100101101110011;
assign LUT_4[37075] = 32'b11111111111111111101111001101011;
assign LUT_4[37076] = 32'b00000000000000000010010011101011;
assign LUT_4[37077] = 32'b11111111111111111011011111100011;
assign LUT_4[37078] = 32'b00000000000000000001101110001111;
assign LUT_4[37079] = 32'b11111111111111111010111010000111;
assign LUT_4[37080] = 32'b11111111111111111110011111100100;
assign LUT_4[37081] = 32'b11111111111111110111101011011100;
assign LUT_4[37082] = 32'b11111111111111111101111010001000;
assign LUT_4[37083] = 32'b11111111111111110111000110000000;
assign LUT_4[37084] = 32'b11111111111111111011100000000000;
assign LUT_4[37085] = 32'b11111111111111110100101011111000;
assign LUT_4[37086] = 32'b11111111111111111010111010100100;
assign LUT_4[37087] = 32'b11111111111111110100000110011100;
assign LUT_4[37088] = 32'b00000000000000000101111100101000;
assign LUT_4[37089] = 32'b11111111111111111111001000100000;
assign LUT_4[37090] = 32'b00000000000000000101010111001100;
assign LUT_4[37091] = 32'b11111111111111111110100011000100;
assign LUT_4[37092] = 32'b00000000000000000010111101000100;
assign LUT_4[37093] = 32'b11111111111111111100001000111100;
assign LUT_4[37094] = 32'b00000000000000000010010111101000;
assign LUT_4[37095] = 32'b11111111111111111011100011100000;
assign LUT_4[37096] = 32'b11111111111111111111001000111101;
assign LUT_4[37097] = 32'b11111111111111111000010100110101;
assign LUT_4[37098] = 32'b11111111111111111110100011100001;
assign LUT_4[37099] = 32'b11111111111111110111101111011001;
assign LUT_4[37100] = 32'b11111111111111111100001001011001;
assign LUT_4[37101] = 32'b11111111111111110101010101010001;
assign LUT_4[37102] = 32'b11111111111111111011100011111101;
assign LUT_4[37103] = 32'b11111111111111110100101111110101;
assign LUT_4[37104] = 32'b00000000000000000011101110010110;
assign LUT_4[37105] = 32'b11111111111111111100111010001110;
assign LUT_4[37106] = 32'b00000000000000000011001000111010;
assign LUT_4[37107] = 32'b11111111111111111100010100110010;
assign LUT_4[37108] = 32'b00000000000000000000101110110010;
assign LUT_4[37109] = 32'b11111111111111111001111010101010;
assign LUT_4[37110] = 32'b00000000000000000000001001010110;
assign LUT_4[37111] = 32'b11111111111111111001010101001110;
assign LUT_4[37112] = 32'b11111111111111111100111010101011;
assign LUT_4[37113] = 32'b11111111111111110110000110100011;
assign LUT_4[37114] = 32'b11111111111111111100010101001111;
assign LUT_4[37115] = 32'b11111111111111110101100001000111;
assign LUT_4[37116] = 32'b11111111111111111001111011000111;
assign LUT_4[37117] = 32'b11111111111111110011000110111111;
assign LUT_4[37118] = 32'b11111111111111111001010101101011;
assign LUT_4[37119] = 32'b11111111111111110010100001100011;
assign LUT_4[37120] = 32'b00000000000000001000011111101000;
assign LUT_4[37121] = 32'b00000000000000000001101011100000;
assign LUT_4[37122] = 32'b00000000000000000111111010001100;
assign LUT_4[37123] = 32'b00000000000000000001000110000100;
assign LUT_4[37124] = 32'b00000000000000000101100000000100;
assign LUT_4[37125] = 32'b11111111111111111110101011111100;
assign LUT_4[37126] = 32'b00000000000000000100111010101000;
assign LUT_4[37127] = 32'b11111111111111111110000110100000;
assign LUT_4[37128] = 32'b00000000000000000001101011111101;
assign LUT_4[37129] = 32'b11111111111111111010110111110101;
assign LUT_4[37130] = 32'b00000000000000000001000110100001;
assign LUT_4[37131] = 32'b11111111111111111010010010011001;
assign LUT_4[37132] = 32'b11111111111111111110101100011001;
assign LUT_4[37133] = 32'b11111111111111110111111000010001;
assign LUT_4[37134] = 32'b11111111111111111110000110111101;
assign LUT_4[37135] = 32'b11111111111111110111010010110101;
assign LUT_4[37136] = 32'b00000000000000000110010001010110;
assign LUT_4[37137] = 32'b11111111111111111111011101001110;
assign LUT_4[37138] = 32'b00000000000000000101101011111010;
assign LUT_4[37139] = 32'b11111111111111111110110111110010;
assign LUT_4[37140] = 32'b00000000000000000011010001110010;
assign LUT_4[37141] = 32'b11111111111111111100011101101010;
assign LUT_4[37142] = 32'b00000000000000000010101100010110;
assign LUT_4[37143] = 32'b11111111111111111011111000001110;
assign LUT_4[37144] = 32'b11111111111111111111011101101011;
assign LUT_4[37145] = 32'b11111111111111111000101001100011;
assign LUT_4[37146] = 32'b11111111111111111110111000001111;
assign LUT_4[37147] = 32'b11111111111111111000000100000111;
assign LUT_4[37148] = 32'b11111111111111111100011110000111;
assign LUT_4[37149] = 32'b11111111111111110101101001111111;
assign LUT_4[37150] = 32'b11111111111111111011111000101011;
assign LUT_4[37151] = 32'b11111111111111110101000100100011;
assign LUT_4[37152] = 32'b00000000000000000110111010101111;
assign LUT_4[37153] = 32'b00000000000000000000000110100111;
assign LUT_4[37154] = 32'b00000000000000000110010101010011;
assign LUT_4[37155] = 32'b11111111111111111111100001001011;
assign LUT_4[37156] = 32'b00000000000000000011111011001011;
assign LUT_4[37157] = 32'b11111111111111111101000111000011;
assign LUT_4[37158] = 32'b00000000000000000011010101101111;
assign LUT_4[37159] = 32'b11111111111111111100100001100111;
assign LUT_4[37160] = 32'b00000000000000000000000111000100;
assign LUT_4[37161] = 32'b11111111111111111001010010111100;
assign LUT_4[37162] = 32'b11111111111111111111100001101000;
assign LUT_4[37163] = 32'b11111111111111111000101101100000;
assign LUT_4[37164] = 32'b11111111111111111101000111100000;
assign LUT_4[37165] = 32'b11111111111111110110010011011000;
assign LUT_4[37166] = 32'b11111111111111111100100010000100;
assign LUT_4[37167] = 32'b11111111111111110101101101111100;
assign LUT_4[37168] = 32'b00000000000000000100101100011101;
assign LUT_4[37169] = 32'b11111111111111111101111000010101;
assign LUT_4[37170] = 32'b00000000000000000100000111000001;
assign LUT_4[37171] = 32'b11111111111111111101010010111001;
assign LUT_4[37172] = 32'b00000000000000000001101100111001;
assign LUT_4[37173] = 32'b11111111111111111010111000110001;
assign LUT_4[37174] = 32'b00000000000000000001000111011101;
assign LUT_4[37175] = 32'b11111111111111111010010011010101;
assign LUT_4[37176] = 32'b11111111111111111101111000110010;
assign LUT_4[37177] = 32'b11111111111111110111000100101010;
assign LUT_4[37178] = 32'b11111111111111111101010011010110;
assign LUT_4[37179] = 32'b11111111111111110110011111001110;
assign LUT_4[37180] = 32'b11111111111111111010111001001110;
assign LUT_4[37181] = 32'b11111111111111110100000101000110;
assign LUT_4[37182] = 32'b11111111111111111010010011110010;
assign LUT_4[37183] = 32'b11111111111111110011011111101010;
assign LUT_4[37184] = 32'b00000000000000001001110110111100;
assign LUT_4[37185] = 32'b00000000000000000011000010110100;
assign LUT_4[37186] = 32'b00000000000000001001010001100000;
assign LUT_4[37187] = 32'b00000000000000000010011101011000;
assign LUT_4[37188] = 32'b00000000000000000110110111011000;
assign LUT_4[37189] = 32'b00000000000000000000000011010000;
assign LUT_4[37190] = 32'b00000000000000000110010001111100;
assign LUT_4[37191] = 32'b11111111111111111111011101110100;
assign LUT_4[37192] = 32'b00000000000000000011000011010001;
assign LUT_4[37193] = 32'b11111111111111111100001111001001;
assign LUT_4[37194] = 32'b00000000000000000010011101110101;
assign LUT_4[37195] = 32'b11111111111111111011101001101101;
assign LUT_4[37196] = 32'b00000000000000000000000011101101;
assign LUT_4[37197] = 32'b11111111111111111001001111100101;
assign LUT_4[37198] = 32'b11111111111111111111011110010001;
assign LUT_4[37199] = 32'b11111111111111111000101010001001;
assign LUT_4[37200] = 32'b00000000000000000111101000101010;
assign LUT_4[37201] = 32'b00000000000000000000110100100010;
assign LUT_4[37202] = 32'b00000000000000000111000011001110;
assign LUT_4[37203] = 32'b00000000000000000000001111000110;
assign LUT_4[37204] = 32'b00000000000000000100101001000110;
assign LUT_4[37205] = 32'b11111111111111111101110100111110;
assign LUT_4[37206] = 32'b00000000000000000100000011101010;
assign LUT_4[37207] = 32'b11111111111111111101001111100010;
assign LUT_4[37208] = 32'b00000000000000000000110100111111;
assign LUT_4[37209] = 32'b11111111111111111010000000110111;
assign LUT_4[37210] = 32'b00000000000000000000001111100011;
assign LUT_4[37211] = 32'b11111111111111111001011011011011;
assign LUT_4[37212] = 32'b11111111111111111101110101011011;
assign LUT_4[37213] = 32'b11111111111111110111000001010011;
assign LUT_4[37214] = 32'b11111111111111111101001111111111;
assign LUT_4[37215] = 32'b11111111111111110110011011110111;
assign LUT_4[37216] = 32'b00000000000000001000010010000011;
assign LUT_4[37217] = 32'b00000000000000000001011101111011;
assign LUT_4[37218] = 32'b00000000000000000111101100100111;
assign LUT_4[37219] = 32'b00000000000000000000111000011111;
assign LUT_4[37220] = 32'b00000000000000000101010010011111;
assign LUT_4[37221] = 32'b11111111111111111110011110010111;
assign LUT_4[37222] = 32'b00000000000000000100101101000011;
assign LUT_4[37223] = 32'b11111111111111111101111000111011;
assign LUT_4[37224] = 32'b00000000000000000001011110011000;
assign LUT_4[37225] = 32'b11111111111111111010101010010000;
assign LUT_4[37226] = 32'b00000000000000000000111000111100;
assign LUT_4[37227] = 32'b11111111111111111010000100110100;
assign LUT_4[37228] = 32'b11111111111111111110011110110100;
assign LUT_4[37229] = 32'b11111111111111110111101010101100;
assign LUT_4[37230] = 32'b11111111111111111101111001011000;
assign LUT_4[37231] = 32'b11111111111111110111000101010000;
assign LUT_4[37232] = 32'b00000000000000000110000011110001;
assign LUT_4[37233] = 32'b11111111111111111111001111101001;
assign LUT_4[37234] = 32'b00000000000000000101011110010101;
assign LUT_4[37235] = 32'b11111111111111111110101010001101;
assign LUT_4[37236] = 32'b00000000000000000011000100001101;
assign LUT_4[37237] = 32'b11111111111111111100010000000101;
assign LUT_4[37238] = 32'b00000000000000000010011110110001;
assign LUT_4[37239] = 32'b11111111111111111011101010101001;
assign LUT_4[37240] = 32'b11111111111111111111010000000110;
assign LUT_4[37241] = 32'b11111111111111111000011011111110;
assign LUT_4[37242] = 32'b11111111111111111110101010101010;
assign LUT_4[37243] = 32'b11111111111111110111110110100010;
assign LUT_4[37244] = 32'b11111111111111111100010000100010;
assign LUT_4[37245] = 32'b11111111111111110101011100011010;
assign LUT_4[37246] = 32'b11111111111111111011101011000110;
assign LUT_4[37247] = 32'b11111111111111110100110110111110;
assign LUT_4[37248] = 32'b00000000000000001011000101110000;
assign LUT_4[37249] = 32'b00000000000000000100010001101000;
assign LUT_4[37250] = 32'b00000000000000001010100000010100;
assign LUT_4[37251] = 32'b00000000000000000011101100001100;
assign LUT_4[37252] = 32'b00000000000000001000000110001100;
assign LUT_4[37253] = 32'b00000000000000000001010010000100;
assign LUT_4[37254] = 32'b00000000000000000111100000110000;
assign LUT_4[37255] = 32'b00000000000000000000101100101000;
assign LUT_4[37256] = 32'b00000000000000000100010010000101;
assign LUT_4[37257] = 32'b11111111111111111101011101111101;
assign LUT_4[37258] = 32'b00000000000000000011101100101001;
assign LUT_4[37259] = 32'b11111111111111111100111000100001;
assign LUT_4[37260] = 32'b00000000000000000001010010100001;
assign LUT_4[37261] = 32'b11111111111111111010011110011001;
assign LUT_4[37262] = 32'b00000000000000000000101101000101;
assign LUT_4[37263] = 32'b11111111111111111001111000111101;
assign LUT_4[37264] = 32'b00000000000000001000110111011110;
assign LUT_4[37265] = 32'b00000000000000000010000011010110;
assign LUT_4[37266] = 32'b00000000000000001000010010000010;
assign LUT_4[37267] = 32'b00000000000000000001011101111010;
assign LUT_4[37268] = 32'b00000000000000000101110111111010;
assign LUT_4[37269] = 32'b11111111111111111111000011110010;
assign LUT_4[37270] = 32'b00000000000000000101010010011110;
assign LUT_4[37271] = 32'b11111111111111111110011110010110;
assign LUT_4[37272] = 32'b00000000000000000010000011110011;
assign LUT_4[37273] = 32'b11111111111111111011001111101011;
assign LUT_4[37274] = 32'b00000000000000000001011110010111;
assign LUT_4[37275] = 32'b11111111111111111010101010001111;
assign LUT_4[37276] = 32'b11111111111111111111000100001111;
assign LUT_4[37277] = 32'b11111111111111111000010000000111;
assign LUT_4[37278] = 32'b11111111111111111110011110110011;
assign LUT_4[37279] = 32'b11111111111111110111101010101011;
assign LUT_4[37280] = 32'b00000000000000001001100000110111;
assign LUT_4[37281] = 32'b00000000000000000010101100101111;
assign LUT_4[37282] = 32'b00000000000000001000111011011011;
assign LUT_4[37283] = 32'b00000000000000000010000111010011;
assign LUT_4[37284] = 32'b00000000000000000110100001010011;
assign LUT_4[37285] = 32'b11111111111111111111101101001011;
assign LUT_4[37286] = 32'b00000000000000000101111011110111;
assign LUT_4[37287] = 32'b11111111111111111111000111101111;
assign LUT_4[37288] = 32'b00000000000000000010101101001100;
assign LUT_4[37289] = 32'b11111111111111111011111001000100;
assign LUT_4[37290] = 32'b00000000000000000010000111110000;
assign LUT_4[37291] = 32'b11111111111111111011010011101000;
assign LUT_4[37292] = 32'b11111111111111111111101101101000;
assign LUT_4[37293] = 32'b11111111111111111000111001100000;
assign LUT_4[37294] = 32'b11111111111111111111001000001100;
assign LUT_4[37295] = 32'b11111111111111111000010100000100;
assign LUT_4[37296] = 32'b00000000000000000111010010100101;
assign LUT_4[37297] = 32'b00000000000000000000011110011101;
assign LUT_4[37298] = 32'b00000000000000000110101101001001;
assign LUT_4[37299] = 32'b11111111111111111111111001000001;
assign LUT_4[37300] = 32'b00000000000000000100010011000001;
assign LUT_4[37301] = 32'b11111111111111111101011110111001;
assign LUT_4[37302] = 32'b00000000000000000011101101100101;
assign LUT_4[37303] = 32'b11111111111111111100111001011101;
assign LUT_4[37304] = 32'b00000000000000000000011110111010;
assign LUT_4[37305] = 32'b11111111111111111001101010110010;
assign LUT_4[37306] = 32'b11111111111111111111111001011110;
assign LUT_4[37307] = 32'b11111111111111111001000101010110;
assign LUT_4[37308] = 32'b11111111111111111101011111010110;
assign LUT_4[37309] = 32'b11111111111111110110101011001110;
assign LUT_4[37310] = 32'b11111111111111111100111001111010;
assign LUT_4[37311] = 32'b11111111111111110110000101110010;
assign LUT_4[37312] = 32'b00000000000000001100011101000100;
assign LUT_4[37313] = 32'b00000000000000000101101000111100;
assign LUT_4[37314] = 32'b00000000000000001011110111101000;
assign LUT_4[37315] = 32'b00000000000000000101000011100000;
assign LUT_4[37316] = 32'b00000000000000001001011101100000;
assign LUT_4[37317] = 32'b00000000000000000010101001011000;
assign LUT_4[37318] = 32'b00000000000000001000111000000100;
assign LUT_4[37319] = 32'b00000000000000000010000011111100;
assign LUT_4[37320] = 32'b00000000000000000101101001011001;
assign LUT_4[37321] = 32'b11111111111111111110110101010001;
assign LUT_4[37322] = 32'b00000000000000000101000011111101;
assign LUT_4[37323] = 32'b11111111111111111110001111110101;
assign LUT_4[37324] = 32'b00000000000000000010101001110101;
assign LUT_4[37325] = 32'b11111111111111111011110101101101;
assign LUT_4[37326] = 32'b00000000000000000010000100011001;
assign LUT_4[37327] = 32'b11111111111111111011010000010001;
assign LUT_4[37328] = 32'b00000000000000001010001110110010;
assign LUT_4[37329] = 32'b00000000000000000011011010101010;
assign LUT_4[37330] = 32'b00000000000000001001101001010110;
assign LUT_4[37331] = 32'b00000000000000000010110101001110;
assign LUT_4[37332] = 32'b00000000000000000111001111001110;
assign LUT_4[37333] = 32'b00000000000000000000011011000110;
assign LUT_4[37334] = 32'b00000000000000000110101001110010;
assign LUT_4[37335] = 32'b11111111111111111111110101101010;
assign LUT_4[37336] = 32'b00000000000000000011011011000111;
assign LUT_4[37337] = 32'b11111111111111111100100110111111;
assign LUT_4[37338] = 32'b00000000000000000010110101101011;
assign LUT_4[37339] = 32'b11111111111111111100000001100011;
assign LUT_4[37340] = 32'b00000000000000000000011011100011;
assign LUT_4[37341] = 32'b11111111111111111001100111011011;
assign LUT_4[37342] = 32'b11111111111111111111110110000111;
assign LUT_4[37343] = 32'b11111111111111111001000001111111;
assign LUT_4[37344] = 32'b00000000000000001010111000001011;
assign LUT_4[37345] = 32'b00000000000000000100000100000011;
assign LUT_4[37346] = 32'b00000000000000001010010010101111;
assign LUT_4[37347] = 32'b00000000000000000011011110100111;
assign LUT_4[37348] = 32'b00000000000000000111111000100111;
assign LUT_4[37349] = 32'b00000000000000000001000100011111;
assign LUT_4[37350] = 32'b00000000000000000111010011001011;
assign LUT_4[37351] = 32'b00000000000000000000011111000011;
assign LUT_4[37352] = 32'b00000000000000000100000100100000;
assign LUT_4[37353] = 32'b11111111111111111101010000011000;
assign LUT_4[37354] = 32'b00000000000000000011011111000100;
assign LUT_4[37355] = 32'b11111111111111111100101010111100;
assign LUT_4[37356] = 32'b00000000000000000001000100111100;
assign LUT_4[37357] = 32'b11111111111111111010010000110100;
assign LUT_4[37358] = 32'b00000000000000000000011111100000;
assign LUT_4[37359] = 32'b11111111111111111001101011011000;
assign LUT_4[37360] = 32'b00000000000000001000101001111001;
assign LUT_4[37361] = 32'b00000000000000000001110101110001;
assign LUT_4[37362] = 32'b00000000000000001000000100011101;
assign LUT_4[37363] = 32'b00000000000000000001010000010101;
assign LUT_4[37364] = 32'b00000000000000000101101010010101;
assign LUT_4[37365] = 32'b11111111111111111110110110001101;
assign LUT_4[37366] = 32'b00000000000000000101000100111001;
assign LUT_4[37367] = 32'b11111111111111111110010000110001;
assign LUT_4[37368] = 32'b00000000000000000001110110001110;
assign LUT_4[37369] = 32'b11111111111111111011000010000110;
assign LUT_4[37370] = 32'b00000000000000000001010000110010;
assign LUT_4[37371] = 32'b11111111111111111010011100101010;
assign LUT_4[37372] = 32'b11111111111111111110110110101010;
assign LUT_4[37373] = 32'b11111111111111111000000010100010;
assign LUT_4[37374] = 32'b11111111111111111110010001001110;
assign LUT_4[37375] = 32'b11111111111111110111011101000110;
assign LUT_4[37376] = 32'b00000000000000000010101000001101;
assign LUT_4[37377] = 32'b11111111111111111011110100000101;
assign LUT_4[37378] = 32'b00000000000000000010000010110001;
assign LUT_4[37379] = 32'b11111111111111111011001110101001;
assign LUT_4[37380] = 32'b11111111111111111111101000101001;
assign LUT_4[37381] = 32'b11111111111111111000110100100001;
assign LUT_4[37382] = 32'b11111111111111111111000011001101;
assign LUT_4[37383] = 32'b11111111111111111000001111000101;
assign LUT_4[37384] = 32'b11111111111111111011110100100010;
assign LUT_4[37385] = 32'b11111111111111110101000000011010;
assign LUT_4[37386] = 32'b11111111111111111011001111000110;
assign LUT_4[37387] = 32'b11111111111111110100011010111110;
assign LUT_4[37388] = 32'b11111111111111111000110100111110;
assign LUT_4[37389] = 32'b11111111111111110010000000110110;
assign LUT_4[37390] = 32'b11111111111111111000001111100010;
assign LUT_4[37391] = 32'b11111111111111110001011011011010;
assign LUT_4[37392] = 32'b00000000000000000000011001111011;
assign LUT_4[37393] = 32'b11111111111111111001100101110011;
assign LUT_4[37394] = 32'b11111111111111111111110100011111;
assign LUT_4[37395] = 32'b11111111111111111001000000010111;
assign LUT_4[37396] = 32'b11111111111111111101011010010111;
assign LUT_4[37397] = 32'b11111111111111110110100110001111;
assign LUT_4[37398] = 32'b11111111111111111100110100111011;
assign LUT_4[37399] = 32'b11111111111111110110000000110011;
assign LUT_4[37400] = 32'b11111111111111111001100110010000;
assign LUT_4[37401] = 32'b11111111111111110010110010001000;
assign LUT_4[37402] = 32'b11111111111111111001000000110100;
assign LUT_4[37403] = 32'b11111111111111110010001100101100;
assign LUT_4[37404] = 32'b11111111111111110110100110101100;
assign LUT_4[37405] = 32'b11111111111111101111110010100100;
assign LUT_4[37406] = 32'b11111111111111110110000001010000;
assign LUT_4[37407] = 32'b11111111111111101111001101001000;
assign LUT_4[37408] = 32'b00000000000000000001000011010100;
assign LUT_4[37409] = 32'b11111111111111111010001111001100;
assign LUT_4[37410] = 32'b00000000000000000000011101111000;
assign LUT_4[37411] = 32'b11111111111111111001101001110000;
assign LUT_4[37412] = 32'b11111111111111111110000011110000;
assign LUT_4[37413] = 32'b11111111111111110111001111101000;
assign LUT_4[37414] = 32'b11111111111111111101011110010100;
assign LUT_4[37415] = 32'b11111111111111110110101010001100;
assign LUT_4[37416] = 32'b11111111111111111010001111101001;
assign LUT_4[37417] = 32'b11111111111111110011011011100001;
assign LUT_4[37418] = 32'b11111111111111111001101010001101;
assign LUT_4[37419] = 32'b11111111111111110010110110000101;
assign LUT_4[37420] = 32'b11111111111111110111010000000101;
assign LUT_4[37421] = 32'b11111111111111110000011011111101;
assign LUT_4[37422] = 32'b11111111111111110110101010101001;
assign LUT_4[37423] = 32'b11111111111111101111110110100001;
assign LUT_4[37424] = 32'b11111111111111111110110101000010;
assign LUT_4[37425] = 32'b11111111111111111000000000111010;
assign LUT_4[37426] = 32'b11111111111111111110001111100110;
assign LUT_4[37427] = 32'b11111111111111110111011011011110;
assign LUT_4[37428] = 32'b11111111111111111011110101011110;
assign LUT_4[37429] = 32'b11111111111111110101000001010110;
assign LUT_4[37430] = 32'b11111111111111111011010000000010;
assign LUT_4[37431] = 32'b11111111111111110100011011111010;
assign LUT_4[37432] = 32'b11111111111111111000000001010111;
assign LUT_4[37433] = 32'b11111111111111110001001101001111;
assign LUT_4[37434] = 32'b11111111111111110111011011111011;
assign LUT_4[37435] = 32'b11111111111111110000100111110011;
assign LUT_4[37436] = 32'b11111111111111110101000001110011;
assign LUT_4[37437] = 32'b11111111111111101110001101101011;
assign LUT_4[37438] = 32'b11111111111111110100011100010111;
assign LUT_4[37439] = 32'b11111111111111101101101000001111;
assign LUT_4[37440] = 32'b00000000000000000011111111100001;
assign LUT_4[37441] = 32'b11111111111111111101001011011001;
assign LUT_4[37442] = 32'b00000000000000000011011010000101;
assign LUT_4[37443] = 32'b11111111111111111100100101111101;
assign LUT_4[37444] = 32'b00000000000000000000111111111101;
assign LUT_4[37445] = 32'b11111111111111111010001011110101;
assign LUT_4[37446] = 32'b00000000000000000000011010100001;
assign LUT_4[37447] = 32'b11111111111111111001100110011001;
assign LUT_4[37448] = 32'b11111111111111111101001011110110;
assign LUT_4[37449] = 32'b11111111111111110110010111101110;
assign LUT_4[37450] = 32'b11111111111111111100100110011010;
assign LUT_4[37451] = 32'b11111111111111110101110010010010;
assign LUT_4[37452] = 32'b11111111111111111010001100010010;
assign LUT_4[37453] = 32'b11111111111111110011011000001010;
assign LUT_4[37454] = 32'b11111111111111111001100110110110;
assign LUT_4[37455] = 32'b11111111111111110010110010101110;
assign LUT_4[37456] = 32'b00000000000000000001110001001111;
assign LUT_4[37457] = 32'b11111111111111111010111101000111;
assign LUT_4[37458] = 32'b00000000000000000001001011110011;
assign LUT_4[37459] = 32'b11111111111111111010010111101011;
assign LUT_4[37460] = 32'b11111111111111111110110001101011;
assign LUT_4[37461] = 32'b11111111111111110111111101100011;
assign LUT_4[37462] = 32'b11111111111111111110001100001111;
assign LUT_4[37463] = 32'b11111111111111110111011000000111;
assign LUT_4[37464] = 32'b11111111111111111010111101100100;
assign LUT_4[37465] = 32'b11111111111111110100001001011100;
assign LUT_4[37466] = 32'b11111111111111111010011000001000;
assign LUT_4[37467] = 32'b11111111111111110011100100000000;
assign LUT_4[37468] = 32'b11111111111111110111111110000000;
assign LUT_4[37469] = 32'b11111111111111110001001001111000;
assign LUT_4[37470] = 32'b11111111111111110111011000100100;
assign LUT_4[37471] = 32'b11111111111111110000100100011100;
assign LUT_4[37472] = 32'b00000000000000000010011010101000;
assign LUT_4[37473] = 32'b11111111111111111011100110100000;
assign LUT_4[37474] = 32'b00000000000000000001110101001100;
assign LUT_4[37475] = 32'b11111111111111111011000001000100;
assign LUT_4[37476] = 32'b11111111111111111111011011000100;
assign LUT_4[37477] = 32'b11111111111111111000100110111100;
assign LUT_4[37478] = 32'b11111111111111111110110101101000;
assign LUT_4[37479] = 32'b11111111111111111000000001100000;
assign LUT_4[37480] = 32'b11111111111111111011100110111101;
assign LUT_4[37481] = 32'b11111111111111110100110010110101;
assign LUT_4[37482] = 32'b11111111111111111011000001100001;
assign LUT_4[37483] = 32'b11111111111111110100001101011001;
assign LUT_4[37484] = 32'b11111111111111111000100111011001;
assign LUT_4[37485] = 32'b11111111111111110001110011010001;
assign LUT_4[37486] = 32'b11111111111111111000000001111101;
assign LUT_4[37487] = 32'b11111111111111110001001101110101;
assign LUT_4[37488] = 32'b00000000000000000000001100010110;
assign LUT_4[37489] = 32'b11111111111111111001011000001110;
assign LUT_4[37490] = 32'b11111111111111111111100110111010;
assign LUT_4[37491] = 32'b11111111111111111000110010110010;
assign LUT_4[37492] = 32'b11111111111111111101001100110010;
assign LUT_4[37493] = 32'b11111111111111110110011000101010;
assign LUT_4[37494] = 32'b11111111111111111100100111010110;
assign LUT_4[37495] = 32'b11111111111111110101110011001110;
assign LUT_4[37496] = 32'b11111111111111111001011000101011;
assign LUT_4[37497] = 32'b11111111111111110010100100100011;
assign LUT_4[37498] = 32'b11111111111111111000110011001111;
assign LUT_4[37499] = 32'b11111111111111110001111111000111;
assign LUT_4[37500] = 32'b11111111111111110110011001000111;
assign LUT_4[37501] = 32'b11111111111111101111100100111111;
assign LUT_4[37502] = 32'b11111111111111110101110011101011;
assign LUT_4[37503] = 32'b11111111111111101110111111100011;
assign LUT_4[37504] = 32'b00000000000000000101001110010101;
assign LUT_4[37505] = 32'b11111111111111111110011010001101;
assign LUT_4[37506] = 32'b00000000000000000100101000111001;
assign LUT_4[37507] = 32'b11111111111111111101110100110001;
assign LUT_4[37508] = 32'b00000000000000000010001110110001;
assign LUT_4[37509] = 32'b11111111111111111011011010101001;
assign LUT_4[37510] = 32'b00000000000000000001101001010101;
assign LUT_4[37511] = 32'b11111111111111111010110101001101;
assign LUT_4[37512] = 32'b11111111111111111110011010101010;
assign LUT_4[37513] = 32'b11111111111111110111100110100010;
assign LUT_4[37514] = 32'b11111111111111111101110101001110;
assign LUT_4[37515] = 32'b11111111111111110111000001000110;
assign LUT_4[37516] = 32'b11111111111111111011011011000110;
assign LUT_4[37517] = 32'b11111111111111110100100110111110;
assign LUT_4[37518] = 32'b11111111111111111010110101101010;
assign LUT_4[37519] = 32'b11111111111111110100000001100010;
assign LUT_4[37520] = 32'b00000000000000000011000000000011;
assign LUT_4[37521] = 32'b11111111111111111100001011111011;
assign LUT_4[37522] = 32'b00000000000000000010011010100111;
assign LUT_4[37523] = 32'b11111111111111111011100110011111;
assign LUT_4[37524] = 32'b00000000000000000000000000011111;
assign LUT_4[37525] = 32'b11111111111111111001001100010111;
assign LUT_4[37526] = 32'b11111111111111111111011011000011;
assign LUT_4[37527] = 32'b11111111111111111000100110111011;
assign LUT_4[37528] = 32'b11111111111111111100001100011000;
assign LUT_4[37529] = 32'b11111111111111110101011000010000;
assign LUT_4[37530] = 32'b11111111111111111011100110111100;
assign LUT_4[37531] = 32'b11111111111111110100110010110100;
assign LUT_4[37532] = 32'b11111111111111111001001100110100;
assign LUT_4[37533] = 32'b11111111111111110010011000101100;
assign LUT_4[37534] = 32'b11111111111111111000100111011000;
assign LUT_4[37535] = 32'b11111111111111110001110011010000;
assign LUT_4[37536] = 32'b00000000000000000011101001011100;
assign LUT_4[37537] = 32'b11111111111111111100110101010100;
assign LUT_4[37538] = 32'b00000000000000000011000100000000;
assign LUT_4[37539] = 32'b11111111111111111100001111111000;
assign LUT_4[37540] = 32'b00000000000000000000101001111000;
assign LUT_4[37541] = 32'b11111111111111111001110101110000;
assign LUT_4[37542] = 32'b00000000000000000000000100011100;
assign LUT_4[37543] = 32'b11111111111111111001010000010100;
assign LUT_4[37544] = 32'b11111111111111111100110101110001;
assign LUT_4[37545] = 32'b11111111111111110110000001101001;
assign LUT_4[37546] = 32'b11111111111111111100010000010101;
assign LUT_4[37547] = 32'b11111111111111110101011100001101;
assign LUT_4[37548] = 32'b11111111111111111001110110001101;
assign LUT_4[37549] = 32'b11111111111111110011000010000101;
assign LUT_4[37550] = 32'b11111111111111111001010000110001;
assign LUT_4[37551] = 32'b11111111111111110010011100101001;
assign LUT_4[37552] = 32'b00000000000000000001011011001010;
assign LUT_4[37553] = 32'b11111111111111111010100111000010;
assign LUT_4[37554] = 32'b00000000000000000000110101101110;
assign LUT_4[37555] = 32'b11111111111111111010000001100110;
assign LUT_4[37556] = 32'b11111111111111111110011011100110;
assign LUT_4[37557] = 32'b11111111111111110111100111011110;
assign LUT_4[37558] = 32'b11111111111111111101110110001010;
assign LUT_4[37559] = 32'b11111111111111110111000010000010;
assign LUT_4[37560] = 32'b11111111111111111010100111011111;
assign LUT_4[37561] = 32'b11111111111111110011110011010111;
assign LUT_4[37562] = 32'b11111111111111111010000010000011;
assign LUT_4[37563] = 32'b11111111111111110011001101111011;
assign LUT_4[37564] = 32'b11111111111111110111100111111011;
assign LUT_4[37565] = 32'b11111111111111110000110011110011;
assign LUT_4[37566] = 32'b11111111111111110111000010011111;
assign LUT_4[37567] = 32'b11111111111111110000001110010111;
assign LUT_4[37568] = 32'b00000000000000000110100101101001;
assign LUT_4[37569] = 32'b11111111111111111111110001100001;
assign LUT_4[37570] = 32'b00000000000000000110000000001101;
assign LUT_4[37571] = 32'b11111111111111111111001100000101;
assign LUT_4[37572] = 32'b00000000000000000011100110000101;
assign LUT_4[37573] = 32'b11111111111111111100110001111101;
assign LUT_4[37574] = 32'b00000000000000000011000000101001;
assign LUT_4[37575] = 32'b11111111111111111100001100100001;
assign LUT_4[37576] = 32'b11111111111111111111110001111110;
assign LUT_4[37577] = 32'b11111111111111111000111101110110;
assign LUT_4[37578] = 32'b11111111111111111111001100100010;
assign LUT_4[37579] = 32'b11111111111111111000011000011010;
assign LUT_4[37580] = 32'b11111111111111111100110010011010;
assign LUT_4[37581] = 32'b11111111111111110101111110010010;
assign LUT_4[37582] = 32'b11111111111111111100001100111110;
assign LUT_4[37583] = 32'b11111111111111110101011000110110;
assign LUT_4[37584] = 32'b00000000000000000100010111010111;
assign LUT_4[37585] = 32'b11111111111111111101100011001111;
assign LUT_4[37586] = 32'b00000000000000000011110001111011;
assign LUT_4[37587] = 32'b11111111111111111100111101110011;
assign LUT_4[37588] = 32'b00000000000000000001010111110011;
assign LUT_4[37589] = 32'b11111111111111111010100011101011;
assign LUT_4[37590] = 32'b00000000000000000000110010010111;
assign LUT_4[37591] = 32'b11111111111111111001111110001111;
assign LUT_4[37592] = 32'b11111111111111111101100011101100;
assign LUT_4[37593] = 32'b11111111111111110110101111100100;
assign LUT_4[37594] = 32'b11111111111111111100111110010000;
assign LUT_4[37595] = 32'b11111111111111110110001010001000;
assign LUT_4[37596] = 32'b11111111111111111010100100001000;
assign LUT_4[37597] = 32'b11111111111111110011110000000000;
assign LUT_4[37598] = 32'b11111111111111111001111110101100;
assign LUT_4[37599] = 32'b11111111111111110011001010100100;
assign LUT_4[37600] = 32'b00000000000000000101000000110000;
assign LUT_4[37601] = 32'b11111111111111111110001100101000;
assign LUT_4[37602] = 32'b00000000000000000100011011010100;
assign LUT_4[37603] = 32'b11111111111111111101100111001100;
assign LUT_4[37604] = 32'b00000000000000000010000001001100;
assign LUT_4[37605] = 32'b11111111111111111011001101000100;
assign LUT_4[37606] = 32'b00000000000000000001011011110000;
assign LUT_4[37607] = 32'b11111111111111111010100111101000;
assign LUT_4[37608] = 32'b11111111111111111110001101000101;
assign LUT_4[37609] = 32'b11111111111111110111011000111101;
assign LUT_4[37610] = 32'b11111111111111111101100111101001;
assign LUT_4[37611] = 32'b11111111111111110110110011100001;
assign LUT_4[37612] = 32'b11111111111111111011001101100001;
assign LUT_4[37613] = 32'b11111111111111110100011001011001;
assign LUT_4[37614] = 32'b11111111111111111010101000000101;
assign LUT_4[37615] = 32'b11111111111111110011110011111101;
assign LUT_4[37616] = 32'b00000000000000000010110010011110;
assign LUT_4[37617] = 32'b11111111111111111011111110010110;
assign LUT_4[37618] = 32'b00000000000000000010001101000010;
assign LUT_4[37619] = 32'b11111111111111111011011000111010;
assign LUT_4[37620] = 32'b11111111111111111111110010111010;
assign LUT_4[37621] = 32'b11111111111111111000111110110010;
assign LUT_4[37622] = 32'b11111111111111111111001101011110;
assign LUT_4[37623] = 32'b11111111111111111000011001010110;
assign LUT_4[37624] = 32'b11111111111111111011111110110011;
assign LUT_4[37625] = 32'b11111111111111110101001010101011;
assign LUT_4[37626] = 32'b11111111111111111011011001010111;
assign LUT_4[37627] = 32'b11111111111111110100100101001111;
assign LUT_4[37628] = 32'b11111111111111111000111111001111;
assign LUT_4[37629] = 32'b11111111111111110010001011000111;
assign LUT_4[37630] = 32'b11111111111111111000011001110011;
assign LUT_4[37631] = 32'b11111111111111110001100101101011;
assign LUT_4[37632] = 32'b00000000000000000111100011110000;
assign LUT_4[37633] = 32'b00000000000000000000101111101000;
assign LUT_4[37634] = 32'b00000000000000000110111110010100;
assign LUT_4[37635] = 32'b00000000000000000000001010001100;
assign LUT_4[37636] = 32'b00000000000000000100100100001100;
assign LUT_4[37637] = 32'b11111111111111111101110000000100;
assign LUT_4[37638] = 32'b00000000000000000011111110110000;
assign LUT_4[37639] = 32'b11111111111111111101001010101000;
assign LUT_4[37640] = 32'b00000000000000000000110000000101;
assign LUT_4[37641] = 32'b11111111111111111001111011111101;
assign LUT_4[37642] = 32'b00000000000000000000001010101001;
assign LUT_4[37643] = 32'b11111111111111111001010110100001;
assign LUT_4[37644] = 32'b11111111111111111101110000100001;
assign LUT_4[37645] = 32'b11111111111111110110111100011001;
assign LUT_4[37646] = 32'b11111111111111111101001011000101;
assign LUT_4[37647] = 32'b11111111111111110110010110111101;
assign LUT_4[37648] = 32'b00000000000000000101010101011110;
assign LUT_4[37649] = 32'b11111111111111111110100001010110;
assign LUT_4[37650] = 32'b00000000000000000100110000000010;
assign LUT_4[37651] = 32'b11111111111111111101111011111010;
assign LUT_4[37652] = 32'b00000000000000000010010101111010;
assign LUT_4[37653] = 32'b11111111111111111011100001110010;
assign LUT_4[37654] = 32'b00000000000000000001110000011110;
assign LUT_4[37655] = 32'b11111111111111111010111100010110;
assign LUT_4[37656] = 32'b11111111111111111110100001110011;
assign LUT_4[37657] = 32'b11111111111111110111101101101011;
assign LUT_4[37658] = 32'b11111111111111111101111100010111;
assign LUT_4[37659] = 32'b11111111111111110111001000001111;
assign LUT_4[37660] = 32'b11111111111111111011100010001111;
assign LUT_4[37661] = 32'b11111111111111110100101110000111;
assign LUT_4[37662] = 32'b11111111111111111010111100110011;
assign LUT_4[37663] = 32'b11111111111111110100001000101011;
assign LUT_4[37664] = 32'b00000000000000000101111110110111;
assign LUT_4[37665] = 32'b11111111111111111111001010101111;
assign LUT_4[37666] = 32'b00000000000000000101011001011011;
assign LUT_4[37667] = 32'b11111111111111111110100101010011;
assign LUT_4[37668] = 32'b00000000000000000010111111010011;
assign LUT_4[37669] = 32'b11111111111111111100001011001011;
assign LUT_4[37670] = 32'b00000000000000000010011001110111;
assign LUT_4[37671] = 32'b11111111111111111011100101101111;
assign LUT_4[37672] = 32'b11111111111111111111001011001100;
assign LUT_4[37673] = 32'b11111111111111111000010111000100;
assign LUT_4[37674] = 32'b11111111111111111110100101110000;
assign LUT_4[37675] = 32'b11111111111111110111110001101000;
assign LUT_4[37676] = 32'b11111111111111111100001011101000;
assign LUT_4[37677] = 32'b11111111111111110101010111100000;
assign LUT_4[37678] = 32'b11111111111111111011100110001100;
assign LUT_4[37679] = 32'b11111111111111110100110010000100;
assign LUT_4[37680] = 32'b00000000000000000011110000100101;
assign LUT_4[37681] = 32'b11111111111111111100111100011101;
assign LUT_4[37682] = 32'b00000000000000000011001011001001;
assign LUT_4[37683] = 32'b11111111111111111100010111000001;
assign LUT_4[37684] = 32'b00000000000000000000110001000001;
assign LUT_4[37685] = 32'b11111111111111111001111100111001;
assign LUT_4[37686] = 32'b00000000000000000000001011100101;
assign LUT_4[37687] = 32'b11111111111111111001010111011101;
assign LUT_4[37688] = 32'b11111111111111111100111100111010;
assign LUT_4[37689] = 32'b11111111111111110110001000110010;
assign LUT_4[37690] = 32'b11111111111111111100010111011110;
assign LUT_4[37691] = 32'b11111111111111110101100011010110;
assign LUT_4[37692] = 32'b11111111111111111001111101010110;
assign LUT_4[37693] = 32'b11111111111111110011001001001110;
assign LUT_4[37694] = 32'b11111111111111111001010111111010;
assign LUT_4[37695] = 32'b11111111111111110010100011110010;
assign LUT_4[37696] = 32'b00000000000000001000111011000100;
assign LUT_4[37697] = 32'b00000000000000000010000110111100;
assign LUT_4[37698] = 32'b00000000000000001000010101101000;
assign LUT_4[37699] = 32'b00000000000000000001100001100000;
assign LUT_4[37700] = 32'b00000000000000000101111011100000;
assign LUT_4[37701] = 32'b11111111111111111111000111011000;
assign LUT_4[37702] = 32'b00000000000000000101010110000100;
assign LUT_4[37703] = 32'b11111111111111111110100001111100;
assign LUT_4[37704] = 32'b00000000000000000010000111011001;
assign LUT_4[37705] = 32'b11111111111111111011010011010001;
assign LUT_4[37706] = 32'b00000000000000000001100001111101;
assign LUT_4[37707] = 32'b11111111111111111010101101110101;
assign LUT_4[37708] = 32'b11111111111111111111000111110101;
assign LUT_4[37709] = 32'b11111111111111111000010011101101;
assign LUT_4[37710] = 32'b11111111111111111110100010011001;
assign LUT_4[37711] = 32'b11111111111111110111101110010001;
assign LUT_4[37712] = 32'b00000000000000000110101100110010;
assign LUT_4[37713] = 32'b11111111111111111111111000101010;
assign LUT_4[37714] = 32'b00000000000000000110000111010110;
assign LUT_4[37715] = 32'b11111111111111111111010011001110;
assign LUT_4[37716] = 32'b00000000000000000011101101001110;
assign LUT_4[37717] = 32'b11111111111111111100111001000110;
assign LUT_4[37718] = 32'b00000000000000000011000111110010;
assign LUT_4[37719] = 32'b11111111111111111100010011101010;
assign LUT_4[37720] = 32'b11111111111111111111111001000111;
assign LUT_4[37721] = 32'b11111111111111111001000100111111;
assign LUT_4[37722] = 32'b11111111111111111111010011101011;
assign LUT_4[37723] = 32'b11111111111111111000011111100011;
assign LUT_4[37724] = 32'b11111111111111111100111001100011;
assign LUT_4[37725] = 32'b11111111111111110110000101011011;
assign LUT_4[37726] = 32'b11111111111111111100010100000111;
assign LUT_4[37727] = 32'b11111111111111110101011111111111;
assign LUT_4[37728] = 32'b00000000000000000111010110001011;
assign LUT_4[37729] = 32'b00000000000000000000100010000011;
assign LUT_4[37730] = 32'b00000000000000000110110000101111;
assign LUT_4[37731] = 32'b11111111111111111111111100100111;
assign LUT_4[37732] = 32'b00000000000000000100010110100111;
assign LUT_4[37733] = 32'b11111111111111111101100010011111;
assign LUT_4[37734] = 32'b00000000000000000011110001001011;
assign LUT_4[37735] = 32'b11111111111111111100111101000011;
assign LUT_4[37736] = 32'b00000000000000000000100010100000;
assign LUT_4[37737] = 32'b11111111111111111001101110011000;
assign LUT_4[37738] = 32'b11111111111111111111111101000100;
assign LUT_4[37739] = 32'b11111111111111111001001000111100;
assign LUT_4[37740] = 32'b11111111111111111101100010111100;
assign LUT_4[37741] = 32'b11111111111111110110101110110100;
assign LUT_4[37742] = 32'b11111111111111111100111101100000;
assign LUT_4[37743] = 32'b11111111111111110110001001011000;
assign LUT_4[37744] = 32'b00000000000000000101000111111001;
assign LUT_4[37745] = 32'b11111111111111111110010011110001;
assign LUT_4[37746] = 32'b00000000000000000100100010011101;
assign LUT_4[37747] = 32'b11111111111111111101101110010101;
assign LUT_4[37748] = 32'b00000000000000000010001000010101;
assign LUT_4[37749] = 32'b11111111111111111011010100001101;
assign LUT_4[37750] = 32'b00000000000000000001100010111001;
assign LUT_4[37751] = 32'b11111111111111111010101110110001;
assign LUT_4[37752] = 32'b11111111111111111110010100001110;
assign LUT_4[37753] = 32'b11111111111111110111100000000110;
assign LUT_4[37754] = 32'b11111111111111111101101110110010;
assign LUT_4[37755] = 32'b11111111111111110110111010101010;
assign LUT_4[37756] = 32'b11111111111111111011010100101010;
assign LUT_4[37757] = 32'b11111111111111110100100000100010;
assign LUT_4[37758] = 32'b11111111111111111010101111001110;
assign LUT_4[37759] = 32'b11111111111111110011111011000110;
assign LUT_4[37760] = 32'b00000000000000001010001001111000;
assign LUT_4[37761] = 32'b00000000000000000011010101110000;
assign LUT_4[37762] = 32'b00000000000000001001100100011100;
assign LUT_4[37763] = 32'b00000000000000000010110000010100;
assign LUT_4[37764] = 32'b00000000000000000111001010010100;
assign LUT_4[37765] = 32'b00000000000000000000010110001100;
assign LUT_4[37766] = 32'b00000000000000000110100100111000;
assign LUT_4[37767] = 32'b11111111111111111111110000110000;
assign LUT_4[37768] = 32'b00000000000000000011010110001101;
assign LUT_4[37769] = 32'b11111111111111111100100010000101;
assign LUT_4[37770] = 32'b00000000000000000010110000110001;
assign LUT_4[37771] = 32'b11111111111111111011111100101001;
assign LUT_4[37772] = 32'b00000000000000000000010110101001;
assign LUT_4[37773] = 32'b11111111111111111001100010100001;
assign LUT_4[37774] = 32'b11111111111111111111110001001101;
assign LUT_4[37775] = 32'b11111111111111111000111101000101;
assign LUT_4[37776] = 32'b00000000000000000111111011100110;
assign LUT_4[37777] = 32'b00000000000000000001000111011110;
assign LUT_4[37778] = 32'b00000000000000000111010110001010;
assign LUT_4[37779] = 32'b00000000000000000000100010000010;
assign LUT_4[37780] = 32'b00000000000000000100111100000010;
assign LUT_4[37781] = 32'b11111111111111111110000111111010;
assign LUT_4[37782] = 32'b00000000000000000100010110100110;
assign LUT_4[37783] = 32'b11111111111111111101100010011110;
assign LUT_4[37784] = 32'b00000000000000000001000111111011;
assign LUT_4[37785] = 32'b11111111111111111010010011110011;
assign LUT_4[37786] = 32'b00000000000000000000100010011111;
assign LUT_4[37787] = 32'b11111111111111111001101110010111;
assign LUT_4[37788] = 32'b11111111111111111110001000010111;
assign LUT_4[37789] = 32'b11111111111111110111010100001111;
assign LUT_4[37790] = 32'b11111111111111111101100010111011;
assign LUT_4[37791] = 32'b11111111111111110110101110110011;
assign LUT_4[37792] = 32'b00000000000000001000100100111111;
assign LUT_4[37793] = 32'b00000000000000000001110000110111;
assign LUT_4[37794] = 32'b00000000000000000111111111100011;
assign LUT_4[37795] = 32'b00000000000000000001001011011011;
assign LUT_4[37796] = 32'b00000000000000000101100101011011;
assign LUT_4[37797] = 32'b11111111111111111110110001010011;
assign LUT_4[37798] = 32'b00000000000000000100111111111111;
assign LUT_4[37799] = 32'b11111111111111111110001011110111;
assign LUT_4[37800] = 32'b00000000000000000001110001010100;
assign LUT_4[37801] = 32'b11111111111111111010111101001100;
assign LUT_4[37802] = 32'b00000000000000000001001011111000;
assign LUT_4[37803] = 32'b11111111111111111010010111110000;
assign LUT_4[37804] = 32'b11111111111111111110110001110000;
assign LUT_4[37805] = 32'b11111111111111110111111101101000;
assign LUT_4[37806] = 32'b11111111111111111110001100010100;
assign LUT_4[37807] = 32'b11111111111111110111011000001100;
assign LUT_4[37808] = 32'b00000000000000000110010110101101;
assign LUT_4[37809] = 32'b11111111111111111111100010100101;
assign LUT_4[37810] = 32'b00000000000000000101110001010001;
assign LUT_4[37811] = 32'b11111111111111111110111101001001;
assign LUT_4[37812] = 32'b00000000000000000011010111001001;
assign LUT_4[37813] = 32'b11111111111111111100100011000001;
assign LUT_4[37814] = 32'b00000000000000000010110001101101;
assign LUT_4[37815] = 32'b11111111111111111011111101100101;
assign LUT_4[37816] = 32'b11111111111111111111100011000010;
assign LUT_4[37817] = 32'b11111111111111111000101110111010;
assign LUT_4[37818] = 32'b11111111111111111110111101100110;
assign LUT_4[37819] = 32'b11111111111111111000001001011110;
assign LUT_4[37820] = 32'b11111111111111111100100011011110;
assign LUT_4[37821] = 32'b11111111111111110101101111010110;
assign LUT_4[37822] = 32'b11111111111111111011111110000010;
assign LUT_4[37823] = 32'b11111111111111110101001001111010;
assign LUT_4[37824] = 32'b00000000000000001011100001001100;
assign LUT_4[37825] = 32'b00000000000000000100101101000100;
assign LUT_4[37826] = 32'b00000000000000001010111011110000;
assign LUT_4[37827] = 32'b00000000000000000100000111101000;
assign LUT_4[37828] = 32'b00000000000000001000100001101000;
assign LUT_4[37829] = 32'b00000000000000000001101101100000;
assign LUT_4[37830] = 32'b00000000000000000111111100001100;
assign LUT_4[37831] = 32'b00000000000000000001001000000100;
assign LUT_4[37832] = 32'b00000000000000000100101101100001;
assign LUT_4[37833] = 32'b11111111111111111101111001011001;
assign LUT_4[37834] = 32'b00000000000000000100001000000101;
assign LUT_4[37835] = 32'b11111111111111111101010011111101;
assign LUT_4[37836] = 32'b00000000000000000001101101111101;
assign LUT_4[37837] = 32'b11111111111111111010111001110101;
assign LUT_4[37838] = 32'b00000000000000000001001000100001;
assign LUT_4[37839] = 32'b11111111111111111010010100011001;
assign LUT_4[37840] = 32'b00000000000000001001010010111010;
assign LUT_4[37841] = 32'b00000000000000000010011110110010;
assign LUT_4[37842] = 32'b00000000000000001000101101011110;
assign LUT_4[37843] = 32'b00000000000000000001111001010110;
assign LUT_4[37844] = 32'b00000000000000000110010011010110;
assign LUT_4[37845] = 32'b11111111111111111111011111001110;
assign LUT_4[37846] = 32'b00000000000000000101101101111010;
assign LUT_4[37847] = 32'b11111111111111111110111001110010;
assign LUT_4[37848] = 32'b00000000000000000010011111001111;
assign LUT_4[37849] = 32'b11111111111111111011101011000111;
assign LUT_4[37850] = 32'b00000000000000000001111001110011;
assign LUT_4[37851] = 32'b11111111111111111011000101101011;
assign LUT_4[37852] = 32'b11111111111111111111011111101011;
assign LUT_4[37853] = 32'b11111111111111111000101011100011;
assign LUT_4[37854] = 32'b11111111111111111110111010001111;
assign LUT_4[37855] = 32'b11111111111111111000000110000111;
assign LUT_4[37856] = 32'b00000000000000001001111100010011;
assign LUT_4[37857] = 32'b00000000000000000011001000001011;
assign LUT_4[37858] = 32'b00000000000000001001010110110111;
assign LUT_4[37859] = 32'b00000000000000000010100010101111;
assign LUT_4[37860] = 32'b00000000000000000110111100101111;
assign LUT_4[37861] = 32'b00000000000000000000001000100111;
assign LUT_4[37862] = 32'b00000000000000000110010111010011;
assign LUT_4[37863] = 32'b11111111111111111111100011001011;
assign LUT_4[37864] = 32'b00000000000000000011001000101000;
assign LUT_4[37865] = 32'b11111111111111111100010100100000;
assign LUT_4[37866] = 32'b00000000000000000010100011001100;
assign LUT_4[37867] = 32'b11111111111111111011101111000100;
assign LUT_4[37868] = 32'b00000000000000000000001001000100;
assign LUT_4[37869] = 32'b11111111111111111001010100111100;
assign LUT_4[37870] = 32'b11111111111111111111100011101000;
assign LUT_4[37871] = 32'b11111111111111111000101111100000;
assign LUT_4[37872] = 32'b00000000000000000111101110000001;
assign LUT_4[37873] = 32'b00000000000000000000111001111001;
assign LUT_4[37874] = 32'b00000000000000000111001000100101;
assign LUT_4[37875] = 32'b00000000000000000000010100011101;
assign LUT_4[37876] = 32'b00000000000000000100101110011101;
assign LUT_4[37877] = 32'b11111111111111111101111010010101;
assign LUT_4[37878] = 32'b00000000000000000100001001000001;
assign LUT_4[37879] = 32'b11111111111111111101010100111001;
assign LUT_4[37880] = 32'b00000000000000000000111010010110;
assign LUT_4[37881] = 32'b11111111111111111010000110001110;
assign LUT_4[37882] = 32'b00000000000000000000010100111010;
assign LUT_4[37883] = 32'b11111111111111111001100000110010;
assign LUT_4[37884] = 32'b11111111111111111101111010110010;
assign LUT_4[37885] = 32'b11111111111111110111000110101010;
assign LUT_4[37886] = 32'b11111111111111111101010101010110;
assign LUT_4[37887] = 32'b11111111111111110110100001001110;
assign LUT_4[37888] = 32'b00000000000000000101001110100100;
assign LUT_4[37889] = 32'b11111111111111111110011010011100;
assign LUT_4[37890] = 32'b00000000000000000100101001001000;
assign LUT_4[37891] = 32'b11111111111111111101110101000000;
assign LUT_4[37892] = 32'b00000000000000000010001111000000;
assign LUT_4[37893] = 32'b11111111111111111011011010111000;
assign LUT_4[37894] = 32'b00000000000000000001101001100100;
assign LUT_4[37895] = 32'b11111111111111111010110101011100;
assign LUT_4[37896] = 32'b11111111111111111110011010111001;
assign LUT_4[37897] = 32'b11111111111111110111100110110001;
assign LUT_4[37898] = 32'b11111111111111111101110101011101;
assign LUT_4[37899] = 32'b11111111111111110111000001010101;
assign LUT_4[37900] = 32'b11111111111111111011011011010101;
assign LUT_4[37901] = 32'b11111111111111110100100111001101;
assign LUT_4[37902] = 32'b11111111111111111010110101111001;
assign LUT_4[37903] = 32'b11111111111111110100000001110001;
assign LUT_4[37904] = 32'b00000000000000000011000000010010;
assign LUT_4[37905] = 32'b11111111111111111100001100001010;
assign LUT_4[37906] = 32'b00000000000000000010011010110110;
assign LUT_4[37907] = 32'b11111111111111111011100110101110;
assign LUT_4[37908] = 32'b00000000000000000000000000101110;
assign LUT_4[37909] = 32'b11111111111111111001001100100110;
assign LUT_4[37910] = 32'b11111111111111111111011011010010;
assign LUT_4[37911] = 32'b11111111111111111000100111001010;
assign LUT_4[37912] = 32'b11111111111111111100001100100111;
assign LUT_4[37913] = 32'b11111111111111110101011000011111;
assign LUT_4[37914] = 32'b11111111111111111011100111001011;
assign LUT_4[37915] = 32'b11111111111111110100110011000011;
assign LUT_4[37916] = 32'b11111111111111111001001101000011;
assign LUT_4[37917] = 32'b11111111111111110010011000111011;
assign LUT_4[37918] = 32'b11111111111111111000100111100111;
assign LUT_4[37919] = 32'b11111111111111110001110011011111;
assign LUT_4[37920] = 32'b00000000000000000011101001101011;
assign LUT_4[37921] = 32'b11111111111111111100110101100011;
assign LUT_4[37922] = 32'b00000000000000000011000100001111;
assign LUT_4[37923] = 32'b11111111111111111100010000000111;
assign LUT_4[37924] = 32'b00000000000000000000101010000111;
assign LUT_4[37925] = 32'b11111111111111111001110101111111;
assign LUT_4[37926] = 32'b00000000000000000000000100101011;
assign LUT_4[37927] = 32'b11111111111111111001010000100011;
assign LUT_4[37928] = 32'b11111111111111111100110110000000;
assign LUT_4[37929] = 32'b11111111111111110110000001111000;
assign LUT_4[37930] = 32'b11111111111111111100010000100100;
assign LUT_4[37931] = 32'b11111111111111110101011100011100;
assign LUT_4[37932] = 32'b11111111111111111001110110011100;
assign LUT_4[37933] = 32'b11111111111111110011000010010100;
assign LUT_4[37934] = 32'b11111111111111111001010001000000;
assign LUT_4[37935] = 32'b11111111111111110010011100111000;
assign LUT_4[37936] = 32'b00000000000000000001011011011001;
assign LUT_4[37937] = 32'b11111111111111111010100111010001;
assign LUT_4[37938] = 32'b00000000000000000000110101111101;
assign LUT_4[37939] = 32'b11111111111111111010000001110101;
assign LUT_4[37940] = 32'b11111111111111111110011011110101;
assign LUT_4[37941] = 32'b11111111111111110111100111101101;
assign LUT_4[37942] = 32'b11111111111111111101110110011001;
assign LUT_4[37943] = 32'b11111111111111110111000010010001;
assign LUT_4[37944] = 32'b11111111111111111010100111101110;
assign LUT_4[37945] = 32'b11111111111111110011110011100110;
assign LUT_4[37946] = 32'b11111111111111111010000010010010;
assign LUT_4[37947] = 32'b11111111111111110011001110001010;
assign LUT_4[37948] = 32'b11111111111111110111101000001010;
assign LUT_4[37949] = 32'b11111111111111110000110100000010;
assign LUT_4[37950] = 32'b11111111111111110111000010101110;
assign LUT_4[37951] = 32'b11111111111111110000001110100110;
assign LUT_4[37952] = 32'b00000000000000000110100101111000;
assign LUT_4[37953] = 32'b11111111111111111111110001110000;
assign LUT_4[37954] = 32'b00000000000000000110000000011100;
assign LUT_4[37955] = 32'b11111111111111111111001100010100;
assign LUT_4[37956] = 32'b00000000000000000011100110010100;
assign LUT_4[37957] = 32'b11111111111111111100110010001100;
assign LUT_4[37958] = 32'b00000000000000000011000000111000;
assign LUT_4[37959] = 32'b11111111111111111100001100110000;
assign LUT_4[37960] = 32'b11111111111111111111110010001101;
assign LUT_4[37961] = 32'b11111111111111111000111110000101;
assign LUT_4[37962] = 32'b11111111111111111111001100110001;
assign LUT_4[37963] = 32'b11111111111111111000011000101001;
assign LUT_4[37964] = 32'b11111111111111111100110010101001;
assign LUT_4[37965] = 32'b11111111111111110101111110100001;
assign LUT_4[37966] = 32'b11111111111111111100001101001101;
assign LUT_4[37967] = 32'b11111111111111110101011001000101;
assign LUT_4[37968] = 32'b00000000000000000100010111100110;
assign LUT_4[37969] = 32'b11111111111111111101100011011110;
assign LUT_4[37970] = 32'b00000000000000000011110010001010;
assign LUT_4[37971] = 32'b11111111111111111100111110000010;
assign LUT_4[37972] = 32'b00000000000000000001011000000010;
assign LUT_4[37973] = 32'b11111111111111111010100011111010;
assign LUT_4[37974] = 32'b00000000000000000000110010100110;
assign LUT_4[37975] = 32'b11111111111111111001111110011110;
assign LUT_4[37976] = 32'b11111111111111111101100011111011;
assign LUT_4[37977] = 32'b11111111111111110110101111110011;
assign LUT_4[37978] = 32'b11111111111111111100111110011111;
assign LUT_4[37979] = 32'b11111111111111110110001010010111;
assign LUT_4[37980] = 32'b11111111111111111010100100010111;
assign LUT_4[37981] = 32'b11111111111111110011110000001111;
assign LUT_4[37982] = 32'b11111111111111111001111110111011;
assign LUT_4[37983] = 32'b11111111111111110011001010110011;
assign LUT_4[37984] = 32'b00000000000000000101000000111111;
assign LUT_4[37985] = 32'b11111111111111111110001100110111;
assign LUT_4[37986] = 32'b00000000000000000100011011100011;
assign LUT_4[37987] = 32'b11111111111111111101100111011011;
assign LUT_4[37988] = 32'b00000000000000000010000001011011;
assign LUT_4[37989] = 32'b11111111111111111011001101010011;
assign LUT_4[37990] = 32'b00000000000000000001011011111111;
assign LUT_4[37991] = 32'b11111111111111111010100111110111;
assign LUT_4[37992] = 32'b11111111111111111110001101010100;
assign LUT_4[37993] = 32'b11111111111111110111011001001100;
assign LUT_4[37994] = 32'b11111111111111111101100111111000;
assign LUT_4[37995] = 32'b11111111111111110110110011110000;
assign LUT_4[37996] = 32'b11111111111111111011001101110000;
assign LUT_4[37997] = 32'b11111111111111110100011001101000;
assign LUT_4[37998] = 32'b11111111111111111010101000010100;
assign LUT_4[37999] = 32'b11111111111111110011110100001100;
assign LUT_4[38000] = 32'b00000000000000000010110010101101;
assign LUT_4[38001] = 32'b11111111111111111011111110100101;
assign LUT_4[38002] = 32'b00000000000000000010001101010001;
assign LUT_4[38003] = 32'b11111111111111111011011001001001;
assign LUT_4[38004] = 32'b11111111111111111111110011001001;
assign LUT_4[38005] = 32'b11111111111111111000111111000001;
assign LUT_4[38006] = 32'b11111111111111111111001101101101;
assign LUT_4[38007] = 32'b11111111111111111000011001100101;
assign LUT_4[38008] = 32'b11111111111111111011111111000010;
assign LUT_4[38009] = 32'b11111111111111110101001010111010;
assign LUT_4[38010] = 32'b11111111111111111011011001100110;
assign LUT_4[38011] = 32'b11111111111111110100100101011110;
assign LUT_4[38012] = 32'b11111111111111111000111111011110;
assign LUT_4[38013] = 32'b11111111111111110010001011010110;
assign LUT_4[38014] = 32'b11111111111111111000011010000010;
assign LUT_4[38015] = 32'b11111111111111110001100101111010;
assign LUT_4[38016] = 32'b00000000000000000111110100101100;
assign LUT_4[38017] = 32'b00000000000000000001000000100100;
assign LUT_4[38018] = 32'b00000000000000000111001111010000;
assign LUT_4[38019] = 32'b00000000000000000000011011001000;
assign LUT_4[38020] = 32'b00000000000000000100110101001000;
assign LUT_4[38021] = 32'b11111111111111111110000001000000;
assign LUT_4[38022] = 32'b00000000000000000100001111101100;
assign LUT_4[38023] = 32'b11111111111111111101011011100100;
assign LUT_4[38024] = 32'b00000000000000000001000001000001;
assign LUT_4[38025] = 32'b11111111111111111010001100111001;
assign LUT_4[38026] = 32'b00000000000000000000011011100101;
assign LUT_4[38027] = 32'b11111111111111111001100111011101;
assign LUT_4[38028] = 32'b11111111111111111110000001011101;
assign LUT_4[38029] = 32'b11111111111111110111001101010101;
assign LUT_4[38030] = 32'b11111111111111111101011100000001;
assign LUT_4[38031] = 32'b11111111111111110110100111111001;
assign LUT_4[38032] = 32'b00000000000000000101100110011010;
assign LUT_4[38033] = 32'b11111111111111111110110010010010;
assign LUT_4[38034] = 32'b00000000000000000101000000111110;
assign LUT_4[38035] = 32'b11111111111111111110001100110110;
assign LUT_4[38036] = 32'b00000000000000000010100110110110;
assign LUT_4[38037] = 32'b11111111111111111011110010101110;
assign LUT_4[38038] = 32'b00000000000000000010000001011010;
assign LUT_4[38039] = 32'b11111111111111111011001101010010;
assign LUT_4[38040] = 32'b11111111111111111110110010101111;
assign LUT_4[38041] = 32'b11111111111111110111111110100111;
assign LUT_4[38042] = 32'b11111111111111111110001101010011;
assign LUT_4[38043] = 32'b11111111111111110111011001001011;
assign LUT_4[38044] = 32'b11111111111111111011110011001011;
assign LUT_4[38045] = 32'b11111111111111110100111111000011;
assign LUT_4[38046] = 32'b11111111111111111011001101101111;
assign LUT_4[38047] = 32'b11111111111111110100011001100111;
assign LUT_4[38048] = 32'b00000000000000000110001111110011;
assign LUT_4[38049] = 32'b11111111111111111111011011101011;
assign LUT_4[38050] = 32'b00000000000000000101101010010111;
assign LUT_4[38051] = 32'b11111111111111111110110110001111;
assign LUT_4[38052] = 32'b00000000000000000011010000001111;
assign LUT_4[38053] = 32'b11111111111111111100011100000111;
assign LUT_4[38054] = 32'b00000000000000000010101010110011;
assign LUT_4[38055] = 32'b11111111111111111011110110101011;
assign LUT_4[38056] = 32'b11111111111111111111011100001000;
assign LUT_4[38057] = 32'b11111111111111111000101000000000;
assign LUT_4[38058] = 32'b11111111111111111110110110101100;
assign LUT_4[38059] = 32'b11111111111111111000000010100100;
assign LUT_4[38060] = 32'b11111111111111111100011100100100;
assign LUT_4[38061] = 32'b11111111111111110101101000011100;
assign LUT_4[38062] = 32'b11111111111111111011110111001000;
assign LUT_4[38063] = 32'b11111111111111110101000011000000;
assign LUT_4[38064] = 32'b00000000000000000100000001100001;
assign LUT_4[38065] = 32'b11111111111111111101001101011001;
assign LUT_4[38066] = 32'b00000000000000000011011100000101;
assign LUT_4[38067] = 32'b11111111111111111100100111111101;
assign LUT_4[38068] = 32'b00000000000000000001000001111101;
assign LUT_4[38069] = 32'b11111111111111111010001101110101;
assign LUT_4[38070] = 32'b00000000000000000000011100100001;
assign LUT_4[38071] = 32'b11111111111111111001101000011001;
assign LUT_4[38072] = 32'b11111111111111111101001101110110;
assign LUT_4[38073] = 32'b11111111111111110110011001101110;
assign LUT_4[38074] = 32'b11111111111111111100101000011010;
assign LUT_4[38075] = 32'b11111111111111110101110100010010;
assign LUT_4[38076] = 32'b11111111111111111010001110010010;
assign LUT_4[38077] = 32'b11111111111111110011011010001010;
assign LUT_4[38078] = 32'b11111111111111111001101000110110;
assign LUT_4[38079] = 32'b11111111111111110010110100101110;
assign LUT_4[38080] = 32'b00000000000000001001001100000000;
assign LUT_4[38081] = 32'b00000000000000000010010111111000;
assign LUT_4[38082] = 32'b00000000000000001000100110100100;
assign LUT_4[38083] = 32'b00000000000000000001110010011100;
assign LUT_4[38084] = 32'b00000000000000000110001100011100;
assign LUT_4[38085] = 32'b11111111111111111111011000010100;
assign LUT_4[38086] = 32'b00000000000000000101100111000000;
assign LUT_4[38087] = 32'b11111111111111111110110010111000;
assign LUT_4[38088] = 32'b00000000000000000010011000010101;
assign LUT_4[38089] = 32'b11111111111111111011100100001101;
assign LUT_4[38090] = 32'b00000000000000000001110010111001;
assign LUT_4[38091] = 32'b11111111111111111010111110110001;
assign LUT_4[38092] = 32'b11111111111111111111011000110001;
assign LUT_4[38093] = 32'b11111111111111111000100100101001;
assign LUT_4[38094] = 32'b11111111111111111110110011010101;
assign LUT_4[38095] = 32'b11111111111111110111111111001101;
assign LUT_4[38096] = 32'b00000000000000000110111101101110;
assign LUT_4[38097] = 32'b00000000000000000000001001100110;
assign LUT_4[38098] = 32'b00000000000000000110011000010010;
assign LUT_4[38099] = 32'b11111111111111111111100100001010;
assign LUT_4[38100] = 32'b00000000000000000011111110001010;
assign LUT_4[38101] = 32'b11111111111111111101001010000010;
assign LUT_4[38102] = 32'b00000000000000000011011000101110;
assign LUT_4[38103] = 32'b11111111111111111100100100100110;
assign LUT_4[38104] = 32'b00000000000000000000001010000011;
assign LUT_4[38105] = 32'b11111111111111111001010101111011;
assign LUT_4[38106] = 32'b11111111111111111111100100100111;
assign LUT_4[38107] = 32'b11111111111111111000110000011111;
assign LUT_4[38108] = 32'b11111111111111111101001010011111;
assign LUT_4[38109] = 32'b11111111111111110110010110010111;
assign LUT_4[38110] = 32'b11111111111111111100100101000011;
assign LUT_4[38111] = 32'b11111111111111110101110000111011;
assign LUT_4[38112] = 32'b00000000000000000111100111000111;
assign LUT_4[38113] = 32'b00000000000000000000110010111111;
assign LUT_4[38114] = 32'b00000000000000000111000001101011;
assign LUT_4[38115] = 32'b00000000000000000000001101100011;
assign LUT_4[38116] = 32'b00000000000000000100100111100011;
assign LUT_4[38117] = 32'b11111111111111111101110011011011;
assign LUT_4[38118] = 32'b00000000000000000100000010000111;
assign LUT_4[38119] = 32'b11111111111111111101001101111111;
assign LUT_4[38120] = 32'b00000000000000000000110011011100;
assign LUT_4[38121] = 32'b11111111111111111001111111010100;
assign LUT_4[38122] = 32'b00000000000000000000001110000000;
assign LUT_4[38123] = 32'b11111111111111111001011001111000;
assign LUT_4[38124] = 32'b11111111111111111101110011111000;
assign LUT_4[38125] = 32'b11111111111111110110111111110000;
assign LUT_4[38126] = 32'b11111111111111111101001110011100;
assign LUT_4[38127] = 32'b11111111111111110110011010010100;
assign LUT_4[38128] = 32'b00000000000000000101011000110101;
assign LUT_4[38129] = 32'b11111111111111111110100100101101;
assign LUT_4[38130] = 32'b00000000000000000100110011011001;
assign LUT_4[38131] = 32'b11111111111111111101111111010001;
assign LUT_4[38132] = 32'b00000000000000000010011001010001;
assign LUT_4[38133] = 32'b11111111111111111011100101001001;
assign LUT_4[38134] = 32'b00000000000000000001110011110101;
assign LUT_4[38135] = 32'b11111111111111111010111111101101;
assign LUT_4[38136] = 32'b11111111111111111110100101001010;
assign LUT_4[38137] = 32'b11111111111111110111110001000010;
assign LUT_4[38138] = 32'b11111111111111111101111111101110;
assign LUT_4[38139] = 32'b11111111111111110111001011100110;
assign LUT_4[38140] = 32'b11111111111111111011100101100110;
assign LUT_4[38141] = 32'b11111111111111110100110001011110;
assign LUT_4[38142] = 32'b11111111111111111011000000001010;
assign LUT_4[38143] = 32'b11111111111111110100001100000010;
assign LUT_4[38144] = 32'b00000000000000001010001010000111;
assign LUT_4[38145] = 32'b00000000000000000011010101111111;
assign LUT_4[38146] = 32'b00000000000000001001100100101011;
assign LUT_4[38147] = 32'b00000000000000000010110000100011;
assign LUT_4[38148] = 32'b00000000000000000111001010100011;
assign LUT_4[38149] = 32'b00000000000000000000010110011011;
assign LUT_4[38150] = 32'b00000000000000000110100101000111;
assign LUT_4[38151] = 32'b11111111111111111111110000111111;
assign LUT_4[38152] = 32'b00000000000000000011010110011100;
assign LUT_4[38153] = 32'b11111111111111111100100010010100;
assign LUT_4[38154] = 32'b00000000000000000010110001000000;
assign LUT_4[38155] = 32'b11111111111111111011111100111000;
assign LUT_4[38156] = 32'b00000000000000000000010110111000;
assign LUT_4[38157] = 32'b11111111111111111001100010110000;
assign LUT_4[38158] = 32'b11111111111111111111110001011100;
assign LUT_4[38159] = 32'b11111111111111111000111101010100;
assign LUT_4[38160] = 32'b00000000000000000111111011110101;
assign LUT_4[38161] = 32'b00000000000000000001000111101101;
assign LUT_4[38162] = 32'b00000000000000000111010110011001;
assign LUT_4[38163] = 32'b00000000000000000000100010010001;
assign LUT_4[38164] = 32'b00000000000000000100111100010001;
assign LUT_4[38165] = 32'b11111111111111111110001000001001;
assign LUT_4[38166] = 32'b00000000000000000100010110110101;
assign LUT_4[38167] = 32'b11111111111111111101100010101101;
assign LUT_4[38168] = 32'b00000000000000000001001000001010;
assign LUT_4[38169] = 32'b11111111111111111010010100000010;
assign LUT_4[38170] = 32'b00000000000000000000100010101110;
assign LUT_4[38171] = 32'b11111111111111111001101110100110;
assign LUT_4[38172] = 32'b11111111111111111110001000100110;
assign LUT_4[38173] = 32'b11111111111111110111010100011110;
assign LUT_4[38174] = 32'b11111111111111111101100011001010;
assign LUT_4[38175] = 32'b11111111111111110110101111000010;
assign LUT_4[38176] = 32'b00000000000000001000100101001110;
assign LUT_4[38177] = 32'b00000000000000000001110001000110;
assign LUT_4[38178] = 32'b00000000000000000111111111110010;
assign LUT_4[38179] = 32'b00000000000000000001001011101010;
assign LUT_4[38180] = 32'b00000000000000000101100101101010;
assign LUT_4[38181] = 32'b11111111111111111110110001100010;
assign LUT_4[38182] = 32'b00000000000000000101000000001110;
assign LUT_4[38183] = 32'b11111111111111111110001100000110;
assign LUT_4[38184] = 32'b00000000000000000001110001100011;
assign LUT_4[38185] = 32'b11111111111111111010111101011011;
assign LUT_4[38186] = 32'b00000000000000000001001100000111;
assign LUT_4[38187] = 32'b11111111111111111010010111111111;
assign LUT_4[38188] = 32'b11111111111111111110110001111111;
assign LUT_4[38189] = 32'b11111111111111110111111101110111;
assign LUT_4[38190] = 32'b11111111111111111110001100100011;
assign LUT_4[38191] = 32'b11111111111111110111011000011011;
assign LUT_4[38192] = 32'b00000000000000000110010110111100;
assign LUT_4[38193] = 32'b11111111111111111111100010110100;
assign LUT_4[38194] = 32'b00000000000000000101110001100000;
assign LUT_4[38195] = 32'b11111111111111111110111101011000;
assign LUT_4[38196] = 32'b00000000000000000011010111011000;
assign LUT_4[38197] = 32'b11111111111111111100100011010000;
assign LUT_4[38198] = 32'b00000000000000000010110001111100;
assign LUT_4[38199] = 32'b11111111111111111011111101110100;
assign LUT_4[38200] = 32'b11111111111111111111100011010001;
assign LUT_4[38201] = 32'b11111111111111111000101111001001;
assign LUT_4[38202] = 32'b11111111111111111110111101110101;
assign LUT_4[38203] = 32'b11111111111111111000001001101101;
assign LUT_4[38204] = 32'b11111111111111111100100011101101;
assign LUT_4[38205] = 32'b11111111111111110101101111100101;
assign LUT_4[38206] = 32'b11111111111111111011111110010001;
assign LUT_4[38207] = 32'b11111111111111110101001010001001;
assign LUT_4[38208] = 32'b00000000000000001011100001011011;
assign LUT_4[38209] = 32'b00000000000000000100101101010011;
assign LUT_4[38210] = 32'b00000000000000001010111011111111;
assign LUT_4[38211] = 32'b00000000000000000100000111110111;
assign LUT_4[38212] = 32'b00000000000000001000100001110111;
assign LUT_4[38213] = 32'b00000000000000000001101101101111;
assign LUT_4[38214] = 32'b00000000000000000111111100011011;
assign LUT_4[38215] = 32'b00000000000000000001001000010011;
assign LUT_4[38216] = 32'b00000000000000000100101101110000;
assign LUT_4[38217] = 32'b11111111111111111101111001101000;
assign LUT_4[38218] = 32'b00000000000000000100001000010100;
assign LUT_4[38219] = 32'b11111111111111111101010100001100;
assign LUT_4[38220] = 32'b00000000000000000001101110001100;
assign LUT_4[38221] = 32'b11111111111111111010111010000100;
assign LUT_4[38222] = 32'b00000000000000000001001000110000;
assign LUT_4[38223] = 32'b11111111111111111010010100101000;
assign LUT_4[38224] = 32'b00000000000000001001010011001001;
assign LUT_4[38225] = 32'b00000000000000000010011111000001;
assign LUT_4[38226] = 32'b00000000000000001000101101101101;
assign LUT_4[38227] = 32'b00000000000000000001111001100101;
assign LUT_4[38228] = 32'b00000000000000000110010011100101;
assign LUT_4[38229] = 32'b11111111111111111111011111011101;
assign LUT_4[38230] = 32'b00000000000000000101101110001001;
assign LUT_4[38231] = 32'b11111111111111111110111010000001;
assign LUT_4[38232] = 32'b00000000000000000010011111011110;
assign LUT_4[38233] = 32'b11111111111111111011101011010110;
assign LUT_4[38234] = 32'b00000000000000000001111010000010;
assign LUT_4[38235] = 32'b11111111111111111011000101111010;
assign LUT_4[38236] = 32'b11111111111111111111011111111010;
assign LUT_4[38237] = 32'b11111111111111111000101011110010;
assign LUT_4[38238] = 32'b11111111111111111110111010011110;
assign LUT_4[38239] = 32'b11111111111111111000000110010110;
assign LUT_4[38240] = 32'b00000000000000001001111100100010;
assign LUT_4[38241] = 32'b00000000000000000011001000011010;
assign LUT_4[38242] = 32'b00000000000000001001010111000110;
assign LUT_4[38243] = 32'b00000000000000000010100010111110;
assign LUT_4[38244] = 32'b00000000000000000110111100111110;
assign LUT_4[38245] = 32'b00000000000000000000001000110110;
assign LUT_4[38246] = 32'b00000000000000000110010111100010;
assign LUT_4[38247] = 32'b11111111111111111111100011011010;
assign LUT_4[38248] = 32'b00000000000000000011001000110111;
assign LUT_4[38249] = 32'b11111111111111111100010100101111;
assign LUT_4[38250] = 32'b00000000000000000010100011011011;
assign LUT_4[38251] = 32'b11111111111111111011101111010011;
assign LUT_4[38252] = 32'b00000000000000000000001001010011;
assign LUT_4[38253] = 32'b11111111111111111001010101001011;
assign LUT_4[38254] = 32'b11111111111111111111100011110111;
assign LUT_4[38255] = 32'b11111111111111111000101111101111;
assign LUT_4[38256] = 32'b00000000000000000111101110010000;
assign LUT_4[38257] = 32'b00000000000000000000111010001000;
assign LUT_4[38258] = 32'b00000000000000000111001000110100;
assign LUT_4[38259] = 32'b00000000000000000000010100101100;
assign LUT_4[38260] = 32'b00000000000000000100101110101100;
assign LUT_4[38261] = 32'b11111111111111111101111010100100;
assign LUT_4[38262] = 32'b00000000000000000100001001010000;
assign LUT_4[38263] = 32'b11111111111111111101010101001000;
assign LUT_4[38264] = 32'b00000000000000000000111010100101;
assign LUT_4[38265] = 32'b11111111111111111010000110011101;
assign LUT_4[38266] = 32'b00000000000000000000010101001001;
assign LUT_4[38267] = 32'b11111111111111111001100001000001;
assign LUT_4[38268] = 32'b11111111111111111101111011000001;
assign LUT_4[38269] = 32'b11111111111111110111000110111001;
assign LUT_4[38270] = 32'b11111111111111111101010101100101;
assign LUT_4[38271] = 32'b11111111111111110110100001011101;
assign LUT_4[38272] = 32'b00000000000000001100110000001111;
assign LUT_4[38273] = 32'b00000000000000000101111100000111;
assign LUT_4[38274] = 32'b00000000000000001100001010110011;
assign LUT_4[38275] = 32'b00000000000000000101010110101011;
assign LUT_4[38276] = 32'b00000000000000001001110000101011;
assign LUT_4[38277] = 32'b00000000000000000010111100100011;
assign LUT_4[38278] = 32'b00000000000000001001001011001111;
assign LUT_4[38279] = 32'b00000000000000000010010111000111;
assign LUT_4[38280] = 32'b00000000000000000101111100100100;
assign LUT_4[38281] = 32'b11111111111111111111001000011100;
assign LUT_4[38282] = 32'b00000000000000000101010111001000;
assign LUT_4[38283] = 32'b11111111111111111110100011000000;
assign LUT_4[38284] = 32'b00000000000000000010111101000000;
assign LUT_4[38285] = 32'b11111111111111111100001000111000;
assign LUT_4[38286] = 32'b00000000000000000010010111100100;
assign LUT_4[38287] = 32'b11111111111111111011100011011100;
assign LUT_4[38288] = 32'b00000000000000001010100001111101;
assign LUT_4[38289] = 32'b00000000000000000011101101110101;
assign LUT_4[38290] = 32'b00000000000000001001111100100001;
assign LUT_4[38291] = 32'b00000000000000000011001000011001;
assign LUT_4[38292] = 32'b00000000000000000111100010011001;
assign LUT_4[38293] = 32'b00000000000000000000101110010001;
assign LUT_4[38294] = 32'b00000000000000000110111100111101;
assign LUT_4[38295] = 32'b00000000000000000000001000110101;
assign LUT_4[38296] = 32'b00000000000000000011101110010010;
assign LUT_4[38297] = 32'b11111111111111111100111010001010;
assign LUT_4[38298] = 32'b00000000000000000011001000110110;
assign LUT_4[38299] = 32'b11111111111111111100010100101110;
assign LUT_4[38300] = 32'b00000000000000000000101110101110;
assign LUT_4[38301] = 32'b11111111111111111001111010100110;
assign LUT_4[38302] = 32'b00000000000000000000001001010010;
assign LUT_4[38303] = 32'b11111111111111111001010101001010;
assign LUT_4[38304] = 32'b00000000000000001011001011010110;
assign LUT_4[38305] = 32'b00000000000000000100010111001110;
assign LUT_4[38306] = 32'b00000000000000001010100101111010;
assign LUT_4[38307] = 32'b00000000000000000011110001110010;
assign LUT_4[38308] = 32'b00000000000000001000001011110010;
assign LUT_4[38309] = 32'b00000000000000000001010111101010;
assign LUT_4[38310] = 32'b00000000000000000111100110010110;
assign LUT_4[38311] = 32'b00000000000000000000110010001110;
assign LUT_4[38312] = 32'b00000000000000000100010111101011;
assign LUT_4[38313] = 32'b11111111111111111101100011100011;
assign LUT_4[38314] = 32'b00000000000000000011110010001111;
assign LUT_4[38315] = 32'b11111111111111111100111110000111;
assign LUT_4[38316] = 32'b00000000000000000001011000000111;
assign LUT_4[38317] = 32'b11111111111111111010100011111111;
assign LUT_4[38318] = 32'b00000000000000000000110010101011;
assign LUT_4[38319] = 32'b11111111111111111001111110100011;
assign LUT_4[38320] = 32'b00000000000000001000111101000100;
assign LUT_4[38321] = 32'b00000000000000000010001000111100;
assign LUT_4[38322] = 32'b00000000000000001000010111101000;
assign LUT_4[38323] = 32'b00000000000000000001100011100000;
assign LUT_4[38324] = 32'b00000000000000000101111101100000;
assign LUT_4[38325] = 32'b11111111111111111111001001011000;
assign LUT_4[38326] = 32'b00000000000000000101011000000100;
assign LUT_4[38327] = 32'b11111111111111111110100011111100;
assign LUT_4[38328] = 32'b00000000000000000010001001011001;
assign LUT_4[38329] = 32'b11111111111111111011010101010001;
assign LUT_4[38330] = 32'b00000000000000000001100011111101;
assign LUT_4[38331] = 32'b11111111111111111010101111110101;
assign LUT_4[38332] = 32'b11111111111111111111001001110101;
assign LUT_4[38333] = 32'b11111111111111111000010101101101;
assign LUT_4[38334] = 32'b11111111111111111110100100011001;
assign LUT_4[38335] = 32'b11111111111111110111110000010001;
assign LUT_4[38336] = 32'b00000000000000001110000111100011;
assign LUT_4[38337] = 32'b00000000000000000111010011011011;
assign LUT_4[38338] = 32'b00000000000000001101100010000111;
assign LUT_4[38339] = 32'b00000000000000000110101101111111;
assign LUT_4[38340] = 32'b00000000000000001011000111111111;
assign LUT_4[38341] = 32'b00000000000000000100010011110111;
assign LUT_4[38342] = 32'b00000000000000001010100010100011;
assign LUT_4[38343] = 32'b00000000000000000011101110011011;
assign LUT_4[38344] = 32'b00000000000000000111010011111000;
assign LUT_4[38345] = 32'b00000000000000000000011111110000;
assign LUT_4[38346] = 32'b00000000000000000110101110011100;
assign LUT_4[38347] = 32'b11111111111111111111111010010100;
assign LUT_4[38348] = 32'b00000000000000000100010100010100;
assign LUT_4[38349] = 32'b11111111111111111101100000001100;
assign LUT_4[38350] = 32'b00000000000000000011101110111000;
assign LUT_4[38351] = 32'b11111111111111111100111010110000;
assign LUT_4[38352] = 32'b00000000000000001011111001010001;
assign LUT_4[38353] = 32'b00000000000000000101000101001001;
assign LUT_4[38354] = 32'b00000000000000001011010011110101;
assign LUT_4[38355] = 32'b00000000000000000100011111101101;
assign LUT_4[38356] = 32'b00000000000000001000111001101101;
assign LUT_4[38357] = 32'b00000000000000000010000101100101;
assign LUT_4[38358] = 32'b00000000000000001000010100010001;
assign LUT_4[38359] = 32'b00000000000000000001100000001001;
assign LUT_4[38360] = 32'b00000000000000000101000101100110;
assign LUT_4[38361] = 32'b11111111111111111110010001011110;
assign LUT_4[38362] = 32'b00000000000000000100100000001010;
assign LUT_4[38363] = 32'b11111111111111111101101100000010;
assign LUT_4[38364] = 32'b00000000000000000010000110000010;
assign LUT_4[38365] = 32'b11111111111111111011010001111010;
assign LUT_4[38366] = 32'b00000000000000000001100000100110;
assign LUT_4[38367] = 32'b11111111111111111010101100011110;
assign LUT_4[38368] = 32'b00000000000000001100100010101010;
assign LUT_4[38369] = 32'b00000000000000000101101110100010;
assign LUT_4[38370] = 32'b00000000000000001011111101001110;
assign LUT_4[38371] = 32'b00000000000000000101001001000110;
assign LUT_4[38372] = 32'b00000000000000001001100011000110;
assign LUT_4[38373] = 32'b00000000000000000010101110111110;
assign LUT_4[38374] = 32'b00000000000000001000111101101010;
assign LUT_4[38375] = 32'b00000000000000000010001001100010;
assign LUT_4[38376] = 32'b00000000000000000101101110111111;
assign LUT_4[38377] = 32'b11111111111111111110111010110111;
assign LUT_4[38378] = 32'b00000000000000000101001001100011;
assign LUT_4[38379] = 32'b11111111111111111110010101011011;
assign LUT_4[38380] = 32'b00000000000000000010101111011011;
assign LUT_4[38381] = 32'b11111111111111111011111011010011;
assign LUT_4[38382] = 32'b00000000000000000010001001111111;
assign LUT_4[38383] = 32'b11111111111111111011010101110111;
assign LUT_4[38384] = 32'b00000000000000001010010100011000;
assign LUT_4[38385] = 32'b00000000000000000011100000010000;
assign LUT_4[38386] = 32'b00000000000000001001101110111100;
assign LUT_4[38387] = 32'b00000000000000000010111010110100;
assign LUT_4[38388] = 32'b00000000000000000111010100110100;
assign LUT_4[38389] = 32'b00000000000000000000100000101100;
assign LUT_4[38390] = 32'b00000000000000000110101111011000;
assign LUT_4[38391] = 32'b11111111111111111111111011010000;
assign LUT_4[38392] = 32'b00000000000000000011100000101101;
assign LUT_4[38393] = 32'b11111111111111111100101100100101;
assign LUT_4[38394] = 32'b00000000000000000010111011010001;
assign LUT_4[38395] = 32'b11111111111111111100000111001001;
assign LUT_4[38396] = 32'b00000000000000000000100001001001;
assign LUT_4[38397] = 32'b11111111111111111001101101000001;
assign LUT_4[38398] = 32'b11111111111111111111111011101101;
assign LUT_4[38399] = 32'b11111111111111111001000111100101;
assign LUT_4[38400] = 32'b00000000000000000100010010101100;
assign LUT_4[38401] = 32'b11111111111111111101011110100100;
assign LUT_4[38402] = 32'b00000000000000000011101101010000;
assign LUT_4[38403] = 32'b11111111111111111100111001001000;
assign LUT_4[38404] = 32'b00000000000000000001010011001000;
assign LUT_4[38405] = 32'b11111111111111111010011111000000;
assign LUT_4[38406] = 32'b00000000000000000000101101101100;
assign LUT_4[38407] = 32'b11111111111111111001111001100100;
assign LUT_4[38408] = 32'b11111111111111111101011111000001;
assign LUT_4[38409] = 32'b11111111111111110110101010111001;
assign LUT_4[38410] = 32'b11111111111111111100111001100101;
assign LUT_4[38411] = 32'b11111111111111110110000101011101;
assign LUT_4[38412] = 32'b11111111111111111010011111011101;
assign LUT_4[38413] = 32'b11111111111111110011101011010101;
assign LUT_4[38414] = 32'b11111111111111111001111010000001;
assign LUT_4[38415] = 32'b11111111111111110011000101111001;
assign LUT_4[38416] = 32'b00000000000000000010000100011010;
assign LUT_4[38417] = 32'b11111111111111111011010000010010;
assign LUT_4[38418] = 32'b00000000000000000001011110111110;
assign LUT_4[38419] = 32'b11111111111111111010101010110110;
assign LUT_4[38420] = 32'b11111111111111111111000100110110;
assign LUT_4[38421] = 32'b11111111111111111000010000101110;
assign LUT_4[38422] = 32'b11111111111111111110011111011010;
assign LUT_4[38423] = 32'b11111111111111110111101011010010;
assign LUT_4[38424] = 32'b11111111111111111011010000101111;
assign LUT_4[38425] = 32'b11111111111111110100011100100111;
assign LUT_4[38426] = 32'b11111111111111111010101011010011;
assign LUT_4[38427] = 32'b11111111111111110011110111001011;
assign LUT_4[38428] = 32'b11111111111111111000010001001011;
assign LUT_4[38429] = 32'b11111111111111110001011101000011;
assign LUT_4[38430] = 32'b11111111111111110111101011101111;
assign LUT_4[38431] = 32'b11111111111111110000110111100111;
assign LUT_4[38432] = 32'b00000000000000000010101101110011;
assign LUT_4[38433] = 32'b11111111111111111011111001101011;
assign LUT_4[38434] = 32'b00000000000000000010001000010111;
assign LUT_4[38435] = 32'b11111111111111111011010100001111;
assign LUT_4[38436] = 32'b11111111111111111111101110001111;
assign LUT_4[38437] = 32'b11111111111111111000111010000111;
assign LUT_4[38438] = 32'b11111111111111111111001000110011;
assign LUT_4[38439] = 32'b11111111111111111000010100101011;
assign LUT_4[38440] = 32'b11111111111111111011111010001000;
assign LUT_4[38441] = 32'b11111111111111110101000110000000;
assign LUT_4[38442] = 32'b11111111111111111011010100101100;
assign LUT_4[38443] = 32'b11111111111111110100100000100100;
assign LUT_4[38444] = 32'b11111111111111111000111010100100;
assign LUT_4[38445] = 32'b11111111111111110010000110011100;
assign LUT_4[38446] = 32'b11111111111111111000010101001000;
assign LUT_4[38447] = 32'b11111111111111110001100001000000;
assign LUT_4[38448] = 32'b00000000000000000000011111100001;
assign LUT_4[38449] = 32'b11111111111111111001101011011001;
assign LUT_4[38450] = 32'b11111111111111111111111010000101;
assign LUT_4[38451] = 32'b11111111111111111001000101111101;
assign LUT_4[38452] = 32'b11111111111111111101011111111101;
assign LUT_4[38453] = 32'b11111111111111110110101011110101;
assign LUT_4[38454] = 32'b11111111111111111100111010100001;
assign LUT_4[38455] = 32'b11111111111111110110000110011001;
assign LUT_4[38456] = 32'b11111111111111111001101011110110;
assign LUT_4[38457] = 32'b11111111111111110010110111101110;
assign LUT_4[38458] = 32'b11111111111111111001000110011010;
assign LUT_4[38459] = 32'b11111111111111110010010010010010;
assign LUT_4[38460] = 32'b11111111111111110110101100010010;
assign LUT_4[38461] = 32'b11111111111111101111111000001010;
assign LUT_4[38462] = 32'b11111111111111110110000110110110;
assign LUT_4[38463] = 32'b11111111111111101111010010101110;
assign LUT_4[38464] = 32'b00000000000000000101101010000000;
assign LUT_4[38465] = 32'b11111111111111111110110101111000;
assign LUT_4[38466] = 32'b00000000000000000101000100100100;
assign LUT_4[38467] = 32'b11111111111111111110010000011100;
assign LUT_4[38468] = 32'b00000000000000000010101010011100;
assign LUT_4[38469] = 32'b11111111111111111011110110010100;
assign LUT_4[38470] = 32'b00000000000000000010000101000000;
assign LUT_4[38471] = 32'b11111111111111111011010000111000;
assign LUT_4[38472] = 32'b11111111111111111110110110010101;
assign LUT_4[38473] = 32'b11111111111111111000000010001101;
assign LUT_4[38474] = 32'b11111111111111111110010000111001;
assign LUT_4[38475] = 32'b11111111111111110111011100110001;
assign LUT_4[38476] = 32'b11111111111111111011110110110001;
assign LUT_4[38477] = 32'b11111111111111110101000010101001;
assign LUT_4[38478] = 32'b11111111111111111011010001010101;
assign LUT_4[38479] = 32'b11111111111111110100011101001101;
assign LUT_4[38480] = 32'b00000000000000000011011011101110;
assign LUT_4[38481] = 32'b11111111111111111100100111100110;
assign LUT_4[38482] = 32'b00000000000000000010110110010010;
assign LUT_4[38483] = 32'b11111111111111111100000010001010;
assign LUT_4[38484] = 32'b00000000000000000000011100001010;
assign LUT_4[38485] = 32'b11111111111111111001101000000010;
assign LUT_4[38486] = 32'b11111111111111111111110110101110;
assign LUT_4[38487] = 32'b11111111111111111001000010100110;
assign LUT_4[38488] = 32'b11111111111111111100101000000011;
assign LUT_4[38489] = 32'b11111111111111110101110011111011;
assign LUT_4[38490] = 32'b11111111111111111100000010100111;
assign LUT_4[38491] = 32'b11111111111111110101001110011111;
assign LUT_4[38492] = 32'b11111111111111111001101000011111;
assign LUT_4[38493] = 32'b11111111111111110010110100010111;
assign LUT_4[38494] = 32'b11111111111111111001000011000011;
assign LUT_4[38495] = 32'b11111111111111110010001110111011;
assign LUT_4[38496] = 32'b00000000000000000100000101000111;
assign LUT_4[38497] = 32'b11111111111111111101010000111111;
assign LUT_4[38498] = 32'b00000000000000000011011111101011;
assign LUT_4[38499] = 32'b11111111111111111100101011100011;
assign LUT_4[38500] = 32'b00000000000000000001000101100011;
assign LUT_4[38501] = 32'b11111111111111111010010001011011;
assign LUT_4[38502] = 32'b00000000000000000000100000000111;
assign LUT_4[38503] = 32'b11111111111111111001101011111111;
assign LUT_4[38504] = 32'b11111111111111111101010001011100;
assign LUT_4[38505] = 32'b11111111111111110110011101010100;
assign LUT_4[38506] = 32'b11111111111111111100101100000000;
assign LUT_4[38507] = 32'b11111111111111110101110111111000;
assign LUT_4[38508] = 32'b11111111111111111010010001111000;
assign LUT_4[38509] = 32'b11111111111111110011011101110000;
assign LUT_4[38510] = 32'b11111111111111111001101100011100;
assign LUT_4[38511] = 32'b11111111111111110010111000010100;
assign LUT_4[38512] = 32'b00000000000000000001110110110101;
assign LUT_4[38513] = 32'b11111111111111111011000010101101;
assign LUT_4[38514] = 32'b00000000000000000001010001011001;
assign LUT_4[38515] = 32'b11111111111111111010011101010001;
assign LUT_4[38516] = 32'b11111111111111111110110111010001;
assign LUT_4[38517] = 32'b11111111111111111000000011001001;
assign LUT_4[38518] = 32'b11111111111111111110010001110101;
assign LUT_4[38519] = 32'b11111111111111110111011101101101;
assign LUT_4[38520] = 32'b11111111111111111011000011001010;
assign LUT_4[38521] = 32'b11111111111111110100001111000010;
assign LUT_4[38522] = 32'b11111111111111111010011101101110;
assign LUT_4[38523] = 32'b11111111111111110011101001100110;
assign LUT_4[38524] = 32'b11111111111111111000000011100110;
assign LUT_4[38525] = 32'b11111111111111110001001111011110;
assign LUT_4[38526] = 32'b11111111111111110111011110001010;
assign LUT_4[38527] = 32'b11111111111111110000101010000010;
assign LUT_4[38528] = 32'b00000000000000000110111000110100;
assign LUT_4[38529] = 32'b00000000000000000000000100101100;
assign LUT_4[38530] = 32'b00000000000000000110010011011000;
assign LUT_4[38531] = 32'b11111111111111111111011111010000;
assign LUT_4[38532] = 32'b00000000000000000011111001010000;
assign LUT_4[38533] = 32'b11111111111111111101000101001000;
assign LUT_4[38534] = 32'b00000000000000000011010011110100;
assign LUT_4[38535] = 32'b11111111111111111100011111101100;
assign LUT_4[38536] = 32'b00000000000000000000000101001001;
assign LUT_4[38537] = 32'b11111111111111111001010001000001;
assign LUT_4[38538] = 32'b11111111111111111111011111101101;
assign LUT_4[38539] = 32'b11111111111111111000101011100101;
assign LUT_4[38540] = 32'b11111111111111111101000101100101;
assign LUT_4[38541] = 32'b11111111111111110110010001011101;
assign LUT_4[38542] = 32'b11111111111111111100100000001001;
assign LUT_4[38543] = 32'b11111111111111110101101100000001;
assign LUT_4[38544] = 32'b00000000000000000100101010100010;
assign LUT_4[38545] = 32'b11111111111111111101110110011010;
assign LUT_4[38546] = 32'b00000000000000000100000101000110;
assign LUT_4[38547] = 32'b11111111111111111101010000111110;
assign LUT_4[38548] = 32'b00000000000000000001101010111110;
assign LUT_4[38549] = 32'b11111111111111111010110110110110;
assign LUT_4[38550] = 32'b00000000000000000001000101100010;
assign LUT_4[38551] = 32'b11111111111111111010010001011010;
assign LUT_4[38552] = 32'b11111111111111111101110110110111;
assign LUT_4[38553] = 32'b11111111111111110111000010101111;
assign LUT_4[38554] = 32'b11111111111111111101010001011011;
assign LUT_4[38555] = 32'b11111111111111110110011101010011;
assign LUT_4[38556] = 32'b11111111111111111010110111010011;
assign LUT_4[38557] = 32'b11111111111111110100000011001011;
assign LUT_4[38558] = 32'b11111111111111111010010001110111;
assign LUT_4[38559] = 32'b11111111111111110011011101101111;
assign LUT_4[38560] = 32'b00000000000000000101010011111011;
assign LUT_4[38561] = 32'b11111111111111111110011111110011;
assign LUT_4[38562] = 32'b00000000000000000100101110011111;
assign LUT_4[38563] = 32'b11111111111111111101111010010111;
assign LUT_4[38564] = 32'b00000000000000000010010100010111;
assign LUT_4[38565] = 32'b11111111111111111011100000001111;
assign LUT_4[38566] = 32'b00000000000000000001101110111011;
assign LUT_4[38567] = 32'b11111111111111111010111010110011;
assign LUT_4[38568] = 32'b11111111111111111110100000010000;
assign LUT_4[38569] = 32'b11111111111111110111101100001000;
assign LUT_4[38570] = 32'b11111111111111111101111010110100;
assign LUT_4[38571] = 32'b11111111111111110111000110101100;
assign LUT_4[38572] = 32'b11111111111111111011100000101100;
assign LUT_4[38573] = 32'b11111111111111110100101100100100;
assign LUT_4[38574] = 32'b11111111111111111010111011010000;
assign LUT_4[38575] = 32'b11111111111111110100000111001000;
assign LUT_4[38576] = 32'b00000000000000000011000101101001;
assign LUT_4[38577] = 32'b11111111111111111100010001100001;
assign LUT_4[38578] = 32'b00000000000000000010100000001101;
assign LUT_4[38579] = 32'b11111111111111111011101100000101;
assign LUT_4[38580] = 32'b00000000000000000000000110000101;
assign LUT_4[38581] = 32'b11111111111111111001010001111101;
assign LUT_4[38582] = 32'b11111111111111111111100000101001;
assign LUT_4[38583] = 32'b11111111111111111000101100100001;
assign LUT_4[38584] = 32'b11111111111111111100010001111110;
assign LUT_4[38585] = 32'b11111111111111110101011101110110;
assign LUT_4[38586] = 32'b11111111111111111011101100100010;
assign LUT_4[38587] = 32'b11111111111111110100111000011010;
assign LUT_4[38588] = 32'b11111111111111111001010010011010;
assign LUT_4[38589] = 32'b11111111111111110010011110010010;
assign LUT_4[38590] = 32'b11111111111111111000101100111110;
assign LUT_4[38591] = 32'b11111111111111110001111000110110;
assign LUT_4[38592] = 32'b00000000000000001000010000001000;
assign LUT_4[38593] = 32'b00000000000000000001011100000000;
assign LUT_4[38594] = 32'b00000000000000000111101010101100;
assign LUT_4[38595] = 32'b00000000000000000000110110100100;
assign LUT_4[38596] = 32'b00000000000000000101010000100100;
assign LUT_4[38597] = 32'b11111111111111111110011100011100;
assign LUT_4[38598] = 32'b00000000000000000100101011001000;
assign LUT_4[38599] = 32'b11111111111111111101110111000000;
assign LUT_4[38600] = 32'b00000000000000000001011100011101;
assign LUT_4[38601] = 32'b11111111111111111010101000010101;
assign LUT_4[38602] = 32'b00000000000000000000110111000001;
assign LUT_4[38603] = 32'b11111111111111111010000010111001;
assign LUT_4[38604] = 32'b11111111111111111110011100111001;
assign LUT_4[38605] = 32'b11111111111111110111101000110001;
assign LUT_4[38606] = 32'b11111111111111111101110111011101;
assign LUT_4[38607] = 32'b11111111111111110111000011010101;
assign LUT_4[38608] = 32'b00000000000000000110000001110110;
assign LUT_4[38609] = 32'b11111111111111111111001101101110;
assign LUT_4[38610] = 32'b00000000000000000101011100011010;
assign LUT_4[38611] = 32'b11111111111111111110101000010010;
assign LUT_4[38612] = 32'b00000000000000000011000010010010;
assign LUT_4[38613] = 32'b11111111111111111100001110001010;
assign LUT_4[38614] = 32'b00000000000000000010011100110110;
assign LUT_4[38615] = 32'b11111111111111111011101000101110;
assign LUT_4[38616] = 32'b11111111111111111111001110001011;
assign LUT_4[38617] = 32'b11111111111111111000011010000011;
assign LUT_4[38618] = 32'b11111111111111111110101000101111;
assign LUT_4[38619] = 32'b11111111111111110111110100100111;
assign LUT_4[38620] = 32'b11111111111111111100001110100111;
assign LUT_4[38621] = 32'b11111111111111110101011010011111;
assign LUT_4[38622] = 32'b11111111111111111011101001001011;
assign LUT_4[38623] = 32'b11111111111111110100110101000011;
assign LUT_4[38624] = 32'b00000000000000000110101011001111;
assign LUT_4[38625] = 32'b11111111111111111111110111000111;
assign LUT_4[38626] = 32'b00000000000000000110000101110011;
assign LUT_4[38627] = 32'b11111111111111111111010001101011;
assign LUT_4[38628] = 32'b00000000000000000011101011101011;
assign LUT_4[38629] = 32'b11111111111111111100110111100011;
assign LUT_4[38630] = 32'b00000000000000000011000110001111;
assign LUT_4[38631] = 32'b11111111111111111100010010000111;
assign LUT_4[38632] = 32'b11111111111111111111110111100100;
assign LUT_4[38633] = 32'b11111111111111111001000011011100;
assign LUT_4[38634] = 32'b11111111111111111111010010001000;
assign LUT_4[38635] = 32'b11111111111111111000011110000000;
assign LUT_4[38636] = 32'b11111111111111111100111000000000;
assign LUT_4[38637] = 32'b11111111111111110110000011111000;
assign LUT_4[38638] = 32'b11111111111111111100010010100100;
assign LUT_4[38639] = 32'b11111111111111110101011110011100;
assign LUT_4[38640] = 32'b00000000000000000100011100111101;
assign LUT_4[38641] = 32'b11111111111111111101101000110101;
assign LUT_4[38642] = 32'b00000000000000000011110111100001;
assign LUT_4[38643] = 32'b11111111111111111101000011011001;
assign LUT_4[38644] = 32'b00000000000000000001011101011001;
assign LUT_4[38645] = 32'b11111111111111111010101001010001;
assign LUT_4[38646] = 32'b00000000000000000000110111111101;
assign LUT_4[38647] = 32'b11111111111111111010000011110101;
assign LUT_4[38648] = 32'b11111111111111111101101001010010;
assign LUT_4[38649] = 32'b11111111111111110110110101001010;
assign LUT_4[38650] = 32'b11111111111111111101000011110110;
assign LUT_4[38651] = 32'b11111111111111110110001111101110;
assign LUT_4[38652] = 32'b11111111111111111010101001101110;
assign LUT_4[38653] = 32'b11111111111111110011110101100110;
assign LUT_4[38654] = 32'b11111111111111111010000100010010;
assign LUT_4[38655] = 32'b11111111111111110011010000001010;
assign LUT_4[38656] = 32'b00000000000000001001001110001111;
assign LUT_4[38657] = 32'b00000000000000000010011010000111;
assign LUT_4[38658] = 32'b00000000000000001000101000110011;
assign LUT_4[38659] = 32'b00000000000000000001110100101011;
assign LUT_4[38660] = 32'b00000000000000000110001110101011;
assign LUT_4[38661] = 32'b11111111111111111111011010100011;
assign LUT_4[38662] = 32'b00000000000000000101101001001111;
assign LUT_4[38663] = 32'b11111111111111111110110101000111;
assign LUT_4[38664] = 32'b00000000000000000010011010100100;
assign LUT_4[38665] = 32'b11111111111111111011100110011100;
assign LUT_4[38666] = 32'b00000000000000000001110101001000;
assign LUT_4[38667] = 32'b11111111111111111011000001000000;
assign LUT_4[38668] = 32'b11111111111111111111011011000000;
assign LUT_4[38669] = 32'b11111111111111111000100110111000;
assign LUT_4[38670] = 32'b11111111111111111110110101100100;
assign LUT_4[38671] = 32'b11111111111111111000000001011100;
assign LUT_4[38672] = 32'b00000000000000000110111111111101;
assign LUT_4[38673] = 32'b00000000000000000000001011110101;
assign LUT_4[38674] = 32'b00000000000000000110011010100001;
assign LUT_4[38675] = 32'b11111111111111111111100110011001;
assign LUT_4[38676] = 32'b00000000000000000100000000011001;
assign LUT_4[38677] = 32'b11111111111111111101001100010001;
assign LUT_4[38678] = 32'b00000000000000000011011010111101;
assign LUT_4[38679] = 32'b11111111111111111100100110110101;
assign LUT_4[38680] = 32'b00000000000000000000001100010010;
assign LUT_4[38681] = 32'b11111111111111111001011000001010;
assign LUT_4[38682] = 32'b11111111111111111111100110110110;
assign LUT_4[38683] = 32'b11111111111111111000110010101110;
assign LUT_4[38684] = 32'b11111111111111111101001100101110;
assign LUT_4[38685] = 32'b11111111111111110110011000100110;
assign LUT_4[38686] = 32'b11111111111111111100100111010010;
assign LUT_4[38687] = 32'b11111111111111110101110011001010;
assign LUT_4[38688] = 32'b00000000000000000111101001010110;
assign LUT_4[38689] = 32'b00000000000000000000110101001110;
assign LUT_4[38690] = 32'b00000000000000000111000011111010;
assign LUT_4[38691] = 32'b00000000000000000000001111110010;
assign LUT_4[38692] = 32'b00000000000000000100101001110010;
assign LUT_4[38693] = 32'b11111111111111111101110101101010;
assign LUT_4[38694] = 32'b00000000000000000100000100010110;
assign LUT_4[38695] = 32'b11111111111111111101010000001110;
assign LUT_4[38696] = 32'b00000000000000000000110101101011;
assign LUT_4[38697] = 32'b11111111111111111010000001100011;
assign LUT_4[38698] = 32'b00000000000000000000010000001111;
assign LUT_4[38699] = 32'b11111111111111111001011100000111;
assign LUT_4[38700] = 32'b11111111111111111101110110000111;
assign LUT_4[38701] = 32'b11111111111111110111000001111111;
assign LUT_4[38702] = 32'b11111111111111111101010000101011;
assign LUT_4[38703] = 32'b11111111111111110110011100100011;
assign LUT_4[38704] = 32'b00000000000000000101011011000100;
assign LUT_4[38705] = 32'b11111111111111111110100110111100;
assign LUT_4[38706] = 32'b00000000000000000100110101101000;
assign LUT_4[38707] = 32'b11111111111111111110000001100000;
assign LUT_4[38708] = 32'b00000000000000000010011011100000;
assign LUT_4[38709] = 32'b11111111111111111011100111011000;
assign LUT_4[38710] = 32'b00000000000000000001110110000100;
assign LUT_4[38711] = 32'b11111111111111111011000001111100;
assign LUT_4[38712] = 32'b11111111111111111110100111011001;
assign LUT_4[38713] = 32'b11111111111111110111110011010001;
assign LUT_4[38714] = 32'b11111111111111111110000001111101;
assign LUT_4[38715] = 32'b11111111111111110111001101110101;
assign LUT_4[38716] = 32'b11111111111111111011100111110101;
assign LUT_4[38717] = 32'b11111111111111110100110011101101;
assign LUT_4[38718] = 32'b11111111111111111011000010011001;
assign LUT_4[38719] = 32'b11111111111111110100001110010001;
assign LUT_4[38720] = 32'b00000000000000001010100101100011;
assign LUT_4[38721] = 32'b00000000000000000011110001011011;
assign LUT_4[38722] = 32'b00000000000000001010000000000111;
assign LUT_4[38723] = 32'b00000000000000000011001011111111;
assign LUT_4[38724] = 32'b00000000000000000111100101111111;
assign LUT_4[38725] = 32'b00000000000000000000110001110111;
assign LUT_4[38726] = 32'b00000000000000000111000000100011;
assign LUT_4[38727] = 32'b00000000000000000000001100011011;
assign LUT_4[38728] = 32'b00000000000000000011110001111000;
assign LUT_4[38729] = 32'b11111111111111111100111101110000;
assign LUT_4[38730] = 32'b00000000000000000011001100011100;
assign LUT_4[38731] = 32'b11111111111111111100011000010100;
assign LUT_4[38732] = 32'b00000000000000000000110010010100;
assign LUT_4[38733] = 32'b11111111111111111001111110001100;
assign LUT_4[38734] = 32'b00000000000000000000001100111000;
assign LUT_4[38735] = 32'b11111111111111111001011000110000;
assign LUT_4[38736] = 32'b00000000000000001000010111010001;
assign LUT_4[38737] = 32'b00000000000000000001100011001001;
assign LUT_4[38738] = 32'b00000000000000000111110001110101;
assign LUT_4[38739] = 32'b00000000000000000000111101101101;
assign LUT_4[38740] = 32'b00000000000000000101010111101101;
assign LUT_4[38741] = 32'b11111111111111111110100011100101;
assign LUT_4[38742] = 32'b00000000000000000100110010010001;
assign LUT_4[38743] = 32'b11111111111111111101111110001001;
assign LUT_4[38744] = 32'b00000000000000000001100011100110;
assign LUT_4[38745] = 32'b11111111111111111010101111011110;
assign LUT_4[38746] = 32'b00000000000000000000111110001010;
assign LUT_4[38747] = 32'b11111111111111111010001010000010;
assign LUT_4[38748] = 32'b11111111111111111110100100000010;
assign LUT_4[38749] = 32'b11111111111111110111101111111010;
assign LUT_4[38750] = 32'b11111111111111111101111110100110;
assign LUT_4[38751] = 32'b11111111111111110111001010011110;
assign LUT_4[38752] = 32'b00000000000000001001000000101010;
assign LUT_4[38753] = 32'b00000000000000000010001100100010;
assign LUT_4[38754] = 32'b00000000000000001000011011001110;
assign LUT_4[38755] = 32'b00000000000000000001100111000110;
assign LUT_4[38756] = 32'b00000000000000000110000001000110;
assign LUT_4[38757] = 32'b11111111111111111111001100111110;
assign LUT_4[38758] = 32'b00000000000000000101011011101010;
assign LUT_4[38759] = 32'b11111111111111111110100111100010;
assign LUT_4[38760] = 32'b00000000000000000010001100111111;
assign LUT_4[38761] = 32'b11111111111111111011011000110111;
assign LUT_4[38762] = 32'b00000000000000000001100111100011;
assign LUT_4[38763] = 32'b11111111111111111010110011011011;
assign LUT_4[38764] = 32'b11111111111111111111001101011011;
assign LUT_4[38765] = 32'b11111111111111111000011001010011;
assign LUT_4[38766] = 32'b11111111111111111110100111111111;
assign LUT_4[38767] = 32'b11111111111111110111110011110111;
assign LUT_4[38768] = 32'b00000000000000000110110010011000;
assign LUT_4[38769] = 32'b11111111111111111111111110010000;
assign LUT_4[38770] = 32'b00000000000000000110001100111100;
assign LUT_4[38771] = 32'b11111111111111111111011000110100;
assign LUT_4[38772] = 32'b00000000000000000011110010110100;
assign LUT_4[38773] = 32'b11111111111111111100111110101100;
assign LUT_4[38774] = 32'b00000000000000000011001101011000;
assign LUT_4[38775] = 32'b11111111111111111100011001010000;
assign LUT_4[38776] = 32'b11111111111111111111111110101101;
assign LUT_4[38777] = 32'b11111111111111111001001010100101;
assign LUT_4[38778] = 32'b11111111111111111111011001010001;
assign LUT_4[38779] = 32'b11111111111111111000100101001001;
assign LUT_4[38780] = 32'b11111111111111111100111111001001;
assign LUT_4[38781] = 32'b11111111111111110110001011000001;
assign LUT_4[38782] = 32'b11111111111111111100011001101101;
assign LUT_4[38783] = 32'b11111111111111110101100101100101;
assign LUT_4[38784] = 32'b00000000000000001011110100010111;
assign LUT_4[38785] = 32'b00000000000000000101000000001111;
assign LUT_4[38786] = 32'b00000000000000001011001110111011;
assign LUT_4[38787] = 32'b00000000000000000100011010110011;
assign LUT_4[38788] = 32'b00000000000000001000110100110011;
assign LUT_4[38789] = 32'b00000000000000000010000000101011;
assign LUT_4[38790] = 32'b00000000000000001000001111010111;
assign LUT_4[38791] = 32'b00000000000000000001011011001111;
assign LUT_4[38792] = 32'b00000000000000000101000000101100;
assign LUT_4[38793] = 32'b11111111111111111110001100100100;
assign LUT_4[38794] = 32'b00000000000000000100011011010000;
assign LUT_4[38795] = 32'b11111111111111111101100111001000;
assign LUT_4[38796] = 32'b00000000000000000010000001001000;
assign LUT_4[38797] = 32'b11111111111111111011001101000000;
assign LUT_4[38798] = 32'b00000000000000000001011011101100;
assign LUT_4[38799] = 32'b11111111111111111010100111100100;
assign LUT_4[38800] = 32'b00000000000000001001100110000101;
assign LUT_4[38801] = 32'b00000000000000000010110001111101;
assign LUT_4[38802] = 32'b00000000000000001001000000101001;
assign LUT_4[38803] = 32'b00000000000000000010001100100001;
assign LUT_4[38804] = 32'b00000000000000000110100110100001;
assign LUT_4[38805] = 32'b11111111111111111111110010011001;
assign LUT_4[38806] = 32'b00000000000000000110000001000101;
assign LUT_4[38807] = 32'b11111111111111111111001100111101;
assign LUT_4[38808] = 32'b00000000000000000010110010011010;
assign LUT_4[38809] = 32'b11111111111111111011111110010010;
assign LUT_4[38810] = 32'b00000000000000000010001100111110;
assign LUT_4[38811] = 32'b11111111111111111011011000110110;
assign LUT_4[38812] = 32'b11111111111111111111110010110110;
assign LUT_4[38813] = 32'b11111111111111111000111110101110;
assign LUT_4[38814] = 32'b11111111111111111111001101011010;
assign LUT_4[38815] = 32'b11111111111111111000011001010010;
assign LUT_4[38816] = 32'b00000000000000001010001111011110;
assign LUT_4[38817] = 32'b00000000000000000011011011010110;
assign LUT_4[38818] = 32'b00000000000000001001101010000010;
assign LUT_4[38819] = 32'b00000000000000000010110101111010;
assign LUT_4[38820] = 32'b00000000000000000111001111111010;
assign LUT_4[38821] = 32'b00000000000000000000011011110010;
assign LUT_4[38822] = 32'b00000000000000000110101010011110;
assign LUT_4[38823] = 32'b11111111111111111111110110010110;
assign LUT_4[38824] = 32'b00000000000000000011011011110011;
assign LUT_4[38825] = 32'b11111111111111111100100111101011;
assign LUT_4[38826] = 32'b00000000000000000010110110010111;
assign LUT_4[38827] = 32'b11111111111111111100000010001111;
assign LUT_4[38828] = 32'b00000000000000000000011100001111;
assign LUT_4[38829] = 32'b11111111111111111001101000000111;
assign LUT_4[38830] = 32'b11111111111111111111110110110011;
assign LUT_4[38831] = 32'b11111111111111111001000010101011;
assign LUT_4[38832] = 32'b00000000000000001000000001001100;
assign LUT_4[38833] = 32'b00000000000000000001001101000100;
assign LUT_4[38834] = 32'b00000000000000000111011011110000;
assign LUT_4[38835] = 32'b00000000000000000000100111101000;
assign LUT_4[38836] = 32'b00000000000000000101000001101000;
assign LUT_4[38837] = 32'b11111111111111111110001101100000;
assign LUT_4[38838] = 32'b00000000000000000100011100001100;
assign LUT_4[38839] = 32'b11111111111111111101101000000100;
assign LUT_4[38840] = 32'b00000000000000000001001101100001;
assign LUT_4[38841] = 32'b11111111111111111010011001011001;
assign LUT_4[38842] = 32'b00000000000000000000101000000101;
assign LUT_4[38843] = 32'b11111111111111111001110011111101;
assign LUT_4[38844] = 32'b11111111111111111110001101111101;
assign LUT_4[38845] = 32'b11111111111111110111011001110101;
assign LUT_4[38846] = 32'b11111111111111111101101000100001;
assign LUT_4[38847] = 32'b11111111111111110110110100011001;
assign LUT_4[38848] = 32'b00000000000000001101001011101011;
assign LUT_4[38849] = 32'b00000000000000000110010111100011;
assign LUT_4[38850] = 32'b00000000000000001100100110001111;
assign LUT_4[38851] = 32'b00000000000000000101110010000111;
assign LUT_4[38852] = 32'b00000000000000001010001100000111;
assign LUT_4[38853] = 32'b00000000000000000011010111111111;
assign LUT_4[38854] = 32'b00000000000000001001100110101011;
assign LUT_4[38855] = 32'b00000000000000000010110010100011;
assign LUT_4[38856] = 32'b00000000000000000110011000000000;
assign LUT_4[38857] = 32'b11111111111111111111100011111000;
assign LUT_4[38858] = 32'b00000000000000000101110010100100;
assign LUT_4[38859] = 32'b11111111111111111110111110011100;
assign LUT_4[38860] = 32'b00000000000000000011011000011100;
assign LUT_4[38861] = 32'b11111111111111111100100100010100;
assign LUT_4[38862] = 32'b00000000000000000010110011000000;
assign LUT_4[38863] = 32'b11111111111111111011111110111000;
assign LUT_4[38864] = 32'b00000000000000001010111101011001;
assign LUT_4[38865] = 32'b00000000000000000100001001010001;
assign LUT_4[38866] = 32'b00000000000000001010010111111101;
assign LUT_4[38867] = 32'b00000000000000000011100011110101;
assign LUT_4[38868] = 32'b00000000000000000111111101110101;
assign LUT_4[38869] = 32'b00000000000000000001001001101101;
assign LUT_4[38870] = 32'b00000000000000000111011000011001;
assign LUT_4[38871] = 32'b00000000000000000000100100010001;
assign LUT_4[38872] = 32'b00000000000000000100001001101110;
assign LUT_4[38873] = 32'b11111111111111111101010101100110;
assign LUT_4[38874] = 32'b00000000000000000011100100010010;
assign LUT_4[38875] = 32'b11111111111111111100110000001010;
assign LUT_4[38876] = 32'b00000000000000000001001010001010;
assign LUT_4[38877] = 32'b11111111111111111010010110000010;
assign LUT_4[38878] = 32'b00000000000000000000100100101110;
assign LUT_4[38879] = 32'b11111111111111111001110000100110;
assign LUT_4[38880] = 32'b00000000000000001011100110110010;
assign LUT_4[38881] = 32'b00000000000000000100110010101010;
assign LUT_4[38882] = 32'b00000000000000001011000001010110;
assign LUT_4[38883] = 32'b00000000000000000100001101001110;
assign LUT_4[38884] = 32'b00000000000000001000100111001110;
assign LUT_4[38885] = 32'b00000000000000000001110011000110;
assign LUT_4[38886] = 32'b00000000000000001000000001110010;
assign LUT_4[38887] = 32'b00000000000000000001001101101010;
assign LUT_4[38888] = 32'b00000000000000000100110011000111;
assign LUT_4[38889] = 32'b11111111111111111101111110111111;
assign LUT_4[38890] = 32'b00000000000000000100001101101011;
assign LUT_4[38891] = 32'b11111111111111111101011001100011;
assign LUT_4[38892] = 32'b00000000000000000001110011100011;
assign LUT_4[38893] = 32'b11111111111111111010111111011011;
assign LUT_4[38894] = 32'b00000000000000000001001110000111;
assign LUT_4[38895] = 32'b11111111111111111010011001111111;
assign LUT_4[38896] = 32'b00000000000000001001011000100000;
assign LUT_4[38897] = 32'b00000000000000000010100100011000;
assign LUT_4[38898] = 32'b00000000000000001000110011000100;
assign LUT_4[38899] = 32'b00000000000000000001111110111100;
assign LUT_4[38900] = 32'b00000000000000000110011000111100;
assign LUT_4[38901] = 32'b11111111111111111111100100110100;
assign LUT_4[38902] = 32'b00000000000000000101110011100000;
assign LUT_4[38903] = 32'b11111111111111111110111111011000;
assign LUT_4[38904] = 32'b00000000000000000010100100110101;
assign LUT_4[38905] = 32'b11111111111111111011110000101101;
assign LUT_4[38906] = 32'b00000000000000000001111111011001;
assign LUT_4[38907] = 32'b11111111111111111011001011010001;
assign LUT_4[38908] = 32'b11111111111111111111100101010001;
assign LUT_4[38909] = 32'b11111111111111111000110001001001;
assign LUT_4[38910] = 32'b11111111111111111110111111110101;
assign LUT_4[38911] = 32'b11111111111111111000001011101101;
assign LUT_4[38912] = 32'b11111111111111111111000011001111;
assign LUT_4[38913] = 32'b11111111111111111000001111000111;
assign LUT_4[38914] = 32'b11111111111111111110011101110011;
assign LUT_4[38915] = 32'b11111111111111110111101001101011;
assign LUT_4[38916] = 32'b11111111111111111100000011101011;
assign LUT_4[38917] = 32'b11111111111111110101001111100011;
assign LUT_4[38918] = 32'b11111111111111111011011110001111;
assign LUT_4[38919] = 32'b11111111111111110100101010000111;
assign LUT_4[38920] = 32'b11111111111111111000001111100100;
assign LUT_4[38921] = 32'b11111111111111110001011011011100;
assign LUT_4[38922] = 32'b11111111111111110111101010001000;
assign LUT_4[38923] = 32'b11111111111111110000110110000000;
assign LUT_4[38924] = 32'b11111111111111110101010000000000;
assign LUT_4[38925] = 32'b11111111111111101110011011111000;
assign LUT_4[38926] = 32'b11111111111111110100101010100100;
assign LUT_4[38927] = 32'b11111111111111101101110110011100;
assign LUT_4[38928] = 32'b11111111111111111100110100111101;
assign LUT_4[38929] = 32'b11111111111111110110000000110101;
assign LUT_4[38930] = 32'b11111111111111111100001111100001;
assign LUT_4[38931] = 32'b11111111111111110101011011011001;
assign LUT_4[38932] = 32'b11111111111111111001110101011001;
assign LUT_4[38933] = 32'b11111111111111110011000001010001;
assign LUT_4[38934] = 32'b11111111111111111001001111111101;
assign LUT_4[38935] = 32'b11111111111111110010011011110101;
assign LUT_4[38936] = 32'b11111111111111110110000001010010;
assign LUT_4[38937] = 32'b11111111111111101111001101001010;
assign LUT_4[38938] = 32'b11111111111111110101011011110110;
assign LUT_4[38939] = 32'b11111111111111101110100111101110;
assign LUT_4[38940] = 32'b11111111111111110011000001101110;
assign LUT_4[38941] = 32'b11111111111111101100001101100110;
assign LUT_4[38942] = 32'b11111111111111110010011100010010;
assign LUT_4[38943] = 32'b11111111111111101011101000001010;
assign LUT_4[38944] = 32'b11111111111111111101011110010110;
assign LUT_4[38945] = 32'b11111111111111110110101010001110;
assign LUT_4[38946] = 32'b11111111111111111100111000111010;
assign LUT_4[38947] = 32'b11111111111111110110000100110010;
assign LUT_4[38948] = 32'b11111111111111111010011110110010;
assign LUT_4[38949] = 32'b11111111111111110011101010101010;
assign LUT_4[38950] = 32'b11111111111111111001111001010110;
assign LUT_4[38951] = 32'b11111111111111110011000101001110;
assign LUT_4[38952] = 32'b11111111111111110110101010101011;
assign LUT_4[38953] = 32'b11111111111111101111110110100011;
assign LUT_4[38954] = 32'b11111111111111110110000101001111;
assign LUT_4[38955] = 32'b11111111111111101111010001000111;
assign LUT_4[38956] = 32'b11111111111111110011101011000111;
assign LUT_4[38957] = 32'b11111111111111101100110110111111;
assign LUT_4[38958] = 32'b11111111111111110011000101101011;
assign LUT_4[38959] = 32'b11111111111111101100010001100011;
assign LUT_4[38960] = 32'b11111111111111111011010000000100;
assign LUT_4[38961] = 32'b11111111111111110100011011111100;
assign LUT_4[38962] = 32'b11111111111111111010101010101000;
assign LUT_4[38963] = 32'b11111111111111110011110110100000;
assign LUT_4[38964] = 32'b11111111111111111000010000100000;
assign LUT_4[38965] = 32'b11111111111111110001011100011000;
assign LUT_4[38966] = 32'b11111111111111110111101011000100;
assign LUT_4[38967] = 32'b11111111111111110000110110111100;
assign LUT_4[38968] = 32'b11111111111111110100011100011001;
assign LUT_4[38969] = 32'b11111111111111101101101000010001;
assign LUT_4[38970] = 32'b11111111111111110011110110111101;
assign LUT_4[38971] = 32'b11111111111111101101000010110101;
assign LUT_4[38972] = 32'b11111111111111110001011100110101;
assign LUT_4[38973] = 32'b11111111111111101010101000101101;
assign LUT_4[38974] = 32'b11111111111111110000110111011001;
assign LUT_4[38975] = 32'b11111111111111101010000011010001;
assign LUT_4[38976] = 32'b00000000000000000000011010100011;
assign LUT_4[38977] = 32'b11111111111111111001100110011011;
assign LUT_4[38978] = 32'b11111111111111111111110101000111;
assign LUT_4[38979] = 32'b11111111111111111001000000111111;
assign LUT_4[38980] = 32'b11111111111111111101011010111111;
assign LUT_4[38981] = 32'b11111111111111110110100110110111;
assign LUT_4[38982] = 32'b11111111111111111100110101100011;
assign LUT_4[38983] = 32'b11111111111111110110000001011011;
assign LUT_4[38984] = 32'b11111111111111111001100110111000;
assign LUT_4[38985] = 32'b11111111111111110010110010110000;
assign LUT_4[38986] = 32'b11111111111111111001000001011100;
assign LUT_4[38987] = 32'b11111111111111110010001101010100;
assign LUT_4[38988] = 32'b11111111111111110110100111010100;
assign LUT_4[38989] = 32'b11111111111111101111110011001100;
assign LUT_4[38990] = 32'b11111111111111110110000001111000;
assign LUT_4[38991] = 32'b11111111111111101111001101110000;
assign LUT_4[38992] = 32'b11111111111111111110001100010001;
assign LUT_4[38993] = 32'b11111111111111110111011000001001;
assign LUT_4[38994] = 32'b11111111111111111101100110110101;
assign LUT_4[38995] = 32'b11111111111111110110110010101101;
assign LUT_4[38996] = 32'b11111111111111111011001100101101;
assign LUT_4[38997] = 32'b11111111111111110100011000100101;
assign LUT_4[38998] = 32'b11111111111111111010100111010001;
assign LUT_4[38999] = 32'b11111111111111110011110011001001;
assign LUT_4[39000] = 32'b11111111111111110111011000100110;
assign LUT_4[39001] = 32'b11111111111111110000100100011110;
assign LUT_4[39002] = 32'b11111111111111110110110011001010;
assign LUT_4[39003] = 32'b11111111111111101111111111000010;
assign LUT_4[39004] = 32'b11111111111111110100011001000010;
assign LUT_4[39005] = 32'b11111111111111101101100100111010;
assign LUT_4[39006] = 32'b11111111111111110011110011100110;
assign LUT_4[39007] = 32'b11111111111111101100111111011110;
assign LUT_4[39008] = 32'b11111111111111111110110101101010;
assign LUT_4[39009] = 32'b11111111111111111000000001100010;
assign LUT_4[39010] = 32'b11111111111111111110010000001110;
assign LUT_4[39011] = 32'b11111111111111110111011100000110;
assign LUT_4[39012] = 32'b11111111111111111011110110000110;
assign LUT_4[39013] = 32'b11111111111111110101000001111110;
assign LUT_4[39014] = 32'b11111111111111111011010000101010;
assign LUT_4[39015] = 32'b11111111111111110100011100100010;
assign LUT_4[39016] = 32'b11111111111111111000000001111111;
assign LUT_4[39017] = 32'b11111111111111110001001101110111;
assign LUT_4[39018] = 32'b11111111111111110111011100100011;
assign LUT_4[39019] = 32'b11111111111111110000101000011011;
assign LUT_4[39020] = 32'b11111111111111110101000010011011;
assign LUT_4[39021] = 32'b11111111111111101110001110010011;
assign LUT_4[39022] = 32'b11111111111111110100011100111111;
assign LUT_4[39023] = 32'b11111111111111101101101000110111;
assign LUT_4[39024] = 32'b11111111111111111100100111011000;
assign LUT_4[39025] = 32'b11111111111111110101110011010000;
assign LUT_4[39026] = 32'b11111111111111111100000001111100;
assign LUT_4[39027] = 32'b11111111111111110101001101110100;
assign LUT_4[39028] = 32'b11111111111111111001100111110100;
assign LUT_4[39029] = 32'b11111111111111110010110011101100;
assign LUT_4[39030] = 32'b11111111111111111001000010011000;
assign LUT_4[39031] = 32'b11111111111111110010001110010000;
assign LUT_4[39032] = 32'b11111111111111110101110011101101;
assign LUT_4[39033] = 32'b11111111111111101110111111100101;
assign LUT_4[39034] = 32'b11111111111111110101001110010001;
assign LUT_4[39035] = 32'b11111111111111101110011010001001;
assign LUT_4[39036] = 32'b11111111111111110010110100001001;
assign LUT_4[39037] = 32'b11111111111111101100000000000001;
assign LUT_4[39038] = 32'b11111111111111110010001110101101;
assign LUT_4[39039] = 32'b11111111111111101011011010100101;
assign LUT_4[39040] = 32'b00000000000000000001101001010111;
assign LUT_4[39041] = 32'b11111111111111111010110101001111;
assign LUT_4[39042] = 32'b00000000000000000001000011111011;
assign LUT_4[39043] = 32'b11111111111111111010001111110011;
assign LUT_4[39044] = 32'b11111111111111111110101001110011;
assign LUT_4[39045] = 32'b11111111111111110111110101101011;
assign LUT_4[39046] = 32'b11111111111111111110000100010111;
assign LUT_4[39047] = 32'b11111111111111110111010000001111;
assign LUT_4[39048] = 32'b11111111111111111010110101101100;
assign LUT_4[39049] = 32'b11111111111111110100000001100100;
assign LUT_4[39050] = 32'b11111111111111111010010000010000;
assign LUT_4[39051] = 32'b11111111111111110011011100001000;
assign LUT_4[39052] = 32'b11111111111111110111110110001000;
assign LUT_4[39053] = 32'b11111111111111110001000010000000;
assign LUT_4[39054] = 32'b11111111111111110111010000101100;
assign LUT_4[39055] = 32'b11111111111111110000011100100100;
assign LUT_4[39056] = 32'b11111111111111111111011011000101;
assign LUT_4[39057] = 32'b11111111111111111000100110111101;
assign LUT_4[39058] = 32'b11111111111111111110110101101001;
assign LUT_4[39059] = 32'b11111111111111111000000001100001;
assign LUT_4[39060] = 32'b11111111111111111100011011100001;
assign LUT_4[39061] = 32'b11111111111111110101100111011001;
assign LUT_4[39062] = 32'b11111111111111111011110110000101;
assign LUT_4[39063] = 32'b11111111111111110101000001111101;
assign LUT_4[39064] = 32'b11111111111111111000100111011010;
assign LUT_4[39065] = 32'b11111111111111110001110011010010;
assign LUT_4[39066] = 32'b11111111111111111000000001111110;
assign LUT_4[39067] = 32'b11111111111111110001001101110110;
assign LUT_4[39068] = 32'b11111111111111110101100111110110;
assign LUT_4[39069] = 32'b11111111111111101110110011101110;
assign LUT_4[39070] = 32'b11111111111111110101000010011010;
assign LUT_4[39071] = 32'b11111111111111101110001110010010;
assign LUT_4[39072] = 32'b00000000000000000000000100011110;
assign LUT_4[39073] = 32'b11111111111111111001010000010110;
assign LUT_4[39074] = 32'b11111111111111111111011111000010;
assign LUT_4[39075] = 32'b11111111111111111000101010111010;
assign LUT_4[39076] = 32'b11111111111111111101000100111010;
assign LUT_4[39077] = 32'b11111111111111110110010000110010;
assign LUT_4[39078] = 32'b11111111111111111100011111011110;
assign LUT_4[39079] = 32'b11111111111111110101101011010110;
assign LUT_4[39080] = 32'b11111111111111111001010000110011;
assign LUT_4[39081] = 32'b11111111111111110010011100101011;
assign LUT_4[39082] = 32'b11111111111111111000101011010111;
assign LUT_4[39083] = 32'b11111111111111110001110111001111;
assign LUT_4[39084] = 32'b11111111111111110110010001001111;
assign LUT_4[39085] = 32'b11111111111111101111011101000111;
assign LUT_4[39086] = 32'b11111111111111110101101011110011;
assign LUT_4[39087] = 32'b11111111111111101110110111101011;
assign LUT_4[39088] = 32'b11111111111111111101110110001100;
assign LUT_4[39089] = 32'b11111111111111110111000010000100;
assign LUT_4[39090] = 32'b11111111111111111101010000110000;
assign LUT_4[39091] = 32'b11111111111111110110011100101000;
assign LUT_4[39092] = 32'b11111111111111111010110110101000;
assign LUT_4[39093] = 32'b11111111111111110100000010100000;
assign LUT_4[39094] = 32'b11111111111111111010010001001100;
assign LUT_4[39095] = 32'b11111111111111110011011101000100;
assign LUT_4[39096] = 32'b11111111111111110111000010100001;
assign LUT_4[39097] = 32'b11111111111111110000001110011001;
assign LUT_4[39098] = 32'b11111111111111110110011101000101;
assign LUT_4[39099] = 32'b11111111111111101111101000111101;
assign LUT_4[39100] = 32'b11111111111111110100000010111101;
assign LUT_4[39101] = 32'b11111111111111101101001110110101;
assign LUT_4[39102] = 32'b11111111111111110011011101100001;
assign LUT_4[39103] = 32'b11111111111111101100101001011001;
assign LUT_4[39104] = 32'b00000000000000000011000000101011;
assign LUT_4[39105] = 32'b11111111111111111100001100100011;
assign LUT_4[39106] = 32'b00000000000000000010011011001111;
assign LUT_4[39107] = 32'b11111111111111111011100111000111;
assign LUT_4[39108] = 32'b00000000000000000000000001000111;
assign LUT_4[39109] = 32'b11111111111111111001001100111111;
assign LUT_4[39110] = 32'b11111111111111111111011011101011;
assign LUT_4[39111] = 32'b11111111111111111000100111100011;
assign LUT_4[39112] = 32'b11111111111111111100001101000000;
assign LUT_4[39113] = 32'b11111111111111110101011000111000;
assign LUT_4[39114] = 32'b11111111111111111011100111100100;
assign LUT_4[39115] = 32'b11111111111111110100110011011100;
assign LUT_4[39116] = 32'b11111111111111111001001101011100;
assign LUT_4[39117] = 32'b11111111111111110010011001010100;
assign LUT_4[39118] = 32'b11111111111111111000101000000000;
assign LUT_4[39119] = 32'b11111111111111110001110011111000;
assign LUT_4[39120] = 32'b00000000000000000000110010011001;
assign LUT_4[39121] = 32'b11111111111111111001111110010001;
assign LUT_4[39122] = 32'b00000000000000000000001100111101;
assign LUT_4[39123] = 32'b11111111111111111001011000110101;
assign LUT_4[39124] = 32'b11111111111111111101110010110101;
assign LUT_4[39125] = 32'b11111111111111110110111110101101;
assign LUT_4[39126] = 32'b11111111111111111101001101011001;
assign LUT_4[39127] = 32'b11111111111111110110011001010001;
assign LUT_4[39128] = 32'b11111111111111111001111110101110;
assign LUT_4[39129] = 32'b11111111111111110011001010100110;
assign LUT_4[39130] = 32'b11111111111111111001011001010010;
assign LUT_4[39131] = 32'b11111111111111110010100101001010;
assign LUT_4[39132] = 32'b11111111111111110110111111001010;
assign LUT_4[39133] = 32'b11111111111111110000001011000010;
assign LUT_4[39134] = 32'b11111111111111110110011001101110;
assign LUT_4[39135] = 32'b11111111111111101111100101100110;
assign LUT_4[39136] = 32'b00000000000000000001011011110010;
assign LUT_4[39137] = 32'b11111111111111111010100111101010;
assign LUT_4[39138] = 32'b00000000000000000000110110010110;
assign LUT_4[39139] = 32'b11111111111111111010000010001110;
assign LUT_4[39140] = 32'b11111111111111111110011100001110;
assign LUT_4[39141] = 32'b11111111111111110111101000000110;
assign LUT_4[39142] = 32'b11111111111111111101110110110010;
assign LUT_4[39143] = 32'b11111111111111110111000010101010;
assign LUT_4[39144] = 32'b11111111111111111010101000000111;
assign LUT_4[39145] = 32'b11111111111111110011110011111111;
assign LUT_4[39146] = 32'b11111111111111111010000010101011;
assign LUT_4[39147] = 32'b11111111111111110011001110100011;
assign LUT_4[39148] = 32'b11111111111111110111101000100011;
assign LUT_4[39149] = 32'b11111111111111110000110100011011;
assign LUT_4[39150] = 32'b11111111111111110111000011000111;
assign LUT_4[39151] = 32'b11111111111111110000001110111111;
assign LUT_4[39152] = 32'b11111111111111111111001101100000;
assign LUT_4[39153] = 32'b11111111111111111000011001011000;
assign LUT_4[39154] = 32'b11111111111111111110101000000100;
assign LUT_4[39155] = 32'b11111111111111110111110011111100;
assign LUT_4[39156] = 32'b11111111111111111100001101111100;
assign LUT_4[39157] = 32'b11111111111111110101011001110100;
assign LUT_4[39158] = 32'b11111111111111111011101000100000;
assign LUT_4[39159] = 32'b11111111111111110100110100011000;
assign LUT_4[39160] = 32'b11111111111111111000011001110101;
assign LUT_4[39161] = 32'b11111111111111110001100101101101;
assign LUT_4[39162] = 32'b11111111111111110111110100011001;
assign LUT_4[39163] = 32'b11111111111111110001000000010001;
assign LUT_4[39164] = 32'b11111111111111110101011010010001;
assign LUT_4[39165] = 32'b11111111111111101110100110001001;
assign LUT_4[39166] = 32'b11111111111111110100110100110101;
assign LUT_4[39167] = 32'b11111111111111101110000000101101;
assign LUT_4[39168] = 32'b00000000000000000011111110110010;
assign LUT_4[39169] = 32'b11111111111111111101001010101010;
assign LUT_4[39170] = 32'b00000000000000000011011001010110;
assign LUT_4[39171] = 32'b11111111111111111100100101001110;
assign LUT_4[39172] = 32'b00000000000000000000111111001110;
assign LUT_4[39173] = 32'b11111111111111111010001011000110;
assign LUT_4[39174] = 32'b00000000000000000000011001110010;
assign LUT_4[39175] = 32'b11111111111111111001100101101010;
assign LUT_4[39176] = 32'b11111111111111111101001011000111;
assign LUT_4[39177] = 32'b11111111111111110110010110111111;
assign LUT_4[39178] = 32'b11111111111111111100100101101011;
assign LUT_4[39179] = 32'b11111111111111110101110001100011;
assign LUT_4[39180] = 32'b11111111111111111010001011100011;
assign LUT_4[39181] = 32'b11111111111111110011010111011011;
assign LUT_4[39182] = 32'b11111111111111111001100110000111;
assign LUT_4[39183] = 32'b11111111111111110010110001111111;
assign LUT_4[39184] = 32'b00000000000000000001110000100000;
assign LUT_4[39185] = 32'b11111111111111111010111100011000;
assign LUT_4[39186] = 32'b00000000000000000001001011000100;
assign LUT_4[39187] = 32'b11111111111111111010010110111100;
assign LUT_4[39188] = 32'b11111111111111111110110000111100;
assign LUT_4[39189] = 32'b11111111111111110111111100110100;
assign LUT_4[39190] = 32'b11111111111111111110001011100000;
assign LUT_4[39191] = 32'b11111111111111110111010111011000;
assign LUT_4[39192] = 32'b11111111111111111010111100110101;
assign LUT_4[39193] = 32'b11111111111111110100001000101101;
assign LUT_4[39194] = 32'b11111111111111111010010111011001;
assign LUT_4[39195] = 32'b11111111111111110011100011010001;
assign LUT_4[39196] = 32'b11111111111111110111111101010001;
assign LUT_4[39197] = 32'b11111111111111110001001001001001;
assign LUT_4[39198] = 32'b11111111111111110111010111110101;
assign LUT_4[39199] = 32'b11111111111111110000100011101101;
assign LUT_4[39200] = 32'b00000000000000000010011001111001;
assign LUT_4[39201] = 32'b11111111111111111011100101110001;
assign LUT_4[39202] = 32'b00000000000000000001110100011101;
assign LUT_4[39203] = 32'b11111111111111111011000000010101;
assign LUT_4[39204] = 32'b11111111111111111111011010010101;
assign LUT_4[39205] = 32'b11111111111111111000100110001101;
assign LUT_4[39206] = 32'b11111111111111111110110100111001;
assign LUT_4[39207] = 32'b11111111111111111000000000110001;
assign LUT_4[39208] = 32'b11111111111111111011100110001110;
assign LUT_4[39209] = 32'b11111111111111110100110010000110;
assign LUT_4[39210] = 32'b11111111111111111011000000110010;
assign LUT_4[39211] = 32'b11111111111111110100001100101010;
assign LUT_4[39212] = 32'b11111111111111111000100110101010;
assign LUT_4[39213] = 32'b11111111111111110001110010100010;
assign LUT_4[39214] = 32'b11111111111111111000000001001110;
assign LUT_4[39215] = 32'b11111111111111110001001101000110;
assign LUT_4[39216] = 32'b00000000000000000000001011100111;
assign LUT_4[39217] = 32'b11111111111111111001010111011111;
assign LUT_4[39218] = 32'b11111111111111111111100110001011;
assign LUT_4[39219] = 32'b11111111111111111000110010000011;
assign LUT_4[39220] = 32'b11111111111111111101001100000011;
assign LUT_4[39221] = 32'b11111111111111110110010111111011;
assign LUT_4[39222] = 32'b11111111111111111100100110100111;
assign LUT_4[39223] = 32'b11111111111111110101110010011111;
assign LUT_4[39224] = 32'b11111111111111111001010111111100;
assign LUT_4[39225] = 32'b11111111111111110010100011110100;
assign LUT_4[39226] = 32'b11111111111111111000110010100000;
assign LUT_4[39227] = 32'b11111111111111110001111110011000;
assign LUT_4[39228] = 32'b11111111111111110110011000011000;
assign LUT_4[39229] = 32'b11111111111111101111100100010000;
assign LUT_4[39230] = 32'b11111111111111110101110010111100;
assign LUT_4[39231] = 32'b11111111111111101110111110110100;
assign LUT_4[39232] = 32'b00000000000000000101010110000110;
assign LUT_4[39233] = 32'b11111111111111111110100001111110;
assign LUT_4[39234] = 32'b00000000000000000100110000101010;
assign LUT_4[39235] = 32'b11111111111111111101111100100010;
assign LUT_4[39236] = 32'b00000000000000000010010110100010;
assign LUT_4[39237] = 32'b11111111111111111011100010011010;
assign LUT_4[39238] = 32'b00000000000000000001110001000110;
assign LUT_4[39239] = 32'b11111111111111111010111100111110;
assign LUT_4[39240] = 32'b11111111111111111110100010011011;
assign LUT_4[39241] = 32'b11111111111111110111101110010011;
assign LUT_4[39242] = 32'b11111111111111111101111100111111;
assign LUT_4[39243] = 32'b11111111111111110111001000110111;
assign LUT_4[39244] = 32'b11111111111111111011100010110111;
assign LUT_4[39245] = 32'b11111111111111110100101110101111;
assign LUT_4[39246] = 32'b11111111111111111010111101011011;
assign LUT_4[39247] = 32'b11111111111111110100001001010011;
assign LUT_4[39248] = 32'b00000000000000000011000111110100;
assign LUT_4[39249] = 32'b11111111111111111100010011101100;
assign LUT_4[39250] = 32'b00000000000000000010100010011000;
assign LUT_4[39251] = 32'b11111111111111111011101110010000;
assign LUT_4[39252] = 32'b00000000000000000000001000010000;
assign LUT_4[39253] = 32'b11111111111111111001010100001000;
assign LUT_4[39254] = 32'b11111111111111111111100010110100;
assign LUT_4[39255] = 32'b11111111111111111000101110101100;
assign LUT_4[39256] = 32'b11111111111111111100010100001001;
assign LUT_4[39257] = 32'b11111111111111110101100000000001;
assign LUT_4[39258] = 32'b11111111111111111011101110101101;
assign LUT_4[39259] = 32'b11111111111111110100111010100101;
assign LUT_4[39260] = 32'b11111111111111111001010100100101;
assign LUT_4[39261] = 32'b11111111111111110010100000011101;
assign LUT_4[39262] = 32'b11111111111111111000101111001001;
assign LUT_4[39263] = 32'b11111111111111110001111011000001;
assign LUT_4[39264] = 32'b00000000000000000011110001001101;
assign LUT_4[39265] = 32'b11111111111111111100111101000101;
assign LUT_4[39266] = 32'b00000000000000000011001011110001;
assign LUT_4[39267] = 32'b11111111111111111100010111101001;
assign LUT_4[39268] = 32'b00000000000000000000110001101001;
assign LUT_4[39269] = 32'b11111111111111111001111101100001;
assign LUT_4[39270] = 32'b00000000000000000000001100001101;
assign LUT_4[39271] = 32'b11111111111111111001011000000101;
assign LUT_4[39272] = 32'b11111111111111111100111101100010;
assign LUT_4[39273] = 32'b11111111111111110110001001011010;
assign LUT_4[39274] = 32'b11111111111111111100011000000110;
assign LUT_4[39275] = 32'b11111111111111110101100011111110;
assign LUT_4[39276] = 32'b11111111111111111001111101111110;
assign LUT_4[39277] = 32'b11111111111111110011001001110110;
assign LUT_4[39278] = 32'b11111111111111111001011000100010;
assign LUT_4[39279] = 32'b11111111111111110010100100011010;
assign LUT_4[39280] = 32'b00000000000000000001100010111011;
assign LUT_4[39281] = 32'b11111111111111111010101110110011;
assign LUT_4[39282] = 32'b00000000000000000000111101011111;
assign LUT_4[39283] = 32'b11111111111111111010001001010111;
assign LUT_4[39284] = 32'b11111111111111111110100011010111;
assign LUT_4[39285] = 32'b11111111111111110111101111001111;
assign LUT_4[39286] = 32'b11111111111111111101111101111011;
assign LUT_4[39287] = 32'b11111111111111110111001001110011;
assign LUT_4[39288] = 32'b11111111111111111010101111010000;
assign LUT_4[39289] = 32'b11111111111111110011111011001000;
assign LUT_4[39290] = 32'b11111111111111111010001001110100;
assign LUT_4[39291] = 32'b11111111111111110011010101101100;
assign LUT_4[39292] = 32'b11111111111111110111101111101100;
assign LUT_4[39293] = 32'b11111111111111110000111011100100;
assign LUT_4[39294] = 32'b11111111111111110111001010010000;
assign LUT_4[39295] = 32'b11111111111111110000010110001000;
assign LUT_4[39296] = 32'b00000000000000000110100100111010;
assign LUT_4[39297] = 32'b11111111111111111111110000110010;
assign LUT_4[39298] = 32'b00000000000000000101111111011110;
assign LUT_4[39299] = 32'b11111111111111111111001011010110;
assign LUT_4[39300] = 32'b00000000000000000011100101010110;
assign LUT_4[39301] = 32'b11111111111111111100110001001110;
assign LUT_4[39302] = 32'b00000000000000000010111111111010;
assign LUT_4[39303] = 32'b11111111111111111100001011110010;
assign LUT_4[39304] = 32'b11111111111111111111110001001111;
assign LUT_4[39305] = 32'b11111111111111111000111101000111;
assign LUT_4[39306] = 32'b11111111111111111111001011110011;
assign LUT_4[39307] = 32'b11111111111111111000010111101011;
assign LUT_4[39308] = 32'b11111111111111111100110001101011;
assign LUT_4[39309] = 32'b11111111111111110101111101100011;
assign LUT_4[39310] = 32'b11111111111111111100001100001111;
assign LUT_4[39311] = 32'b11111111111111110101011000000111;
assign LUT_4[39312] = 32'b00000000000000000100010110101000;
assign LUT_4[39313] = 32'b11111111111111111101100010100000;
assign LUT_4[39314] = 32'b00000000000000000011110001001100;
assign LUT_4[39315] = 32'b11111111111111111100111101000100;
assign LUT_4[39316] = 32'b00000000000000000001010111000100;
assign LUT_4[39317] = 32'b11111111111111111010100010111100;
assign LUT_4[39318] = 32'b00000000000000000000110001101000;
assign LUT_4[39319] = 32'b11111111111111111001111101100000;
assign LUT_4[39320] = 32'b11111111111111111101100010111101;
assign LUT_4[39321] = 32'b11111111111111110110101110110101;
assign LUT_4[39322] = 32'b11111111111111111100111101100001;
assign LUT_4[39323] = 32'b11111111111111110110001001011001;
assign LUT_4[39324] = 32'b11111111111111111010100011011001;
assign LUT_4[39325] = 32'b11111111111111110011101111010001;
assign LUT_4[39326] = 32'b11111111111111111001111101111101;
assign LUT_4[39327] = 32'b11111111111111110011001001110101;
assign LUT_4[39328] = 32'b00000000000000000101000000000001;
assign LUT_4[39329] = 32'b11111111111111111110001011111001;
assign LUT_4[39330] = 32'b00000000000000000100011010100101;
assign LUT_4[39331] = 32'b11111111111111111101100110011101;
assign LUT_4[39332] = 32'b00000000000000000010000000011101;
assign LUT_4[39333] = 32'b11111111111111111011001100010101;
assign LUT_4[39334] = 32'b00000000000000000001011011000001;
assign LUT_4[39335] = 32'b11111111111111111010100110111001;
assign LUT_4[39336] = 32'b11111111111111111110001100010110;
assign LUT_4[39337] = 32'b11111111111111110111011000001110;
assign LUT_4[39338] = 32'b11111111111111111101100110111010;
assign LUT_4[39339] = 32'b11111111111111110110110010110010;
assign LUT_4[39340] = 32'b11111111111111111011001100110010;
assign LUT_4[39341] = 32'b11111111111111110100011000101010;
assign LUT_4[39342] = 32'b11111111111111111010100111010110;
assign LUT_4[39343] = 32'b11111111111111110011110011001110;
assign LUT_4[39344] = 32'b00000000000000000010110001101111;
assign LUT_4[39345] = 32'b11111111111111111011111101100111;
assign LUT_4[39346] = 32'b00000000000000000010001100010011;
assign LUT_4[39347] = 32'b11111111111111111011011000001011;
assign LUT_4[39348] = 32'b11111111111111111111110010001011;
assign LUT_4[39349] = 32'b11111111111111111000111110000011;
assign LUT_4[39350] = 32'b11111111111111111111001100101111;
assign LUT_4[39351] = 32'b11111111111111111000011000100111;
assign LUT_4[39352] = 32'b11111111111111111011111110000100;
assign LUT_4[39353] = 32'b11111111111111110101001001111100;
assign LUT_4[39354] = 32'b11111111111111111011011000101000;
assign LUT_4[39355] = 32'b11111111111111110100100100100000;
assign LUT_4[39356] = 32'b11111111111111111000111110100000;
assign LUT_4[39357] = 32'b11111111111111110010001010011000;
assign LUT_4[39358] = 32'b11111111111111111000011001000100;
assign LUT_4[39359] = 32'b11111111111111110001100100111100;
assign LUT_4[39360] = 32'b00000000000000000111111100001110;
assign LUT_4[39361] = 32'b00000000000000000001001000000110;
assign LUT_4[39362] = 32'b00000000000000000111010110110010;
assign LUT_4[39363] = 32'b00000000000000000000100010101010;
assign LUT_4[39364] = 32'b00000000000000000100111100101010;
assign LUT_4[39365] = 32'b11111111111111111110001000100010;
assign LUT_4[39366] = 32'b00000000000000000100010111001110;
assign LUT_4[39367] = 32'b11111111111111111101100011000110;
assign LUT_4[39368] = 32'b00000000000000000001001000100011;
assign LUT_4[39369] = 32'b11111111111111111010010100011011;
assign LUT_4[39370] = 32'b00000000000000000000100011000111;
assign LUT_4[39371] = 32'b11111111111111111001101110111111;
assign LUT_4[39372] = 32'b11111111111111111110001000111111;
assign LUT_4[39373] = 32'b11111111111111110111010100110111;
assign LUT_4[39374] = 32'b11111111111111111101100011100011;
assign LUT_4[39375] = 32'b11111111111111110110101111011011;
assign LUT_4[39376] = 32'b00000000000000000101101101111100;
assign LUT_4[39377] = 32'b11111111111111111110111001110100;
assign LUT_4[39378] = 32'b00000000000000000101001000100000;
assign LUT_4[39379] = 32'b11111111111111111110010100011000;
assign LUT_4[39380] = 32'b00000000000000000010101110011000;
assign LUT_4[39381] = 32'b11111111111111111011111010010000;
assign LUT_4[39382] = 32'b00000000000000000010001000111100;
assign LUT_4[39383] = 32'b11111111111111111011010100110100;
assign LUT_4[39384] = 32'b11111111111111111110111010010001;
assign LUT_4[39385] = 32'b11111111111111111000000110001001;
assign LUT_4[39386] = 32'b11111111111111111110010100110101;
assign LUT_4[39387] = 32'b11111111111111110111100000101101;
assign LUT_4[39388] = 32'b11111111111111111011111010101101;
assign LUT_4[39389] = 32'b11111111111111110101000110100101;
assign LUT_4[39390] = 32'b11111111111111111011010101010001;
assign LUT_4[39391] = 32'b11111111111111110100100001001001;
assign LUT_4[39392] = 32'b00000000000000000110010111010101;
assign LUT_4[39393] = 32'b11111111111111111111100011001101;
assign LUT_4[39394] = 32'b00000000000000000101110001111001;
assign LUT_4[39395] = 32'b11111111111111111110111101110001;
assign LUT_4[39396] = 32'b00000000000000000011010111110001;
assign LUT_4[39397] = 32'b11111111111111111100100011101001;
assign LUT_4[39398] = 32'b00000000000000000010110010010101;
assign LUT_4[39399] = 32'b11111111111111111011111110001101;
assign LUT_4[39400] = 32'b11111111111111111111100011101010;
assign LUT_4[39401] = 32'b11111111111111111000101111100010;
assign LUT_4[39402] = 32'b11111111111111111110111110001110;
assign LUT_4[39403] = 32'b11111111111111111000001010000110;
assign LUT_4[39404] = 32'b11111111111111111100100100000110;
assign LUT_4[39405] = 32'b11111111111111110101101111111110;
assign LUT_4[39406] = 32'b11111111111111111011111110101010;
assign LUT_4[39407] = 32'b11111111111111110101001010100010;
assign LUT_4[39408] = 32'b00000000000000000100001001000011;
assign LUT_4[39409] = 32'b11111111111111111101010100111011;
assign LUT_4[39410] = 32'b00000000000000000011100011100111;
assign LUT_4[39411] = 32'b11111111111111111100101111011111;
assign LUT_4[39412] = 32'b00000000000000000001001001011111;
assign LUT_4[39413] = 32'b11111111111111111010010101010111;
assign LUT_4[39414] = 32'b00000000000000000000100100000011;
assign LUT_4[39415] = 32'b11111111111111111001101111111011;
assign LUT_4[39416] = 32'b11111111111111111101010101011000;
assign LUT_4[39417] = 32'b11111111111111110110100001010000;
assign LUT_4[39418] = 32'b11111111111111111100101111111100;
assign LUT_4[39419] = 32'b11111111111111110101111011110100;
assign LUT_4[39420] = 32'b11111111111111111010010101110100;
assign LUT_4[39421] = 32'b11111111111111110011100001101100;
assign LUT_4[39422] = 32'b11111111111111111001110000011000;
assign LUT_4[39423] = 32'b11111111111111110010111100010000;
assign LUT_4[39424] = 32'b11111111111111111110000111010111;
assign LUT_4[39425] = 32'b11111111111111110111010011001111;
assign LUT_4[39426] = 32'b11111111111111111101100001111011;
assign LUT_4[39427] = 32'b11111111111111110110101101110011;
assign LUT_4[39428] = 32'b11111111111111111011000111110011;
assign LUT_4[39429] = 32'b11111111111111110100010011101011;
assign LUT_4[39430] = 32'b11111111111111111010100010010111;
assign LUT_4[39431] = 32'b11111111111111110011101110001111;
assign LUT_4[39432] = 32'b11111111111111110111010011101100;
assign LUT_4[39433] = 32'b11111111111111110000011111100100;
assign LUT_4[39434] = 32'b11111111111111110110101110010000;
assign LUT_4[39435] = 32'b11111111111111101111111010001000;
assign LUT_4[39436] = 32'b11111111111111110100010100001000;
assign LUT_4[39437] = 32'b11111111111111101101100000000000;
assign LUT_4[39438] = 32'b11111111111111110011101110101100;
assign LUT_4[39439] = 32'b11111111111111101100111010100100;
assign LUT_4[39440] = 32'b11111111111111111011111001000101;
assign LUT_4[39441] = 32'b11111111111111110101000100111101;
assign LUT_4[39442] = 32'b11111111111111111011010011101001;
assign LUT_4[39443] = 32'b11111111111111110100011111100001;
assign LUT_4[39444] = 32'b11111111111111111000111001100001;
assign LUT_4[39445] = 32'b11111111111111110010000101011001;
assign LUT_4[39446] = 32'b11111111111111111000010100000101;
assign LUT_4[39447] = 32'b11111111111111110001011111111101;
assign LUT_4[39448] = 32'b11111111111111110101000101011010;
assign LUT_4[39449] = 32'b11111111111111101110010001010010;
assign LUT_4[39450] = 32'b11111111111111110100011111111110;
assign LUT_4[39451] = 32'b11111111111111101101101011110110;
assign LUT_4[39452] = 32'b11111111111111110010000101110110;
assign LUT_4[39453] = 32'b11111111111111101011010001101110;
assign LUT_4[39454] = 32'b11111111111111110001100000011010;
assign LUT_4[39455] = 32'b11111111111111101010101100010010;
assign LUT_4[39456] = 32'b11111111111111111100100010011110;
assign LUT_4[39457] = 32'b11111111111111110101101110010110;
assign LUT_4[39458] = 32'b11111111111111111011111101000010;
assign LUT_4[39459] = 32'b11111111111111110101001000111010;
assign LUT_4[39460] = 32'b11111111111111111001100010111010;
assign LUT_4[39461] = 32'b11111111111111110010101110110010;
assign LUT_4[39462] = 32'b11111111111111111000111101011110;
assign LUT_4[39463] = 32'b11111111111111110010001001010110;
assign LUT_4[39464] = 32'b11111111111111110101101110110011;
assign LUT_4[39465] = 32'b11111111111111101110111010101011;
assign LUT_4[39466] = 32'b11111111111111110101001001010111;
assign LUT_4[39467] = 32'b11111111111111101110010101001111;
assign LUT_4[39468] = 32'b11111111111111110010101111001111;
assign LUT_4[39469] = 32'b11111111111111101011111011000111;
assign LUT_4[39470] = 32'b11111111111111110010001001110011;
assign LUT_4[39471] = 32'b11111111111111101011010101101011;
assign LUT_4[39472] = 32'b11111111111111111010010100001100;
assign LUT_4[39473] = 32'b11111111111111110011100000000100;
assign LUT_4[39474] = 32'b11111111111111111001101110110000;
assign LUT_4[39475] = 32'b11111111111111110010111010101000;
assign LUT_4[39476] = 32'b11111111111111110111010100101000;
assign LUT_4[39477] = 32'b11111111111111110000100000100000;
assign LUT_4[39478] = 32'b11111111111111110110101111001100;
assign LUT_4[39479] = 32'b11111111111111101111111011000100;
assign LUT_4[39480] = 32'b11111111111111110011100000100001;
assign LUT_4[39481] = 32'b11111111111111101100101100011001;
assign LUT_4[39482] = 32'b11111111111111110010111011000101;
assign LUT_4[39483] = 32'b11111111111111101100000110111101;
assign LUT_4[39484] = 32'b11111111111111110000100000111101;
assign LUT_4[39485] = 32'b11111111111111101001101100110101;
assign LUT_4[39486] = 32'b11111111111111101111111011100001;
assign LUT_4[39487] = 32'b11111111111111101001000111011001;
assign LUT_4[39488] = 32'b11111111111111111111011110101011;
assign LUT_4[39489] = 32'b11111111111111111000101010100011;
assign LUT_4[39490] = 32'b11111111111111111110111001001111;
assign LUT_4[39491] = 32'b11111111111111111000000101000111;
assign LUT_4[39492] = 32'b11111111111111111100011111000111;
assign LUT_4[39493] = 32'b11111111111111110101101010111111;
assign LUT_4[39494] = 32'b11111111111111111011111001101011;
assign LUT_4[39495] = 32'b11111111111111110101000101100011;
assign LUT_4[39496] = 32'b11111111111111111000101011000000;
assign LUT_4[39497] = 32'b11111111111111110001110110111000;
assign LUT_4[39498] = 32'b11111111111111111000000101100100;
assign LUT_4[39499] = 32'b11111111111111110001010001011100;
assign LUT_4[39500] = 32'b11111111111111110101101011011100;
assign LUT_4[39501] = 32'b11111111111111101110110111010100;
assign LUT_4[39502] = 32'b11111111111111110101000110000000;
assign LUT_4[39503] = 32'b11111111111111101110010001111000;
assign LUT_4[39504] = 32'b11111111111111111101010000011001;
assign LUT_4[39505] = 32'b11111111111111110110011100010001;
assign LUT_4[39506] = 32'b11111111111111111100101010111101;
assign LUT_4[39507] = 32'b11111111111111110101110110110101;
assign LUT_4[39508] = 32'b11111111111111111010010000110101;
assign LUT_4[39509] = 32'b11111111111111110011011100101101;
assign LUT_4[39510] = 32'b11111111111111111001101011011001;
assign LUT_4[39511] = 32'b11111111111111110010110111010001;
assign LUT_4[39512] = 32'b11111111111111110110011100101110;
assign LUT_4[39513] = 32'b11111111111111101111101000100110;
assign LUT_4[39514] = 32'b11111111111111110101110111010010;
assign LUT_4[39515] = 32'b11111111111111101111000011001010;
assign LUT_4[39516] = 32'b11111111111111110011011101001010;
assign LUT_4[39517] = 32'b11111111111111101100101001000010;
assign LUT_4[39518] = 32'b11111111111111110010110111101110;
assign LUT_4[39519] = 32'b11111111111111101100000011100110;
assign LUT_4[39520] = 32'b11111111111111111101111001110010;
assign LUT_4[39521] = 32'b11111111111111110111000101101010;
assign LUT_4[39522] = 32'b11111111111111111101010100010110;
assign LUT_4[39523] = 32'b11111111111111110110100000001110;
assign LUT_4[39524] = 32'b11111111111111111010111010001110;
assign LUT_4[39525] = 32'b11111111111111110100000110000110;
assign LUT_4[39526] = 32'b11111111111111111010010100110010;
assign LUT_4[39527] = 32'b11111111111111110011100000101010;
assign LUT_4[39528] = 32'b11111111111111110111000110000111;
assign LUT_4[39529] = 32'b11111111111111110000010001111111;
assign LUT_4[39530] = 32'b11111111111111110110100000101011;
assign LUT_4[39531] = 32'b11111111111111101111101100100011;
assign LUT_4[39532] = 32'b11111111111111110100000110100011;
assign LUT_4[39533] = 32'b11111111111111101101010010011011;
assign LUT_4[39534] = 32'b11111111111111110011100001000111;
assign LUT_4[39535] = 32'b11111111111111101100101100111111;
assign LUT_4[39536] = 32'b11111111111111111011101011100000;
assign LUT_4[39537] = 32'b11111111111111110100110111011000;
assign LUT_4[39538] = 32'b11111111111111111011000110000100;
assign LUT_4[39539] = 32'b11111111111111110100010001111100;
assign LUT_4[39540] = 32'b11111111111111111000101011111100;
assign LUT_4[39541] = 32'b11111111111111110001110111110100;
assign LUT_4[39542] = 32'b11111111111111111000000110100000;
assign LUT_4[39543] = 32'b11111111111111110001010010011000;
assign LUT_4[39544] = 32'b11111111111111110100110111110101;
assign LUT_4[39545] = 32'b11111111111111101110000011101101;
assign LUT_4[39546] = 32'b11111111111111110100010010011001;
assign LUT_4[39547] = 32'b11111111111111101101011110010001;
assign LUT_4[39548] = 32'b11111111111111110001111000010001;
assign LUT_4[39549] = 32'b11111111111111101011000100001001;
assign LUT_4[39550] = 32'b11111111111111110001010010110101;
assign LUT_4[39551] = 32'b11111111111111101010011110101101;
assign LUT_4[39552] = 32'b00000000000000000000101101011111;
assign LUT_4[39553] = 32'b11111111111111111001111001010111;
assign LUT_4[39554] = 32'b00000000000000000000001000000011;
assign LUT_4[39555] = 32'b11111111111111111001010011111011;
assign LUT_4[39556] = 32'b11111111111111111101101101111011;
assign LUT_4[39557] = 32'b11111111111111110110111001110011;
assign LUT_4[39558] = 32'b11111111111111111101001000011111;
assign LUT_4[39559] = 32'b11111111111111110110010100010111;
assign LUT_4[39560] = 32'b11111111111111111001111001110100;
assign LUT_4[39561] = 32'b11111111111111110011000101101100;
assign LUT_4[39562] = 32'b11111111111111111001010100011000;
assign LUT_4[39563] = 32'b11111111111111110010100000010000;
assign LUT_4[39564] = 32'b11111111111111110110111010010000;
assign LUT_4[39565] = 32'b11111111111111110000000110001000;
assign LUT_4[39566] = 32'b11111111111111110110010100110100;
assign LUT_4[39567] = 32'b11111111111111101111100000101100;
assign LUT_4[39568] = 32'b11111111111111111110011111001101;
assign LUT_4[39569] = 32'b11111111111111110111101011000101;
assign LUT_4[39570] = 32'b11111111111111111101111001110001;
assign LUT_4[39571] = 32'b11111111111111110111000101101001;
assign LUT_4[39572] = 32'b11111111111111111011011111101001;
assign LUT_4[39573] = 32'b11111111111111110100101011100001;
assign LUT_4[39574] = 32'b11111111111111111010111010001101;
assign LUT_4[39575] = 32'b11111111111111110100000110000101;
assign LUT_4[39576] = 32'b11111111111111110111101011100010;
assign LUT_4[39577] = 32'b11111111111111110000110111011010;
assign LUT_4[39578] = 32'b11111111111111110111000110000110;
assign LUT_4[39579] = 32'b11111111111111110000010001111110;
assign LUT_4[39580] = 32'b11111111111111110100101011111110;
assign LUT_4[39581] = 32'b11111111111111101101110111110110;
assign LUT_4[39582] = 32'b11111111111111110100000110100010;
assign LUT_4[39583] = 32'b11111111111111101101010010011010;
assign LUT_4[39584] = 32'b11111111111111111111001000100110;
assign LUT_4[39585] = 32'b11111111111111111000010100011110;
assign LUT_4[39586] = 32'b11111111111111111110100011001010;
assign LUT_4[39587] = 32'b11111111111111110111101111000010;
assign LUT_4[39588] = 32'b11111111111111111100001001000010;
assign LUT_4[39589] = 32'b11111111111111110101010100111010;
assign LUT_4[39590] = 32'b11111111111111111011100011100110;
assign LUT_4[39591] = 32'b11111111111111110100101111011110;
assign LUT_4[39592] = 32'b11111111111111111000010100111011;
assign LUT_4[39593] = 32'b11111111111111110001100000110011;
assign LUT_4[39594] = 32'b11111111111111110111101111011111;
assign LUT_4[39595] = 32'b11111111111111110000111011010111;
assign LUT_4[39596] = 32'b11111111111111110101010101010111;
assign LUT_4[39597] = 32'b11111111111111101110100001001111;
assign LUT_4[39598] = 32'b11111111111111110100101111111011;
assign LUT_4[39599] = 32'b11111111111111101101111011110011;
assign LUT_4[39600] = 32'b11111111111111111100111010010100;
assign LUT_4[39601] = 32'b11111111111111110110000110001100;
assign LUT_4[39602] = 32'b11111111111111111100010100111000;
assign LUT_4[39603] = 32'b11111111111111110101100000110000;
assign LUT_4[39604] = 32'b11111111111111111001111010110000;
assign LUT_4[39605] = 32'b11111111111111110011000110101000;
assign LUT_4[39606] = 32'b11111111111111111001010101010100;
assign LUT_4[39607] = 32'b11111111111111110010100001001100;
assign LUT_4[39608] = 32'b11111111111111110110000110101001;
assign LUT_4[39609] = 32'b11111111111111101111010010100001;
assign LUT_4[39610] = 32'b11111111111111110101100001001101;
assign LUT_4[39611] = 32'b11111111111111101110101101000101;
assign LUT_4[39612] = 32'b11111111111111110011000111000101;
assign LUT_4[39613] = 32'b11111111111111101100010010111101;
assign LUT_4[39614] = 32'b11111111111111110010100001101001;
assign LUT_4[39615] = 32'b11111111111111101011101101100001;
assign LUT_4[39616] = 32'b00000000000000000010000100110011;
assign LUT_4[39617] = 32'b11111111111111111011010000101011;
assign LUT_4[39618] = 32'b00000000000000000001011111010111;
assign LUT_4[39619] = 32'b11111111111111111010101011001111;
assign LUT_4[39620] = 32'b11111111111111111111000101001111;
assign LUT_4[39621] = 32'b11111111111111111000010001000111;
assign LUT_4[39622] = 32'b11111111111111111110011111110011;
assign LUT_4[39623] = 32'b11111111111111110111101011101011;
assign LUT_4[39624] = 32'b11111111111111111011010001001000;
assign LUT_4[39625] = 32'b11111111111111110100011101000000;
assign LUT_4[39626] = 32'b11111111111111111010101011101100;
assign LUT_4[39627] = 32'b11111111111111110011110111100100;
assign LUT_4[39628] = 32'b11111111111111111000010001100100;
assign LUT_4[39629] = 32'b11111111111111110001011101011100;
assign LUT_4[39630] = 32'b11111111111111110111101100001000;
assign LUT_4[39631] = 32'b11111111111111110000111000000000;
assign LUT_4[39632] = 32'b11111111111111111111110110100001;
assign LUT_4[39633] = 32'b11111111111111111001000010011001;
assign LUT_4[39634] = 32'b11111111111111111111010001000101;
assign LUT_4[39635] = 32'b11111111111111111000011100111101;
assign LUT_4[39636] = 32'b11111111111111111100110110111101;
assign LUT_4[39637] = 32'b11111111111111110110000010110101;
assign LUT_4[39638] = 32'b11111111111111111100010001100001;
assign LUT_4[39639] = 32'b11111111111111110101011101011001;
assign LUT_4[39640] = 32'b11111111111111111001000010110110;
assign LUT_4[39641] = 32'b11111111111111110010001110101110;
assign LUT_4[39642] = 32'b11111111111111111000011101011010;
assign LUT_4[39643] = 32'b11111111111111110001101001010010;
assign LUT_4[39644] = 32'b11111111111111110110000011010010;
assign LUT_4[39645] = 32'b11111111111111101111001111001010;
assign LUT_4[39646] = 32'b11111111111111110101011101110110;
assign LUT_4[39647] = 32'b11111111111111101110101001101110;
assign LUT_4[39648] = 32'b00000000000000000000011111111010;
assign LUT_4[39649] = 32'b11111111111111111001101011110010;
assign LUT_4[39650] = 32'b11111111111111111111111010011110;
assign LUT_4[39651] = 32'b11111111111111111001000110010110;
assign LUT_4[39652] = 32'b11111111111111111101100000010110;
assign LUT_4[39653] = 32'b11111111111111110110101100001110;
assign LUT_4[39654] = 32'b11111111111111111100111010111010;
assign LUT_4[39655] = 32'b11111111111111110110000110110010;
assign LUT_4[39656] = 32'b11111111111111111001101100001111;
assign LUT_4[39657] = 32'b11111111111111110010111000000111;
assign LUT_4[39658] = 32'b11111111111111111001000110110011;
assign LUT_4[39659] = 32'b11111111111111110010010010101011;
assign LUT_4[39660] = 32'b11111111111111110110101100101011;
assign LUT_4[39661] = 32'b11111111111111101111111000100011;
assign LUT_4[39662] = 32'b11111111111111110110000111001111;
assign LUT_4[39663] = 32'b11111111111111101111010011000111;
assign LUT_4[39664] = 32'b11111111111111111110010001101000;
assign LUT_4[39665] = 32'b11111111111111110111011101100000;
assign LUT_4[39666] = 32'b11111111111111111101101100001100;
assign LUT_4[39667] = 32'b11111111111111110110111000000100;
assign LUT_4[39668] = 32'b11111111111111111011010010000100;
assign LUT_4[39669] = 32'b11111111111111110100011101111100;
assign LUT_4[39670] = 32'b11111111111111111010101100101000;
assign LUT_4[39671] = 32'b11111111111111110011111000100000;
assign LUT_4[39672] = 32'b11111111111111110111011101111101;
assign LUT_4[39673] = 32'b11111111111111110000101001110101;
assign LUT_4[39674] = 32'b11111111111111110110111000100001;
assign LUT_4[39675] = 32'b11111111111111110000000100011001;
assign LUT_4[39676] = 32'b11111111111111110100011110011001;
assign LUT_4[39677] = 32'b11111111111111101101101010010001;
assign LUT_4[39678] = 32'b11111111111111110011111000111101;
assign LUT_4[39679] = 32'b11111111111111101101000100110101;
assign LUT_4[39680] = 32'b00000000000000000011000010111010;
assign LUT_4[39681] = 32'b11111111111111111100001110110010;
assign LUT_4[39682] = 32'b00000000000000000010011101011110;
assign LUT_4[39683] = 32'b11111111111111111011101001010110;
assign LUT_4[39684] = 32'b00000000000000000000000011010110;
assign LUT_4[39685] = 32'b11111111111111111001001111001110;
assign LUT_4[39686] = 32'b11111111111111111111011101111010;
assign LUT_4[39687] = 32'b11111111111111111000101001110010;
assign LUT_4[39688] = 32'b11111111111111111100001111001111;
assign LUT_4[39689] = 32'b11111111111111110101011011000111;
assign LUT_4[39690] = 32'b11111111111111111011101001110011;
assign LUT_4[39691] = 32'b11111111111111110100110101101011;
assign LUT_4[39692] = 32'b11111111111111111001001111101011;
assign LUT_4[39693] = 32'b11111111111111110010011011100011;
assign LUT_4[39694] = 32'b11111111111111111000101010001111;
assign LUT_4[39695] = 32'b11111111111111110001110110000111;
assign LUT_4[39696] = 32'b00000000000000000000110100101000;
assign LUT_4[39697] = 32'b11111111111111111010000000100000;
assign LUT_4[39698] = 32'b00000000000000000000001111001100;
assign LUT_4[39699] = 32'b11111111111111111001011011000100;
assign LUT_4[39700] = 32'b11111111111111111101110101000100;
assign LUT_4[39701] = 32'b11111111111111110111000000111100;
assign LUT_4[39702] = 32'b11111111111111111101001111101000;
assign LUT_4[39703] = 32'b11111111111111110110011011100000;
assign LUT_4[39704] = 32'b11111111111111111010000000111101;
assign LUT_4[39705] = 32'b11111111111111110011001100110101;
assign LUT_4[39706] = 32'b11111111111111111001011011100001;
assign LUT_4[39707] = 32'b11111111111111110010100111011001;
assign LUT_4[39708] = 32'b11111111111111110111000001011001;
assign LUT_4[39709] = 32'b11111111111111110000001101010001;
assign LUT_4[39710] = 32'b11111111111111110110011011111101;
assign LUT_4[39711] = 32'b11111111111111101111100111110101;
assign LUT_4[39712] = 32'b00000000000000000001011110000001;
assign LUT_4[39713] = 32'b11111111111111111010101001111001;
assign LUT_4[39714] = 32'b00000000000000000000111000100101;
assign LUT_4[39715] = 32'b11111111111111111010000100011101;
assign LUT_4[39716] = 32'b11111111111111111110011110011101;
assign LUT_4[39717] = 32'b11111111111111110111101010010101;
assign LUT_4[39718] = 32'b11111111111111111101111001000001;
assign LUT_4[39719] = 32'b11111111111111110111000100111001;
assign LUT_4[39720] = 32'b11111111111111111010101010010110;
assign LUT_4[39721] = 32'b11111111111111110011110110001110;
assign LUT_4[39722] = 32'b11111111111111111010000100111010;
assign LUT_4[39723] = 32'b11111111111111110011010000110010;
assign LUT_4[39724] = 32'b11111111111111110111101010110010;
assign LUT_4[39725] = 32'b11111111111111110000110110101010;
assign LUT_4[39726] = 32'b11111111111111110111000101010110;
assign LUT_4[39727] = 32'b11111111111111110000010001001110;
assign LUT_4[39728] = 32'b11111111111111111111001111101111;
assign LUT_4[39729] = 32'b11111111111111111000011011100111;
assign LUT_4[39730] = 32'b11111111111111111110101010010011;
assign LUT_4[39731] = 32'b11111111111111110111110110001011;
assign LUT_4[39732] = 32'b11111111111111111100010000001011;
assign LUT_4[39733] = 32'b11111111111111110101011100000011;
assign LUT_4[39734] = 32'b11111111111111111011101010101111;
assign LUT_4[39735] = 32'b11111111111111110100110110100111;
assign LUT_4[39736] = 32'b11111111111111111000011100000100;
assign LUT_4[39737] = 32'b11111111111111110001100111111100;
assign LUT_4[39738] = 32'b11111111111111110111110110101000;
assign LUT_4[39739] = 32'b11111111111111110001000010100000;
assign LUT_4[39740] = 32'b11111111111111110101011100100000;
assign LUT_4[39741] = 32'b11111111111111101110101000011000;
assign LUT_4[39742] = 32'b11111111111111110100110111000100;
assign LUT_4[39743] = 32'b11111111111111101110000010111100;
assign LUT_4[39744] = 32'b00000000000000000100011010001110;
assign LUT_4[39745] = 32'b11111111111111111101100110000110;
assign LUT_4[39746] = 32'b00000000000000000011110100110010;
assign LUT_4[39747] = 32'b11111111111111111101000000101010;
assign LUT_4[39748] = 32'b00000000000000000001011010101010;
assign LUT_4[39749] = 32'b11111111111111111010100110100010;
assign LUT_4[39750] = 32'b00000000000000000000110101001110;
assign LUT_4[39751] = 32'b11111111111111111010000001000110;
assign LUT_4[39752] = 32'b11111111111111111101100110100011;
assign LUT_4[39753] = 32'b11111111111111110110110010011011;
assign LUT_4[39754] = 32'b11111111111111111101000001000111;
assign LUT_4[39755] = 32'b11111111111111110110001100111111;
assign LUT_4[39756] = 32'b11111111111111111010100110111111;
assign LUT_4[39757] = 32'b11111111111111110011110010110111;
assign LUT_4[39758] = 32'b11111111111111111010000001100011;
assign LUT_4[39759] = 32'b11111111111111110011001101011011;
assign LUT_4[39760] = 32'b00000000000000000010001011111100;
assign LUT_4[39761] = 32'b11111111111111111011010111110100;
assign LUT_4[39762] = 32'b00000000000000000001100110100000;
assign LUT_4[39763] = 32'b11111111111111111010110010011000;
assign LUT_4[39764] = 32'b11111111111111111111001100011000;
assign LUT_4[39765] = 32'b11111111111111111000011000010000;
assign LUT_4[39766] = 32'b11111111111111111110100110111100;
assign LUT_4[39767] = 32'b11111111111111110111110010110100;
assign LUT_4[39768] = 32'b11111111111111111011011000010001;
assign LUT_4[39769] = 32'b11111111111111110100100100001001;
assign LUT_4[39770] = 32'b11111111111111111010110010110101;
assign LUT_4[39771] = 32'b11111111111111110011111110101101;
assign LUT_4[39772] = 32'b11111111111111111000011000101101;
assign LUT_4[39773] = 32'b11111111111111110001100100100101;
assign LUT_4[39774] = 32'b11111111111111110111110011010001;
assign LUT_4[39775] = 32'b11111111111111110000111111001001;
assign LUT_4[39776] = 32'b00000000000000000010110101010101;
assign LUT_4[39777] = 32'b11111111111111111100000001001101;
assign LUT_4[39778] = 32'b00000000000000000010001111111001;
assign LUT_4[39779] = 32'b11111111111111111011011011110001;
assign LUT_4[39780] = 32'b11111111111111111111110101110001;
assign LUT_4[39781] = 32'b11111111111111111001000001101001;
assign LUT_4[39782] = 32'b11111111111111111111010000010101;
assign LUT_4[39783] = 32'b11111111111111111000011100001101;
assign LUT_4[39784] = 32'b11111111111111111100000001101010;
assign LUT_4[39785] = 32'b11111111111111110101001101100010;
assign LUT_4[39786] = 32'b11111111111111111011011100001110;
assign LUT_4[39787] = 32'b11111111111111110100101000000110;
assign LUT_4[39788] = 32'b11111111111111111001000010000110;
assign LUT_4[39789] = 32'b11111111111111110010001101111110;
assign LUT_4[39790] = 32'b11111111111111111000011100101010;
assign LUT_4[39791] = 32'b11111111111111110001101000100010;
assign LUT_4[39792] = 32'b00000000000000000000100111000011;
assign LUT_4[39793] = 32'b11111111111111111001110010111011;
assign LUT_4[39794] = 32'b00000000000000000000000001100111;
assign LUT_4[39795] = 32'b11111111111111111001001101011111;
assign LUT_4[39796] = 32'b11111111111111111101100111011111;
assign LUT_4[39797] = 32'b11111111111111110110110011010111;
assign LUT_4[39798] = 32'b11111111111111111101000010000011;
assign LUT_4[39799] = 32'b11111111111111110110001101111011;
assign LUT_4[39800] = 32'b11111111111111111001110011011000;
assign LUT_4[39801] = 32'b11111111111111110010111111010000;
assign LUT_4[39802] = 32'b11111111111111111001001101111100;
assign LUT_4[39803] = 32'b11111111111111110010011001110100;
assign LUT_4[39804] = 32'b11111111111111110110110011110100;
assign LUT_4[39805] = 32'b11111111111111101111111111101100;
assign LUT_4[39806] = 32'b11111111111111110110001110011000;
assign LUT_4[39807] = 32'b11111111111111101111011010010000;
assign LUT_4[39808] = 32'b00000000000000000101101001000010;
assign LUT_4[39809] = 32'b11111111111111111110110100111010;
assign LUT_4[39810] = 32'b00000000000000000101000011100110;
assign LUT_4[39811] = 32'b11111111111111111110001111011110;
assign LUT_4[39812] = 32'b00000000000000000010101001011110;
assign LUT_4[39813] = 32'b11111111111111111011110101010110;
assign LUT_4[39814] = 32'b00000000000000000010000100000010;
assign LUT_4[39815] = 32'b11111111111111111011001111111010;
assign LUT_4[39816] = 32'b11111111111111111110110101010111;
assign LUT_4[39817] = 32'b11111111111111111000000001001111;
assign LUT_4[39818] = 32'b11111111111111111110001111111011;
assign LUT_4[39819] = 32'b11111111111111110111011011110011;
assign LUT_4[39820] = 32'b11111111111111111011110101110011;
assign LUT_4[39821] = 32'b11111111111111110101000001101011;
assign LUT_4[39822] = 32'b11111111111111111011010000010111;
assign LUT_4[39823] = 32'b11111111111111110100011100001111;
assign LUT_4[39824] = 32'b00000000000000000011011010110000;
assign LUT_4[39825] = 32'b11111111111111111100100110101000;
assign LUT_4[39826] = 32'b00000000000000000010110101010100;
assign LUT_4[39827] = 32'b11111111111111111100000001001100;
assign LUT_4[39828] = 32'b00000000000000000000011011001100;
assign LUT_4[39829] = 32'b11111111111111111001100111000100;
assign LUT_4[39830] = 32'b11111111111111111111110101110000;
assign LUT_4[39831] = 32'b11111111111111111001000001101000;
assign LUT_4[39832] = 32'b11111111111111111100100111000101;
assign LUT_4[39833] = 32'b11111111111111110101110010111101;
assign LUT_4[39834] = 32'b11111111111111111100000001101001;
assign LUT_4[39835] = 32'b11111111111111110101001101100001;
assign LUT_4[39836] = 32'b11111111111111111001100111100001;
assign LUT_4[39837] = 32'b11111111111111110010110011011001;
assign LUT_4[39838] = 32'b11111111111111111001000010000101;
assign LUT_4[39839] = 32'b11111111111111110010001101111101;
assign LUT_4[39840] = 32'b00000000000000000100000100001001;
assign LUT_4[39841] = 32'b11111111111111111101010000000001;
assign LUT_4[39842] = 32'b00000000000000000011011110101101;
assign LUT_4[39843] = 32'b11111111111111111100101010100101;
assign LUT_4[39844] = 32'b00000000000000000001000100100101;
assign LUT_4[39845] = 32'b11111111111111111010010000011101;
assign LUT_4[39846] = 32'b00000000000000000000011111001001;
assign LUT_4[39847] = 32'b11111111111111111001101011000001;
assign LUT_4[39848] = 32'b11111111111111111101010000011110;
assign LUT_4[39849] = 32'b11111111111111110110011100010110;
assign LUT_4[39850] = 32'b11111111111111111100101011000010;
assign LUT_4[39851] = 32'b11111111111111110101110110111010;
assign LUT_4[39852] = 32'b11111111111111111010010000111010;
assign LUT_4[39853] = 32'b11111111111111110011011100110010;
assign LUT_4[39854] = 32'b11111111111111111001101011011110;
assign LUT_4[39855] = 32'b11111111111111110010110111010110;
assign LUT_4[39856] = 32'b00000000000000000001110101110111;
assign LUT_4[39857] = 32'b11111111111111111011000001101111;
assign LUT_4[39858] = 32'b00000000000000000001010000011011;
assign LUT_4[39859] = 32'b11111111111111111010011100010011;
assign LUT_4[39860] = 32'b11111111111111111110110110010011;
assign LUT_4[39861] = 32'b11111111111111111000000010001011;
assign LUT_4[39862] = 32'b11111111111111111110010000110111;
assign LUT_4[39863] = 32'b11111111111111110111011100101111;
assign LUT_4[39864] = 32'b11111111111111111011000010001100;
assign LUT_4[39865] = 32'b11111111111111110100001110000100;
assign LUT_4[39866] = 32'b11111111111111111010011100110000;
assign LUT_4[39867] = 32'b11111111111111110011101000101000;
assign LUT_4[39868] = 32'b11111111111111111000000010101000;
assign LUT_4[39869] = 32'b11111111111111110001001110100000;
assign LUT_4[39870] = 32'b11111111111111110111011101001100;
assign LUT_4[39871] = 32'b11111111111111110000101001000100;
assign LUT_4[39872] = 32'b00000000000000000111000000010110;
assign LUT_4[39873] = 32'b00000000000000000000001100001110;
assign LUT_4[39874] = 32'b00000000000000000110011010111010;
assign LUT_4[39875] = 32'b11111111111111111111100110110010;
assign LUT_4[39876] = 32'b00000000000000000100000000110010;
assign LUT_4[39877] = 32'b11111111111111111101001100101010;
assign LUT_4[39878] = 32'b00000000000000000011011011010110;
assign LUT_4[39879] = 32'b11111111111111111100100111001110;
assign LUT_4[39880] = 32'b00000000000000000000001100101011;
assign LUT_4[39881] = 32'b11111111111111111001011000100011;
assign LUT_4[39882] = 32'b11111111111111111111100111001111;
assign LUT_4[39883] = 32'b11111111111111111000110011000111;
assign LUT_4[39884] = 32'b11111111111111111101001101000111;
assign LUT_4[39885] = 32'b11111111111111110110011000111111;
assign LUT_4[39886] = 32'b11111111111111111100100111101011;
assign LUT_4[39887] = 32'b11111111111111110101110011100011;
assign LUT_4[39888] = 32'b00000000000000000100110010000100;
assign LUT_4[39889] = 32'b11111111111111111101111101111100;
assign LUT_4[39890] = 32'b00000000000000000100001100101000;
assign LUT_4[39891] = 32'b11111111111111111101011000100000;
assign LUT_4[39892] = 32'b00000000000000000001110010100000;
assign LUT_4[39893] = 32'b11111111111111111010111110011000;
assign LUT_4[39894] = 32'b00000000000000000001001101000100;
assign LUT_4[39895] = 32'b11111111111111111010011000111100;
assign LUT_4[39896] = 32'b11111111111111111101111110011001;
assign LUT_4[39897] = 32'b11111111111111110111001010010001;
assign LUT_4[39898] = 32'b11111111111111111101011000111101;
assign LUT_4[39899] = 32'b11111111111111110110100100110101;
assign LUT_4[39900] = 32'b11111111111111111010111110110101;
assign LUT_4[39901] = 32'b11111111111111110100001010101101;
assign LUT_4[39902] = 32'b11111111111111111010011001011001;
assign LUT_4[39903] = 32'b11111111111111110011100101010001;
assign LUT_4[39904] = 32'b00000000000000000101011011011101;
assign LUT_4[39905] = 32'b11111111111111111110100111010101;
assign LUT_4[39906] = 32'b00000000000000000100110110000001;
assign LUT_4[39907] = 32'b11111111111111111110000001111001;
assign LUT_4[39908] = 32'b00000000000000000010011011111001;
assign LUT_4[39909] = 32'b11111111111111111011100111110001;
assign LUT_4[39910] = 32'b00000000000000000001110110011101;
assign LUT_4[39911] = 32'b11111111111111111011000010010101;
assign LUT_4[39912] = 32'b11111111111111111110100111110010;
assign LUT_4[39913] = 32'b11111111111111110111110011101010;
assign LUT_4[39914] = 32'b11111111111111111110000010010110;
assign LUT_4[39915] = 32'b11111111111111110111001110001110;
assign LUT_4[39916] = 32'b11111111111111111011101000001110;
assign LUT_4[39917] = 32'b11111111111111110100110100000110;
assign LUT_4[39918] = 32'b11111111111111111011000010110010;
assign LUT_4[39919] = 32'b11111111111111110100001110101010;
assign LUT_4[39920] = 32'b00000000000000000011001101001011;
assign LUT_4[39921] = 32'b11111111111111111100011001000011;
assign LUT_4[39922] = 32'b00000000000000000010100111101111;
assign LUT_4[39923] = 32'b11111111111111111011110011100111;
assign LUT_4[39924] = 32'b00000000000000000000001101100111;
assign LUT_4[39925] = 32'b11111111111111111001011001011111;
assign LUT_4[39926] = 32'b11111111111111111111101000001011;
assign LUT_4[39927] = 32'b11111111111111111000110100000011;
assign LUT_4[39928] = 32'b11111111111111111100011001100000;
assign LUT_4[39929] = 32'b11111111111111110101100101011000;
assign LUT_4[39930] = 32'b11111111111111111011110100000100;
assign LUT_4[39931] = 32'b11111111111111110100111111111100;
assign LUT_4[39932] = 32'b11111111111111111001011001111100;
assign LUT_4[39933] = 32'b11111111111111110010100101110100;
assign LUT_4[39934] = 32'b11111111111111111000110100100000;
assign LUT_4[39935] = 32'b11111111111111110010000000011000;
assign LUT_4[39936] = 32'b00000000000000000000101101101110;
assign LUT_4[39937] = 32'b11111111111111111001111001100110;
assign LUT_4[39938] = 32'b00000000000000000000001000010010;
assign LUT_4[39939] = 32'b11111111111111111001010100001010;
assign LUT_4[39940] = 32'b11111111111111111101101110001010;
assign LUT_4[39941] = 32'b11111111111111110110111010000010;
assign LUT_4[39942] = 32'b11111111111111111101001000101110;
assign LUT_4[39943] = 32'b11111111111111110110010100100110;
assign LUT_4[39944] = 32'b11111111111111111001111010000011;
assign LUT_4[39945] = 32'b11111111111111110011000101111011;
assign LUT_4[39946] = 32'b11111111111111111001010100100111;
assign LUT_4[39947] = 32'b11111111111111110010100000011111;
assign LUT_4[39948] = 32'b11111111111111110110111010011111;
assign LUT_4[39949] = 32'b11111111111111110000000110010111;
assign LUT_4[39950] = 32'b11111111111111110110010101000011;
assign LUT_4[39951] = 32'b11111111111111101111100000111011;
assign LUT_4[39952] = 32'b11111111111111111110011111011100;
assign LUT_4[39953] = 32'b11111111111111110111101011010100;
assign LUT_4[39954] = 32'b11111111111111111101111010000000;
assign LUT_4[39955] = 32'b11111111111111110111000101111000;
assign LUT_4[39956] = 32'b11111111111111111011011111111000;
assign LUT_4[39957] = 32'b11111111111111110100101011110000;
assign LUT_4[39958] = 32'b11111111111111111010111010011100;
assign LUT_4[39959] = 32'b11111111111111110100000110010100;
assign LUT_4[39960] = 32'b11111111111111110111101011110001;
assign LUT_4[39961] = 32'b11111111111111110000110111101001;
assign LUT_4[39962] = 32'b11111111111111110111000110010101;
assign LUT_4[39963] = 32'b11111111111111110000010010001101;
assign LUT_4[39964] = 32'b11111111111111110100101100001101;
assign LUT_4[39965] = 32'b11111111111111101101111000000101;
assign LUT_4[39966] = 32'b11111111111111110100000110110001;
assign LUT_4[39967] = 32'b11111111111111101101010010101001;
assign LUT_4[39968] = 32'b11111111111111111111001000110101;
assign LUT_4[39969] = 32'b11111111111111111000010100101101;
assign LUT_4[39970] = 32'b11111111111111111110100011011001;
assign LUT_4[39971] = 32'b11111111111111110111101111010001;
assign LUT_4[39972] = 32'b11111111111111111100001001010001;
assign LUT_4[39973] = 32'b11111111111111110101010101001001;
assign LUT_4[39974] = 32'b11111111111111111011100011110101;
assign LUT_4[39975] = 32'b11111111111111110100101111101101;
assign LUT_4[39976] = 32'b11111111111111111000010101001010;
assign LUT_4[39977] = 32'b11111111111111110001100001000010;
assign LUT_4[39978] = 32'b11111111111111110111101111101110;
assign LUT_4[39979] = 32'b11111111111111110000111011100110;
assign LUT_4[39980] = 32'b11111111111111110101010101100110;
assign LUT_4[39981] = 32'b11111111111111101110100001011110;
assign LUT_4[39982] = 32'b11111111111111110100110000001010;
assign LUT_4[39983] = 32'b11111111111111101101111100000010;
assign LUT_4[39984] = 32'b11111111111111111100111010100011;
assign LUT_4[39985] = 32'b11111111111111110110000110011011;
assign LUT_4[39986] = 32'b11111111111111111100010101000111;
assign LUT_4[39987] = 32'b11111111111111110101100000111111;
assign LUT_4[39988] = 32'b11111111111111111001111010111111;
assign LUT_4[39989] = 32'b11111111111111110011000110110111;
assign LUT_4[39990] = 32'b11111111111111111001010101100011;
assign LUT_4[39991] = 32'b11111111111111110010100001011011;
assign LUT_4[39992] = 32'b11111111111111110110000110111000;
assign LUT_4[39993] = 32'b11111111111111101111010010110000;
assign LUT_4[39994] = 32'b11111111111111110101100001011100;
assign LUT_4[39995] = 32'b11111111111111101110101101010100;
assign LUT_4[39996] = 32'b11111111111111110011000111010100;
assign LUT_4[39997] = 32'b11111111111111101100010011001100;
assign LUT_4[39998] = 32'b11111111111111110010100001111000;
assign LUT_4[39999] = 32'b11111111111111101011101101110000;
assign LUT_4[40000] = 32'b00000000000000000010000101000010;
assign LUT_4[40001] = 32'b11111111111111111011010000111010;
assign LUT_4[40002] = 32'b00000000000000000001011111100110;
assign LUT_4[40003] = 32'b11111111111111111010101011011110;
assign LUT_4[40004] = 32'b11111111111111111111000101011110;
assign LUT_4[40005] = 32'b11111111111111111000010001010110;
assign LUT_4[40006] = 32'b11111111111111111110100000000010;
assign LUT_4[40007] = 32'b11111111111111110111101011111010;
assign LUT_4[40008] = 32'b11111111111111111011010001010111;
assign LUT_4[40009] = 32'b11111111111111110100011101001111;
assign LUT_4[40010] = 32'b11111111111111111010101011111011;
assign LUT_4[40011] = 32'b11111111111111110011110111110011;
assign LUT_4[40012] = 32'b11111111111111111000010001110011;
assign LUT_4[40013] = 32'b11111111111111110001011101101011;
assign LUT_4[40014] = 32'b11111111111111110111101100010111;
assign LUT_4[40015] = 32'b11111111111111110000111000001111;
assign LUT_4[40016] = 32'b11111111111111111111110110110000;
assign LUT_4[40017] = 32'b11111111111111111001000010101000;
assign LUT_4[40018] = 32'b11111111111111111111010001010100;
assign LUT_4[40019] = 32'b11111111111111111000011101001100;
assign LUT_4[40020] = 32'b11111111111111111100110111001100;
assign LUT_4[40021] = 32'b11111111111111110110000011000100;
assign LUT_4[40022] = 32'b11111111111111111100010001110000;
assign LUT_4[40023] = 32'b11111111111111110101011101101000;
assign LUT_4[40024] = 32'b11111111111111111001000011000101;
assign LUT_4[40025] = 32'b11111111111111110010001110111101;
assign LUT_4[40026] = 32'b11111111111111111000011101101001;
assign LUT_4[40027] = 32'b11111111111111110001101001100001;
assign LUT_4[40028] = 32'b11111111111111110110000011100001;
assign LUT_4[40029] = 32'b11111111111111101111001111011001;
assign LUT_4[40030] = 32'b11111111111111110101011110000101;
assign LUT_4[40031] = 32'b11111111111111101110101001111101;
assign LUT_4[40032] = 32'b00000000000000000000100000001001;
assign LUT_4[40033] = 32'b11111111111111111001101100000001;
assign LUT_4[40034] = 32'b11111111111111111111111010101101;
assign LUT_4[40035] = 32'b11111111111111111001000110100101;
assign LUT_4[40036] = 32'b11111111111111111101100000100101;
assign LUT_4[40037] = 32'b11111111111111110110101100011101;
assign LUT_4[40038] = 32'b11111111111111111100111011001001;
assign LUT_4[40039] = 32'b11111111111111110110000111000001;
assign LUT_4[40040] = 32'b11111111111111111001101100011110;
assign LUT_4[40041] = 32'b11111111111111110010111000010110;
assign LUT_4[40042] = 32'b11111111111111111001000111000010;
assign LUT_4[40043] = 32'b11111111111111110010010010111010;
assign LUT_4[40044] = 32'b11111111111111110110101100111010;
assign LUT_4[40045] = 32'b11111111111111101111111000110010;
assign LUT_4[40046] = 32'b11111111111111110110000111011110;
assign LUT_4[40047] = 32'b11111111111111101111010011010110;
assign LUT_4[40048] = 32'b11111111111111111110010001110111;
assign LUT_4[40049] = 32'b11111111111111110111011101101111;
assign LUT_4[40050] = 32'b11111111111111111101101100011011;
assign LUT_4[40051] = 32'b11111111111111110110111000010011;
assign LUT_4[40052] = 32'b11111111111111111011010010010011;
assign LUT_4[40053] = 32'b11111111111111110100011110001011;
assign LUT_4[40054] = 32'b11111111111111111010101100110111;
assign LUT_4[40055] = 32'b11111111111111110011111000101111;
assign LUT_4[40056] = 32'b11111111111111110111011110001100;
assign LUT_4[40057] = 32'b11111111111111110000101010000100;
assign LUT_4[40058] = 32'b11111111111111110110111000110000;
assign LUT_4[40059] = 32'b11111111111111110000000100101000;
assign LUT_4[40060] = 32'b11111111111111110100011110101000;
assign LUT_4[40061] = 32'b11111111111111101101101010100000;
assign LUT_4[40062] = 32'b11111111111111110011111001001100;
assign LUT_4[40063] = 32'b11111111111111101101000101000100;
assign LUT_4[40064] = 32'b00000000000000000011010011110110;
assign LUT_4[40065] = 32'b11111111111111111100011111101110;
assign LUT_4[40066] = 32'b00000000000000000010101110011010;
assign LUT_4[40067] = 32'b11111111111111111011111010010010;
assign LUT_4[40068] = 32'b00000000000000000000010100010010;
assign LUT_4[40069] = 32'b11111111111111111001100000001010;
assign LUT_4[40070] = 32'b11111111111111111111101110110110;
assign LUT_4[40071] = 32'b11111111111111111000111010101110;
assign LUT_4[40072] = 32'b11111111111111111100100000001011;
assign LUT_4[40073] = 32'b11111111111111110101101100000011;
assign LUT_4[40074] = 32'b11111111111111111011111010101111;
assign LUT_4[40075] = 32'b11111111111111110101000110100111;
assign LUT_4[40076] = 32'b11111111111111111001100000100111;
assign LUT_4[40077] = 32'b11111111111111110010101100011111;
assign LUT_4[40078] = 32'b11111111111111111000111011001011;
assign LUT_4[40079] = 32'b11111111111111110010000111000011;
assign LUT_4[40080] = 32'b00000000000000000001000101100100;
assign LUT_4[40081] = 32'b11111111111111111010010001011100;
assign LUT_4[40082] = 32'b00000000000000000000100000001000;
assign LUT_4[40083] = 32'b11111111111111111001101100000000;
assign LUT_4[40084] = 32'b11111111111111111110000110000000;
assign LUT_4[40085] = 32'b11111111111111110111010001111000;
assign LUT_4[40086] = 32'b11111111111111111101100000100100;
assign LUT_4[40087] = 32'b11111111111111110110101100011100;
assign LUT_4[40088] = 32'b11111111111111111010010001111001;
assign LUT_4[40089] = 32'b11111111111111110011011101110001;
assign LUT_4[40090] = 32'b11111111111111111001101100011101;
assign LUT_4[40091] = 32'b11111111111111110010111000010101;
assign LUT_4[40092] = 32'b11111111111111110111010010010101;
assign LUT_4[40093] = 32'b11111111111111110000011110001101;
assign LUT_4[40094] = 32'b11111111111111110110101100111001;
assign LUT_4[40095] = 32'b11111111111111101111111000110001;
assign LUT_4[40096] = 32'b00000000000000000001101110111101;
assign LUT_4[40097] = 32'b11111111111111111010111010110101;
assign LUT_4[40098] = 32'b00000000000000000001001001100001;
assign LUT_4[40099] = 32'b11111111111111111010010101011001;
assign LUT_4[40100] = 32'b11111111111111111110101111011001;
assign LUT_4[40101] = 32'b11111111111111110111111011010001;
assign LUT_4[40102] = 32'b11111111111111111110001001111101;
assign LUT_4[40103] = 32'b11111111111111110111010101110101;
assign LUT_4[40104] = 32'b11111111111111111010111011010010;
assign LUT_4[40105] = 32'b11111111111111110100000111001010;
assign LUT_4[40106] = 32'b11111111111111111010010101110110;
assign LUT_4[40107] = 32'b11111111111111110011100001101110;
assign LUT_4[40108] = 32'b11111111111111110111111011101110;
assign LUT_4[40109] = 32'b11111111111111110001000111100110;
assign LUT_4[40110] = 32'b11111111111111110111010110010010;
assign LUT_4[40111] = 32'b11111111111111110000100010001010;
assign LUT_4[40112] = 32'b11111111111111111111100000101011;
assign LUT_4[40113] = 32'b11111111111111111000101100100011;
assign LUT_4[40114] = 32'b11111111111111111110111011001111;
assign LUT_4[40115] = 32'b11111111111111111000000111000111;
assign LUT_4[40116] = 32'b11111111111111111100100001000111;
assign LUT_4[40117] = 32'b11111111111111110101101100111111;
assign LUT_4[40118] = 32'b11111111111111111011111011101011;
assign LUT_4[40119] = 32'b11111111111111110101000111100011;
assign LUT_4[40120] = 32'b11111111111111111000101101000000;
assign LUT_4[40121] = 32'b11111111111111110001111000111000;
assign LUT_4[40122] = 32'b11111111111111111000000111100100;
assign LUT_4[40123] = 32'b11111111111111110001010011011100;
assign LUT_4[40124] = 32'b11111111111111110101101101011100;
assign LUT_4[40125] = 32'b11111111111111101110111001010100;
assign LUT_4[40126] = 32'b11111111111111110101001000000000;
assign LUT_4[40127] = 32'b11111111111111101110010011111000;
assign LUT_4[40128] = 32'b00000000000000000100101011001010;
assign LUT_4[40129] = 32'b11111111111111111101110111000010;
assign LUT_4[40130] = 32'b00000000000000000100000101101110;
assign LUT_4[40131] = 32'b11111111111111111101010001100110;
assign LUT_4[40132] = 32'b00000000000000000001101011100110;
assign LUT_4[40133] = 32'b11111111111111111010110111011110;
assign LUT_4[40134] = 32'b00000000000000000001000110001010;
assign LUT_4[40135] = 32'b11111111111111111010010010000010;
assign LUT_4[40136] = 32'b11111111111111111101110111011111;
assign LUT_4[40137] = 32'b11111111111111110111000011010111;
assign LUT_4[40138] = 32'b11111111111111111101010010000011;
assign LUT_4[40139] = 32'b11111111111111110110011101111011;
assign LUT_4[40140] = 32'b11111111111111111010110111111011;
assign LUT_4[40141] = 32'b11111111111111110100000011110011;
assign LUT_4[40142] = 32'b11111111111111111010010010011111;
assign LUT_4[40143] = 32'b11111111111111110011011110010111;
assign LUT_4[40144] = 32'b00000000000000000010011100111000;
assign LUT_4[40145] = 32'b11111111111111111011101000110000;
assign LUT_4[40146] = 32'b00000000000000000001110111011100;
assign LUT_4[40147] = 32'b11111111111111111011000011010100;
assign LUT_4[40148] = 32'b11111111111111111111011101010100;
assign LUT_4[40149] = 32'b11111111111111111000101001001100;
assign LUT_4[40150] = 32'b11111111111111111110110111111000;
assign LUT_4[40151] = 32'b11111111111111111000000011110000;
assign LUT_4[40152] = 32'b11111111111111111011101001001101;
assign LUT_4[40153] = 32'b11111111111111110100110101000101;
assign LUT_4[40154] = 32'b11111111111111111011000011110001;
assign LUT_4[40155] = 32'b11111111111111110100001111101001;
assign LUT_4[40156] = 32'b11111111111111111000101001101001;
assign LUT_4[40157] = 32'b11111111111111110001110101100001;
assign LUT_4[40158] = 32'b11111111111111111000000100001101;
assign LUT_4[40159] = 32'b11111111111111110001010000000101;
assign LUT_4[40160] = 32'b00000000000000000011000110010001;
assign LUT_4[40161] = 32'b11111111111111111100010010001001;
assign LUT_4[40162] = 32'b00000000000000000010100000110101;
assign LUT_4[40163] = 32'b11111111111111111011101100101101;
assign LUT_4[40164] = 32'b00000000000000000000000110101101;
assign LUT_4[40165] = 32'b11111111111111111001010010100101;
assign LUT_4[40166] = 32'b11111111111111111111100001010001;
assign LUT_4[40167] = 32'b11111111111111111000101101001001;
assign LUT_4[40168] = 32'b11111111111111111100010010100110;
assign LUT_4[40169] = 32'b11111111111111110101011110011110;
assign LUT_4[40170] = 32'b11111111111111111011101101001010;
assign LUT_4[40171] = 32'b11111111111111110100111001000010;
assign LUT_4[40172] = 32'b11111111111111111001010011000010;
assign LUT_4[40173] = 32'b11111111111111110010011110111010;
assign LUT_4[40174] = 32'b11111111111111111000101101100110;
assign LUT_4[40175] = 32'b11111111111111110001111001011110;
assign LUT_4[40176] = 32'b00000000000000000000110111111111;
assign LUT_4[40177] = 32'b11111111111111111010000011110111;
assign LUT_4[40178] = 32'b00000000000000000000010010100011;
assign LUT_4[40179] = 32'b11111111111111111001011110011011;
assign LUT_4[40180] = 32'b11111111111111111101111000011011;
assign LUT_4[40181] = 32'b11111111111111110111000100010011;
assign LUT_4[40182] = 32'b11111111111111111101010010111111;
assign LUT_4[40183] = 32'b11111111111111110110011110110111;
assign LUT_4[40184] = 32'b11111111111111111010000100010100;
assign LUT_4[40185] = 32'b11111111111111110011010000001100;
assign LUT_4[40186] = 32'b11111111111111111001011110111000;
assign LUT_4[40187] = 32'b11111111111111110010101010110000;
assign LUT_4[40188] = 32'b11111111111111110111000100110000;
assign LUT_4[40189] = 32'b11111111111111110000010000101000;
assign LUT_4[40190] = 32'b11111111111111110110011111010100;
assign LUT_4[40191] = 32'b11111111111111101111101011001100;
assign LUT_4[40192] = 32'b00000000000000000101101001010001;
assign LUT_4[40193] = 32'b11111111111111111110110101001001;
assign LUT_4[40194] = 32'b00000000000000000101000011110101;
assign LUT_4[40195] = 32'b11111111111111111110001111101101;
assign LUT_4[40196] = 32'b00000000000000000010101001101101;
assign LUT_4[40197] = 32'b11111111111111111011110101100101;
assign LUT_4[40198] = 32'b00000000000000000010000100010001;
assign LUT_4[40199] = 32'b11111111111111111011010000001001;
assign LUT_4[40200] = 32'b11111111111111111110110101100110;
assign LUT_4[40201] = 32'b11111111111111111000000001011110;
assign LUT_4[40202] = 32'b11111111111111111110010000001010;
assign LUT_4[40203] = 32'b11111111111111110111011100000010;
assign LUT_4[40204] = 32'b11111111111111111011110110000010;
assign LUT_4[40205] = 32'b11111111111111110101000001111010;
assign LUT_4[40206] = 32'b11111111111111111011010000100110;
assign LUT_4[40207] = 32'b11111111111111110100011100011110;
assign LUT_4[40208] = 32'b00000000000000000011011010111111;
assign LUT_4[40209] = 32'b11111111111111111100100110110111;
assign LUT_4[40210] = 32'b00000000000000000010110101100011;
assign LUT_4[40211] = 32'b11111111111111111100000001011011;
assign LUT_4[40212] = 32'b00000000000000000000011011011011;
assign LUT_4[40213] = 32'b11111111111111111001100111010011;
assign LUT_4[40214] = 32'b11111111111111111111110101111111;
assign LUT_4[40215] = 32'b11111111111111111001000001110111;
assign LUT_4[40216] = 32'b11111111111111111100100111010100;
assign LUT_4[40217] = 32'b11111111111111110101110011001100;
assign LUT_4[40218] = 32'b11111111111111111100000001111000;
assign LUT_4[40219] = 32'b11111111111111110101001101110000;
assign LUT_4[40220] = 32'b11111111111111111001100111110000;
assign LUT_4[40221] = 32'b11111111111111110010110011101000;
assign LUT_4[40222] = 32'b11111111111111111001000010010100;
assign LUT_4[40223] = 32'b11111111111111110010001110001100;
assign LUT_4[40224] = 32'b00000000000000000100000100011000;
assign LUT_4[40225] = 32'b11111111111111111101010000010000;
assign LUT_4[40226] = 32'b00000000000000000011011110111100;
assign LUT_4[40227] = 32'b11111111111111111100101010110100;
assign LUT_4[40228] = 32'b00000000000000000001000100110100;
assign LUT_4[40229] = 32'b11111111111111111010010000101100;
assign LUT_4[40230] = 32'b00000000000000000000011111011000;
assign LUT_4[40231] = 32'b11111111111111111001101011010000;
assign LUT_4[40232] = 32'b11111111111111111101010000101101;
assign LUT_4[40233] = 32'b11111111111111110110011100100101;
assign LUT_4[40234] = 32'b11111111111111111100101011010001;
assign LUT_4[40235] = 32'b11111111111111110101110111001001;
assign LUT_4[40236] = 32'b11111111111111111010010001001001;
assign LUT_4[40237] = 32'b11111111111111110011011101000001;
assign LUT_4[40238] = 32'b11111111111111111001101011101101;
assign LUT_4[40239] = 32'b11111111111111110010110111100101;
assign LUT_4[40240] = 32'b00000000000000000001110110000110;
assign LUT_4[40241] = 32'b11111111111111111011000001111110;
assign LUT_4[40242] = 32'b00000000000000000001010000101010;
assign LUT_4[40243] = 32'b11111111111111111010011100100010;
assign LUT_4[40244] = 32'b11111111111111111110110110100010;
assign LUT_4[40245] = 32'b11111111111111111000000010011010;
assign LUT_4[40246] = 32'b11111111111111111110010001000110;
assign LUT_4[40247] = 32'b11111111111111110111011100111110;
assign LUT_4[40248] = 32'b11111111111111111011000010011011;
assign LUT_4[40249] = 32'b11111111111111110100001110010011;
assign LUT_4[40250] = 32'b11111111111111111010011100111111;
assign LUT_4[40251] = 32'b11111111111111110011101000110111;
assign LUT_4[40252] = 32'b11111111111111111000000010110111;
assign LUT_4[40253] = 32'b11111111111111110001001110101111;
assign LUT_4[40254] = 32'b11111111111111110111011101011011;
assign LUT_4[40255] = 32'b11111111111111110000101001010011;
assign LUT_4[40256] = 32'b00000000000000000111000000100101;
assign LUT_4[40257] = 32'b00000000000000000000001100011101;
assign LUT_4[40258] = 32'b00000000000000000110011011001001;
assign LUT_4[40259] = 32'b11111111111111111111100111000001;
assign LUT_4[40260] = 32'b00000000000000000100000001000001;
assign LUT_4[40261] = 32'b11111111111111111101001100111001;
assign LUT_4[40262] = 32'b00000000000000000011011011100101;
assign LUT_4[40263] = 32'b11111111111111111100100111011101;
assign LUT_4[40264] = 32'b00000000000000000000001100111010;
assign LUT_4[40265] = 32'b11111111111111111001011000110010;
assign LUT_4[40266] = 32'b11111111111111111111100111011110;
assign LUT_4[40267] = 32'b11111111111111111000110011010110;
assign LUT_4[40268] = 32'b11111111111111111101001101010110;
assign LUT_4[40269] = 32'b11111111111111110110011001001110;
assign LUT_4[40270] = 32'b11111111111111111100100111111010;
assign LUT_4[40271] = 32'b11111111111111110101110011110010;
assign LUT_4[40272] = 32'b00000000000000000100110010010011;
assign LUT_4[40273] = 32'b11111111111111111101111110001011;
assign LUT_4[40274] = 32'b00000000000000000100001100110111;
assign LUT_4[40275] = 32'b11111111111111111101011000101111;
assign LUT_4[40276] = 32'b00000000000000000001110010101111;
assign LUT_4[40277] = 32'b11111111111111111010111110100111;
assign LUT_4[40278] = 32'b00000000000000000001001101010011;
assign LUT_4[40279] = 32'b11111111111111111010011001001011;
assign LUT_4[40280] = 32'b11111111111111111101111110101000;
assign LUT_4[40281] = 32'b11111111111111110111001010100000;
assign LUT_4[40282] = 32'b11111111111111111101011001001100;
assign LUT_4[40283] = 32'b11111111111111110110100101000100;
assign LUT_4[40284] = 32'b11111111111111111010111111000100;
assign LUT_4[40285] = 32'b11111111111111110100001010111100;
assign LUT_4[40286] = 32'b11111111111111111010011001101000;
assign LUT_4[40287] = 32'b11111111111111110011100101100000;
assign LUT_4[40288] = 32'b00000000000000000101011011101100;
assign LUT_4[40289] = 32'b11111111111111111110100111100100;
assign LUT_4[40290] = 32'b00000000000000000100110110010000;
assign LUT_4[40291] = 32'b11111111111111111110000010001000;
assign LUT_4[40292] = 32'b00000000000000000010011100001000;
assign LUT_4[40293] = 32'b11111111111111111011101000000000;
assign LUT_4[40294] = 32'b00000000000000000001110110101100;
assign LUT_4[40295] = 32'b11111111111111111011000010100100;
assign LUT_4[40296] = 32'b11111111111111111110101000000001;
assign LUT_4[40297] = 32'b11111111111111110111110011111001;
assign LUT_4[40298] = 32'b11111111111111111110000010100101;
assign LUT_4[40299] = 32'b11111111111111110111001110011101;
assign LUT_4[40300] = 32'b11111111111111111011101000011101;
assign LUT_4[40301] = 32'b11111111111111110100110100010101;
assign LUT_4[40302] = 32'b11111111111111111011000011000001;
assign LUT_4[40303] = 32'b11111111111111110100001110111001;
assign LUT_4[40304] = 32'b00000000000000000011001101011010;
assign LUT_4[40305] = 32'b11111111111111111100011001010010;
assign LUT_4[40306] = 32'b00000000000000000010100111111110;
assign LUT_4[40307] = 32'b11111111111111111011110011110110;
assign LUT_4[40308] = 32'b00000000000000000000001101110110;
assign LUT_4[40309] = 32'b11111111111111111001011001101110;
assign LUT_4[40310] = 32'b11111111111111111111101000011010;
assign LUT_4[40311] = 32'b11111111111111111000110100010010;
assign LUT_4[40312] = 32'b11111111111111111100011001101111;
assign LUT_4[40313] = 32'b11111111111111110101100101100111;
assign LUT_4[40314] = 32'b11111111111111111011110100010011;
assign LUT_4[40315] = 32'b11111111111111110101000000001011;
assign LUT_4[40316] = 32'b11111111111111111001011010001011;
assign LUT_4[40317] = 32'b11111111111111110010100110000011;
assign LUT_4[40318] = 32'b11111111111111111000110100101111;
assign LUT_4[40319] = 32'b11111111111111110010000000100111;
assign LUT_4[40320] = 32'b00000000000000001000001111011001;
assign LUT_4[40321] = 32'b00000000000000000001011011010001;
assign LUT_4[40322] = 32'b00000000000000000111101001111101;
assign LUT_4[40323] = 32'b00000000000000000000110101110101;
assign LUT_4[40324] = 32'b00000000000000000101001111110101;
assign LUT_4[40325] = 32'b11111111111111111110011011101101;
assign LUT_4[40326] = 32'b00000000000000000100101010011001;
assign LUT_4[40327] = 32'b11111111111111111101110110010001;
assign LUT_4[40328] = 32'b00000000000000000001011011101110;
assign LUT_4[40329] = 32'b11111111111111111010100111100110;
assign LUT_4[40330] = 32'b00000000000000000000110110010010;
assign LUT_4[40331] = 32'b11111111111111111010000010001010;
assign LUT_4[40332] = 32'b11111111111111111110011100001010;
assign LUT_4[40333] = 32'b11111111111111110111101000000010;
assign LUT_4[40334] = 32'b11111111111111111101110110101110;
assign LUT_4[40335] = 32'b11111111111111110111000010100110;
assign LUT_4[40336] = 32'b00000000000000000110000001000111;
assign LUT_4[40337] = 32'b11111111111111111111001100111111;
assign LUT_4[40338] = 32'b00000000000000000101011011101011;
assign LUT_4[40339] = 32'b11111111111111111110100111100011;
assign LUT_4[40340] = 32'b00000000000000000011000001100011;
assign LUT_4[40341] = 32'b11111111111111111100001101011011;
assign LUT_4[40342] = 32'b00000000000000000010011100000111;
assign LUT_4[40343] = 32'b11111111111111111011100111111111;
assign LUT_4[40344] = 32'b11111111111111111111001101011100;
assign LUT_4[40345] = 32'b11111111111111111000011001010100;
assign LUT_4[40346] = 32'b11111111111111111110101000000000;
assign LUT_4[40347] = 32'b11111111111111110111110011111000;
assign LUT_4[40348] = 32'b11111111111111111100001101111000;
assign LUT_4[40349] = 32'b11111111111111110101011001110000;
assign LUT_4[40350] = 32'b11111111111111111011101000011100;
assign LUT_4[40351] = 32'b11111111111111110100110100010100;
assign LUT_4[40352] = 32'b00000000000000000110101010100000;
assign LUT_4[40353] = 32'b11111111111111111111110110011000;
assign LUT_4[40354] = 32'b00000000000000000110000101000100;
assign LUT_4[40355] = 32'b11111111111111111111010000111100;
assign LUT_4[40356] = 32'b00000000000000000011101010111100;
assign LUT_4[40357] = 32'b11111111111111111100110110110100;
assign LUT_4[40358] = 32'b00000000000000000011000101100000;
assign LUT_4[40359] = 32'b11111111111111111100010001011000;
assign LUT_4[40360] = 32'b11111111111111111111110110110101;
assign LUT_4[40361] = 32'b11111111111111111001000010101101;
assign LUT_4[40362] = 32'b11111111111111111111010001011001;
assign LUT_4[40363] = 32'b11111111111111111000011101010001;
assign LUT_4[40364] = 32'b11111111111111111100110111010001;
assign LUT_4[40365] = 32'b11111111111111110110000011001001;
assign LUT_4[40366] = 32'b11111111111111111100010001110101;
assign LUT_4[40367] = 32'b11111111111111110101011101101101;
assign LUT_4[40368] = 32'b00000000000000000100011100001110;
assign LUT_4[40369] = 32'b11111111111111111101101000000110;
assign LUT_4[40370] = 32'b00000000000000000011110110110010;
assign LUT_4[40371] = 32'b11111111111111111101000010101010;
assign LUT_4[40372] = 32'b00000000000000000001011100101010;
assign LUT_4[40373] = 32'b11111111111111111010101000100010;
assign LUT_4[40374] = 32'b00000000000000000000110111001110;
assign LUT_4[40375] = 32'b11111111111111111010000011000110;
assign LUT_4[40376] = 32'b11111111111111111101101000100011;
assign LUT_4[40377] = 32'b11111111111111110110110100011011;
assign LUT_4[40378] = 32'b11111111111111111101000011000111;
assign LUT_4[40379] = 32'b11111111111111110110001110111111;
assign LUT_4[40380] = 32'b11111111111111111010101000111111;
assign LUT_4[40381] = 32'b11111111111111110011110100110111;
assign LUT_4[40382] = 32'b11111111111111111010000011100011;
assign LUT_4[40383] = 32'b11111111111111110011001111011011;
assign LUT_4[40384] = 32'b00000000000000001001100110101101;
assign LUT_4[40385] = 32'b00000000000000000010110010100101;
assign LUT_4[40386] = 32'b00000000000000001001000001010001;
assign LUT_4[40387] = 32'b00000000000000000010001101001001;
assign LUT_4[40388] = 32'b00000000000000000110100111001001;
assign LUT_4[40389] = 32'b11111111111111111111110011000001;
assign LUT_4[40390] = 32'b00000000000000000110000001101101;
assign LUT_4[40391] = 32'b11111111111111111111001101100101;
assign LUT_4[40392] = 32'b00000000000000000010110011000010;
assign LUT_4[40393] = 32'b11111111111111111011111110111010;
assign LUT_4[40394] = 32'b00000000000000000010001101100110;
assign LUT_4[40395] = 32'b11111111111111111011011001011110;
assign LUT_4[40396] = 32'b11111111111111111111110011011110;
assign LUT_4[40397] = 32'b11111111111111111000111111010110;
assign LUT_4[40398] = 32'b11111111111111111111001110000010;
assign LUT_4[40399] = 32'b11111111111111111000011001111010;
assign LUT_4[40400] = 32'b00000000000000000111011000011011;
assign LUT_4[40401] = 32'b00000000000000000000100100010011;
assign LUT_4[40402] = 32'b00000000000000000110110010111111;
assign LUT_4[40403] = 32'b11111111111111111111111110110111;
assign LUT_4[40404] = 32'b00000000000000000100011000110111;
assign LUT_4[40405] = 32'b11111111111111111101100100101111;
assign LUT_4[40406] = 32'b00000000000000000011110011011011;
assign LUT_4[40407] = 32'b11111111111111111100111111010011;
assign LUT_4[40408] = 32'b00000000000000000000100100110000;
assign LUT_4[40409] = 32'b11111111111111111001110000101000;
assign LUT_4[40410] = 32'b11111111111111111111111111010100;
assign LUT_4[40411] = 32'b11111111111111111001001011001100;
assign LUT_4[40412] = 32'b11111111111111111101100101001100;
assign LUT_4[40413] = 32'b11111111111111110110110001000100;
assign LUT_4[40414] = 32'b11111111111111111100111111110000;
assign LUT_4[40415] = 32'b11111111111111110110001011101000;
assign LUT_4[40416] = 32'b00000000000000001000000001110100;
assign LUT_4[40417] = 32'b00000000000000000001001101101100;
assign LUT_4[40418] = 32'b00000000000000000111011100011000;
assign LUT_4[40419] = 32'b00000000000000000000101000010000;
assign LUT_4[40420] = 32'b00000000000000000101000010010000;
assign LUT_4[40421] = 32'b11111111111111111110001110001000;
assign LUT_4[40422] = 32'b00000000000000000100011100110100;
assign LUT_4[40423] = 32'b11111111111111111101101000101100;
assign LUT_4[40424] = 32'b00000000000000000001001110001001;
assign LUT_4[40425] = 32'b11111111111111111010011010000001;
assign LUT_4[40426] = 32'b00000000000000000000101000101101;
assign LUT_4[40427] = 32'b11111111111111111001110100100101;
assign LUT_4[40428] = 32'b11111111111111111110001110100101;
assign LUT_4[40429] = 32'b11111111111111110111011010011101;
assign LUT_4[40430] = 32'b11111111111111111101101001001001;
assign LUT_4[40431] = 32'b11111111111111110110110101000001;
assign LUT_4[40432] = 32'b00000000000000000101110011100010;
assign LUT_4[40433] = 32'b11111111111111111110111111011010;
assign LUT_4[40434] = 32'b00000000000000000101001110000110;
assign LUT_4[40435] = 32'b11111111111111111110011001111110;
assign LUT_4[40436] = 32'b00000000000000000010110011111110;
assign LUT_4[40437] = 32'b11111111111111111011111111110110;
assign LUT_4[40438] = 32'b00000000000000000010001110100010;
assign LUT_4[40439] = 32'b11111111111111111011011010011010;
assign LUT_4[40440] = 32'b11111111111111111110111111110111;
assign LUT_4[40441] = 32'b11111111111111111000001011101111;
assign LUT_4[40442] = 32'b11111111111111111110011010011011;
assign LUT_4[40443] = 32'b11111111111111110111100110010011;
assign LUT_4[40444] = 32'b11111111111111111100000000010011;
assign LUT_4[40445] = 32'b11111111111111110101001100001011;
assign LUT_4[40446] = 32'b11111111111111111011011010110111;
assign LUT_4[40447] = 32'b11111111111111110100100110101111;
assign LUT_4[40448] = 32'b11111111111111111111110001110110;
assign LUT_4[40449] = 32'b11111111111111111000111101101110;
assign LUT_4[40450] = 32'b11111111111111111111001100011010;
assign LUT_4[40451] = 32'b11111111111111111000011000010010;
assign LUT_4[40452] = 32'b11111111111111111100110010010010;
assign LUT_4[40453] = 32'b11111111111111110101111110001010;
assign LUT_4[40454] = 32'b11111111111111111100001100110110;
assign LUT_4[40455] = 32'b11111111111111110101011000101110;
assign LUT_4[40456] = 32'b11111111111111111000111110001011;
assign LUT_4[40457] = 32'b11111111111111110010001010000011;
assign LUT_4[40458] = 32'b11111111111111111000011000101111;
assign LUT_4[40459] = 32'b11111111111111110001100100100111;
assign LUT_4[40460] = 32'b11111111111111110101111110100111;
assign LUT_4[40461] = 32'b11111111111111101111001010011111;
assign LUT_4[40462] = 32'b11111111111111110101011001001011;
assign LUT_4[40463] = 32'b11111111111111101110100101000011;
assign LUT_4[40464] = 32'b11111111111111111101100011100100;
assign LUT_4[40465] = 32'b11111111111111110110101111011100;
assign LUT_4[40466] = 32'b11111111111111111100111110001000;
assign LUT_4[40467] = 32'b11111111111111110110001010000000;
assign LUT_4[40468] = 32'b11111111111111111010100100000000;
assign LUT_4[40469] = 32'b11111111111111110011101111111000;
assign LUT_4[40470] = 32'b11111111111111111001111110100100;
assign LUT_4[40471] = 32'b11111111111111110011001010011100;
assign LUT_4[40472] = 32'b11111111111111110110101111111001;
assign LUT_4[40473] = 32'b11111111111111101111111011110001;
assign LUT_4[40474] = 32'b11111111111111110110001010011101;
assign LUT_4[40475] = 32'b11111111111111101111010110010101;
assign LUT_4[40476] = 32'b11111111111111110011110000010101;
assign LUT_4[40477] = 32'b11111111111111101100111100001101;
assign LUT_4[40478] = 32'b11111111111111110011001010111001;
assign LUT_4[40479] = 32'b11111111111111101100010110110001;
assign LUT_4[40480] = 32'b11111111111111111110001100111101;
assign LUT_4[40481] = 32'b11111111111111110111011000110101;
assign LUT_4[40482] = 32'b11111111111111111101100111100001;
assign LUT_4[40483] = 32'b11111111111111110110110011011001;
assign LUT_4[40484] = 32'b11111111111111111011001101011001;
assign LUT_4[40485] = 32'b11111111111111110100011001010001;
assign LUT_4[40486] = 32'b11111111111111111010100111111101;
assign LUT_4[40487] = 32'b11111111111111110011110011110101;
assign LUT_4[40488] = 32'b11111111111111110111011001010010;
assign LUT_4[40489] = 32'b11111111111111110000100101001010;
assign LUT_4[40490] = 32'b11111111111111110110110011110110;
assign LUT_4[40491] = 32'b11111111111111101111111111101110;
assign LUT_4[40492] = 32'b11111111111111110100011001101110;
assign LUT_4[40493] = 32'b11111111111111101101100101100110;
assign LUT_4[40494] = 32'b11111111111111110011110100010010;
assign LUT_4[40495] = 32'b11111111111111101101000000001010;
assign LUT_4[40496] = 32'b11111111111111111011111110101011;
assign LUT_4[40497] = 32'b11111111111111110101001010100011;
assign LUT_4[40498] = 32'b11111111111111111011011001001111;
assign LUT_4[40499] = 32'b11111111111111110100100101000111;
assign LUT_4[40500] = 32'b11111111111111111000111111000111;
assign LUT_4[40501] = 32'b11111111111111110010001010111111;
assign LUT_4[40502] = 32'b11111111111111111000011001101011;
assign LUT_4[40503] = 32'b11111111111111110001100101100011;
assign LUT_4[40504] = 32'b11111111111111110101001011000000;
assign LUT_4[40505] = 32'b11111111111111101110010110111000;
assign LUT_4[40506] = 32'b11111111111111110100100101100100;
assign LUT_4[40507] = 32'b11111111111111101101110001011100;
assign LUT_4[40508] = 32'b11111111111111110010001011011100;
assign LUT_4[40509] = 32'b11111111111111101011010111010100;
assign LUT_4[40510] = 32'b11111111111111110001100110000000;
assign LUT_4[40511] = 32'b11111111111111101010110001111000;
assign LUT_4[40512] = 32'b00000000000000000001001001001010;
assign LUT_4[40513] = 32'b11111111111111111010010101000010;
assign LUT_4[40514] = 32'b00000000000000000000100011101110;
assign LUT_4[40515] = 32'b11111111111111111001101111100110;
assign LUT_4[40516] = 32'b11111111111111111110001001100110;
assign LUT_4[40517] = 32'b11111111111111110111010101011110;
assign LUT_4[40518] = 32'b11111111111111111101100100001010;
assign LUT_4[40519] = 32'b11111111111111110110110000000010;
assign LUT_4[40520] = 32'b11111111111111111010010101011111;
assign LUT_4[40521] = 32'b11111111111111110011100001010111;
assign LUT_4[40522] = 32'b11111111111111111001110000000011;
assign LUT_4[40523] = 32'b11111111111111110010111011111011;
assign LUT_4[40524] = 32'b11111111111111110111010101111011;
assign LUT_4[40525] = 32'b11111111111111110000100001110011;
assign LUT_4[40526] = 32'b11111111111111110110110000011111;
assign LUT_4[40527] = 32'b11111111111111101111111100010111;
assign LUT_4[40528] = 32'b11111111111111111110111010111000;
assign LUT_4[40529] = 32'b11111111111111111000000110110000;
assign LUT_4[40530] = 32'b11111111111111111110010101011100;
assign LUT_4[40531] = 32'b11111111111111110111100001010100;
assign LUT_4[40532] = 32'b11111111111111111011111011010100;
assign LUT_4[40533] = 32'b11111111111111110101000111001100;
assign LUT_4[40534] = 32'b11111111111111111011010101111000;
assign LUT_4[40535] = 32'b11111111111111110100100001110000;
assign LUT_4[40536] = 32'b11111111111111111000000111001101;
assign LUT_4[40537] = 32'b11111111111111110001010011000101;
assign LUT_4[40538] = 32'b11111111111111110111100001110001;
assign LUT_4[40539] = 32'b11111111111111110000101101101001;
assign LUT_4[40540] = 32'b11111111111111110101000111101001;
assign LUT_4[40541] = 32'b11111111111111101110010011100001;
assign LUT_4[40542] = 32'b11111111111111110100100010001101;
assign LUT_4[40543] = 32'b11111111111111101101101110000101;
assign LUT_4[40544] = 32'b11111111111111111111100100010001;
assign LUT_4[40545] = 32'b11111111111111111000110000001001;
assign LUT_4[40546] = 32'b11111111111111111110111110110101;
assign LUT_4[40547] = 32'b11111111111111111000001010101101;
assign LUT_4[40548] = 32'b11111111111111111100100100101101;
assign LUT_4[40549] = 32'b11111111111111110101110000100101;
assign LUT_4[40550] = 32'b11111111111111111011111111010001;
assign LUT_4[40551] = 32'b11111111111111110101001011001001;
assign LUT_4[40552] = 32'b11111111111111111000110000100110;
assign LUT_4[40553] = 32'b11111111111111110001111100011110;
assign LUT_4[40554] = 32'b11111111111111111000001011001010;
assign LUT_4[40555] = 32'b11111111111111110001010111000010;
assign LUT_4[40556] = 32'b11111111111111110101110001000010;
assign LUT_4[40557] = 32'b11111111111111101110111100111010;
assign LUT_4[40558] = 32'b11111111111111110101001011100110;
assign LUT_4[40559] = 32'b11111111111111101110010111011110;
assign LUT_4[40560] = 32'b11111111111111111101010101111111;
assign LUT_4[40561] = 32'b11111111111111110110100001110111;
assign LUT_4[40562] = 32'b11111111111111111100110000100011;
assign LUT_4[40563] = 32'b11111111111111110101111100011011;
assign LUT_4[40564] = 32'b11111111111111111010010110011011;
assign LUT_4[40565] = 32'b11111111111111110011100010010011;
assign LUT_4[40566] = 32'b11111111111111111001110000111111;
assign LUT_4[40567] = 32'b11111111111111110010111100110111;
assign LUT_4[40568] = 32'b11111111111111110110100010010100;
assign LUT_4[40569] = 32'b11111111111111101111101110001100;
assign LUT_4[40570] = 32'b11111111111111110101111100111000;
assign LUT_4[40571] = 32'b11111111111111101111001000110000;
assign LUT_4[40572] = 32'b11111111111111110011100010110000;
assign LUT_4[40573] = 32'b11111111111111101100101110101000;
assign LUT_4[40574] = 32'b11111111111111110010111101010100;
assign LUT_4[40575] = 32'b11111111111111101100001001001100;
assign LUT_4[40576] = 32'b00000000000000000010010111111110;
assign LUT_4[40577] = 32'b11111111111111111011100011110110;
assign LUT_4[40578] = 32'b00000000000000000001110010100010;
assign LUT_4[40579] = 32'b11111111111111111010111110011010;
assign LUT_4[40580] = 32'b11111111111111111111011000011010;
assign LUT_4[40581] = 32'b11111111111111111000100100010010;
assign LUT_4[40582] = 32'b11111111111111111110110010111110;
assign LUT_4[40583] = 32'b11111111111111110111111110110110;
assign LUT_4[40584] = 32'b11111111111111111011100100010011;
assign LUT_4[40585] = 32'b11111111111111110100110000001011;
assign LUT_4[40586] = 32'b11111111111111111010111110110111;
assign LUT_4[40587] = 32'b11111111111111110100001010101111;
assign LUT_4[40588] = 32'b11111111111111111000100100101111;
assign LUT_4[40589] = 32'b11111111111111110001110000100111;
assign LUT_4[40590] = 32'b11111111111111110111111111010011;
assign LUT_4[40591] = 32'b11111111111111110001001011001011;
assign LUT_4[40592] = 32'b00000000000000000000001001101100;
assign LUT_4[40593] = 32'b11111111111111111001010101100100;
assign LUT_4[40594] = 32'b11111111111111111111100100010000;
assign LUT_4[40595] = 32'b11111111111111111000110000001000;
assign LUT_4[40596] = 32'b11111111111111111101001010001000;
assign LUT_4[40597] = 32'b11111111111111110110010110000000;
assign LUT_4[40598] = 32'b11111111111111111100100100101100;
assign LUT_4[40599] = 32'b11111111111111110101110000100100;
assign LUT_4[40600] = 32'b11111111111111111001010110000001;
assign LUT_4[40601] = 32'b11111111111111110010100001111001;
assign LUT_4[40602] = 32'b11111111111111111000110000100101;
assign LUT_4[40603] = 32'b11111111111111110001111100011101;
assign LUT_4[40604] = 32'b11111111111111110110010110011101;
assign LUT_4[40605] = 32'b11111111111111101111100010010101;
assign LUT_4[40606] = 32'b11111111111111110101110001000001;
assign LUT_4[40607] = 32'b11111111111111101110111100111001;
assign LUT_4[40608] = 32'b00000000000000000000110011000101;
assign LUT_4[40609] = 32'b11111111111111111001111110111101;
assign LUT_4[40610] = 32'b00000000000000000000001101101001;
assign LUT_4[40611] = 32'b11111111111111111001011001100001;
assign LUT_4[40612] = 32'b11111111111111111101110011100001;
assign LUT_4[40613] = 32'b11111111111111110110111111011001;
assign LUT_4[40614] = 32'b11111111111111111101001110000101;
assign LUT_4[40615] = 32'b11111111111111110110011001111101;
assign LUT_4[40616] = 32'b11111111111111111001111111011010;
assign LUT_4[40617] = 32'b11111111111111110011001011010010;
assign LUT_4[40618] = 32'b11111111111111111001011001111110;
assign LUT_4[40619] = 32'b11111111111111110010100101110110;
assign LUT_4[40620] = 32'b11111111111111110110111111110110;
assign LUT_4[40621] = 32'b11111111111111110000001011101110;
assign LUT_4[40622] = 32'b11111111111111110110011010011010;
assign LUT_4[40623] = 32'b11111111111111101111100110010010;
assign LUT_4[40624] = 32'b11111111111111111110100100110011;
assign LUT_4[40625] = 32'b11111111111111110111110000101011;
assign LUT_4[40626] = 32'b11111111111111111101111111010111;
assign LUT_4[40627] = 32'b11111111111111110111001011001111;
assign LUT_4[40628] = 32'b11111111111111111011100101001111;
assign LUT_4[40629] = 32'b11111111111111110100110001000111;
assign LUT_4[40630] = 32'b11111111111111111010111111110011;
assign LUT_4[40631] = 32'b11111111111111110100001011101011;
assign LUT_4[40632] = 32'b11111111111111110111110001001000;
assign LUT_4[40633] = 32'b11111111111111110000111101000000;
assign LUT_4[40634] = 32'b11111111111111110111001011101100;
assign LUT_4[40635] = 32'b11111111111111110000010111100100;
assign LUT_4[40636] = 32'b11111111111111110100110001100100;
assign LUT_4[40637] = 32'b11111111111111101101111101011100;
assign LUT_4[40638] = 32'b11111111111111110100001100001000;
assign LUT_4[40639] = 32'b11111111111111101101011000000000;
assign LUT_4[40640] = 32'b00000000000000000011101111010010;
assign LUT_4[40641] = 32'b11111111111111111100111011001010;
assign LUT_4[40642] = 32'b00000000000000000011001001110110;
assign LUT_4[40643] = 32'b11111111111111111100010101101110;
assign LUT_4[40644] = 32'b00000000000000000000101111101110;
assign LUT_4[40645] = 32'b11111111111111111001111011100110;
assign LUT_4[40646] = 32'b00000000000000000000001010010010;
assign LUT_4[40647] = 32'b11111111111111111001010110001010;
assign LUT_4[40648] = 32'b11111111111111111100111011100111;
assign LUT_4[40649] = 32'b11111111111111110110000111011111;
assign LUT_4[40650] = 32'b11111111111111111100010110001011;
assign LUT_4[40651] = 32'b11111111111111110101100010000011;
assign LUT_4[40652] = 32'b11111111111111111001111100000011;
assign LUT_4[40653] = 32'b11111111111111110011000111111011;
assign LUT_4[40654] = 32'b11111111111111111001010110100111;
assign LUT_4[40655] = 32'b11111111111111110010100010011111;
assign LUT_4[40656] = 32'b00000000000000000001100001000000;
assign LUT_4[40657] = 32'b11111111111111111010101100111000;
assign LUT_4[40658] = 32'b00000000000000000000111011100100;
assign LUT_4[40659] = 32'b11111111111111111010000111011100;
assign LUT_4[40660] = 32'b11111111111111111110100001011100;
assign LUT_4[40661] = 32'b11111111111111110111101101010100;
assign LUT_4[40662] = 32'b11111111111111111101111100000000;
assign LUT_4[40663] = 32'b11111111111111110111000111111000;
assign LUT_4[40664] = 32'b11111111111111111010101101010101;
assign LUT_4[40665] = 32'b11111111111111110011111001001101;
assign LUT_4[40666] = 32'b11111111111111111010000111111001;
assign LUT_4[40667] = 32'b11111111111111110011010011110001;
assign LUT_4[40668] = 32'b11111111111111110111101101110001;
assign LUT_4[40669] = 32'b11111111111111110000111001101001;
assign LUT_4[40670] = 32'b11111111111111110111001000010101;
assign LUT_4[40671] = 32'b11111111111111110000010100001101;
assign LUT_4[40672] = 32'b00000000000000000010001010011001;
assign LUT_4[40673] = 32'b11111111111111111011010110010001;
assign LUT_4[40674] = 32'b00000000000000000001100100111101;
assign LUT_4[40675] = 32'b11111111111111111010110000110101;
assign LUT_4[40676] = 32'b11111111111111111111001010110101;
assign LUT_4[40677] = 32'b11111111111111111000010110101101;
assign LUT_4[40678] = 32'b11111111111111111110100101011001;
assign LUT_4[40679] = 32'b11111111111111110111110001010001;
assign LUT_4[40680] = 32'b11111111111111111011010110101110;
assign LUT_4[40681] = 32'b11111111111111110100100010100110;
assign LUT_4[40682] = 32'b11111111111111111010110001010010;
assign LUT_4[40683] = 32'b11111111111111110011111101001010;
assign LUT_4[40684] = 32'b11111111111111111000010111001010;
assign LUT_4[40685] = 32'b11111111111111110001100011000010;
assign LUT_4[40686] = 32'b11111111111111110111110001101110;
assign LUT_4[40687] = 32'b11111111111111110000111101100110;
assign LUT_4[40688] = 32'b11111111111111111111111100000111;
assign LUT_4[40689] = 32'b11111111111111111001000111111111;
assign LUT_4[40690] = 32'b11111111111111111111010110101011;
assign LUT_4[40691] = 32'b11111111111111111000100010100011;
assign LUT_4[40692] = 32'b11111111111111111100111100100011;
assign LUT_4[40693] = 32'b11111111111111110110001000011011;
assign LUT_4[40694] = 32'b11111111111111111100010111000111;
assign LUT_4[40695] = 32'b11111111111111110101100010111111;
assign LUT_4[40696] = 32'b11111111111111111001001000011100;
assign LUT_4[40697] = 32'b11111111111111110010010100010100;
assign LUT_4[40698] = 32'b11111111111111111000100011000000;
assign LUT_4[40699] = 32'b11111111111111110001101110111000;
assign LUT_4[40700] = 32'b11111111111111110110001000111000;
assign LUT_4[40701] = 32'b11111111111111101111010100110000;
assign LUT_4[40702] = 32'b11111111111111110101100011011100;
assign LUT_4[40703] = 32'b11111111111111101110101111010100;
assign LUT_4[40704] = 32'b00000000000000000100101101011001;
assign LUT_4[40705] = 32'b11111111111111111101111001010001;
assign LUT_4[40706] = 32'b00000000000000000100000111111101;
assign LUT_4[40707] = 32'b11111111111111111101010011110101;
assign LUT_4[40708] = 32'b00000000000000000001101101110101;
assign LUT_4[40709] = 32'b11111111111111111010111001101101;
assign LUT_4[40710] = 32'b00000000000000000001001000011001;
assign LUT_4[40711] = 32'b11111111111111111010010100010001;
assign LUT_4[40712] = 32'b11111111111111111101111001101110;
assign LUT_4[40713] = 32'b11111111111111110111000101100110;
assign LUT_4[40714] = 32'b11111111111111111101010100010010;
assign LUT_4[40715] = 32'b11111111111111110110100000001010;
assign LUT_4[40716] = 32'b11111111111111111010111010001010;
assign LUT_4[40717] = 32'b11111111111111110100000110000010;
assign LUT_4[40718] = 32'b11111111111111111010010100101110;
assign LUT_4[40719] = 32'b11111111111111110011100000100110;
assign LUT_4[40720] = 32'b00000000000000000010011111000111;
assign LUT_4[40721] = 32'b11111111111111111011101010111111;
assign LUT_4[40722] = 32'b00000000000000000001111001101011;
assign LUT_4[40723] = 32'b11111111111111111011000101100011;
assign LUT_4[40724] = 32'b11111111111111111111011111100011;
assign LUT_4[40725] = 32'b11111111111111111000101011011011;
assign LUT_4[40726] = 32'b11111111111111111110111010000111;
assign LUT_4[40727] = 32'b11111111111111111000000101111111;
assign LUT_4[40728] = 32'b11111111111111111011101011011100;
assign LUT_4[40729] = 32'b11111111111111110100110111010100;
assign LUT_4[40730] = 32'b11111111111111111011000110000000;
assign LUT_4[40731] = 32'b11111111111111110100010001111000;
assign LUT_4[40732] = 32'b11111111111111111000101011111000;
assign LUT_4[40733] = 32'b11111111111111110001110111110000;
assign LUT_4[40734] = 32'b11111111111111111000000110011100;
assign LUT_4[40735] = 32'b11111111111111110001010010010100;
assign LUT_4[40736] = 32'b00000000000000000011001000100000;
assign LUT_4[40737] = 32'b11111111111111111100010100011000;
assign LUT_4[40738] = 32'b00000000000000000010100011000100;
assign LUT_4[40739] = 32'b11111111111111111011101110111100;
assign LUT_4[40740] = 32'b00000000000000000000001000111100;
assign LUT_4[40741] = 32'b11111111111111111001010100110100;
assign LUT_4[40742] = 32'b11111111111111111111100011100000;
assign LUT_4[40743] = 32'b11111111111111111000101111011000;
assign LUT_4[40744] = 32'b11111111111111111100010100110101;
assign LUT_4[40745] = 32'b11111111111111110101100000101101;
assign LUT_4[40746] = 32'b11111111111111111011101111011001;
assign LUT_4[40747] = 32'b11111111111111110100111011010001;
assign LUT_4[40748] = 32'b11111111111111111001010101010001;
assign LUT_4[40749] = 32'b11111111111111110010100001001001;
assign LUT_4[40750] = 32'b11111111111111111000101111110101;
assign LUT_4[40751] = 32'b11111111111111110001111011101101;
assign LUT_4[40752] = 32'b00000000000000000000111010001110;
assign LUT_4[40753] = 32'b11111111111111111010000110000110;
assign LUT_4[40754] = 32'b00000000000000000000010100110010;
assign LUT_4[40755] = 32'b11111111111111111001100000101010;
assign LUT_4[40756] = 32'b11111111111111111101111010101010;
assign LUT_4[40757] = 32'b11111111111111110111000110100010;
assign LUT_4[40758] = 32'b11111111111111111101010101001110;
assign LUT_4[40759] = 32'b11111111111111110110100001000110;
assign LUT_4[40760] = 32'b11111111111111111010000110100011;
assign LUT_4[40761] = 32'b11111111111111110011010010011011;
assign LUT_4[40762] = 32'b11111111111111111001100001000111;
assign LUT_4[40763] = 32'b11111111111111110010101100111111;
assign LUT_4[40764] = 32'b11111111111111110111000110111111;
assign LUT_4[40765] = 32'b11111111111111110000010010110111;
assign LUT_4[40766] = 32'b11111111111111110110100001100011;
assign LUT_4[40767] = 32'b11111111111111101111101101011011;
assign LUT_4[40768] = 32'b00000000000000000110000100101101;
assign LUT_4[40769] = 32'b11111111111111111111010000100101;
assign LUT_4[40770] = 32'b00000000000000000101011111010001;
assign LUT_4[40771] = 32'b11111111111111111110101011001001;
assign LUT_4[40772] = 32'b00000000000000000011000101001001;
assign LUT_4[40773] = 32'b11111111111111111100010001000001;
assign LUT_4[40774] = 32'b00000000000000000010011111101101;
assign LUT_4[40775] = 32'b11111111111111111011101011100101;
assign LUT_4[40776] = 32'b11111111111111111111010001000010;
assign LUT_4[40777] = 32'b11111111111111111000011100111010;
assign LUT_4[40778] = 32'b11111111111111111110101011100110;
assign LUT_4[40779] = 32'b11111111111111110111110111011110;
assign LUT_4[40780] = 32'b11111111111111111100010001011110;
assign LUT_4[40781] = 32'b11111111111111110101011101010110;
assign LUT_4[40782] = 32'b11111111111111111011101100000010;
assign LUT_4[40783] = 32'b11111111111111110100110111111010;
assign LUT_4[40784] = 32'b00000000000000000011110110011011;
assign LUT_4[40785] = 32'b11111111111111111101000010010011;
assign LUT_4[40786] = 32'b00000000000000000011010000111111;
assign LUT_4[40787] = 32'b11111111111111111100011100110111;
assign LUT_4[40788] = 32'b00000000000000000000110110110111;
assign LUT_4[40789] = 32'b11111111111111111010000010101111;
assign LUT_4[40790] = 32'b00000000000000000000010001011011;
assign LUT_4[40791] = 32'b11111111111111111001011101010011;
assign LUT_4[40792] = 32'b11111111111111111101000010110000;
assign LUT_4[40793] = 32'b11111111111111110110001110101000;
assign LUT_4[40794] = 32'b11111111111111111100011101010100;
assign LUT_4[40795] = 32'b11111111111111110101101001001100;
assign LUT_4[40796] = 32'b11111111111111111010000011001100;
assign LUT_4[40797] = 32'b11111111111111110011001111000100;
assign LUT_4[40798] = 32'b11111111111111111001011101110000;
assign LUT_4[40799] = 32'b11111111111111110010101001101000;
assign LUT_4[40800] = 32'b00000000000000000100011111110100;
assign LUT_4[40801] = 32'b11111111111111111101101011101100;
assign LUT_4[40802] = 32'b00000000000000000011111010011000;
assign LUT_4[40803] = 32'b11111111111111111101000110010000;
assign LUT_4[40804] = 32'b00000000000000000001100000010000;
assign LUT_4[40805] = 32'b11111111111111111010101100001000;
assign LUT_4[40806] = 32'b00000000000000000000111010110100;
assign LUT_4[40807] = 32'b11111111111111111010000110101100;
assign LUT_4[40808] = 32'b11111111111111111101101100001001;
assign LUT_4[40809] = 32'b11111111111111110110111000000001;
assign LUT_4[40810] = 32'b11111111111111111101000110101101;
assign LUT_4[40811] = 32'b11111111111111110110010010100101;
assign LUT_4[40812] = 32'b11111111111111111010101100100101;
assign LUT_4[40813] = 32'b11111111111111110011111000011101;
assign LUT_4[40814] = 32'b11111111111111111010000111001001;
assign LUT_4[40815] = 32'b11111111111111110011010011000001;
assign LUT_4[40816] = 32'b00000000000000000010010001100010;
assign LUT_4[40817] = 32'b11111111111111111011011101011010;
assign LUT_4[40818] = 32'b00000000000000000001101100000110;
assign LUT_4[40819] = 32'b11111111111111111010110111111110;
assign LUT_4[40820] = 32'b11111111111111111111010001111110;
assign LUT_4[40821] = 32'b11111111111111111000011101110110;
assign LUT_4[40822] = 32'b11111111111111111110101100100010;
assign LUT_4[40823] = 32'b11111111111111110111111000011010;
assign LUT_4[40824] = 32'b11111111111111111011011101110111;
assign LUT_4[40825] = 32'b11111111111111110100101001101111;
assign LUT_4[40826] = 32'b11111111111111111010111000011011;
assign LUT_4[40827] = 32'b11111111111111110100000100010011;
assign LUT_4[40828] = 32'b11111111111111111000011110010011;
assign LUT_4[40829] = 32'b11111111111111110001101010001011;
assign LUT_4[40830] = 32'b11111111111111110111111000110111;
assign LUT_4[40831] = 32'b11111111111111110001000100101111;
assign LUT_4[40832] = 32'b00000000000000000111010011100001;
assign LUT_4[40833] = 32'b00000000000000000000011111011001;
assign LUT_4[40834] = 32'b00000000000000000110101110000101;
assign LUT_4[40835] = 32'b11111111111111111111111001111101;
assign LUT_4[40836] = 32'b00000000000000000100010011111101;
assign LUT_4[40837] = 32'b11111111111111111101011111110101;
assign LUT_4[40838] = 32'b00000000000000000011101110100001;
assign LUT_4[40839] = 32'b11111111111111111100111010011001;
assign LUT_4[40840] = 32'b00000000000000000000011111110110;
assign LUT_4[40841] = 32'b11111111111111111001101011101110;
assign LUT_4[40842] = 32'b11111111111111111111111010011010;
assign LUT_4[40843] = 32'b11111111111111111001000110010010;
assign LUT_4[40844] = 32'b11111111111111111101100000010010;
assign LUT_4[40845] = 32'b11111111111111110110101100001010;
assign LUT_4[40846] = 32'b11111111111111111100111010110110;
assign LUT_4[40847] = 32'b11111111111111110110000110101110;
assign LUT_4[40848] = 32'b00000000000000000101000101001111;
assign LUT_4[40849] = 32'b11111111111111111110010001000111;
assign LUT_4[40850] = 32'b00000000000000000100011111110011;
assign LUT_4[40851] = 32'b11111111111111111101101011101011;
assign LUT_4[40852] = 32'b00000000000000000010000101101011;
assign LUT_4[40853] = 32'b11111111111111111011010001100011;
assign LUT_4[40854] = 32'b00000000000000000001100000001111;
assign LUT_4[40855] = 32'b11111111111111111010101100000111;
assign LUT_4[40856] = 32'b11111111111111111110010001100100;
assign LUT_4[40857] = 32'b11111111111111110111011101011100;
assign LUT_4[40858] = 32'b11111111111111111101101100001000;
assign LUT_4[40859] = 32'b11111111111111110110111000000000;
assign LUT_4[40860] = 32'b11111111111111111011010010000000;
assign LUT_4[40861] = 32'b11111111111111110100011101111000;
assign LUT_4[40862] = 32'b11111111111111111010101100100100;
assign LUT_4[40863] = 32'b11111111111111110011111000011100;
assign LUT_4[40864] = 32'b00000000000000000101101110101000;
assign LUT_4[40865] = 32'b11111111111111111110111010100000;
assign LUT_4[40866] = 32'b00000000000000000101001001001100;
assign LUT_4[40867] = 32'b11111111111111111110010101000100;
assign LUT_4[40868] = 32'b00000000000000000010101111000100;
assign LUT_4[40869] = 32'b11111111111111111011111010111100;
assign LUT_4[40870] = 32'b00000000000000000010001001101000;
assign LUT_4[40871] = 32'b11111111111111111011010101100000;
assign LUT_4[40872] = 32'b11111111111111111110111010111101;
assign LUT_4[40873] = 32'b11111111111111111000000110110101;
assign LUT_4[40874] = 32'b11111111111111111110010101100001;
assign LUT_4[40875] = 32'b11111111111111110111100001011001;
assign LUT_4[40876] = 32'b11111111111111111011111011011001;
assign LUT_4[40877] = 32'b11111111111111110101000111010001;
assign LUT_4[40878] = 32'b11111111111111111011010101111101;
assign LUT_4[40879] = 32'b11111111111111110100100001110101;
assign LUT_4[40880] = 32'b00000000000000000011100000010110;
assign LUT_4[40881] = 32'b11111111111111111100101100001110;
assign LUT_4[40882] = 32'b00000000000000000010111010111010;
assign LUT_4[40883] = 32'b11111111111111111100000110110010;
assign LUT_4[40884] = 32'b00000000000000000000100000110010;
assign LUT_4[40885] = 32'b11111111111111111001101100101010;
assign LUT_4[40886] = 32'b11111111111111111111111011010110;
assign LUT_4[40887] = 32'b11111111111111111001000111001110;
assign LUT_4[40888] = 32'b11111111111111111100101100101011;
assign LUT_4[40889] = 32'b11111111111111110101111000100011;
assign LUT_4[40890] = 32'b11111111111111111100000111001111;
assign LUT_4[40891] = 32'b11111111111111110101010011000111;
assign LUT_4[40892] = 32'b11111111111111111001101101000111;
assign LUT_4[40893] = 32'b11111111111111110010111000111111;
assign LUT_4[40894] = 32'b11111111111111111001000111101011;
assign LUT_4[40895] = 32'b11111111111111110010010011100011;
assign LUT_4[40896] = 32'b00000000000000001000101010110101;
assign LUT_4[40897] = 32'b00000000000000000001110110101101;
assign LUT_4[40898] = 32'b00000000000000001000000101011001;
assign LUT_4[40899] = 32'b00000000000000000001010001010001;
assign LUT_4[40900] = 32'b00000000000000000101101011010001;
assign LUT_4[40901] = 32'b11111111111111111110110111001001;
assign LUT_4[40902] = 32'b00000000000000000101000101110101;
assign LUT_4[40903] = 32'b11111111111111111110010001101101;
assign LUT_4[40904] = 32'b00000000000000000001110111001010;
assign LUT_4[40905] = 32'b11111111111111111011000011000010;
assign LUT_4[40906] = 32'b00000000000000000001010001101110;
assign LUT_4[40907] = 32'b11111111111111111010011101100110;
assign LUT_4[40908] = 32'b11111111111111111110110111100110;
assign LUT_4[40909] = 32'b11111111111111111000000011011110;
assign LUT_4[40910] = 32'b11111111111111111110010010001010;
assign LUT_4[40911] = 32'b11111111111111110111011110000010;
assign LUT_4[40912] = 32'b00000000000000000110011100100011;
assign LUT_4[40913] = 32'b11111111111111111111101000011011;
assign LUT_4[40914] = 32'b00000000000000000101110111000111;
assign LUT_4[40915] = 32'b11111111111111111111000010111111;
assign LUT_4[40916] = 32'b00000000000000000011011100111111;
assign LUT_4[40917] = 32'b11111111111111111100101000110111;
assign LUT_4[40918] = 32'b00000000000000000010110111100011;
assign LUT_4[40919] = 32'b11111111111111111100000011011011;
assign LUT_4[40920] = 32'b11111111111111111111101000111000;
assign LUT_4[40921] = 32'b11111111111111111000110100110000;
assign LUT_4[40922] = 32'b11111111111111111111000011011100;
assign LUT_4[40923] = 32'b11111111111111111000001111010100;
assign LUT_4[40924] = 32'b11111111111111111100101001010100;
assign LUT_4[40925] = 32'b11111111111111110101110101001100;
assign LUT_4[40926] = 32'b11111111111111111100000011111000;
assign LUT_4[40927] = 32'b11111111111111110101001111110000;
assign LUT_4[40928] = 32'b00000000000000000111000101111100;
assign LUT_4[40929] = 32'b00000000000000000000010001110100;
assign LUT_4[40930] = 32'b00000000000000000110100000100000;
assign LUT_4[40931] = 32'b11111111111111111111101100011000;
assign LUT_4[40932] = 32'b00000000000000000100000110011000;
assign LUT_4[40933] = 32'b11111111111111111101010010010000;
assign LUT_4[40934] = 32'b00000000000000000011100000111100;
assign LUT_4[40935] = 32'b11111111111111111100101100110100;
assign LUT_4[40936] = 32'b00000000000000000000010010010001;
assign LUT_4[40937] = 32'b11111111111111111001011110001001;
assign LUT_4[40938] = 32'b11111111111111111111101100110101;
assign LUT_4[40939] = 32'b11111111111111111000111000101101;
assign LUT_4[40940] = 32'b11111111111111111101010010101101;
assign LUT_4[40941] = 32'b11111111111111110110011110100101;
assign LUT_4[40942] = 32'b11111111111111111100101101010001;
assign LUT_4[40943] = 32'b11111111111111110101111001001001;
assign LUT_4[40944] = 32'b00000000000000000100110111101010;
assign LUT_4[40945] = 32'b11111111111111111110000011100010;
assign LUT_4[40946] = 32'b00000000000000000100010010001110;
assign LUT_4[40947] = 32'b11111111111111111101011110000110;
assign LUT_4[40948] = 32'b00000000000000000001111000000110;
assign LUT_4[40949] = 32'b11111111111111111011000011111110;
assign LUT_4[40950] = 32'b00000000000000000001010010101010;
assign LUT_4[40951] = 32'b11111111111111111010011110100010;
assign LUT_4[40952] = 32'b11111111111111111110000011111111;
assign LUT_4[40953] = 32'b11111111111111110111001111110111;
assign LUT_4[40954] = 32'b11111111111111111101011110100011;
assign LUT_4[40955] = 32'b11111111111111110110101010011011;
assign LUT_4[40956] = 32'b11111111111111111011000100011011;
assign LUT_4[40957] = 32'b11111111111111110100010000010011;
assign LUT_4[40958] = 32'b11111111111111111010011110111111;
assign LUT_4[40959] = 32'b11111111111111110011101010110111;
assign LUT_4[40960] = 32'b00000000000000001101100011100000;
assign LUT_4[40961] = 32'b00000000000000000110101111011000;
assign LUT_4[40962] = 32'b00000000000000001100111110000100;
assign LUT_4[40963] = 32'b00000000000000000110001001111100;
assign LUT_4[40964] = 32'b00000000000000001010100011111100;
assign LUT_4[40965] = 32'b00000000000000000011101111110100;
assign LUT_4[40966] = 32'b00000000000000001001111110100000;
assign LUT_4[40967] = 32'b00000000000000000011001010011000;
assign LUT_4[40968] = 32'b00000000000000000110101111110101;
assign LUT_4[40969] = 32'b11111111111111111111111011101101;
assign LUT_4[40970] = 32'b00000000000000000110001010011001;
assign LUT_4[40971] = 32'b11111111111111111111010110010001;
assign LUT_4[40972] = 32'b00000000000000000011110000010001;
assign LUT_4[40973] = 32'b11111111111111111100111100001001;
assign LUT_4[40974] = 32'b00000000000000000011001010110101;
assign LUT_4[40975] = 32'b11111111111111111100010110101101;
assign LUT_4[40976] = 32'b00000000000000001011010101001110;
assign LUT_4[40977] = 32'b00000000000000000100100001000110;
assign LUT_4[40978] = 32'b00000000000000001010101111110010;
assign LUT_4[40979] = 32'b00000000000000000011111011101010;
assign LUT_4[40980] = 32'b00000000000000001000010101101010;
assign LUT_4[40981] = 32'b00000000000000000001100001100010;
assign LUT_4[40982] = 32'b00000000000000000111110000001110;
assign LUT_4[40983] = 32'b00000000000000000000111100000110;
assign LUT_4[40984] = 32'b00000000000000000100100001100011;
assign LUT_4[40985] = 32'b11111111111111111101101101011011;
assign LUT_4[40986] = 32'b00000000000000000011111100000111;
assign LUT_4[40987] = 32'b11111111111111111101000111111111;
assign LUT_4[40988] = 32'b00000000000000000001100001111111;
assign LUT_4[40989] = 32'b11111111111111111010101101110111;
assign LUT_4[40990] = 32'b00000000000000000000111100100011;
assign LUT_4[40991] = 32'b11111111111111111010001000011011;
assign LUT_4[40992] = 32'b00000000000000001011111110100111;
assign LUT_4[40993] = 32'b00000000000000000101001010011111;
assign LUT_4[40994] = 32'b00000000000000001011011001001011;
assign LUT_4[40995] = 32'b00000000000000000100100101000011;
assign LUT_4[40996] = 32'b00000000000000001000111111000011;
assign LUT_4[40997] = 32'b00000000000000000010001010111011;
assign LUT_4[40998] = 32'b00000000000000001000011001100111;
assign LUT_4[40999] = 32'b00000000000000000001100101011111;
assign LUT_4[41000] = 32'b00000000000000000101001010111100;
assign LUT_4[41001] = 32'b11111111111111111110010110110100;
assign LUT_4[41002] = 32'b00000000000000000100100101100000;
assign LUT_4[41003] = 32'b11111111111111111101110001011000;
assign LUT_4[41004] = 32'b00000000000000000010001011011000;
assign LUT_4[41005] = 32'b11111111111111111011010111010000;
assign LUT_4[41006] = 32'b00000000000000000001100101111100;
assign LUT_4[41007] = 32'b11111111111111111010110001110100;
assign LUT_4[41008] = 32'b00000000000000001001110000010101;
assign LUT_4[41009] = 32'b00000000000000000010111100001101;
assign LUT_4[41010] = 32'b00000000000000001001001010111001;
assign LUT_4[41011] = 32'b00000000000000000010010110110001;
assign LUT_4[41012] = 32'b00000000000000000110110000110001;
assign LUT_4[41013] = 32'b11111111111111111111111100101001;
assign LUT_4[41014] = 32'b00000000000000000110001011010101;
assign LUT_4[41015] = 32'b11111111111111111111010111001101;
assign LUT_4[41016] = 32'b00000000000000000010111100101010;
assign LUT_4[41017] = 32'b11111111111111111100001000100010;
assign LUT_4[41018] = 32'b00000000000000000010010111001110;
assign LUT_4[41019] = 32'b11111111111111111011100011000110;
assign LUT_4[41020] = 32'b11111111111111111111111101000110;
assign LUT_4[41021] = 32'b11111111111111111001001000111110;
assign LUT_4[41022] = 32'b11111111111111111111010111101010;
assign LUT_4[41023] = 32'b11111111111111111000100011100010;
assign LUT_4[41024] = 32'b00000000000000001110111010110100;
assign LUT_4[41025] = 32'b00000000000000001000000110101100;
assign LUT_4[41026] = 32'b00000000000000001110010101011000;
assign LUT_4[41027] = 32'b00000000000000000111100001010000;
assign LUT_4[41028] = 32'b00000000000000001011111011010000;
assign LUT_4[41029] = 32'b00000000000000000101000111001000;
assign LUT_4[41030] = 32'b00000000000000001011010101110100;
assign LUT_4[41031] = 32'b00000000000000000100100001101100;
assign LUT_4[41032] = 32'b00000000000000001000000111001001;
assign LUT_4[41033] = 32'b00000000000000000001010011000001;
assign LUT_4[41034] = 32'b00000000000000000111100001101101;
assign LUT_4[41035] = 32'b00000000000000000000101101100101;
assign LUT_4[41036] = 32'b00000000000000000101000111100101;
assign LUT_4[41037] = 32'b11111111111111111110010011011101;
assign LUT_4[41038] = 32'b00000000000000000100100010001001;
assign LUT_4[41039] = 32'b11111111111111111101101110000001;
assign LUT_4[41040] = 32'b00000000000000001100101100100010;
assign LUT_4[41041] = 32'b00000000000000000101111000011010;
assign LUT_4[41042] = 32'b00000000000000001100000111000110;
assign LUT_4[41043] = 32'b00000000000000000101010010111110;
assign LUT_4[41044] = 32'b00000000000000001001101100111110;
assign LUT_4[41045] = 32'b00000000000000000010111000110110;
assign LUT_4[41046] = 32'b00000000000000001001000111100010;
assign LUT_4[41047] = 32'b00000000000000000010010011011010;
assign LUT_4[41048] = 32'b00000000000000000101111000110111;
assign LUT_4[41049] = 32'b11111111111111111111000100101111;
assign LUT_4[41050] = 32'b00000000000000000101010011011011;
assign LUT_4[41051] = 32'b11111111111111111110011111010011;
assign LUT_4[41052] = 32'b00000000000000000010111001010011;
assign LUT_4[41053] = 32'b11111111111111111100000101001011;
assign LUT_4[41054] = 32'b00000000000000000010010011110111;
assign LUT_4[41055] = 32'b11111111111111111011011111101111;
assign LUT_4[41056] = 32'b00000000000000001101010101111011;
assign LUT_4[41057] = 32'b00000000000000000110100001110011;
assign LUT_4[41058] = 32'b00000000000000001100110000011111;
assign LUT_4[41059] = 32'b00000000000000000101111100010111;
assign LUT_4[41060] = 32'b00000000000000001010010110010111;
assign LUT_4[41061] = 32'b00000000000000000011100010001111;
assign LUT_4[41062] = 32'b00000000000000001001110000111011;
assign LUT_4[41063] = 32'b00000000000000000010111100110011;
assign LUT_4[41064] = 32'b00000000000000000110100010010000;
assign LUT_4[41065] = 32'b11111111111111111111101110001000;
assign LUT_4[41066] = 32'b00000000000000000101111100110100;
assign LUT_4[41067] = 32'b11111111111111111111001000101100;
assign LUT_4[41068] = 32'b00000000000000000011100010101100;
assign LUT_4[41069] = 32'b11111111111111111100101110100100;
assign LUT_4[41070] = 32'b00000000000000000010111101010000;
assign LUT_4[41071] = 32'b11111111111111111100001001001000;
assign LUT_4[41072] = 32'b00000000000000001011000111101001;
assign LUT_4[41073] = 32'b00000000000000000100010011100001;
assign LUT_4[41074] = 32'b00000000000000001010100010001101;
assign LUT_4[41075] = 32'b00000000000000000011101110000101;
assign LUT_4[41076] = 32'b00000000000000001000001000000101;
assign LUT_4[41077] = 32'b00000000000000000001010011111101;
assign LUT_4[41078] = 32'b00000000000000000111100010101001;
assign LUT_4[41079] = 32'b00000000000000000000101110100001;
assign LUT_4[41080] = 32'b00000000000000000100010011111110;
assign LUT_4[41081] = 32'b11111111111111111101011111110110;
assign LUT_4[41082] = 32'b00000000000000000011101110100010;
assign LUT_4[41083] = 32'b11111111111111111100111010011010;
assign LUT_4[41084] = 32'b00000000000000000001010100011010;
assign LUT_4[41085] = 32'b11111111111111111010100000010010;
assign LUT_4[41086] = 32'b00000000000000000000101110111110;
assign LUT_4[41087] = 32'b11111111111111111001111010110110;
assign LUT_4[41088] = 32'b00000000000000010000001001101000;
assign LUT_4[41089] = 32'b00000000000000001001010101100000;
assign LUT_4[41090] = 32'b00000000000000001111100100001100;
assign LUT_4[41091] = 32'b00000000000000001000110000000100;
assign LUT_4[41092] = 32'b00000000000000001101001010000100;
assign LUT_4[41093] = 32'b00000000000000000110010101111100;
assign LUT_4[41094] = 32'b00000000000000001100100100101000;
assign LUT_4[41095] = 32'b00000000000000000101110000100000;
assign LUT_4[41096] = 32'b00000000000000001001010101111101;
assign LUT_4[41097] = 32'b00000000000000000010100001110101;
assign LUT_4[41098] = 32'b00000000000000001000110000100001;
assign LUT_4[41099] = 32'b00000000000000000001111100011001;
assign LUT_4[41100] = 32'b00000000000000000110010110011001;
assign LUT_4[41101] = 32'b11111111111111111111100010010001;
assign LUT_4[41102] = 32'b00000000000000000101110000111101;
assign LUT_4[41103] = 32'b11111111111111111110111100110101;
assign LUT_4[41104] = 32'b00000000000000001101111011010110;
assign LUT_4[41105] = 32'b00000000000000000111000111001110;
assign LUT_4[41106] = 32'b00000000000000001101010101111010;
assign LUT_4[41107] = 32'b00000000000000000110100001110010;
assign LUT_4[41108] = 32'b00000000000000001010111011110010;
assign LUT_4[41109] = 32'b00000000000000000100000111101010;
assign LUT_4[41110] = 32'b00000000000000001010010110010110;
assign LUT_4[41111] = 32'b00000000000000000011100010001110;
assign LUT_4[41112] = 32'b00000000000000000111000111101011;
assign LUT_4[41113] = 32'b00000000000000000000010011100011;
assign LUT_4[41114] = 32'b00000000000000000110100010001111;
assign LUT_4[41115] = 32'b11111111111111111111101110000111;
assign LUT_4[41116] = 32'b00000000000000000100001000000111;
assign LUT_4[41117] = 32'b11111111111111111101010011111111;
assign LUT_4[41118] = 32'b00000000000000000011100010101011;
assign LUT_4[41119] = 32'b11111111111111111100101110100011;
assign LUT_4[41120] = 32'b00000000000000001110100100101111;
assign LUT_4[41121] = 32'b00000000000000000111110000100111;
assign LUT_4[41122] = 32'b00000000000000001101111111010011;
assign LUT_4[41123] = 32'b00000000000000000111001011001011;
assign LUT_4[41124] = 32'b00000000000000001011100101001011;
assign LUT_4[41125] = 32'b00000000000000000100110001000011;
assign LUT_4[41126] = 32'b00000000000000001010111111101111;
assign LUT_4[41127] = 32'b00000000000000000100001011100111;
assign LUT_4[41128] = 32'b00000000000000000111110001000100;
assign LUT_4[41129] = 32'b00000000000000000000111100111100;
assign LUT_4[41130] = 32'b00000000000000000111001011101000;
assign LUT_4[41131] = 32'b00000000000000000000010111100000;
assign LUT_4[41132] = 32'b00000000000000000100110001100000;
assign LUT_4[41133] = 32'b11111111111111111101111101011000;
assign LUT_4[41134] = 32'b00000000000000000100001100000100;
assign LUT_4[41135] = 32'b11111111111111111101010111111100;
assign LUT_4[41136] = 32'b00000000000000001100010110011101;
assign LUT_4[41137] = 32'b00000000000000000101100010010101;
assign LUT_4[41138] = 32'b00000000000000001011110001000001;
assign LUT_4[41139] = 32'b00000000000000000100111100111001;
assign LUT_4[41140] = 32'b00000000000000001001010110111001;
assign LUT_4[41141] = 32'b00000000000000000010100010110001;
assign LUT_4[41142] = 32'b00000000000000001000110001011101;
assign LUT_4[41143] = 32'b00000000000000000001111101010101;
assign LUT_4[41144] = 32'b00000000000000000101100010110010;
assign LUT_4[41145] = 32'b11111111111111111110101110101010;
assign LUT_4[41146] = 32'b00000000000000000100111101010110;
assign LUT_4[41147] = 32'b11111111111111111110001001001110;
assign LUT_4[41148] = 32'b00000000000000000010100011001110;
assign LUT_4[41149] = 32'b11111111111111111011101111000110;
assign LUT_4[41150] = 32'b00000000000000000001111101110010;
assign LUT_4[41151] = 32'b11111111111111111011001001101010;
assign LUT_4[41152] = 32'b00000000000000010001100000111100;
assign LUT_4[41153] = 32'b00000000000000001010101100110100;
assign LUT_4[41154] = 32'b00000000000000010000111011100000;
assign LUT_4[41155] = 32'b00000000000000001010000111011000;
assign LUT_4[41156] = 32'b00000000000000001110100001011000;
assign LUT_4[41157] = 32'b00000000000000000111101101010000;
assign LUT_4[41158] = 32'b00000000000000001101111011111100;
assign LUT_4[41159] = 32'b00000000000000000111000111110100;
assign LUT_4[41160] = 32'b00000000000000001010101101010001;
assign LUT_4[41161] = 32'b00000000000000000011111001001001;
assign LUT_4[41162] = 32'b00000000000000001010000111110101;
assign LUT_4[41163] = 32'b00000000000000000011010011101101;
assign LUT_4[41164] = 32'b00000000000000000111101101101101;
assign LUT_4[41165] = 32'b00000000000000000000111001100101;
assign LUT_4[41166] = 32'b00000000000000000111001000010001;
assign LUT_4[41167] = 32'b00000000000000000000010100001001;
assign LUT_4[41168] = 32'b00000000000000001111010010101010;
assign LUT_4[41169] = 32'b00000000000000001000011110100010;
assign LUT_4[41170] = 32'b00000000000000001110101101001110;
assign LUT_4[41171] = 32'b00000000000000000111111001000110;
assign LUT_4[41172] = 32'b00000000000000001100010011000110;
assign LUT_4[41173] = 32'b00000000000000000101011110111110;
assign LUT_4[41174] = 32'b00000000000000001011101101101010;
assign LUT_4[41175] = 32'b00000000000000000100111001100010;
assign LUT_4[41176] = 32'b00000000000000001000011110111111;
assign LUT_4[41177] = 32'b00000000000000000001101010110111;
assign LUT_4[41178] = 32'b00000000000000000111111001100011;
assign LUT_4[41179] = 32'b00000000000000000001000101011011;
assign LUT_4[41180] = 32'b00000000000000000101011111011011;
assign LUT_4[41181] = 32'b11111111111111111110101011010011;
assign LUT_4[41182] = 32'b00000000000000000100111001111111;
assign LUT_4[41183] = 32'b11111111111111111110000101110111;
assign LUT_4[41184] = 32'b00000000000000001111111100000011;
assign LUT_4[41185] = 32'b00000000000000001001000111111011;
assign LUT_4[41186] = 32'b00000000000000001111010110100111;
assign LUT_4[41187] = 32'b00000000000000001000100010011111;
assign LUT_4[41188] = 32'b00000000000000001100111100011111;
assign LUT_4[41189] = 32'b00000000000000000110001000010111;
assign LUT_4[41190] = 32'b00000000000000001100010111000011;
assign LUT_4[41191] = 32'b00000000000000000101100010111011;
assign LUT_4[41192] = 32'b00000000000000001001001000011000;
assign LUT_4[41193] = 32'b00000000000000000010010100010000;
assign LUT_4[41194] = 32'b00000000000000001000100010111100;
assign LUT_4[41195] = 32'b00000000000000000001101110110100;
assign LUT_4[41196] = 32'b00000000000000000110001000110100;
assign LUT_4[41197] = 32'b11111111111111111111010100101100;
assign LUT_4[41198] = 32'b00000000000000000101100011011000;
assign LUT_4[41199] = 32'b11111111111111111110101111010000;
assign LUT_4[41200] = 32'b00000000000000001101101101110001;
assign LUT_4[41201] = 32'b00000000000000000110111001101001;
assign LUT_4[41202] = 32'b00000000000000001101001000010101;
assign LUT_4[41203] = 32'b00000000000000000110010100001101;
assign LUT_4[41204] = 32'b00000000000000001010101110001101;
assign LUT_4[41205] = 32'b00000000000000000011111010000101;
assign LUT_4[41206] = 32'b00000000000000001010001000110001;
assign LUT_4[41207] = 32'b00000000000000000011010100101001;
assign LUT_4[41208] = 32'b00000000000000000110111010000110;
assign LUT_4[41209] = 32'b00000000000000000000000101111110;
assign LUT_4[41210] = 32'b00000000000000000110010100101010;
assign LUT_4[41211] = 32'b11111111111111111111100000100010;
assign LUT_4[41212] = 32'b00000000000000000011111010100010;
assign LUT_4[41213] = 32'b11111111111111111101000110011010;
assign LUT_4[41214] = 32'b00000000000000000011010101000110;
assign LUT_4[41215] = 32'b11111111111111111100100000111110;
assign LUT_4[41216] = 32'b00000000000000010010011111000011;
assign LUT_4[41217] = 32'b00000000000000001011101010111011;
assign LUT_4[41218] = 32'b00000000000000010001111001100111;
assign LUT_4[41219] = 32'b00000000000000001011000101011111;
assign LUT_4[41220] = 32'b00000000000000001111011111011111;
assign LUT_4[41221] = 32'b00000000000000001000101011010111;
assign LUT_4[41222] = 32'b00000000000000001110111010000011;
assign LUT_4[41223] = 32'b00000000000000001000000101111011;
assign LUT_4[41224] = 32'b00000000000000001011101011011000;
assign LUT_4[41225] = 32'b00000000000000000100110111010000;
assign LUT_4[41226] = 32'b00000000000000001011000101111100;
assign LUT_4[41227] = 32'b00000000000000000100010001110100;
assign LUT_4[41228] = 32'b00000000000000001000101011110100;
assign LUT_4[41229] = 32'b00000000000000000001110111101100;
assign LUT_4[41230] = 32'b00000000000000001000000110011000;
assign LUT_4[41231] = 32'b00000000000000000001010010010000;
assign LUT_4[41232] = 32'b00000000000000010000010000110001;
assign LUT_4[41233] = 32'b00000000000000001001011100101001;
assign LUT_4[41234] = 32'b00000000000000001111101011010101;
assign LUT_4[41235] = 32'b00000000000000001000110111001101;
assign LUT_4[41236] = 32'b00000000000000001101010001001101;
assign LUT_4[41237] = 32'b00000000000000000110011101000101;
assign LUT_4[41238] = 32'b00000000000000001100101011110001;
assign LUT_4[41239] = 32'b00000000000000000101110111101001;
assign LUT_4[41240] = 32'b00000000000000001001011101000110;
assign LUT_4[41241] = 32'b00000000000000000010101000111110;
assign LUT_4[41242] = 32'b00000000000000001000110111101010;
assign LUT_4[41243] = 32'b00000000000000000010000011100010;
assign LUT_4[41244] = 32'b00000000000000000110011101100010;
assign LUT_4[41245] = 32'b11111111111111111111101001011010;
assign LUT_4[41246] = 32'b00000000000000000101111000000110;
assign LUT_4[41247] = 32'b11111111111111111111000011111110;
assign LUT_4[41248] = 32'b00000000000000010000111010001010;
assign LUT_4[41249] = 32'b00000000000000001010000110000010;
assign LUT_4[41250] = 32'b00000000000000010000010100101110;
assign LUT_4[41251] = 32'b00000000000000001001100000100110;
assign LUT_4[41252] = 32'b00000000000000001101111010100110;
assign LUT_4[41253] = 32'b00000000000000000111000110011110;
assign LUT_4[41254] = 32'b00000000000000001101010101001010;
assign LUT_4[41255] = 32'b00000000000000000110100001000010;
assign LUT_4[41256] = 32'b00000000000000001010000110011111;
assign LUT_4[41257] = 32'b00000000000000000011010010010111;
assign LUT_4[41258] = 32'b00000000000000001001100001000011;
assign LUT_4[41259] = 32'b00000000000000000010101100111011;
assign LUT_4[41260] = 32'b00000000000000000111000110111011;
assign LUT_4[41261] = 32'b00000000000000000000010010110011;
assign LUT_4[41262] = 32'b00000000000000000110100001011111;
assign LUT_4[41263] = 32'b11111111111111111111101101010111;
assign LUT_4[41264] = 32'b00000000000000001110101011111000;
assign LUT_4[41265] = 32'b00000000000000000111110111110000;
assign LUT_4[41266] = 32'b00000000000000001110000110011100;
assign LUT_4[41267] = 32'b00000000000000000111010010010100;
assign LUT_4[41268] = 32'b00000000000000001011101100010100;
assign LUT_4[41269] = 32'b00000000000000000100111000001100;
assign LUT_4[41270] = 32'b00000000000000001011000110111000;
assign LUT_4[41271] = 32'b00000000000000000100010010110000;
assign LUT_4[41272] = 32'b00000000000000000111111000001101;
assign LUT_4[41273] = 32'b00000000000000000001000100000101;
assign LUT_4[41274] = 32'b00000000000000000111010010110001;
assign LUT_4[41275] = 32'b00000000000000000000011110101001;
assign LUT_4[41276] = 32'b00000000000000000100111000101001;
assign LUT_4[41277] = 32'b11111111111111111110000100100001;
assign LUT_4[41278] = 32'b00000000000000000100010011001101;
assign LUT_4[41279] = 32'b11111111111111111101011111000101;
assign LUT_4[41280] = 32'b00000000000000010011110110010111;
assign LUT_4[41281] = 32'b00000000000000001101000010001111;
assign LUT_4[41282] = 32'b00000000000000010011010000111011;
assign LUT_4[41283] = 32'b00000000000000001100011100110011;
assign LUT_4[41284] = 32'b00000000000000010000110110110011;
assign LUT_4[41285] = 32'b00000000000000001010000010101011;
assign LUT_4[41286] = 32'b00000000000000010000010001010111;
assign LUT_4[41287] = 32'b00000000000000001001011101001111;
assign LUT_4[41288] = 32'b00000000000000001101000010101100;
assign LUT_4[41289] = 32'b00000000000000000110001110100100;
assign LUT_4[41290] = 32'b00000000000000001100011101010000;
assign LUT_4[41291] = 32'b00000000000000000101101001001000;
assign LUT_4[41292] = 32'b00000000000000001010000011001000;
assign LUT_4[41293] = 32'b00000000000000000011001111000000;
assign LUT_4[41294] = 32'b00000000000000001001011101101100;
assign LUT_4[41295] = 32'b00000000000000000010101001100100;
assign LUT_4[41296] = 32'b00000000000000010001101000000101;
assign LUT_4[41297] = 32'b00000000000000001010110011111101;
assign LUT_4[41298] = 32'b00000000000000010001000010101001;
assign LUT_4[41299] = 32'b00000000000000001010001110100001;
assign LUT_4[41300] = 32'b00000000000000001110101000100001;
assign LUT_4[41301] = 32'b00000000000000000111110100011001;
assign LUT_4[41302] = 32'b00000000000000001110000011000101;
assign LUT_4[41303] = 32'b00000000000000000111001110111101;
assign LUT_4[41304] = 32'b00000000000000001010110100011010;
assign LUT_4[41305] = 32'b00000000000000000100000000010010;
assign LUT_4[41306] = 32'b00000000000000001010001110111110;
assign LUT_4[41307] = 32'b00000000000000000011011010110110;
assign LUT_4[41308] = 32'b00000000000000000111110100110110;
assign LUT_4[41309] = 32'b00000000000000000001000000101110;
assign LUT_4[41310] = 32'b00000000000000000111001111011010;
assign LUT_4[41311] = 32'b00000000000000000000011011010010;
assign LUT_4[41312] = 32'b00000000000000010010010001011110;
assign LUT_4[41313] = 32'b00000000000000001011011101010110;
assign LUT_4[41314] = 32'b00000000000000010001101100000010;
assign LUT_4[41315] = 32'b00000000000000001010110111111010;
assign LUT_4[41316] = 32'b00000000000000001111010001111010;
assign LUT_4[41317] = 32'b00000000000000001000011101110010;
assign LUT_4[41318] = 32'b00000000000000001110101100011110;
assign LUT_4[41319] = 32'b00000000000000000111111000010110;
assign LUT_4[41320] = 32'b00000000000000001011011101110011;
assign LUT_4[41321] = 32'b00000000000000000100101001101011;
assign LUT_4[41322] = 32'b00000000000000001010111000010111;
assign LUT_4[41323] = 32'b00000000000000000100000100001111;
assign LUT_4[41324] = 32'b00000000000000001000011110001111;
assign LUT_4[41325] = 32'b00000000000000000001101010000111;
assign LUT_4[41326] = 32'b00000000000000000111111000110011;
assign LUT_4[41327] = 32'b00000000000000000001000100101011;
assign LUT_4[41328] = 32'b00000000000000010000000011001100;
assign LUT_4[41329] = 32'b00000000000000001001001111000100;
assign LUT_4[41330] = 32'b00000000000000001111011101110000;
assign LUT_4[41331] = 32'b00000000000000001000101001101000;
assign LUT_4[41332] = 32'b00000000000000001101000011101000;
assign LUT_4[41333] = 32'b00000000000000000110001111100000;
assign LUT_4[41334] = 32'b00000000000000001100011110001100;
assign LUT_4[41335] = 32'b00000000000000000101101010000100;
assign LUT_4[41336] = 32'b00000000000000001001001111100001;
assign LUT_4[41337] = 32'b00000000000000000010011011011001;
assign LUT_4[41338] = 32'b00000000000000001000101010000101;
assign LUT_4[41339] = 32'b00000000000000000001110101111101;
assign LUT_4[41340] = 32'b00000000000000000110001111111101;
assign LUT_4[41341] = 32'b11111111111111111111011011110101;
assign LUT_4[41342] = 32'b00000000000000000101101010100001;
assign LUT_4[41343] = 32'b11111111111111111110110110011001;
assign LUT_4[41344] = 32'b00000000000000010101000101001011;
assign LUT_4[41345] = 32'b00000000000000001110010001000011;
assign LUT_4[41346] = 32'b00000000000000010100011111101111;
assign LUT_4[41347] = 32'b00000000000000001101101011100111;
assign LUT_4[41348] = 32'b00000000000000010010000101100111;
assign LUT_4[41349] = 32'b00000000000000001011010001011111;
assign LUT_4[41350] = 32'b00000000000000010001100000001011;
assign LUT_4[41351] = 32'b00000000000000001010101100000011;
assign LUT_4[41352] = 32'b00000000000000001110010001100000;
assign LUT_4[41353] = 32'b00000000000000000111011101011000;
assign LUT_4[41354] = 32'b00000000000000001101101100000100;
assign LUT_4[41355] = 32'b00000000000000000110110111111100;
assign LUT_4[41356] = 32'b00000000000000001011010001111100;
assign LUT_4[41357] = 32'b00000000000000000100011101110100;
assign LUT_4[41358] = 32'b00000000000000001010101100100000;
assign LUT_4[41359] = 32'b00000000000000000011111000011000;
assign LUT_4[41360] = 32'b00000000000000010010110110111001;
assign LUT_4[41361] = 32'b00000000000000001100000010110001;
assign LUT_4[41362] = 32'b00000000000000010010010001011101;
assign LUT_4[41363] = 32'b00000000000000001011011101010101;
assign LUT_4[41364] = 32'b00000000000000001111110111010101;
assign LUT_4[41365] = 32'b00000000000000001001000011001101;
assign LUT_4[41366] = 32'b00000000000000001111010001111001;
assign LUT_4[41367] = 32'b00000000000000001000011101110001;
assign LUT_4[41368] = 32'b00000000000000001100000011001110;
assign LUT_4[41369] = 32'b00000000000000000101001111000110;
assign LUT_4[41370] = 32'b00000000000000001011011101110010;
assign LUT_4[41371] = 32'b00000000000000000100101001101010;
assign LUT_4[41372] = 32'b00000000000000001001000011101010;
assign LUT_4[41373] = 32'b00000000000000000010001111100010;
assign LUT_4[41374] = 32'b00000000000000001000011110001110;
assign LUT_4[41375] = 32'b00000000000000000001101010000110;
assign LUT_4[41376] = 32'b00000000000000010011100000010010;
assign LUT_4[41377] = 32'b00000000000000001100101100001010;
assign LUT_4[41378] = 32'b00000000000000010010111010110110;
assign LUT_4[41379] = 32'b00000000000000001100000110101110;
assign LUT_4[41380] = 32'b00000000000000010000100000101110;
assign LUT_4[41381] = 32'b00000000000000001001101100100110;
assign LUT_4[41382] = 32'b00000000000000001111111011010010;
assign LUT_4[41383] = 32'b00000000000000001001000111001010;
assign LUT_4[41384] = 32'b00000000000000001100101100100111;
assign LUT_4[41385] = 32'b00000000000000000101111000011111;
assign LUT_4[41386] = 32'b00000000000000001100000111001011;
assign LUT_4[41387] = 32'b00000000000000000101010011000011;
assign LUT_4[41388] = 32'b00000000000000001001101101000011;
assign LUT_4[41389] = 32'b00000000000000000010111000111011;
assign LUT_4[41390] = 32'b00000000000000001001000111100111;
assign LUT_4[41391] = 32'b00000000000000000010010011011111;
assign LUT_4[41392] = 32'b00000000000000010001010010000000;
assign LUT_4[41393] = 32'b00000000000000001010011101111000;
assign LUT_4[41394] = 32'b00000000000000010000101100100100;
assign LUT_4[41395] = 32'b00000000000000001001111000011100;
assign LUT_4[41396] = 32'b00000000000000001110010010011100;
assign LUT_4[41397] = 32'b00000000000000000111011110010100;
assign LUT_4[41398] = 32'b00000000000000001101101101000000;
assign LUT_4[41399] = 32'b00000000000000000110111000111000;
assign LUT_4[41400] = 32'b00000000000000001010011110010101;
assign LUT_4[41401] = 32'b00000000000000000011101010001101;
assign LUT_4[41402] = 32'b00000000000000001001111000111001;
assign LUT_4[41403] = 32'b00000000000000000011000100110001;
assign LUT_4[41404] = 32'b00000000000000000111011110110001;
assign LUT_4[41405] = 32'b00000000000000000000101010101001;
assign LUT_4[41406] = 32'b00000000000000000110111001010101;
assign LUT_4[41407] = 32'b00000000000000000000000101001101;
assign LUT_4[41408] = 32'b00000000000000010110011100011111;
assign LUT_4[41409] = 32'b00000000000000001111101000010111;
assign LUT_4[41410] = 32'b00000000000000010101110111000011;
assign LUT_4[41411] = 32'b00000000000000001111000010111011;
assign LUT_4[41412] = 32'b00000000000000010011011100111011;
assign LUT_4[41413] = 32'b00000000000000001100101000110011;
assign LUT_4[41414] = 32'b00000000000000010010110111011111;
assign LUT_4[41415] = 32'b00000000000000001100000011010111;
assign LUT_4[41416] = 32'b00000000000000001111101000110100;
assign LUT_4[41417] = 32'b00000000000000001000110100101100;
assign LUT_4[41418] = 32'b00000000000000001111000011011000;
assign LUT_4[41419] = 32'b00000000000000001000001111010000;
assign LUT_4[41420] = 32'b00000000000000001100101001010000;
assign LUT_4[41421] = 32'b00000000000000000101110101001000;
assign LUT_4[41422] = 32'b00000000000000001100000011110100;
assign LUT_4[41423] = 32'b00000000000000000101001111101100;
assign LUT_4[41424] = 32'b00000000000000010100001110001101;
assign LUT_4[41425] = 32'b00000000000000001101011010000101;
assign LUT_4[41426] = 32'b00000000000000010011101000110001;
assign LUT_4[41427] = 32'b00000000000000001100110100101001;
assign LUT_4[41428] = 32'b00000000000000010001001110101001;
assign LUT_4[41429] = 32'b00000000000000001010011010100001;
assign LUT_4[41430] = 32'b00000000000000010000101001001101;
assign LUT_4[41431] = 32'b00000000000000001001110101000101;
assign LUT_4[41432] = 32'b00000000000000001101011010100010;
assign LUT_4[41433] = 32'b00000000000000000110100110011010;
assign LUT_4[41434] = 32'b00000000000000001100110101000110;
assign LUT_4[41435] = 32'b00000000000000000110000000111110;
assign LUT_4[41436] = 32'b00000000000000001010011010111110;
assign LUT_4[41437] = 32'b00000000000000000011100110110110;
assign LUT_4[41438] = 32'b00000000000000001001110101100010;
assign LUT_4[41439] = 32'b00000000000000000011000001011010;
assign LUT_4[41440] = 32'b00000000000000010100110111100110;
assign LUT_4[41441] = 32'b00000000000000001110000011011110;
assign LUT_4[41442] = 32'b00000000000000010100010010001010;
assign LUT_4[41443] = 32'b00000000000000001101011110000010;
assign LUT_4[41444] = 32'b00000000000000010001111000000010;
assign LUT_4[41445] = 32'b00000000000000001011000011111010;
assign LUT_4[41446] = 32'b00000000000000010001010010100110;
assign LUT_4[41447] = 32'b00000000000000001010011110011110;
assign LUT_4[41448] = 32'b00000000000000001110000011111011;
assign LUT_4[41449] = 32'b00000000000000000111001111110011;
assign LUT_4[41450] = 32'b00000000000000001101011110011111;
assign LUT_4[41451] = 32'b00000000000000000110101010010111;
assign LUT_4[41452] = 32'b00000000000000001011000100010111;
assign LUT_4[41453] = 32'b00000000000000000100010000001111;
assign LUT_4[41454] = 32'b00000000000000001010011110111011;
assign LUT_4[41455] = 32'b00000000000000000011101010110011;
assign LUT_4[41456] = 32'b00000000000000010010101001010100;
assign LUT_4[41457] = 32'b00000000000000001011110101001100;
assign LUT_4[41458] = 32'b00000000000000010010000011111000;
assign LUT_4[41459] = 32'b00000000000000001011001111110000;
assign LUT_4[41460] = 32'b00000000000000001111101001110000;
assign LUT_4[41461] = 32'b00000000000000001000110101101000;
assign LUT_4[41462] = 32'b00000000000000001111000100010100;
assign LUT_4[41463] = 32'b00000000000000001000010000001100;
assign LUT_4[41464] = 32'b00000000000000001011110101101001;
assign LUT_4[41465] = 32'b00000000000000000101000001100001;
assign LUT_4[41466] = 32'b00000000000000001011010000001101;
assign LUT_4[41467] = 32'b00000000000000000100011100000101;
assign LUT_4[41468] = 32'b00000000000000001000110110000101;
assign LUT_4[41469] = 32'b00000000000000000010000001111101;
assign LUT_4[41470] = 32'b00000000000000001000010000101001;
assign LUT_4[41471] = 32'b00000000000000000001011100100001;
assign LUT_4[41472] = 32'b00000000000000001100100111101000;
assign LUT_4[41473] = 32'b00000000000000000101110011100000;
assign LUT_4[41474] = 32'b00000000000000001100000010001100;
assign LUT_4[41475] = 32'b00000000000000000101001110000100;
assign LUT_4[41476] = 32'b00000000000000001001101000000100;
assign LUT_4[41477] = 32'b00000000000000000010110011111100;
assign LUT_4[41478] = 32'b00000000000000001001000010101000;
assign LUT_4[41479] = 32'b00000000000000000010001110100000;
assign LUT_4[41480] = 32'b00000000000000000101110011111101;
assign LUT_4[41481] = 32'b11111111111111111110111111110101;
assign LUT_4[41482] = 32'b00000000000000000101001110100001;
assign LUT_4[41483] = 32'b11111111111111111110011010011001;
assign LUT_4[41484] = 32'b00000000000000000010110100011001;
assign LUT_4[41485] = 32'b11111111111111111100000000010001;
assign LUT_4[41486] = 32'b00000000000000000010001110111101;
assign LUT_4[41487] = 32'b11111111111111111011011010110101;
assign LUT_4[41488] = 32'b00000000000000001010011001010110;
assign LUT_4[41489] = 32'b00000000000000000011100101001110;
assign LUT_4[41490] = 32'b00000000000000001001110011111010;
assign LUT_4[41491] = 32'b00000000000000000010111111110010;
assign LUT_4[41492] = 32'b00000000000000000111011001110010;
assign LUT_4[41493] = 32'b00000000000000000000100101101010;
assign LUT_4[41494] = 32'b00000000000000000110110100010110;
assign LUT_4[41495] = 32'b00000000000000000000000000001110;
assign LUT_4[41496] = 32'b00000000000000000011100101101011;
assign LUT_4[41497] = 32'b11111111111111111100110001100011;
assign LUT_4[41498] = 32'b00000000000000000011000000001111;
assign LUT_4[41499] = 32'b11111111111111111100001100000111;
assign LUT_4[41500] = 32'b00000000000000000000100110000111;
assign LUT_4[41501] = 32'b11111111111111111001110001111111;
assign LUT_4[41502] = 32'b00000000000000000000000000101011;
assign LUT_4[41503] = 32'b11111111111111111001001100100011;
assign LUT_4[41504] = 32'b00000000000000001011000010101111;
assign LUT_4[41505] = 32'b00000000000000000100001110100111;
assign LUT_4[41506] = 32'b00000000000000001010011101010011;
assign LUT_4[41507] = 32'b00000000000000000011101001001011;
assign LUT_4[41508] = 32'b00000000000000001000000011001011;
assign LUT_4[41509] = 32'b00000000000000000001001111000011;
assign LUT_4[41510] = 32'b00000000000000000111011101101111;
assign LUT_4[41511] = 32'b00000000000000000000101001100111;
assign LUT_4[41512] = 32'b00000000000000000100001111000100;
assign LUT_4[41513] = 32'b11111111111111111101011010111100;
assign LUT_4[41514] = 32'b00000000000000000011101001101000;
assign LUT_4[41515] = 32'b11111111111111111100110101100000;
assign LUT_4[41516] = 32'b00000000000000000001001111100000;
assign LUT_4[41517] = 32'b11111111111111111010011011011000;
assign LUT_4[41518] = 32'b00000000000000000000101010000100;
assign LUT_4[41519] = 32'b11111111111111111001110101111100;
assign LUT_4[41520] = 32'b00000000000000001000110100011101;
assign LUT_4[41521] = 32'b00000000000000000010000000010101;
assign LUT_4[41522] = 32'b00000000000000001000001111000001;
assign LUT_4[41523] = 32'b00000000000000000001011010111001;
assign LUT_4[41524] = 32'b00000000000000000101110100111001;
assign LUT_4[41525] = 32'b11111111111111111111000000110001;
assign LUT_4[41526] = 32'b00000000000000000101001111011101;
assign LUT_4[41527] = 32'b11111111111111111110011011010101;
assign LUT_4[41528] = 32'b00000000000000000010000000110010;
assign LUT_4[41529] = 32'b11111111111111111011001100101010;
assign LUT_4[41530] = 32'b00000000000000000001011011010110;
assign LUT_4[41531] = 32'b11111111111111111010100111001110;
assign LUT_4[41532] = 32'b11111111111111111111000001001110;
assign LUT_4[41533] = 32'b11111111111111111000001101000110;
assign LUT_4[41534] = 32'b11111111111111111110011011110010;
assign LUT_4[41535] = 32'b11111111111111110111100111101010;
assign LUT_4[41536] = 32'b00000000000000001101111110111100;
assign LUT_4[41537] = 32'b00000000000000000111001010110100;
assign LUT_4[41538] = 32'b00000000000000001101011001100000;
assign LUT_4[41539] = 32'b00000000000000000110100101011000;
assign LUT_4[41540] = 32'b00000000000000001010111111011000;
assign LUT_4[41541] = 32'b00000000000000000100001011010000;
assign LUT_4[41542] = 32'b00000000000000001010011001111100;
assign LUT_4[41543] = 32'b00000000000000000011100101110100;
assign LUT_4[41544] = 32'b00000000000000000111001011010001;
assign LUT_4[41545] = 32'b00000000000000000000010111001001;
assign LUT_4[41546] = 32'b00000000000000000110100101110101;
assign LUT_4[41547] = 32'b11111111111111111111110001101101;
assign LUT_4[41548] = 32'b00000000000000000100001011101101;
assign LUT_4[41549] = 32'b11111111111111111101010111100101;
assign LUT_4[41550] = 32'b00000000000000000011100110010001;
assign LUT_4[41551] = 32'b11111111111111111100110010001001;
assign LUT_4[41552] = 32'b00000000000000001011110000101010;
assign LUT_4[41553] = 32'b00000000000000000100111100100010;
assign LUT_4[41554] = 32'b00000000000000001011001011001110;
assign LUT_4[41555] = 32'b00000000000000000100010111000110;
assign LUT_4[41556] = 32'b00000000000000001000110001000110;
assign LUT_4[41557] = 32'b00000000000000000001111100111110;
assign LUT_4[41558] = 32'b00000000000000001000001011101010;
assign LUT_4[41559] = 32'b00000000000000000001010111100010;
assign LUT_4[41560] = 32'b00000000000000000100111100111111;
assign LUT_4[41561] = 32'b11111111111111111110001000110111;
assign LUT_4[41562] = 32'b00000000000000000100010111100011;
assign LUT_4[41563] = 32'b11111111111111111101100011011011;
assign LUT_4[41564] = 32'b00000000000000000001111101011011;
assign LUT_4[41565] = 32'b11111111111111111011001001010011;
assign LUT_4[41566] = 32'b00000000000000000001010111111111;
assign LUT_4[41567] = 32'b11111111111111111010100011110111;
assign LUT_4[41568] = 32'b00000000000000001100011010000011;
assign LUT_4[41569] = 32'b00000000000000000101100101111011;
assign LUT_4[41570] = 32'b00000000000000001011110100100111;
assign LUT_4[41571] = 32'b00000000000000000101000000011111;
assign LUT_4[41572] = 32'b00000000000000001001011010011111;
assign LUT_4[41573] = 32'b00000000000000000010100110010111;
assign LUT_4[41574] = 32'b00000000000000001000110101000011;
assign LUT_4[41575] = 32'b00000000000000000010000000111011;
assign LUT_4[41576] = 32'b00000000000000000101100110011000;
assign LUT_4[41577] = 32'b11111111111111111110110010010000;
assign LUT_4[41578] = 32'b00000000000000000101000000111100;
assign LUT_4[41579] = 32'b11111111111111111110001100110100;
assign LUT_4[41580] = 32'b00000000000000000010100110110100;
assign LUT_4[41581] = 32'b11111111111111111011110010101100;
assign LUT_4[41582] = 32'b00000000000000000010000001011000;
assign LUT_4[41583] = 32'b11111111111111111011001101010000;
assign LUT_4[41584] = 32'b00000000000000001010001011110001;
assign LUT_4[41585] = 32'b00000000000000000011010111101001;
assign LUT_4[41586] = 32'b00000000000000001001100110010101;
assign LUT_4[41587] = 32'b00000000000000000010110010001101;
assign LUT_4[41588] = 32'b00000000000000000111001100001101;
assign LUT_4[41589] = 32'b00000000000000000000011000000101;
assign LUT_4[41590] = 32'b00000000000000000110100110110001;
assign LUT_4[41591] = 32'b11111111111111111111110010101001;
assign LUT_4[41592] = 32'b00000000000000000011011000000110;
assign LUT_4[41593] = 32'b11111111111111111100100011111110;
assign LUT_4[41594] = 32'b00000000000000000010110010101010;
assign LUT_4[41595] = 32'b11111111111111111011111110100010;
assign LUT_4[41596] = 32'b00000000000000000000011000100010;
assign LUT_4[41597] = 32'b11111111111111111001100100011010;
assign LUT_4[41598] = 32'b11111111111111111111110011000110;
assign LUT_4[41599] = 32'b11111111111111111000111110111110;
assign LUT_4[41600] = 32'b00000000000000001111001101110000;
assign LUT_4[41601] = 32'b00000000000000001000011001101000;
assign LUT_4[41602] = 32'b00000000000000001110101000010100;
assign LUT_4[41603] = 32'b00000000000000000111110100001100;
assign LUT_4[41604] = 32'b00000000000000001100001110001100;
assign LUT_4[41605] = 32'b00000000000000000101011010000100;
assign LUT_4[41606] = 32'b00000000000000001011101000110000;
assign LUT_4[41607] = 32'b00000000000000000100110100101000;
assign LUT_4[41608] = 32'b00000000000000001000011010000101;
assign LUT_4[41609] = 32'b00000000000000000001100101111101;
assign LUT_4[41610] = 32'b00000000000000000111110100101001;
assign LUT_4[41611] = 32'b00000000000000000001000000100001;
assign LUT_4[41612] = 32'b00000000000000000101011010100001;
assign LUT_4[41613] = 32'b11111111111111111110100110011001;
assign LUT_4[41614] = 32'b00000000000000000100110101000101;
assign LUT_4[41615] = 32'b11111111111111111110000000111101;
assign LUT_4[41616] = 32'b00000000000000001100111111011110;
assign LUT_4[41617] = 32'b00000000000000000110001011010110;
assign LUT_4[41618] = 32'b00000000000000001100011010000010;
assign LUT_4[41619] = 32'b00000000000000000101100101111010;
assign LUT_4[41620] = 32'b00000000000000001001111111111010;
assign LUT_4[41621] = 32'b00000000000000000011001011110010;
assign LUT_4[41622] = 32'b00000000000000001001011010011110;
assign LUT_4[41623] = 32'b00000000000000000010100110010110;
assign LUT_4[41624] = 32'b00000000000000000110001011110011;
assign LUT_4[41625] = 32'b11111111111111111111010111101011;
assign LUT_4[41626] = 32'b00000000000000000101100110010111;
assign LUT_4[41627] = 32'b11111111111111111110110010001111;
assign LUT_4[41628] = 32'b00000000000000000011001100001111;
assign LUT_4[41629] = 32'b11111111111111111100011000000111;
assign LUT_4[41630] = 32'b00000000000000000010100110110011;
assign LUT_4[41631] = 32'b11111111111111111011110010101011;
assign LUT_4[41632] = 32'b00000000000000001101101000110111;
assign LUT_4[41633] = 32'b00000000000000000110110100101111;
assign LUT_4[41634] = 32'b00000000000000001101000011011011;
assign LUT_4[41635] = 32'b00000000000000000110001111010011;
assign LUT_4[41636] = 32'b00000000000000001010101001010011;
assign LUT_4[41637] = 32'b00000000000000000011110101001011;
assign LUT_4[41638] = 32'b00000000000000001010000011110111;
assign LUT_4[41639] = 32'b00000000000000000011001111101111;
assign LUT_4[41640] = 32'b00000000000000000110110101001100;
assign LUT_4[41641] = 32'b00000000000000000000000001000100;
assign LUT_4[41642] = 32'b00000000000000000110001111110000;
assign LUT_4[41643] = 32'b11111111111111111111011011101000;
assign LUT_4[41644] = 32'b00000000000000000011110101101000;
assign LUT_4[41645] = 32'b11111111111111111101000001100000;
assign LUT_4[41646] = 32'b00000000000000000011010000001100;
assign LUT_4[41647] = 32'b11111111111111111100011100000100;
assign LUT_4[41648] = 32'b00000000000000001011011010100101;
assign LUT_4[41649] = 32'b00000000000000000100100110011101;
assign LUT_4[41650] = 32'b00000000000000001010110101001001;
assign LUT_4[41651] = 32'b00000000000000000100000001000001;
assign LUT_4[41652] = 32'b00000000000000001000011011000001;
assign LUT_4[41653] = 32'b00000000000000000001100110111001;
assign LUT_4[41654] = 32'b00000000000000000111110101100101;
assign LUT_4[41655] = 32'b00000000000000000001000001011101;
assign LUT_4[41656] = 32'b00000000000000000100100110111010;
assign LUT_4[41657] = 32'b11111111111111111101110010110010;
assign LUT_4[41658] = 32'b00000000000000000100000001011110;
assign LUT_4[41659] = 32'b11111111111111111101001101010110;
assign LUT_4[41660] = 32'b00000000000000000001100111010110;
assign LUT_4[41661] = 32'b11111111111111111010110011001110;
assign LUT_4[41662] = 32'b00000000000000000001000001111010;
assign LUT_4[41663] = 32'b11111111111111111010001101110010;
assign LUT_4[41664] = 32'b00000000000000010000100101000100;
assign LUT_4[41665] = 32'b00000000000000001001110000111100;
assign LUT_4[41666] = 32'b00000000000000001111111111101000;
assign LUT_4[41667] = 32'b00000000000000001001001011100000;
assign LUT_4[41668] = 32'b00000000000000001101100101100000;
assign LUT_4[41669] = 32'b00000000000000000110110001011000;
assign LUT_4[41670] = 32'b00000000000000001101000000000100;
assign LUT_4[41671] = 32'b00000000000000000110001011111100;
assign LUT_4[41672] = 32'b00000000000000001001110001011001;
assign LUT_4[41673] = 32'b00000000000000000010111101010001;
assign LUT_4[41674] = 32'b00000000000000001001001011111101;
assign LUT_4[41675] = 32'b00000000000000000010010111110101;
assign LUT_4[41676] = 32'b00000000000000000110110001110101;
assign LUT_4[41677] = 32'b11111111111111111111111101101101;
assign LUT_4[41678] = 32'b00000000000000000110001100011001;
assign LUT_4[41679] = 32'b11111111111111111111011000010001;
assign LUT_4[41680] = 32'b00000000000000001110010110110010;
assign LUT_4[41681] = 32'b00000000000000000111100010101010;
assign LUT_4[41682] = 32'b00000000000000001101110001010110;
assign LUT_4[41683] = 32'b00000000000000000110111101001110;
assign LUT_4[41684] = 32'b00000000000000001011010111001110;
assign LUT_4[41685] = 32'b00000000000000000100100011000110;
assign LUT_4[41686] = 32'b00000000000000001010110001110010;
assign LUT_4[41687] = 32'b00000000000000000011111101101010;
assign LUT_4[41688] = 32'b00000000000000000111100011000111;
assign LUT_4[41689] = 32'b00000000000000000000101110111111;
assign LUT_4[41690] = 32'b00000000000000000110111101101011;
assign LUT_4[41691] = 32'b00000000000000000000001001100011;
assign LUT_4[41692] = 32'b00000000000000000100100011100011;
assign LUT_4[41693] = 32'b11111111111111111101101111011011;
assign LUT_4[41694] = 32'b00000000000000000011111110000111;
assign LUT_4[41695] = 32'b11111111111111111101001001111111;
assign LUT_4[41696] = 32'b00000000000000001111000000001011;
assign LUT_4[41697] = 32'b00000000000000001000001100000011;
assign LUT_4[41698] = 32'b00000000000000001110011010101111;
assign LUT_4[41699] = 32'b00000000000000000111100110100111;
assign LUT_4[41700] = 32'b00000000000000001100000000100111;
assign LUT_4[41701] = 32'b00000000000000000101001100011111;
assign LUT_4[41702] = 32'b00000000000000001011011011001011;
assign LUT_4[41703] = 32'b00000000000000000100100111000011;
assign LUT_4[41704] = 32'b00000000000000001000001100100000;
assign LUT_4[41705] = 32'b00000000000000000001011000011000;
assign LUT_4[41706] = 32'b00000000000000000111100111000100;
assign LUT_4[41707] = 32'b00000000000000000000110010111100;
assign LUT_4[41708] = 32'b00000000000000000101001100111100;
assign LUT_4[41709] = 32'b11111111111111111110011000110100;
assign LUT_4[41710] = 32'b00000000000000000100100111100000;
assign LUT_4[41711] = 32'b11111111111111111101110011011000;
assign LUT_4[41712] = 32'b00000000000000001100110001111001;
assign LUT_4[41713] = 32'b00000000000000000101111101110001;
assign LUT_4[41714] = 32'b00000000000000001100001100011101;
assign LUT_4[41715] = 32'b00000000000000000101011000010101;
assign LUT_4[41716] = 32'b00000000000000001001110010010101;
assign LUT_4[41717] = 32'b00000000000000000010111110001101;
assign LUT_4[41718] = 32'b00000000000000001001001100111001;
assign LUT_4[41719] = 32'b00000000000000000010011000110001;
assign LUT_4[41720] = 32'b00000000000000000101111110001110;
assign LUT_4[41721] = 32'b11111111111111111111001010000110;
assign LUT_4[41722] = 32'b00000000000000000101011000110010;
assign LUT_4[41723] = 32'b11111111111111111110100100101010;
assign LUT_4[41724] = 32'b00000000000000000010111110101010;
assign LUT_4[41725] = 32'b11111111111111111100001010100010;
assign LUT_4[41726] = 32'b00000000000000000010011001001110;
assign LUT_4[41727] = 32'b11111111111111111011100101000110;
assign LUT_4[41728] = 32'b00000000000000010001100011001011;
assign LUT_4[41729] = 32'b00000000000000001010101111000011;
assign LUT_4[41730] = 32'b00000000000000010000111101101111;
assign LUT_4[41731] = 32'b00000000000000001010001001100111;
assign LUT_4[41732] = 32'b00000000000000001110100011100111;
assign LUT_4[41733] = 32'b00000000000000000111101111011111;
assign LUT_4[41734] = 32'b00000000000000001101111110001011;
assign LUT_4[41735] = 32'b00000000000000000111001010000011;
assign LUT_4[41736] = 32'b00000000000000001010101111100000;
assign LUT_4[41737] = 32'b00000000000000000011111011011000;
assign LUT_4[41738] = 32'b00000000000000001010001010000100;
assign LUT_4[41739] = 32'b00000000000000000011010101111100;
assign LUT_4[41740] = 32'b00000000000000000111101111111100;
assign LUT_4[41741] = 32'b00000000000000000000111011110100;
assign LUT_4[41742] = 32'b00000000000000000111001010100000;
assign LUT_4[41743] = 32'b00000000000000000000010110011000;
assign LUT_4[41744] = 32'b00000000000000001111010100111001;
assign LUT_4[41745] = 32'b00000000000000001000100000110001;
assign LUT_4[41746] = 32'b00000000000000001110101111011101;
assign LUT_4[41747] = 32'b00000000000000000111111011010101;
assign LUT_4[41748] = 32'b00000000000000001100010101010101;
assign LUT_4[41749] = 32'b00000000000000000101100001001101;
assign LUT_4[41750] = 32'b00000000000000001011101111111001;
assign LUT_4[41751] = 32'b00000000000000000100111011110001;
assign LUT_4[41752] = 32'b00000000000000001000100001001110;
assign LUT_4[41753] = 32'b00000000000000000001101101000110;
assign LUT_4[41754] = 32'b00000000000000000111111011110010;
assign LUT_4[41755] = 32'b00000000000000000001000111101010;
assign LUT_4[41756] = 32'b00000000000000000101100001101010;
assign LUT_4[41757] = 32'b11111111111111111110101101100010;
assign LUT_4[41758] = 32'b00000000000000000100111100001110;
assign LUT_4[41759] = 32'b11111111111111111110001000000110;
assign LUT_4[41760] = 32'b00000000000000001111111110010010;
assign LUT_4[41761] = 32'b00000000000000001001001010001010;
assign LUT_4[41762] = 32'b00000000000000001111011000110110;
assign LUT_4[41763] = 32'b00000000000000001000100100101110;
assign LUT_4[41764] = 32'b00000000000000001100111110101110;
assign LUT_4[41765] = 32'b00000000000000000110001010100110;
assign LUT_4[41766] = 32'b00000000000000001100011001010010;
assign LUT_4[41767] = 32'b00000000000000000101100101001010;
assign LUT_4[41768] = 32'b00000000000000001001001010100111;
assign LUT_4[41769] = 32'b00000000000000000010010110011111;
assign LUT_4[41770] = 32'b00000000000000001000100101001011;
assign LUT_4[41771] = 32'b00000000000000000001110001000011;
assign LUT_4[41772] = 32'b00000000000000000110001011000011;
assign LUT_4[41773] = 32'b11111111111111111111010110111011;
assign LUT_4[41774] = 32'b00000000000000000101100101100111;
assign LUT_4[41775] = 32'b11111111111111111110110001011111;
assign LUT_4[41776] = 32'b00000000000000001101110000000000;
assign LUT_4[41777] = 32'b00000000000000000110111011111000;
assign LUT_4[41778] = 32'b00000000000000001101001010100100;
assign LUT_4[41779] = 32'b00000000000000000110010110011100;
assign LUT_4[41780] = 32'b00000000000000001010110000011100;
assign LUT_4[41781] = 32'b00000000000000000011111100010100;
assign LUT_4[41782] = 32'b00000000000000001010001011000000;
assign LUT_4[41783] = 32'b00000000000000000011010110111000;
assign LUT_4[41784] = 32'b00000000000000000110111100010101;
assign LUT_4[41785] = 32'b00000000000000000000001000001101;
assign LUT_4[41786] = 32'b00000000000000000110010110111001;
assign LUT_4[41787] = 32'b11111111111111111111100010110001;
assign LUT_4[41788] = 32'b00000000000000000011111100110001;
assign LUT_4[41789] = 32'b11111111111111111101001000101001;
assign LUT_4[41790] = 32'b00000000000000000011010111010101;
assign LUT_4[41791] = 32'b11111111111111111100100011001101;
assign LUT_4[41792] = 32'b00000000000000010010111010011111;
assign LUT_4[41793] = 32'b00000000000000001100000110010111;
assign LUT_4[41794] = 32'b00000000000000010010010101000011;
assign LUT_4[41795] = 32'b00000000000000001011100000111011;
assign LUT_4[41796] = 32'b00000000000000001111111010111011;
assign LUT_4[41797] = 32'b00000000000000001001000110110011;
assign LUT_4[41798] = 32'b00000000000000001111010101011111;
assign LUT_4[41799] = 32'b00000000000000001000100001010111;
assign LUT_4[41800] = 32'b00000000000000001100000110110100;
assign LUT_4[41801] = 32'b00000000000000000101010010101100;
assign LUT_4[41802] = 32'b00000000000000001011100001011000;
assign LUT_4[41803] = 32'b00000000000000000100101101010000;
assign LUT_4[41804] = 32'b00000000000000001001000111010000;
assign LUT_4[41805] = 32'b00000000000000000010010011001000;
assign LUT_4[41806] = 32'b00000000000000001000100001110100;
assign LUT_4[41807] = 32'b00000000000000000001101101101100;
assign LUT_4[41808] = 32'b00000000000000010000101100001101;
assign LUT_4[41809] = 32'b00000000000000001001111000000101;
assign LUT_4[41810] = 32'b00000000000000010000000110110001;
assign LUT_4[41811] = 32'b00000000000000001001010010101001;
assign LUT_4[41812] = 32'b00000000000000001101101100101001;
assign LUT_4[41813] = 32'b00000000000000000110111000100001;
assign LUT_4[41814] = 32'b00000000000000001101000111001101;
assign LUT_4[41815] = 32'b00000000000000000110010011000101;
assign LUT_4[41816] = 32'b00000000000000001001111000100010;
assign LUT_4[41817] = 32'b00000000000000000011000100011010;
assign LUT_4[41818] = 32'b00000000000000001001010011000110;
assign LUT_4[41819] = 32'b00000000000000000010011110111110;
assign LUT_4[41820] = 32'b00000000000000000110111000111110;
assign LUT_4[41821] = 32'b00000000000000000000000100110110;
assign LUT_4[41822] = 32'b00000000000000000110010011100010;
assign LUT_4[41823] = 32'b11111111111111111111011111011010;
assign LUT_4[41824] = 32'b00000000000000010001010101100110;
assign LUT_4[41825] = 32'b00000000000000001010100001011110;
assign LUT_4[41826] = 32'b00000000000000010000110000001010;
assign LUT_4[41827] = 32'b00000000000000001001111100000010;
assign LUT_4[41828] = 32'b00000000000000001110010110000010;
assign LUT_4[41829] = 32'b00000000000000000111100001111010;
assign LUT_4[41830] = 32'b00000000000000001101110000100110;
assign LUT_4[41831] = 32'b00000000000000000110111100011110;
assign LUT_4[41832] = 32'b00000000000000001010100001111011;
assign LUT_4[41833] = 32'b00000000000000000011101101110011;
assign LUT_4[41834] = 32'b00000000000000001001111100011111;
assign LUT_4[41835] = 32'b00000000000000000011001000010111;
assign LUT_4[41836] = 32'b00000000000000000111100010010111;
assign LUT_4[41837] = 32'b00000000000000000000101110001111;
assign LUT_4[41838] = 32'b00000000000000000110111100111011;
assign LUT_4[41839] = 32'b00000000000000000000001000110011;
assign LUT_4[41840] = 32'b00000000000000001111000111010100;
assign LUT_4[41841] = 32'b00000000000000001000010011001100;
assign LUT_4[41842] = 32'b00000000000000001110100001111000;
assign LUT_4[41843] = 32'b00000000000000000111101101110000;
assign LUT_4[41844] = 32'b00000000000000001100000111110000;
assign LUT_4[41845] = 32'b00000000000000000101010011101000;
assign LUT_4[41846] = 32'b00000000000000001011100010010100;
assign LUT_4[41847] = 32'b00000000000000000100101110001100;
assign LUT_4[41848] = 32'b00000000000000001000010011101001;
assign LUT_4[41849] = 32'b00000000000000000001011111100001;
assign LUT_4[41850] = 32'b00000000000000000111101110001101;
assign LUT_4[41851] = 32'b00000000000000000000111010000101;
assign LUT_4[41852] = 32'b00000000000000000101010100000101;
assign LUT_4[41853] = 32'b11111111111111111110011111111101;
assign LUT_4[41854] = 32'b00000000000000000100101110101001;
assign LUT_4[41855] = 32'b11111111111111111101111010100001;
assign LUT_4[41856] = 32'b00000000000000010100001001010011;
assign LUT_4[41857] = 32'b00000000000000001101010101001011;
assign LUT_4[41858] = 32'b00000000000000010011100011110111;
assign LUT_4[41859] = 32'b00000000000000001100101111101111;
assign LUT_4[41860] = 32'b00000000000000010001001001101111;
assign LUT_4[41861] = 32'b00000000000000001010010101100111;
assign LUT_4[41862] = 32'b00000000000000010000100100010011;
assign LUT_4[41863] = 32'b00000000000000001001110000001011;
assign LUT_4[41864] = 32'b00000000000000001101010101101000;
assign LUT_4[41865] = 32'b00000000000000000110100001100000;
assign LUT_4[41866] = 32'b00000000000000001100110000001100;
assign LUT_4[41867] = 32'b00000000000000000101111100000100;
assign LUT_4[41868] = 32'b00000000000000001010010110000100;
assign LUT_4[41869] = 32'b00000000000000000011100001111100;
assign LUT_4[41870] = 32'b00000000000000001001110000101000;
assign LUT_4[41871] = 32'b00000000000000000010111100100000;
assign LUT_4[41872] = 32'b00000000000000010001111011000001;
assign LUT_4[41873] = 32'b00000000000000001011000110111001;
assign LUT_4[41874] = 32'b00000000000000010001010101100101;
assign LUT_4[41875] = 32'b00000000000000001010100001011101;
assign LUT_4[41876] = 32'b00000000000000001110111011011101;
assign LUT_4[41877] = 32'b00000000000000001000000111010101;
assign LUT_4[41878] = 32'b00000000000000001110010110000001;
assign LUT_4[41879] = 32'b00000000000000000111100001111001;
assign LUT_4[41880] = 32'b00000000000000001011000111010110;
assign LUT_4[41881] = 32'b00000000000000000100010011001110;
assign LUT_4[41882] = 32'b00000000000000001010100001111010;
assign LUT_4[41883] = 32'b00000000000000000011101101110010;
assign LUT_4[41884] = 32'b00000000000000001000000111110010;
assign LUT_4[41885] = 32'b00000000000000000001010011101010;
assign LUT_4[41886] = 32'b00000000000000000111100010010110;
assign LUT_4[41887] = 32'b00000000000000000000101110001110;
assign LUT_4[41888] = 32'b00000000000000010010100100011010;
assign LUT_4[41889] = 32'b00000000000000001011110000010010;
assign LUT_4[41890] = 32'b00000000000000010001111110111110;
assign LUT_4[41891] = 32'b00000000000000001011001010110110;
assign LUT_4[41892] = 32'b00000000000000001111100100110110;
assign LUT_4[41893] = 32'b00000000000000001000110000101110;
assign LUT_4[41894] = 32'b00000000000000001110111111011010;
assign LUT_4[41895] = 32'b00000000000000001000001011010010;
assign LUT_4[41896] = 32'b00000000000000001011110000101111;
assign LUT_4[41897] = 32'b00000000000000000100111100100111;
assign LUT_4[41898] = 32'b00000000000000001011001011010011;
assign LUT_4[41899] = 32'b00000000000000000100010111001011;
assign LUT_4[41900] = 32'b00000000000000001000110001001011;
assign LUT_4[41901] = 32'b00000000000000000001111101000011;
assign LUT_4[41902] = 32'b00000000000000001000001011101111;
assign LUT_4[41903] = 32'b00000000000000000001010111100111;
assign LUT_4[41904] = 32'b00000000000000010000010110001000;
assign LUT_4[41905] = 32'b00000000000000001001100010000000;
assign LUT_4[41906] = 32'b00000000000000001111110000101100;
assign LUT_4[41907] = 32'b00000000000000001000111100100100;
assign LUT_4[41908] = 32'b00000000000000001101010110100100;
assign LUT_4[41909] = 32'b00000000000000000110100010011100;
assign LUT_4[41910] = 32'b00000000000000001100110001001000;
assign LUT_4[41911] = 32'b00000000000000000101111101000000;
assign LUT_4[41912] = 32'b00000000000000001001100010011101;
assign LUT_4[41913] = 32'b00000000000000000010101110010101;
assign LUT_4[41914] = 32'b00000000000000001000111101000001;
assign LUT_4[41915] = 32'b00000000000000000010001000111001;
assign LUT_4[41916] = 32'b00000000000000000110100010111001;
assign LUT_4[41917] = 32'b11111111111111111111101110110001;
assign LUT_4[41918] = 32'b00000000000000000101111101011101;
assign LUT_4[41919] = 32'b11111111111111111111001001010101;
assign LUT_4[41920] = 32'b00000000000000010101100000100111;
assign LUT_4[41921] = 32'b00000000000000001110101100011111;
assign LUT_4[41922] = 32'b00000000000000010100111011001011;
assign LUT_4[41923] = 32'b00000000000000001110000111000011;
assign LUT_4[41924] = 32'b00000000000000010010100001000011;
assign LUT_4[41925] = 32'b00000000000000001011101100111011;
assign LUT_4[41926] = 32'b00000000000000010001111011100111;
assign LUT_4[41927] = 32'b00000000000000001011000111011111;
assign LUT_4[41928] = 32'b00000000000000001110101100111100;
assign LUT_4[41929] = 32'b00000000000000000111111000110100;
assign LUT_4[41930] = 32'b00000000000000001110000111100000;
assign LUT_4[41931] = 32'b00000000000000000111010011011000;
assign LUT_4[41932] = 32'b00000000000000001011101101011000;
assign LUT_4[41933] = 32'b00000000000000000100111001010000;
assign LUT_4[41934] = 32'b00000000000000001011000111111100;
assign LUT_4[41935] = 32'b00000000000000000100010011110100;
assign LUT_4[41936] = 32'b00000000000000010011010010010101;
assign LUT_4[41937] = 32'b00000000000000001100011110001101;
assign LUT_4[41938] = 32'b00000000000000010010101100111001;
assign LUT_4[41939] = 32'b00000000000000001011111000110001;
assign LUT_4[41940] = 32'b00000000000000010000010010110001;
assign LUT_4[41941] = 32'b00000000000000001001011110101001;
assign LUT_4[41942] = 32'b00000000000000001111101101010101;
assign LUT_4[41943] = 32'b00000000000000001000111001001101;
assign LUT_4[41944] = 32'b00000000000000001100011110101010;
assign LUT_4[41945] = 32'b00000000000000000101101010100010;
assign LUT_4[41946] = 32'b00000000000000001011111001001110;
assign LUT_4[41947] = 32'b00000000000000000101000101000110;
assign LUT_4[41948] = 32'b00000000000000001001011111000110;
assign LUT_4[41949] = 32'b00000000000000000010101010111110;
assign LUT_4[41950] = 32'b00000000000000001000111001101010;
assign LUT_4[41951] = 32'b00000000000000000010000101100010;
assign LUT_4[41952] = 32'b00000000000000010011111011101110;
assign LUT_4[41953] = 32'b00000000000000001101000111100110;
assign LUT_4[41954] = 32'b00000000000000010011010110010010;
assign LUT_4[41955] = 32'b00000000000000001100100010001010;
assign LUT_4[41956] = 32'b00000000000000010000111100001010;
assign LUT_4[41957] = 32'b00000000000000001010001000000010;
assign LUT_4[41958] = 32'b00000000000000010000010110101110;
assign LUT_4[41959] = 32'b00000000000000001001100010100110;
assign LUT_4[41960] = 32'b00000000000000001101001000000011;
assign LUT_4[41961] = 32'b00000000000000000110010011111011;
assign LUT_4[41962] = 32'b00000000000000001100100010100111;
assign LUT_4[41963] = 32'b00000000000000000101101110011111;
assign LUT_4[41964] = 32'b00000000000000001010001000011111;
assign LUT_4[41965] = 32'b00000000000000000011010100010111;
assign LUT_4[41966] = 32'b00000000000000001001100011000011;
assign LUT_4[41967] = 32'b00000000000000000010101110111011;
assign LUT_4[41968] = 32'b00000000000000010001101101011100;
assign LUT_4[41969] = 32'b00000000000000001010111001010100;
assign LUT_4[41970] = 32'b00000000000000010001001000000000;
assign LUT_4[41971] = 32'b00000000000000001010010011111000;
assign LUT_4[41972] = 32'b00000000000000001110101101111000;
assign LUT_4[41973] = 32'b00000000000000000111111001110000;
assign LUT_4[41974] = 32'b00000000000000001110001000011100;
assign LUT_4[41975] = 32'b00000000000000000111010100010100;
assign LUT_4[41976] = 32'b00000000000000001010111001110001;
assign LUT_4[41977] = 32'b00000000000000000100000101101001;
assign LUT_4[41978] = 32'b00000000000000001010010100010101;
assign LUT_4[41979] = 32'b00000000000000000011100000001101;
assign LUT_4[41980] = 32'b00000000000000000111111010001101;
assign LUT_4[41981] = 32'b00000000000000000001000110000101;
assign LUT_4[41982] = 32'b00000000000000000111010100110001;
assign LUT_4[41983] = 32'b00000000000000000000100000101001;
assign LUT_4[41984] = 32'b00000000000000001111001101111111;
assign LUT_4[41985] = 32'b00000000000000001000011001110111;
assign LUT_4[41986] = 32'b00000000000000001110101000100011;
assign LUT_4[41987] = 32'b00000000000000000111110100011011;
assign LUT_4[41988] = 32'b00000000000000001100001110011011;
assign LUT_4[41989] = 32'b00000000000000000101011010010011;
assign LUT_4[41990] = 32'b00000000000000001011101000111111;
assign LUT_4[41991] = 32'b00000000000000000100110100110111;
assign LUT_4[41992] = 32'b00000000000000001000011010010100;
assign LUT_4[41993] = 32'b00000000000000000001100110001100;
assign LUT_4[41994] = 32'b00000000000000000111110100111000;
assign LUT_4[41995] = 32'b00000000000000000001000000110000;
assign LUT_4[41996] = 32'b00000000000000000101011010110000;
assign LUT_4[41997] = 32'b11111111111111111110100110101000;
assign LUT_4[41998] = 32'b00000000000000000100110101010100;
assign LUT_4[41999] = 32'b11111111111111111110000001001100;
assign LUT_4[42000] = 32'b00000000000000001100111111101101;
assign LUT_4[42001] = 32'b00000000000000000110001011100101;
assign LUT_4[42002] = 32'b00000000000000001100011010010001;
assign LUT_4[42003] = 32'b00000000000000000101100110001001;
assign LUT_4[42004] = 32'b00000000000000001010000000001001;
assign LUT_4[42005] = 32'b00000000000000000011001100000001;
assign LUT_4[42006] = 32'b00000000000000001001011010101101;
assign LUT_4[42007] = 32'b00000000000000000010100110100101;
assign LUT_4[42008] = 32'b00000000000000000110001100000010;
assign LUT_4[42009] = 32'b11111111111111111111010111111010;
assign LUT_4[42010] = 32'b00000000000000000101100110100110;
assign LUT_4[42011] = 32'b11111111111111111110110010011110;
assign LUT_4[42012] = 32'b00000000000000000011001100011110;
assign LUT_4[42013] = 32'b11111111111111111100011000010110;
assign LUT_4[42014] = 32'b00000000000000000010100111000010;
assign LUT_4[42015] = 32'b11111111111111111011110010111010;
assign LUT_4[42016] = 32'b00000000000000001101101001000110;
assign LUT_4[42017] = 32'b00000000000000000110110100111110;
assign LUT_4[42018] = 32'b00000000000000001101000011101010;
assign LUT_4[42019] = 32'b00000000000000000110001111100010;
assign LUT_4[42020] = 32'b00000000000000001010101001100010;
assign LUT_4[42021] = 32'b00000000000000000011110101011010;
assign LUT_4[42022] = 32'b00000000000000001010000100000110;
assign LUT_4[42023] = 32'b00000000000000000011001111111110;
assign LUT_4[42024] = 32'b00000000000000000110110101011011;
assign LUT_4[42025] = 32'b00000000000000000000000001010011;
assign LUT_4[42026] = 32'b00000000000000000110001111111111;
assign LUT_4[42027] = 32'b11111111111111111111011011110111;
assign LUT_4[42028] = 32'b00000000000000000011110101110111;
assign LUT_4[42029] = 32'b11111111111111111101000001101111;
assign LUT_4[42030] = 32'b00000000000000000011010000011011;
assign LUT_4[42031] = 32'b11111111111111111100011100010011;
assign LUT_4[42032] = 32'b00000000000000001011011010110100;
assign LUT_4[42033] = 32'b00000000000000000100100110101100;
assign LUT_4[42034] = 32'b00000000000000001010110101011000;
assign LUT_4[42035] = 32'b00000000000000000100000001010000;
assign LUT_4[42036] = 32'b00000000000000001000011011010000;
assign LUT_4[42037] = 32'b00000000000000000001100111001000;
assign LUT_4[42038] = 32'b00000000000000000111110101110100;
assign LUT_4[42039] = 32'b00000000000000000001000001101100;
assign LUT_4[42040] = 32'b00000000000000000100100111001001;
assign LUT_4[42041] = 32'b11111111111111111101110011000001;
assign LUT_4[42042] = 32'b00000000000000000100000001101101;
assign LUT_4[42043] = 32'b11111111111111111101001101100101;
assign LUT_4[42044] = 32'b00000000000000000001100111100101;
assign LUT_4[42045] = 32'b11111111111111111010110011011101;
assign LUT_4[42046] = 32'b00000000000000000001000010001001;
assign LUT_4[42047] = 32'b11111111111111111010001110000001;
assign LUT_4[42048] = 32'b00000000000000010000100101010011;
assign LUT_4[42049] = 32'b00000000000000001001110001001011;
assign LUT_4[42050] = 32'b00000000000000001111111111110111;
assign LUT_4[42051] = 32'b00000000000000001001001011101111;
assign LUT_4[42052] = 32'b00000000000000001101100101101111;
assign LUT_4[42053] = 32'b00000000000000000110110001100111;
assign LUT_4[42054] = 32'b00000000000000001101000000010011;
assign LUT_4[42055] = 32'b00000000000000000110001100001011;
assign LUT_4[42056] = 32'b00000000000000001001110001101000;
assign LUT_4[42057] = 32'b00000000000000000010111101100000;
assign LUT_4[42058] = 32'b00000000000000001001001100001100;
assign LUT_4[42059] = 32'b00000000000000000010011000000100;
assign LUT_4[42060] = 32'b00000000000000000110110010000100;
assign LUT_4[42061] = 32'b11111111111111111111111101111100;
assign LUT_4[42062] = 32'b00000000000000000110001100101000;
assign LUT_4[42063] = 32'b11111111111111111111011000100000;
assign LUT_4[42064] = 32'b00000000000000001110010111000001;
assign LUT_4[42065] = 32'b00000000000000000111100010111001;
assign LUT_4[42066] = 32'b00000000000000001101110001100101;
assign LUT_4[42067] = 32'b00000000000000000110111101011101;
assign LUT_4[42068] = 32'b00000000000000001011010111011101;
assign LUT_4[42069] = 32'b00000000000000000100100011010101;
assign LUT_4[42070] = 32'b00000000000000001010110010000001;
assign LUT_4[42071] = 32'b00000000000000000011111101111001;
assign LUT_4[42072] = 32'b00000000000000000111100011010110;
assign LUT_4[42073] = 32'b00000000000000000000101111001110;
assign LUT_4[42074] = 32'b00000000000000000110111101111010;
assign LUT_4[42075] = 32'b00000000000000000000001001110010;
assign LUT_4[42076] = 32'b00000000000000000100100011110010;
assign LUT_4[42077] = 32'b11111111111111111101101111101010;
assign LUT_4[42078] = 32'b00000000000000000011111110010110;
assign LUT_4[42079] = 32'b11111111111111111101001010001110;
assign LUT_4[42080] = 32'b00000000000000001111000000011010;
assign LUT_4[42081] = 32'b00000000000000001000001100010010;
assign LUT_4[42082] = 32'b00000000000000001110011010111110;
assign LUT_4[42083] = 32'b00000000000000000111100110110110;
assign LUT_4[42084] = 32'b00000000000000001100000000110110;
assign LUT_4[42085] = 32'b00000000000000000101001100101110;
assign LUT_4[42086] = 32'b00000000000000001011011011011010;
assign LUT_4[42087] = 32'b00000000000000000100100111010010;
assign LUT_4[42088] = 32'b00000000000000001000001100101111;
assign LUT_4[42089] = 32'b00000000000000000001011000100111;
assign LUT_4[42090] = 32'b00000000000000000111100111010011;
assign LUT_4[42091] = 32'b00000000000000000000110011001011;
assign LUT_4[42092] = 32'b00000000000000000101001101001011;
assign LUT_4[42093] = 32'b11111111111111111110011001000011;
assign LUT_4[42094] = 32'b00000000000000000100100111101111;
assign LUT_4[42095] = 32'b11111111111111111101110011100111;
assign LUT_4[42096] = 32'b00000000000000001100110010001000;
assign LUT_4[42097] = 32'b00000000000000000101111110000000;
assign LUT_4[42098] = 32'b00000000000000001100001100101100;
assign LUT_4[42099] = 32'b00000000000000000101011000100100;
assign LUT_4[42100] = 32'b00000000000000001001110010100100;
assign LUT_4[42101] = 32'b00000000000000000010111110011100;
assign LUT_4[42102] = 32'b00000000000000001001001101001000;
assign LUT_4[42103] = 32'b00000000000000000010011001000000;
assign LUT_4[42104] = 32'b00000000000000000101111110011101;
assign LUT_4[42105] = 32'b11111111111111111111001010010101;
assign LUT_4[42106] = 32'b00000000000000000101011001000001;
assign LUT_4[42107] = 32'b11111111111111111110100100111001;
assign LUT_4[42108] = 32'b00000000000000000010111110111001;
assign LUT_4[42109] = 32'b11111111111111111100001010110001;
assign LUT_4[42110] = 32'b00000000000000000010011001011101;
assign LUT_4[42111] = 32'b11111111111111111011100101010101;
assign LUT_4[42112] = 32'b00000000000000010001110100000111;
assign LUT_4[42113] = 32'b00000000000000001010111111111111;
assign LUT_4[42114] = 32'b00000000000000010001001110101011;
assign LUT_4[42115] = 32'b00000000000000001010011010100011;
assign LUT_4[42116] = 32'b00000000000000001110110100100011;
assign LUT_4[42117] = 32'b00000000000000001000000000011011;
assign LUT_4[42118] = 32'b00000000000000001110001111000111;
assign LUT_4[42119] = 32'b00000000000000000111011010111111;
assign LUT_4[42120] = 32'b00000000000000001011000000011100;
assign LUT_4[42121] = 32'b00000000000000000100001100010100;
assign LUT_4[42122] = 32'b00000000000000001010011011000000;
assign LUT_4[42123] = 32'b00000000000000000011100110111000;
assign LUT_4[42124] = 32'b00000000000000001000000000111000;
assign LUT_4[42125] = 32'b00000000000000000001001100110000;
assign LUT_4[42126] = 32'b00000000000000000111011011011100;
assign LUT_4[42127] = 32'b00000000000000000000100111010100;
assign LUT_4[42128] = 32'b00000000000000001111100101110101;
assign LUT_4[42129] = 32'b00000000000000001000110001101101;
assign LUT_4[42130] = 32'b00000000000000001111000000011001;
assign LUT_4[42131] = 32'b00000000000000001000001100010001;
assign LUT_4[42132] = 32'b00000000000000001100100110010001;
assign LUT_4[42133] = 32'b00000000000000000101110010001001;
assign LUT_4[42134] = 32'b00000000000000001100000000110101;
assign LUT_4[42135] = 32'b00000000000000000101001100101101;
assign LUT_4[42136] = 32'b00000000000000001000110010001010;
assign LUT_4[42137] = 32'b00000000000000000001111110000010;
assign LUT_4[42138] = 32'b00000000000000001000001100101110;
assign LUT_4[42139] = 32'b00000000000000000001011000100110;
assign LUT_4[42140] = 32'b00000000000000000101110010100110;
assign LUT_4[42141] = 32'b11111111111111111110111110011110;
assign LUT_4[42142] = 32'b00000000000000000101001101001010;
assign LUT_4[42143] = 32'b11111111111111111110011001000010;
assign LUT_4[42144] = 32'b00000000000000010000001111001110;
assign LUT_4[42145] = 32'b00000000000000001001011011000110;
assign LUT_4[42146] = 32'b00000000000000001111101001110010;
assign LUT_4[42147] = 32'b00000000000000001000110101101010;
assign LUT_4[42148] = 32'b00000000000000001101001111101010;
assign LUT_4[42149] = 32'b00000000000000000110011011100010;
assign LUT_4[42150] = 32'b00000000000000001100101010001110;
assign LUT_4[42151] = 32'b00000000000000000101110110000110;
assign LUT_4[42152] = 32'b00000000000000001001011011100011;
assign LUT_4[42153] = 32'b00000000000000000010100111011011;
assign LUT_4[42154] = 32'b00000000000000001000110110000111;
assign LUT_4[42155] = 32'b00000000000000000010000001111111;
assign LUT_4[42156] = 32'b00000000000000000110011011111111;
assign LUT_4[42157] = 32'b11111111111111111111100111110111;
assign LUT_4[42158] = 32'b00000000000000000101110110100011;
assign LUT_4[42159] = 32'b11111111111111111111000010011011;
assign LUT_4[42160] = 32'b00000000000000001110000000111100;
assign LUT_4[42161] = 32'b00000000000000000111001100110100;
assign LUT_4[42162] = 32'b00000000000000001101011011100000;
assign LUT_4[42163] = 32'b00000000000000000110100111011000;
assign LUT_4[42164] = 32'b00000000000000001011000001011000;
assign LUT_4[42165] = 32'b00000000000000000100001101010000;
assign LUT_4[42166] = 32'b00000000000000001010011011111100;
assign LUT_4[42167] = 32'b00000000000000000011100111110100;
assign LUT_4[42168] = 32'b00000000000000000111001101010001;
assign LUT_4[42169] = 32'b00000000000000000000011001001001;
assign LUT_4[42170] = 32'b00000000000000000110100111110101;
assign LUT_4[42171] = 32'b11111111111111111111110011101101;
assign LUT_4[42172] = 32'b00000000000000000100001101101101;
assign LUT_4[42173] = 32'b11111111111111111101011001100101;
assign LUT_4[42174] = 32'b00000000000000000011101000010001;
assign LUT_4[42175] = 32'b11111111111111111100110100001001;
assign LUT_4[42176] = 32'b00000000000000010011001011011011;
assign LUT_4[42177] = 32'b00000000000000001100010111010011;
assign LUT_4[42178] = 32'b00000000000000010010100101111111;
assign LUT_4[42179] = 32'b00000000000000001011110001110111;
assign LUT_4[42180] = 32'b00000000000000010000001011110111;
assign LUT_4[42181] = 32'b00000000000000001001010111101111;
assign LUT_4[42182] = 32'b00000000000000001111100110011011;
assign LUT_4[42183] = 32'b00000000000000001000110010010011;
assign LUT_4[42184] = 32'b00000000000000001100010111110000;
assign LUT_4[42185] = 32'b00000000000000000101100011101000;
assign LUT_4[42186] = 32'b00000000000000001011110010010100;
assign LUT_4[42187] = 32'b00000000000000000100111110001100;
assign LUT_4[42188] = 32'b00000000000000001001011000001100;
assign LUT_4[42189] = 32'b00000000000000000010100100000100;
assign LUT_4[42190] = 32'b00000000000000001000110010110000;
assign LUT_4[42191] = 32'b00000000000000000001111110101000;
assign LUT_4[42192] = 32'b00000000000000010000111101001001;
assign LUT_4[42193] = 32'b00000000000000001010001001000001;
assign LUT_4[42194] = 32'b00000000000000010000010111101101;
assign LUT_4[42195] = 32'b00000000000000001001100011100101;
assign LUT_4[42196] = 32'b00000000000000001101111101100101;
assign LUT_4[42197] = 32'b00000000000000000111001001011101;
assign LUT_4[42198] = 32'b00000000000000001101011000001001;
assign LUT_4[42199] = 32'b00000000000000000110100100000001;
assign LUT_4[42200] = 32'b00000000000000001010001001011110;
assign LUT_4[42201] = 32'b00000000000000000011010101010110;
assign LUT_4[42202] = 32'b00000000000000001001100100000010;
assign LUT_4[42203] = 32'b00000000000000000010101111111010;
assign LUT_4[42204] = 32'b00000000000000000111001001111010;
assign LUT_4[42205] = 32'b00000000000000000000010101110010;
assign LUT_4[42206] = 32'b00000000000000000110100100011110;
assign LUT_4[42207] = 32'b11111111111111111111110000010110;
assign LUT_4[42208] = 32'b00000000000000010001100110100010;
assign LUT_4[42209] = 32'b00000000000000001010110010011010;
assign LUT_4[42210] = 32'b00000000000000010001000001000110;
assign LUT_4[42211] = 32'b00000000000000001010001100111110;
assign LUT_4[42212] = 32'b00000000000000001110100110111110;
assign LUT_4[42213] = 32'b00000000000000000111110010110110;
assign LUT_4[42214] = 32'b00000000000000001110000001100010;
assign LUT_4[42215] = 32'b00000000000000000111001101011010;
assign LUT_4[42216] = 32'b00000000000000001010110010110111;
assign LUT_4[42217] = 32'b00000000000000000011111110101111;
assign LUT_4[42218] = 32'b00000000000000001010001101011011;
assign LUT_4[42219] = 32'b00000000000000000011011001010011;
assign LUT_4[42220] = 32'b00000000000000000111110011010011;
assign LUT_4[42221] = 32'b00000000000000000000111111001011;
assign LUT_4[42222] = 32'b00000000000000000111001101110111;
assign LUT_4[42223] = 32'b00000000000000000000011001101111;
assign LUT_4[42224] = 32'b00000000000000001111011000010000;
assign LUT_4[42225] = 32'b00000000000000001000100100001000;
assign LUT_4[42226] = 32'b00000000000000001110110010110100;
assign LUT_4[42227] = 32'b00000000000000000111111110101100;
assign LUT_4[42228] = 32'b00000000000000001100011000101100;
assign LUT_4[42229] = 32'b00000000000000000101100100100100;
assign LUT_4[42230] = 32'b00000000000000001011110011010000;
assign LUT_4[42231] = 32'b00000000000000000100111111001000;
assign LUT_4[42232] = 32'b00000000000000001000100100100101;
assign LUT_4[42233] = 32'b00000000000000000001110000011101;
assign LUT_4[42234] = 32'b00000000000000000111111111001001;
assign LUT_4[42235] = 32'b00000000000000000001001011000001;
assign LUT_4[42236] = 32'b00000000000000000101100101000001;
assign LUT_4[42237] = 32'b11111111111111111110110000111001;
assign LUT_4[42238] = 32'b00000000000000000100111111100101;
assign LUT_4[42239] = 32'b11111111111111111110001011011101;
assign LUT_4[42240] = 32'b00000000000000010100001001100010;
assign LUT_4[42241] = 32'b00000000000000001101010101011010;
assign LUT_4[42242] = 32'b00000000000000010011100100000110;
assign LUT_4[42243] = 32'b00000000000000001100101111111110;
assign LUT_4[42244] = 32'b00000000000000010001001001111110;
assign LUT_4[42245] = 32'b00000000000000001010010101110110;
assign LUT_4[42246] = 32'b00000000000000010000100100100010;
assign LUT_4[42247] = 32'b00000000000000001001110000011010;
assign LUT_4[42248] = 32'b00000000000000001101010101110111;
assign LUT_4[42249] = 32'b00000000000000000110100001101111;
assign LUT_4[42250] = 32'b00000000000000001100110000011011;
assign LUT_4[42251] = 32'b00000000000000000101111100010011;
assign LUT_4[42252] = 32'b00000000000000001010010110010011;
assign LUT_4[42253] = 32'b00000000000000000011100010001011;
assign LUT_4[42254] = 32'b00000000000000001001110000110111;
assign LUT_4[42255] = 32'b00000000000000000010111100101111;
assign LUT_4[42256] = 32'b00000000000000010001111011010000;
assign LUT_4[42257] = 32'b00000000000000001011000111001000;
assign LUT_4[42258] = 32'b00000000000000010001010101110100;
assign LUT_4[42259] = 32'b00000000000000001010100001101100;
assign LUT_4[42260] = 32'b00000000000000001110111011101100;
assign LUT_4[42261] = 32'b00000000000000001000000111100100;
assign LUT_4[42262] = 32'b00000000000000001110010110010000;
assign LUT_4[42263] = 32'b00000000000000000111100010001000;
assign LUT_4[42264] = 32'b00000000000000001011000111100101;
assign LUT_4[42265] = 32'b00000000000000000100010011011101;
assign LUT_4[42266] = 32'b00000000000000001010100010001001;
assign LUT_4[42267] = 32'b00000000000000000011101110000001;
assign LUT_4[42268] = 32'b00000000000000001000001000000001;
assign LUT_4[42269] = 32'b00000000000000000001010011111001;
assign LUT_4[42270] = 32'b00000000000000000111100010100101;
assign LUT_4[42271] = 32'b00000000000000000000101110011101;
assign LUT_4[42272] = 32'b00000000000000010010100100101001;
assign LUT_4[42273] = 32'b00000000000000001011110000100001;
assign LUT_4[42274] = 32'b00000000000000010001111111001101;
assign LUT_4[42275] = 32'b00000000000000001011001011000101;
assign LUT_4[42276] = 32'b00000000000000001111100101000101;
assign LUT_4[42277] = 32'b00000000000000001000110000111101;
assign LUT_4[42278] = 32'b00000000000000001110111111101001;
assign LUT_4[42279] = 32'b00000000000000001000001011100001;
assign LUT_4[42280] = 32'b00000000000000001011110000111110;
assign LUT_4[42281] = 32'b00000000000000000100111100110110;
assign LUT_4[42282] = 32'b00000000000000001011001011100010;
assign LUT_4[42283] = 32'b00000000000000000100010111011010;
assign LUT_4[42284] = 32'b00000000000000001000110001011010;
assign LUT_4[42285] = 32'b00000000000000000001111101010010;
assign LUT_4[42286] = 32'b00000000000000001000001011111110;
assign LUT_4[42287] = 32'b00000000000000000001010111110110;
assign LUT_4[42288] = 32'b00000000000000010000010110010111;
assign LUT_4[42289] = 32'b00000000000000001001100010001111;
assign LUT_4[42290] = 32'b00000000000000001111110000111011;
assign LUT_4[42291] = 32'b00000000000000001000111100110011;
assign LUT_4[42292] = 32'b00000000000000001101010110110011;
assign LUT_4[42293] = 32'b00000000000000000110100010101011;
assign LUT_4[42294] = 32'b00000000000000001100110001010111;
assign LUT_4[42295] = 32'b00000000000000000101111101001111;
assign LUT_4[42296] = 32'b00000000000000001001100010101100;
assign LUT_4[42297] = 32'b00000000000000000010101110100100;
assign LUT_4[42298] = 32'b00000000000000001000111101010000;
assign LUT_4[42299] = 32'b00000000000000000010001001001000;
assign LUT_4[42300] = 32'b00000000000000000110100011001000;
assign LUT_4[42301] = 32'b11111111111111111111101111000000;
assign LUT_4[42302] = 32'b00000000000000000101111101101100;
assign LUT_4[42303] = 32'b11111111111111111111001001100100;
assign LUT_4[42304] = 32'b00000000000000010101100000110110;
assign LUT_4[42305] = 32'b00000000000000001110101100101110;
assign LUT_4[42306] = 32'b00000000000000010100111011011010;
assign LUT_4[42307] = 32'b00000000000000001110000111010010;
assign LUT_4[42308] = 32'b00000000000000010010100001010010;
assign LUT_4[42309] = 32'b00000000000000001011101101001010;
assign LUT_4[42310] = 32'b00000000000000010001111011110110;
assign LUT_4[42311] = 32'b00000000000000001011000111101110;
assign LUT_4[42312] = 32'b00000000000000001110101101001011;
assign LUT_4[42313] = 32'b00000000000000000111111001000011;
assign LUT_4[42314] = 32'b00000000000000001110000111101111;
assign LUT_4[42315] = 32'b00000000000000000111010011100111;
assign LUT_4[42316] = 32'b00000000000000001011101101100111;
assign LUT_4[42317] = 32'b00000000000000000100111001011111;
assign LUT_4[42318] = 32'b00000000000000001011001000001011;
assign LUT_4[42319] = 32'b00000000000000000100010100000011;
assign LUT_4[42320] = 32'b00000000000000010011010010100100;
assign LUT_4[42321] = 32'b00000000000000001100011110011100;
assign LUT_4[42322] = 32'b00000000000000010010101101001000;
assign LUT_4[42323] = 32'b00000000000000001011111001000000;
assign LUT_4[42324] = 32'b00000000000000010000010011000000;
assign LUT_4[42325] = 32'b00000000000000001001011110111000;
assign LUT_4[42326] = 32'b00000000000000001111101101100100;
assign LUT_4[42327] = 32'b00000000000000001000111001011100;
assign LUT_4[42328] = 32'b00000000000000001100011110111001;
assign LUT_4[42329] = 32'b00000000000000000101101010110001;
assign LUT_4[42330] = 32'b00000000000000001011111001011101;
assign LUT_4[42331] = 32'b00000000000000000101000101010101;
assign LUT_4[42332] = 32'b00000000000000001001011111010101;
assign LUT_4[42333] = 32'b00000000000000000010101011001101;
assign LUT_4[42334] = 32'b00000000000000001000111001111001;
assign LUT_4[42335] = 32'b00000000000000000010000101110001;
assign LUT_4[42336] = 32'b00000000000000010011111011111101;
assign LUT_4[42337] = 32'b00000000000000001101000111110101;
assign LUT_4[42338] = 32'b00000000000000010011010110100001;
assign LUT_4[42339] = 32'b00000000000000001100100010011001;
assign LUT_4[42340] = 32'b00000000000000010000111100011001;
assign LUT_4[42341] = 32'b00000000000000001010001000010001;
assign LUT_4[42342] = 32'b00000000000000010000010110111101;
assign LUT_4[42343] = 32'b00000000000000001001100010110101;
assign LUT_4[42344] = 32'b00000000000000001101001000010010;
assign LUT_4[42345] = 32'b00000000000000000110010100001010;
assign LUT_4[42346] = 32'b00000000000000001100100010110110;
assign LUT_4[42347] = 32'b00000000000000000101101110101110;
assign LUT_4[42348] = 32'b00000000000000001010001000101110;
assign LUT_4[42349] = 32'b00000000000000000011010100100110;
assign LUT_4[42350] = 32'b00000000000000001001100011010010;
assign LUT_4[42351] = 32'b00000000000000000010101111001010;
assign LUT_4[42352] = 32'b00000000000000010001101101101011;
assign LUT_4[42353] = 32'b00000000000000001010111001100011;
assign LUT_4[42354] = 32'b00000000000000010001001000001111;
assign LUT_4[42355] = 32'b00000000000000001010010100000111;
assign LUT_4[42356] = 32'b00000000000000001110101110000111;
assign LUT_4[42357] = 32'b00000000000000000111111001111111;
assign LUT_4[42358] = 32'b00000000000000001110001000101011;
assign LUT_4[42359] = 32'b00000000000000000111010100100011;
assign LUT_4[42360] = 32'b00000000000000001010111010000000;
assign LUT_4[42361] = 32'b00000000000000000100000101111000;
assign LUT_4[42362] = 32'b00000000000000001010010100100100;
assign LUT_4[42363] = 32'b00000000000000000011100000011100;
assign LUT_4[42364] = 32'b00000000000000000111111010011100;
assign LUT_4[42365] = 32'b00000000000000000001000110010100;
assign LUT_4[42366] = 32'b00000000000000000111010101000000;
assign LUT_4[42367] = 32'b00000000000000000000100000111000;
assign LUT_4[42368] = 32'b00000000000000010110101111101010;
assign LUT_4[42369] = 32'b00000000000000001111111011100010;
assign LUT_4[42370] = 32'b00000000000000010110001010001110;
assign LUT_4[42371] = 32'b00000000000000001111010110000110;
assign LUT_4[42372] = 32'b00000000000000010011110000000110;
assign LUT_4[42373] = 32'b00000000000000001100111011111110;
assign LUT_4[42374] = 32'b00000000000000010011001010101010;
assign LUT_4[42375] = 32'b00000000000000001100010110100010;
assign LUT_4[42376] = 32'b00000000000000001111111011111111;
assign LUT_4[42377] = 32'b00000000000000001001000111110111;
assign LUT_4[42378] = 32'b00000000000000001111010110100011;
assign LUT_4[42379] = 32'b00000000000000001000100010011011;
assign LUT_4[42380] = 32'b00000000000000001100111100011011;
assign LUT_4[42381] = 32'b00000000000000000110001000010011;
assign LUT_4[42382] = 32'b00000000000000001100010110111111;
assign LUT_4[42383] = 32'b00000000000000000101100010110111;
assign LUT_4[42384] = 32'b00000000000000010100100001011000;
assign LUT_4[42385] = 32'b00000000000000001101101101010000;
assign LUT_4[42386] = 32'b00000000000000010011111011111100;
assign LUT_4[42387] = 32'b00000000000000001101000111110100;
assign LUT_4[42388] = 32'b00000000000000010001100001110100;
assign LUT_4[42389] = 32'b00000000000000001010101101101100;
assign LUT_4[42390] = 32'b00000000000000010000111100011000;
assign LUT_4[42391] = 32'b00000000000000001010001000010000;
assign LUT_4[42392] = 32'b00000000000000001101101101101101;
assign LUT_4[42393] = 32'b00000000000000000110111001100101;
assign LUT_4[42394] = 32'b00000000000000001101001000010001;
assign LUT_4[42395] = 32'b00000000000000000110010100001001;
assign LUT_4[42396] = 32'b00000000000000001010101110001001;
assign LUT_4[42397] = 32'b00000000000000000011111010000001;
assign LUT_4[42398] = 32'b00000000000000001010001000101101;
assign LUT_4[42399] = 32'b00000000000000000011010100100101;
assign LUT_4[42400] = 32'b00000000000000010101001010110001;
assign LUT_4[42401] = 32'b00000000000000001110010110101001;
assign LUT_4[42402] = 32'b00000000000000010100100101010101;
assign LUT_4[42403] = 32'b00000000000000001101110001001101;
assign LUT_4[42404] = 32'b00000000000000010010001011001101;
assign LUT_4[42405] = 32'b00000000000000001011010111000101;
assign LUT_4[42406] = 32'b00000000000000010001100101110001;
assign LUT_4[42407] = 32'b00000000000000001010110001101001;
assign LUT_4[42408] = 32'b00000000000000001110010111000110;
assign LUT_4[42409] = 32'b00000000000000000111100010111110;
assign LUT_4[42410] = 32'b00000000000000001101110001101010;
assign LUT_4[42411] = 32'b00000000000000000110111101100010;
assign LUT_4[42412] = 32'b00000000000000001011010111100010;
assign LUT_4[42413] = 32'b00000000000000000100100011011010;
assign LUT_4[42414] = 32'b00000000000000001010110010000110;
assign LUT_4[42415] = 32'b00000000000000000011111101111110;
assign LUT_4[42416] = 32'b00000000000000010010111100011111;
assign LUT_4[42417] = 32'b00000000000000001100001000010111;
assign LUT_4[42418] = 32'b00000000000000010010010111000011;
assign LUT_4[42419] = 32'b00000000000000001011100010111011;
assign LUT_4[42420] = 32'b00000000000000001111111100111011;
assign LUT_4[42421] = 32'b00000000000000001001001000110011;
assign LUT_4[42422] = 32'b00000000000000001111010111011111;
assign LUT_4[42423] = 32'b00000000000000001000100011010111;
assign LUT_4[42424] = 32'b00000000000000001100001000110100;
assign LUT_4[42425] = 32'b00000000000000000101010100101100;
assign LUT_4[42426] = 32'b00000000000000001011100011011000;
assign LUT_4[42427] = 32'b00000000000000000100101111010000;
assign LUT_4[42428] = 32'b00000000000000001001001001010000;
assign LUT_4[42429] = 32'b00000000000000000010010101001000;
assign LUT_4[42430] = 32'b00000000000000001000100011110100;
assign LUT_4[42431] = 32'b00000000000000000001101111101100;
assign LUT_4[42432] = 32'b00000000000000011000000110111110;
assign LUT_4[42433] = 32'b00000000000000010001010010110110;
assign LUT_4[42434] = 32'b00000000000000010111100001100010;
assign LUT_4[42435] = 32'b00000000000000010000101101011010;
assign LUT_4[42436] = 32'b00000000000000010101000111011010;
assign LUT_4[42437] = 32'b00000000000000001110010011010010;
assign LUT_4[42438] = 32'b00000000000000010100100001111110;
assign LUT_4[42439] = 32'b00000000000000001101101101110110;
assign LUT_4[42440] = 32'b00000000000000010001010011010011;
assign LUT_4[42441] = 32'b00000000000000001010011111001011;
assign LUT_4[42442] = 32'b00000000000000010000101101110111;
assign LUT_4[42443] = 32'b00000000000000001001111001101111;
assign LUT_4[42444] = 32'b00000000000000001110010011101111;
assign LUT_4[42445] = 32'b00000000000000000111011111100111;
assign LUT_4[42446] = 32'b00000000000000001101101110010011;
assign LUT_4[42447] = 32'b00000000000000000110111010001011;
assign LUT_4[42448] = 32'b00000000000000010101111000101100;
assign LUT_4[42449] = 32'b00000000000000001111000100100100;
assign LUT_4[42450] = 32'b00000000000000010101010011010000;
assign LUT_4[42451] = 32'b00000000000000001110011111001000;
assign LUT_4[42452] = 32'b00000000000000010010111001001000;
assign LUT_4[42453] = 32'b00000000000000001100000101000000;
assign LUT_4[42454] = 32'b00000000000000010010010011101100;
assign LUT_4[42455] = 32'b00000000000000001011011111100100;
assign LUT_4[42456] = 32'b00000000000000001111000101000001;
assign LUT_4[42457] = 32'b00000000000000001000010000111001;
assign LUT_4[42458] = 32'b00000000000000001110011111100101;
assign LUT_4[42459] = 32'b00000000000000000111101011011101;
assign LUT_4[42460] = 32'b00000000000000001100000101011101;
assign LUT_4[42461] = 32'b00000000000000000101010001010101;
assign LUT_4[42462] = 32'b00000000000000001011100000000001;
assign LUT_4[42463] = 32'b00000000000000000100101011111001;
assign LUT_4[42464] = 32'b00000000000000010110100010000101;
assign LUT_4[42465] = 32'b00000000000000001111101101111101;
assign LUT_4[42466] = 32'b00000000000000010101111100101001;
assign LUT_4[42467] = 32'b00000000000000001111001000100001;
assign LUT_4[42468] = 32'b00000000000000010011100010100001;
assign LUT_4[42469] = 32'b00000000000000001100101110011001;
assign LUT_4[42470] = 32'b00000000000000010010111101000101;
assign LUT_4[42471] = 32'b00000000000000001100001000111101;
assign LUT_4[42472] = 32'b00000000000000001111101110011010;
assign LUT_4[42473] = 32'b00000000000000001000111010010010;
assign LUT_4[42474] = 32'b00000000000000001111001000111110;
assign LUT_4[42475] = 32'b00000000000000001000010100110110;
assign LUT_4[42476] = 32'b00000000000000001100101110110110;
assign LUT_4[42477] = 32'b00000000000000000101111010101110;
assign LUT_4[42478] = 32'b00000000000000001100001001011010;
assign LUT_4[42479] = 32'b00000000000000000101010101010010;
assign LUT_4[42480] = 32'b00000000000000010100010011110011;
assign LUT_4[42481] = 32'b00000000000000001101011111101011;
assign LUT_4[42482] = 32'b00000000000000010011101110010111;
assign LUT_4[42483] = 32'b00000000000000001100111010001111;
assign LUT_4[42484] = 32'b00000000000000010001010100001111;
assign LUT_4[42485] = 32'b00000000000000001010100000000111;
assign LUT_4[42486] = 32'b00000000000000010000101110110011;
assign LUT_4[42487] = 32'b00000000000000001001111010101011;
assign LUT_4[42488] = 32'b00000000000000001101100000001000;
assign LUT_4[42489] = 32'b00000000000000000110101100000000;
assign LUT_4[42490] = 32'b00000000000000001100111010101100;
assign LUT_4[42491] = 32'b00000000000000000110000110100100;
assign LUT_4[42492] = 32'b00000000000000001010100000100100;
assign LUT_4[42493] = 32'b00000000000000000011101100011100;
assign LUT_4[42494] = 32'b00000000000000001001111011001000;
assign LUT_4[42495] = 32'b00000000000000000011000111000000;
assign LUT_4[42496] = 32'b00000000000000001110010010000111;
assign LUT_4[42497] = 32'b00000000000000000111011101111111;
assign LUT_4[42498] = 32'b00000000000000001101101100101011;
assign LUT_4[42499] = 32'b00000000000000000110111000100011;
assign LUT_4[42500] = 32'b00000000000000001011010010100011;
assign LUT_4[42501] = 32'b00000000000000000100011110011011;
assign LUT_4[42502] = 32'b00000000000000001010101101000111;
assign LUT_4[42503] = 32'b00000000000000000011111000111111;
assign LUT_4[42504] = 32'b00000000000000000111011110011100;
assign LUT_4[42505] = 32'b00000000000000000000101010010100;
assign LUT_4[42506] = 32'b00000000000000000110111001000000;
assign LUT_4[42507] = 32'b00000000000000000000000100111000;
assign LUT_4[42508] = 32'b00000000000000000100011110111000;
assign LUT_4[42509] = 32'b11111111111111111101101010110000;
assign LUT_4[42510] = 32'b00000000000000000011111001011100;
assign LUT_4[42511] = 32'b11111111111111111101000101010100;
assign LUT_4[42512] = 32'b00000000000000001100000011110101;
assign LUT_4[42513] = 32'b00000000000000000101001111101101;
assign LUT_4[42514] = 32'b00000000000000001011011110011001;
assign LUT_4[42515] = 32'b00000000000000000100101010010001;
assign LUT_4[42516] = 32'b00000000000000001001000100010001;
assign LUT_4[42517] = 32'b00000000000000000010010000001001;
assign LUT_4[42518] = 32'b00000000000000001000011110110101;
assign LUT_4[42519] = 32'b00000000000000000001101010101101;
assign LUT_4[42520] = 32'b00000000000000000101010000001010;
assign LUT_4[42521] = 32'b11111111111111111110011100000010;
assign LUT_4[42522] = 32'b00000000000000000100101010101110;
assign LUT_4[42523] = 32'b11111111111111111101110110100110;
assign LUT_4[42524] = 32'b00000000000000000010010000100110;
assign LUT_4[42525] = 32'b11111111111111111011011100011110;
assign LUT_4[42526] = 32'b00000000000000000001101011001010;
assign LUT_4[42527] = 32'b11111111111111111010110111000010;
assign LUT_4[42528] = 32'b00000000000000001100101101001110;
assign LUT_4[42529] = 32'b00000000000000000101111001000110;
assign LUT_4[42530] = 32'b00000000000000001100000111110010;
assign LUT_4[42531] = 32'b00000000000000000101010011101010;
assign LUT_4[42532] = 32'b00000000000000001001101101101010;
assign LUT_4[42533] = 32'b00000000000000000010111001100010;
assign LUT_4[42534] = 32'b00000000000000001001001000001110;
assign LUT_4[42535] = 32'b00000000000000000010010100000110;
assign LUT_4[42536] = 32'b00000000000000000101111001100011;
assign LUT_4[42537] = 32'b11111111111111111111000101011011;
assign LUT_4[42538] = 32'b00000000000000000101010100000111;
assign LUT_4[42539] = 32'b11111111111111111110011111111111;
assign LUT_4[42540] = 32'b00000000000000000010111001111111;
assign LUT_4[42541] = 32'b11111111111111111100000101110111;
assign LUT_4[42542] = 32'b00000000000000000010010100100011;
assign LUT_4[42543] = 32'b11111111111111111011100000011011;
assign LUT_4[42544] = 32'b00000000000000001010011110111100;
assign LUT_4[42545] = 32'b00000000000000000011101010110100;
assign LUT_4[42546] = 32'b00000000000000001001111001100000;
assign LUT_4[42547] = 32'b00000000000000000011000101011000;
assign LUT_4[42548] = 32'b00000000000000000111011111011000;
assign LUT_4[42549] = 32'b00000000000000000000101011010000;
assign LUT_4[42550] = 32'b00000000000000000110111001111100;
assign LUT_4[42551] = 32'b00000000000000000000000101110100;
assign LUT_4[42552] = 32'b00000000000000000011101011010001;
assign LUT_4[42553] = 32'b11111111111111111100110111001001;
assign LUT_4[42554] = 32'b00000000000000000011000101110101;
assign LUT_4[42555] = 32'b11111111111111111100010001101101;
assign LUT_4[42556] = 32'b00000000000000000000101011101101;
assign LUT_4[42557] = 32'b11111111111111111001110111100101;
assign LUT_4[42558] = 32'b00000000000000000000000110010001;
assign LUT_4[42559] = 32'b11111111111111111001010010001001;
assign LUT_4[42560] = 32'b00000000000000001111101001011011;
assign LUT_4[42561] = 32'b00000000000000001000110101010011;
assign LUT_4[42562] = 32'b00000000000000001111000011111111;
assign LUT_4[42563] = 32'b00000000000000001000001111110111;
assign LUT_4[42564] = 32'b00000000000000001100101001110111;
assign LUT_4[42565] = 32'b00000000000000000101110101101111;
assign LUT_4[42566] = 32'b00000000000000001100000100011011;
assign LUT_4[42567] = 32'b00000000000000000101010000010011;
assign LUT_4[42568] = 32'b00000000000000001000110101110000;
assign LUT_4[42569] = 32'b00000000000000000010000001101000;
assign LUT_4[42570] = 32'b00000000000000001000010000010100;
assign LUT_4[42571] = 32'b00000000000000000001011100001100;
assign LUT_4[42572] = 32'b00000000000000000101110110001100;
assign LUT_4[42573] = 32'b11111111111111111111000010000100;
assign LUT_4[42574] = 32'b00000000000000000101010000110000;
assign LUT_4[42575] = 32'b11111111111111111110011100101000;
assign LUT_4[42576] = 32'b00000000000000001101011011001001;
assign LUT_4[42577] = 32'b00000000000000000110100111000001;
assign LUT_4[42578] = 32'b00000000000000001100110101101101;
assign LUT_4[42579] = 32'b00000000000000000110000001100101;
assign LUT_4[42580] = 32'b00000000000000001010011011100101;
assign LUT_4[42581] = 32'b00000000000000000011100111011101;
assign LUT_4[42582] = 32'b00000000000000001001110110001001;
assign LUT_4[42583] = 32'b00000000000000000011000010000001;
assign LUT_4[42584] = 32'b00000000000000000110100111011110;
assign LUT_4[42585] = 32'b11111111111111111111110011010110;
assign LUT_4[42586] = 32'b00000000000000000110000010000010;
assign LUT_4[42587] = 32'b11111111111111111111001101111010;
assign LUT_4[42588] = 32'b00000000000000000011100111111010;
assign LUT_4[42589] = 32'b11111111111111111100110011110010;
assign LUT_4[42590] = 32'b00000000000000000011000010011110;
assign LUT_4[42591] = 32'b11111111111111111100001110010110;
assign LUT_4[42592] = 32'b00000000000000001110000100100010;
assign LUT_4[42593] = 32'b00000000000000000111010000011010;
assign LUT_4[42594] = 32'b00000000000000001101011111000110;
assign LUT_4[42595] = 32'b00000000000000000110101010111110;
assign LUT_4[42596] = 32'b00000000000000001011000100111110;
assign LUT_4[42597] = 32'b00000000000000000100010000110110;
assign LUT_4[42598] = 32'b00000000000000001010011111100010;
assign LUT_4[42599] = 32'b00000000000000000011101011011010;
assign LUT_4[42600] = 32'b00000000000000000111010000110111;
assign LUT_4[42601] = 32'b00000000000000000000011100101111;
assign LUT_4[42602] = 32'b00000000000000000110101011011011;
assign LUT_4[42603] = 32'b11111111111111111111110111010011;
assign LUT_4[42604] = 32'b00000000000000000100010001010011;
assign LUT_4[42605] = 32'b11111111111111111101011101001011;
assign LUT_4[42606] = 32'b00000000000000000011101011110111;
assign LUT_4[42607] = 32'b11111111111111111100110111101111;
assign LUT_4[42608] = 32'b00000000000000001011110110010000;
assign LUT_4[42609] = 32'b00000000000000000101000010001000;
assign LUT_4[42610] = 32'b00000000000000001011010000110100;
assign LUT_4[42611] = 32'b00000000000000000100011100101100;
assign LUT_4[42612] = 32'b00000000000000001000110110101100;
assign LUT_4[42613] = 32'b00000000000000000010000010100100;
assign LUT_4[42614] = 32'b00000000000000001000010001010000;
assign LUT_4[42615] = 32'b00000000000000000001011101001000;
assign LUT_4[42616] = 32'b00000000000000000101000010100101;
assign LUT_4[42617] = 32'b11111111111111111110001110011101;
assign LUT_4[42618] = 32'b00000000000000000100011101001001;
assign LUT_4[42619] = 32'b11111111111111111101101001000001;
assign LUT_4[42620] = 32'b00000000000000000010000011000001;
assign LUT_4[42621] = 32'b11111111111111111011001110111001;
assign LUT_4[42622] = 32'b00000000000000000001011101100101;
assign LUT_4[42623] = 32'b11111111111111111010101001011101;
assign LUT_4[42624] = 32'b00000000000000010000111000001111;
assign LUT_4[42625] = 32'b00000000000000001010000100000111;
assign LUT_4[42626] = 32'b00000000000000010000010010110011;
assign LUT_4[42627] = 32'b00000000000000001001011110101011;
assign LUT_4[42628] = 32'b00000000000000001101111000101011;
assign LUT_4[42629] = 32'b00000000000000000111000100100011;
assign LUT_4[42630] = 32'b00000000000000001101010011001111;
assign LUT_4[42631] = 32'b00000000000000000110011111000111;
assign LUT_4[42632] = 32'b00000000000000001010000100100100;
assign LUT_4[42633] = 32'b00000000000000000011010000011100;
assign LUT_4[42634] = 32'b00000000000000001001011111001000;
assign LUT_4[42635] = 32'b00000000000000000010101011000000;
assign LUT_4[42636] = 32'b00000000000000000111000101000000;
assign LUT_4[42637] = 32'b00000000000000000000010000111000;
assign LUT_4[42638] = 32'b00000000000000000110011111100100;
assign LUT_4[42639] = 32'b11111111111111111111101011011100;
assign LUT_4[42640] = 32'b00000000000000001110101001111101;
assign LUT_4[42641] = 32'b00000000000000000111110101110101;
assign LUT_4[42642] = 32'b00000000000000001110000100100001;
assign LUT_4[42643] = 32'b00000000000000000111010000011001;
assign LUT_4[42644] = 32'b00000000000000001011101010011001;
assign LUT_4[42645] = 32'b00000000000000000100110110010001;
assign LUT_4[42646] = 32'b00000000000000001011000100111101;
assign LUT_4[42647] = 32'b00000000000000000100010000110101;
assign LUT_4[42648] = 32'b00000000000000000111110110010010;
assign LUT_4[42649] = 32'b00000000000000000001000010001010;
assign LUT_4[42650] = 32'b00000000000000000111010000110110;
assign LUT_4[42651] = 32'b00000000000000000000011100101110;
assign LUT_4[42652] = 32'b00000000000000000100110110101110;
assign LUT_4[42653] = 32'b11111111111111111110000010100110;
assign LUT_4[42654] = 32'b00000000000000000100010001010010;
assign LUT_4[42655] = 32'b11111111111111111101011101001010;
assign LUT_4[42656] = 32'b00000000000000001111010011010110;
assign LUT_4[42657] = 32'b00000000000000001000011111001110;
assign LUT_4[42658] = 32'b00000000000000001110101101111010;
assign LUT_4[42659] = 32'b00000000000000000111111001110010;
assign LUT_4[42660] = 32'b00000000000000001100010011110010;
assign LUT_4[42661] = 32'b00000000000000000101011111101010;
assign LUT_4[42662] = 32'b00000000000000001011101110010110;
assign LUT_4[42663] = 32'b00000000000000000100111010001110;
assign LUT_4[42664] = 32'b00000000000000001000011111101011;
assign LUT_4[42665] = 32'b00000000000000000001101011100011;
assign LUT_4[42666] = 32'b00000000000000000111111010001111;
assign LUT_4[42667] = 32'b00000000000000000001000110000111;
assign LUT_4[42668] = 32'b00000000000000000101100000000111;
assign LUT_4[42669] = 32'b11111111111111111110101011111111;
assign LUT_4[42670] = 32'b00000000000000000100111010101011;
assign LUT_4[42671] = 32'b11111111111111111110000110100011;
assign LUT_4[42672] = 32'b00000000000000001101000101000100;
assign LUT_4[42673] = 32'b00000000000000000110010000111100;
assign LUT_4[42674] = 32'b00000000000000001100011111101000;
assign LUT_4[42675] = 32'b00000000000000000101101011100000;
assign LUT_4[42676] = 32'b00000000000000001010000101100000;
assign LUT_4[42677] = 32'b00000000000000000011010001011000;
assign LUT_4[42678] = 32'b00000000000000001001100000000100;
assign LUT_4[42679] = 32'b00000000000000000010101011111100;
assign LUT_4[42680] = 32'b00000000000000000110010001011001;
assign LUT_4[42681] = 32'b11111111111111111111011101010001;
assign LUT_4[42682] = 32'b00000000000000000101101011111101;
assign LUT_4[42683] = 32'b11111111111111111110110111110101;
assign LUT_4[42684] = 32'b00000000000000000011010001110101;
assign LUT_4[42685] = 32'b11111111111111111100011101101101;
assign LUT_4[42686] = 32'b00000000000000000010101100011001;
assign LUT_4[42687] = 32'b11111111111111111011111000010001;
assign LUT_4[42688] = 32'b00000000000000010010001111100011;
assign LUT_4[42689] = 32'b00000000000000001011011011011011;
assign LUT_4[42690] = 32'b00000000000000010001101010000111;
assign LUT_4[42691] = 32'b00000000000000001010110101111111;
assign LUT_4[42692] = 32'b00000000000000001111001111111111;
assign LUT_4[42693] = 32'b00000000000000001000011011110111;
assign LUT_4[42694] = 32'b00000000000000001110101010100011;
assign LUT_4[42695] = 32'b00000000000000000111110110011011;
assign LUT_4[42696] = 32'b00000000000000001011011011111000;
assign LUT_4[42697] = 32'b00000000000000000100100111110000;
assign LUT_4[42698] = 32'b00000000000000001010110110011100;
assign LUT_4[42699] = 32'b00000000000000000100000010010100;
assign LUT_4[42700] = 32'b00000000000000001000011100010100;
assign LUT_4[42701] = 32'b00000000000000000001101000001100;
assign LUT_4[42702] = 32'b00000000000000000111110110111000;
assign LUT_4[42703] = 32'b00000000000000000001000010110000;
assign LUT_4[42704] = 32'b00000000000000010000000001010001;
assign LUT_4[42705] = 32'b00000000000000001001001101001001;
assign LUT_4[42706] = 32'b00000000000000001111011011110101;
assign LUT_4[42707] = 32'b00000000000000001000100111101101;
assign LUT_4[42708] = 32'b00000000000000001101000001101101;
assign LUT_4[42709] = 32'b00000000000000000110001101100101;
assign LUT_4[42710] = 32'b00000000000000001100011100010001;
assign LUT_4[42711] = 32'b00000000000000000101101000001001;
assign LUT_4[42712] = 32'b00000000000000001001001101100110;
assign LUT_4[42713] = 32'b00000000000000000010011001011110;
assign LUT_4[42714] = 32'b00000000000000001000101000001010;
assign LUT_4[42715] = 32'b00000000000000000001110100000010;
assign LUT_4[42716] = 32'b00000000000000000110001110000010;
assign LUT_4[42717] = 32'b11111111111111111111011001111010;
assign LUT_4[42718] = 32'b00000000000000000101101000100110;
assign LUT_4[42719] = 32'b11111111111111111110110100011110;
assign LUT_4[42720] = 32'b00000000000000010000101010101010;
assign LUT_4[42721] = 32'b00000000000000001001110110100010;
assign LUT_4[42722] = 32'b00000000000000010000000101001110;
assign LUT_4[42723] = 32'b00000000000000001001010001000110;
assign LUT_4[42724] = 32'b00000000000000001101101011000110;
assign LUT_4[42725] = 32'b00000000000000000110110110111110;
assign LUT_4[42726] = 32'b00000000000000001101000101101010;
assign LUT_4[42727] = 32'b00000000000000000110010001100010;
assign LUT_4[42728] = 32'b00000000000000001001110110111111;
assign LUT_4[42729] = 32'b00000000000000000011000010110111;
assign LUT_4[42730] = 32'b00000000000000001001010001100011;
assign LUT_4[42731] = 32'b00000000000000000010011101011011;
assign LUT_4[42732] = 32'b00000000000000000110110111011011;
assign LUT_4[42733] = 32'b00000000000000000000000011010011;
assign LUT_4[42734] = 32'b00000000000000000110010001111111;
assign LUT_4[42735] = 32'b11111111111111111111011101110111;
assign LUT_4[42736] = 32'b00000000000000001110011100011000;
assign LUT_4[42737] = 32'b00000000000000000111101000010000;
assign LUT_4[42738] = 32'b00000000000000001101110110111100;
assign LUT_4[42739] = 32'b00000000000000000111000010110100;
assign LUT_4[42740] = 32'b00000000000000001011011100110100;
assign LUT_4[42741] = 32'b00000000000000000100101000101100;
assign LUT_4[42742] = 32'b00000000000000001010110111011000;
assign LUT_4[42743] = 32'b00000000000000000100000011010000;
assign LUT_4[42744] = 32'b00000000000000000111101000101101;
assign LUT_4[42745] = 32'b00000000000000000000110100100101;
assign LUT_4[42746] = 32'b00000000000000000111000011010001;
assign LUT_4[42747] = 32'b00000000000000000000001111001001;
assign LUT_4[42748] = 32'b00000000000000000100101001001001;
assign LUT_4[42749] = 32'b11111111111111111101110101000001;
assign LUT_4[42750] = 32'b00000000000000000100000011101101;
assign LUT_4[42751] = 32'b11111111111111111101001111100101;
assign LUT_4[42752] = 32'b00000000000000010011001101101010;
assign LUT_4[42753] = 32'b00000000000000001100011001100010;
assign LUT_4[42754] = 32'b00000000000000010010101000001110;
assign LUT_4[42755] = 32'b00000000000000001011110100000110;
assign LUT_4[42756] = 32'b00000000000000010000001110000110;
assign LUT_4[42757] = 32'b00000000000000001001011001111110;
assign LUT_4[42758] = 32'b00000000000000001111101000101010;
assign LUT_4[42759] = 32'b00000000000000001000110100100010;
assign LUT_4[42760] = 32'b00000000000000001100011001111111;
assign LUT_4[42761] = 32'b00000000000000000101100101110111;
assign LUT_4[42762] = 32'b00000000000000001011110100100011;
assign LUT_4[42763] = 32'b00000000000000000101000000011011;
assign LUT_4[42764] = 32'b00000000000000001001011010011011;
assign LUT_4[42765] = 32'b00000000000000000010100110010011;
assign LUT_4[42766] = 32'b00000000000000001000110100111111;
assign LUT_4[42767] = 32'b00000000000000000010000000110111;
assign LUT_4[42768] = 32'b00000000000000010000111111011000;
assign LUT_4[42769] = 32'b00000000000000001010001011010000;
assign LUT_4[42770] = 32'b00000000000000010000011001111100;
assign LUT_4[42771] = 32'b00000000000000001001100101110100;
assign LUT_4[42772] = 32'b00000000000000001101111111110100;
assign LUT_4[42773] = 32'b00000000000000000111001011101100;
assign LUT_4[42774] = 32'b00000000000000001101011010011000;
assign LUT_4[42775] = 32'b00000000000000000110100110010000;
assign LUT_4[42776] = 32'b00000000000000001010001011101101;
assign LUT_4[42777] = 32'b00000000000000000011010111100101;
assign LUT_4[42778] = 32'b00000000000000001001100110010001;
assign LUT_4[42779] = 32'b00000000000000000010110010001001;
assign LUT_4[42780] = 32'b00000000000000000111001100001001;
assign LUT_4[42781] = 32'b00000000000000000000011000000001;
assign LUT_4[42782] = 32'b00000000000000000110100110101101;
assign LUT_4[42783] = 32'b11111111111111111111110010100101;
assign LUT_4[42784] = 32'b00000000000000010001101000110001;
assign LUT_4[42785] = 32'b00000000000000001010110100101001;
assign LUT_4[42786] = 32'b00000000000000010001000011010101;
assign LUT_4[42787] = 32'b00000000000000001010001111001101;
assign LUT_4[42788] = 32'b00000000000000001110101001001101;
assign LUT_4[42789] = 32'b00000000000000000111110101000101;
assign LUT_4[42790] = 32'b00000000000000001110000011110001;
assign LUT_4[42791] = 32'b00000000000000000111001111101001;
assign LUT_4[42792] = 32'b00000000000000001010110101000110;
assign LUT_4[42793] = 32'b00000000000000000100000000111110;
assign LUT_4[42794] = 32'b00000000000000001010001111101010;
assign LUT_4[42795] = 32'b00000000000000000011011011100010;
assign LUT_4[42796] = 32'b00000000000000000111110101100010;
assign LUT_4[42797] = 32'b00000000000000000001000001011010;
assign LUT_4[42798] = 32'b00000000000000000111010000000110;
assign LUT_4[42799] = 32'b00000000000000000000011011111110;
assign LUT_4[42800] = 32'b00000000000000001111011010011111;
assign LUT_4[42801] = 32'b00000000000000001000100110010111;
assign LUT_4[42802] = 32'b00000000000000001110110101000011;
assign LUT_4[42803] = 32'b00000000000000001000000000111011;
assign LUT_4[42804] = 32'b00000000000000001100011010111011;
assign LUT_4[42805] = 32'b00000000000000000101100110110011;
assign LUT_4[42806] = 32'b00000000000000001011110101011111;
assign LUT_4[42807] = 32'b00000000000000000101000001010111;
assign LUT_4[42808] = 32'b00000000000000001000100110110100;
assign LUT_4[42809] = 32'b00000000000000000001110010101100;
assign LUT_4[42810] = 32'b00000000000000001000000001011000;
assign LUT_4[42811] = 32'b00000000000000000001001101010000;
assign LUT_4[42812] = 32'b00000000000000000101100111010000;
assign LUT_4[42813] = 32'b11111111111111111110110011001000;
assign LUT_4[42814] = 32'b00000000000000000101000001110100;
assign LUT_4[42815] = 32'b11111111111111111110001101101100;
assign LUT_4[42816] = 32'b00000000000000010100100100111110;
assign LUT_4[42817] = 32'b00000000000000001101110000110110;
assign LUT_4[42818] = 32'b00000000000000010011111111100010;
assign LUT_4[42819] = 32'b00000000000000001101001011011010;
assign LUT_4[42820] = 32'b00000000000000010001100101011010;
assign LUT_4[42821] = 32'b00000000000000001010110001010010;
assign LUT_4[42822] = 32'b00000000000000010000111111111110;
assign LUT_4[42823] = 32'b00000000000000001010001011110110;
assign LUT_4[42824] = 32'b00000000000000001101110001010011;
assign LUT_4[42825] = 32'b00000000000000000110111101001011;
assign LUT_4[42826] = 32'b00000000000000001101001011110111;
assign LUT_4[42827] = 32'b00000000000000000110010111101111;
assign LUT_4[42828] = 32'b00000000000000001010110001101111;
assign LUT_4[42829] = 32'b00000000000000000011111101100111;
assign LUT_4[42830] = 32'b00000000000000001010001100010011;
assign LUT_4[42831] = 32'b00000000000000000011011000001011;
assign LUT_4[42832] = 32'b00000000000000010010010110101100;
assign LUT_4[42833] = 32'b00000000000000001011100010100100;
assign LUT_4[42834] = 32'b00000000000000010001110001010000;
assign LUT_4[42835] = 32'b00000000000000001010111101001000;
assign LUT_4[42836] = 32'b00000000000000001111010111001000;
assign LUT_4[42837] = 32'b00000000000000001000100011000000;
assign LUT_4[42838] = 32'b00000000000000001110110001101100;
assign LUT_4[42839] = 32'b00000000000000000111111101100100;
assign LUT_4[42840] = 32'b00000000000000001011100011000001;
assign LUT_4[42841] = 32'b00000000000000000100101110111001;
assign LUT_4[42842] = 32'b00000000000000001010111101100101;
assign LUT_4[42843] = 32'b00000000000000000100001001011101;
assign LUT_4[42844] = 32'b00000000000000001000100011011101;
assign LUT_4[42845] = 32'b00000000000000000001101111010101;
assign LUT_4[42846] = 32'b00000000000000000111111110000001;
assign LUT_4[42847] = 32'b00000000000000000001001001111001;
assign LUT_4[42848] = 32'b00000000000000010011000000000101;
assign LUT_4[42849] = 32'b00000000000000001100001011111101;
assign LUT_4[42850] = 32'b00000000000000010010011010101001;
assign LUT_4[42851] = 32'b00000000000000001011100110100001;
assign LUT_4[42852] = 32'b00000000000000010000000000100001;
assign LUT_4[42853] = 32'b00000000000000001001001100011001;
assign LUT_4[42854] = 32'b00000000000000001111011011000101;
assign LUT_4[42855] = 32'b00000000000000001000100110111101;
assign LUT_4[42856] = 32'b00000000000000001100001100011010;
assign LUT_4[42857] = 32'b00000000000000000101011000010010;
assign LUT_4[42858] = 32'b00000000000000001011100110111110;
assign LUT_4[42859] = 32'b00000000000000000100110010110110;
assign LUT_4[42860] = 32'b00000000000000001001001100110110;
assign LUT_4[42861] = 32'b00000000000000000010011000101110;
assign LUT_4[42862] = 32'b00000000000000001000100111011010;
assign LUT_4[42863] = 32'b00000000000000000001110011010010;
assign LUT_4[42864] = 32'b00000000000000010000110001110011;
assign LUT_4[42865] = 32'b00000000000000001001111101101011;
assign LUT_4[42866] = 32'b00000000000000010000001100010111;
assign LUT_4[42867] = 32'b00000000000000001001011000001111;
assign LUT_4[42868] = 32'b00000000000000001101110010001111;
assign LUT_4[42869] = 32'b00000000000000000110111110000111;
assign LUT_4[42870] = 32'b00000000000000001101001100110011;
assign LUT_4[42871] = 32'b00000000000000000110011000101011;
assign LUT_4[42872] = 32'b00000000000000001001111110001000;
assign LUT_4[42873] = 32'b00000000000000000011001010000000;
assign LUT_4[42874] = 32'b00000000000000001001011000101100;
assign LUT_4[42875] = 32'b00000000000000000010100100100100;
assign LUT_4[42876] = 32'b00000000000000000110111110100100;
assign LUT_4[42877] = 32'b00000000000000000000001010011100;
assign LUT_4[42878] = 32'b00000000000000000110011001001000;
assign LUT_4[42879] = 32'b11111111111111111111100101000000;
assign LUT_4[42880] = 32'b00000000000000010101110011110010;
assign LUT_4[42881] = 32'b00000000000000001110111111101010;
assign LUT_4[42882] = 32'b00000000000000010101001110010110;
assign LUT_4[42883] = 32'b00000000000000001110011010001110;
assign LUT_4[42884] = 32'b00000000000000010010110100001110;
assign LUT_4[42885] = 32'b00000000000000001100000000000110;
assign LUT_4[42886] = 32'b00000000000000010010001110110010;
assign LUT_4[42887] = 32'b00000000000000001011011010101010;
assign LUT_4[42888] = 32'b00000000000000001111000000000111;
assign LUT_4[42889] = 32'b00000000000000001000001011111111;
assign LUT_4[42890] = 32'b00000000000000001110011010101011;
assign LUT_4[42891] = 32'b00000000000000000111100110100011;
assign LUT_4[42892] = 32'b00000000000000001100000000100011;
assign LUT_4[42893] = 32'b00000000000000000101001100011011;
assign LUT_4[42894] = 32'b00000000000000001011011011000111;
assign LUT_4[42895] = 32'b00000000000000000100100110111111;
assign LUT_4[42896] = 32'b00000000000000010011100101100000;
assign LUT_4[42897] = 32'b00000000000000001100110001011000;
assign LUT_4[42898] = 32'b00000000000000010011000000000100;
assign LUT_4[42899] = 32'b00000000000000001100001011111100;
assign LUT_4[42900] = 32'b00000000000000010000100101111100;
assign LUT_4[42901] = 32'b00000000000000001001110001110100;
assign LUT_4[42902] = 32'b00000000000000010000000000100000;
assign LUT_4[42903] = 32'b00000000000000001001001100011000;
assign LUT_4[42904] = 32'b00000000000000001100110001110101;
assign LUT_4[42905] = 32'b00000000000000000101111101101101;
assign LUT_4[42906] = 32'b00000000000000001100001100011001;
assign LUT_4[42907] = 32'b00000000000000000101011000010001;
assign LUT_4[42908] = 32'b00000000000000001001110010010001;
assign LUT_4[42909] = 32'b00000000000000000010111110001001;
assign LUT_4[42910] = 32'b00000000000000001001001100110101;
assign LUT_4[42911] = 32'b00000000000000000010011000101101;
assign LUT_4[42912] = 32'b00000000000000010100001110111001;
assign LUT_4[42913] = 32'b00000000000000001101011010110001;
assign LUT_4[42914] = 32'b00000000000000010011101001011101;
assign LUT_4[42915] = 32'b00000000000000001100110101010101;
assign LUT_4[42916] = 32'b00000000000000010001001111010101;
assign LUT_4[42917] = 32'b00000000000000001010011011001101;
assign LUT_4[42918] = 32'b00000000000000010000101001111001;
assign LUT_4[42919] = 32'b00000000000000001001110101110001;
assign LUT_4[42920] = 32'b00000000000000001101011011001110;
assign LUT_4[42921] = 32'b00000000000000000110100111000110;
assign LUT_4[42922] = 32'b00000000000000001100110101110010;
assign LUT_4[42923] = 32'b00000000000000000110000001101010;
assign LUT_4[42924] = 32'b00000000000000001010011011101010;
assign LUT_4[42925] = 32'b00000000000000000011100111100010;
assign LUT_4[42926] = 32'b00000000000000001001110110001110;
assign LUT_4[42927] = 32'b00000000000000000011000010000110;
assign LUT_4[42928] = 32'b00000000000000010010000000100111;
assign LUT_4[42929] = 32'b00000000000000001011001100011111;
assign LUT_4[42930] = 32'b00000000000000010001011011001011;
assign LUT_4[42931] = 32'b00000000000000001010100111000011;
assign LUT_4[42932] = 32'b00000000000000001111000001000011;
assign LUT_4[42933] = 32'b00000000000000001000001100111011;
assign LUT_4[42934] = 32'b00000000000000001110011011100111;
assign LUT_4[42935] = 32'b00000000000000000111100111011111;
assign LUT_4[42936] = 32'b00000000000000001011001100111100;
assign LUT_4[42937] = 32'b00000000000000000100011000110100;
assign LUT_4[42938] = 32'b00000000000000001010100111100000;
assign LUT_4[42939] = 32'b00000000000000000011110011011000;
assign LUT_4[42940] = 32'b00000000000000001000001101011000;
assign LUT_4[42941] = 32'b00000000000000000001011001010000;
assign LUT_4[42942] = 32'b00000000000000000111100111111100;
assign LUT_4[42943] = 32'b00000000000000000000110011110100;
assign LUT_4[42944] = 32'b00000000000000010111001011000110;
assign LUT_4[42945] = 32'b00000000000000010000010110111110;
assign LUT_4[42946] = 32'b00000000000000010110100101101010;
assign LUT_4[42947] = 32'b00000000000000001111110001100010;
assign LUT_4[42948] = 32'b00000000000000010100001011100010;
assign LUT_4[42949] = 32'b00000000000000001101010111011010;
assign LUT_4[42950] = 32'b00000000000000010011100110000110;
assign LUT_4[42951] = 32'b00000000000000001100110001111110;
assign LUT_4[42952] = 32'b00000000000000010000010111011011;
assign LUT_4[42953] = 32'b00000000000000001001100011010011;
assign LUT_4[42954] = 32'b00000000000000001111110001111111;
assign LUT_4[42955] = 32'b00000000000000001000111101110111;
assign LUT_4[42956] = 32'b00000000000000001101010111110111;
assign LUT_4[42957] = 32'b00000000000000000110100011101111;
assign LUT_4[42958] = 32'b00000000000000001100110010011011;
assign LUT_4[42959] = 32'b00000000000000000101111110010011;
assign LUT_4[42960] = 32'b00000000000000010100111100110100;
assign LUT_4[42961] = 32'b00000000000000001110001000101100;
assign LUT_4[42962] = 32'b00000000000000010100010111011000;
assign LUT_4[42963] = 32'b00000000000000001101100011010000;
assign LUT_4[42964] = 32'b00000000000000010001111101010000;
assign LUT_4[42965] = 32'b00000000000000001011001001001000;
assign LUT_4[42966] = 32'b00000000000000010001010111110100;
assign LUT_4[42967] = 32'b00000000000000001010100011101100;
assign LUT_4[42968] = 32'b00000000000000001110001001001001;
assign LUT_4[42969] = 32'b00000000000000000111010101000001;
assign LUT_4[42970] = 32'b00000000000000001101100011101101;
assign LUT_4[42971] = 32'b00000000000000000110101111100101;
assign LUT_4[42972] = 32'b00000000000000001011001001100101;
assign LUT_4[42973] = 32'b00000000000000000100010101011101;
assign LUT_4[42974] = 32'b00000000000000001010100100001001;
assign LUT_4[42975] = 32'b00000000000000000011110000000001;
assign LUT_4[42976] = 32'b00000000000000010101100110001101;
assign LUT_4[42977] = 32'b00000000000000001110110010000101;
assign LUT_4[42978] = 32'b00000000000000010101000000110001;
assign LUT_4[42979] = 32'b00000000000000001110001100101001;
assign LUT_4[42980] = 32'b00000000000000010010100110101001;
assign LUT_4[42981] = 32'b00000000000000001011110010100001;
assign LUT_4[42982] = 32'b00000000000000010010000001001101;
assign LUT_4[42983] = 32'b00000000000000001011001101000101;
assign LUT_4[42984] = 32'b00000000000000001110110010100010;
assign LUT_4[42985] = 32'b00000000000000000111111110011010;
assign LUT_4[42986] = 32'b00000000000000001110001101000110;
assign LUT_4[42987] = 32'b00000000000000000111011000111110;
assign LUT_4[42988] = 32'b00000000000000001011110010111110;
assign LUT_4[42989] = 32'b00000000000000000100111110110110;
assign LUT_4[42990] = 32'b00000000000000001011001101100010;
assign LUT_4[42991] = 32'b00000000000000000100011001011010;
assign LUT_4[42992] = 32'b00000000000000010011010111111011;
assign LUT_4[42993] = 32'b00000000000000001100100011110011;
assign LUT_4[42994] = 32'b00000000000000010010110010011111;
assign LUT_4[42995] = 32'b00000000000000001011111110010111;
assign LUT_4[42996] = 32'b00000000000000010000011000010111;
assign LUT_4[42997] = 32'b00000000000000001001100100001111;
assign LUT_4[42998] = 32'b00000000000000001111110010111011;
assign LUT_4[42999] = 32'b00000000000000001000111110110011;
assign LUT_4[43000] = 32'b00000000000000001100100100010000;
assign LUT_4[43001] = 32'b00000000000000000101110000001000;
assign LUT_4[43002] = 32'b00000000000000001011111110110100;
assign LUT_4[43003] = 32'b00000000000000000101001010101100;
assign LUT_4[43004] = 32'b00000000000000001001100100101100;
assign LUT_4[43005] = 32'b00000000000000000010110000100100;
assign LUT_4[43006] = 32'b00000000000000001000111111010000;
assign LUT_4[43007] = 32'b00000000000000000010001011001000;
assign LUT_4[43008] = 32'b00000000000000001001000010101010;
assign LUT_4[43009] = 32'b00000000000000000010001110100010;
assign LUT_4[43010] = 32'b00000000000000001000011101001110;
assign LUT_4[43011] = 32'b00000000000000000001101001000110;
assign LUT_4[43012] = 32'b00000000000000000110000011000110;
assign LUT_4[43013] = 32'b11111111111111111111001110111110;
assign LUT_4[43014] = 32'b00000000000000000101011101101010;
assign LUT_4[43015] = 32'b11111111111111111110101001100010;
assign LUT_4[43016] = 32'b00000000000000000010001110111111;
assign LUT_4[43017] = 32'b11111111111111111011011010110111;
assign LUT_4[43018] = 32'b00000000000000000001101001100011;
assign LUT_4[43019] = 32'b11111111111111111010110101011011;
assign LUT_4[43020] = 32'b11111111111111111111001111011011;
assign LUT_4[43021] = 32'b11111111111111111000011011010011;
assign LUT_4[43022] = 32'b11111111111111111110101001111111;
assign LUT_4[43023] = 32'b11111111111111110111110101110111;
assign LUT_4[43024] = 32'b00000000000000000110110100011000;
assign LUT_4[43025] = 32'b00000000000000000000000000010000;
assign LUT_4[43026] = 32'b00000000000000000110001110111100;
assign LUT_4[43027] = 32'b11111111111111111111011010110100;
assign LUT_4[43028] = 32'b00000000000000000011110100110100;
assign LUT_4[43029] = 32'b11111111111111111101000000101100;
assign LUT_4[43030] = 32'b00000000000000000011001111011000;
assign LUT_4[43031] = 32'b11111111111111111100011011010000;
assign LUT_4[43032] = 32'b00000000000000000000000000101101;
assign LUT_4[43033] = 32'b11111111111111111001001100100101;
assign LUT_4[43034] = 32'b11111111111111111111011011010001;
assign LUT_4[43035] = 32'b11111111111111111000100111001001;
assign LUT_4[43036] = 32'b11111111111111111101000001001001;
assign LUT_4[43037] = 32'b11111111111111110110001101000001;
assign LUT_4[43038] = 32'b11111111111111111100011011101101;
assign LUT_4[43039] = 32'b11111111111111110101100111100101;
assign LUT_4[43040] = 32'b00000000000000000111011101110001;
assign LUT_4[43041] = 32'b00000000000000000000101001101001;
assign LUT_4[43042] = 32'b00000000000000000110111000010101;
assign LUT_4[43043] = 32'b00000000000000000000000100001101;
assign LUT_4[43044] = 32'b00000000000000000100011110001101;
assign LUT_4[43045] = 32'b11111111111111111101101010000101;
assign LUT_4[43046] = 32'b00000000000000000011111000110001;
assign LUT_4[43047] = 32'b11111111111111111101000100101001;
assign LUT_4[43048] = 32'b00000000000000000000101010000110;
assign LUT_4[43049] = 32'b11111111111111111001110101111110;
assign LUT_4[43050] = 32'b00000000000000000000000100101010;
assign LUT_4[43051] = 32'b11111111111111111001010000100010;
assign LUT_4[43052] = 32'b11111111111111111101101010100010;
assign LUT_4[43053] = 32'b11111111111111110110110110011010;
assign LUT_4[43054] = 32'b11111111111111111101000101000110;
assign LUT_4[43055] = 32'b11111111111111110110010000111110;
assign LUT_4[43056] = 32'b00000000000000000101001111011111;
assign LUT_4[43057] = 32'b11111111111111111110011011010111;
assign LUT_4[43058] = 32'b00000000000000000100101010000011;
assign LUT_4[43059] = 32'b11111111111111111101110101111011;
assign LUT_4[43060] = 32'b00000000000000000010001111111011;
assign LUT_4[43061] = 32'b11111111111111111011011011110011;
assign LUT_4[43062] = 32'b00000000000000000001101010011111;
assign LUT_4[43063] = 32'b11111111111111111010110110010111;
assign LUT_4[43064] = 32'b11111111111111111110011011110100;
assign LUT_4[43065] = 32'b11111111111111110111100111101100;
assign LUT_4[43066] = 32'b11111111111111111101110110011000;
assign LUT_4[43067] = 32'b11111111111111110111000010010000;
assign LUT_4[43068] = 32'b11111111111111111011011100010000;
assign LUT_4[43069] = 32'b11111111111111110100101000001000;
assign LUT_4[43070] = 32'b11111111111111111010110110110100;
assign LUT_4[43071] = 32'b11111111111111110100000010101100;
assign LUT_4[43072] = 32'b00000000000000001010011001111110;
assign LUT_4[43073] = 32'b00000000000000000011100101110110;
assign LUT_4[43074] = 32'b00000000000000001001110100100010;
assign LUT_4[43075] = 32'b00000000000000000011000000011010;
assign LUT_4[43076] = 32'b00000000000000000111011010011010;
assign LUT_4[43077] = 32'b00000000000000000000100110010010;
assign LUT_4[43078] = 32'b00000000000000000110110100111110;
assign LUT_4[43079] = 32'b00000000000000000000000000110110;
assign LUT_4[43080] = 32'b00000000000000000011100110010011;
assign LUT_4[43081] = 32'b11111111111111111100110010001011;
assign LUT_4[43082] = 32'b00000000000000000011000000110111;
assign LUT_4[43083] = 32'b11111111111111111100001100101111;
assign LUT_4[43084] = 32'b00000000000000000000100110101111;
assign LUT_4[43085] = 32'b11111111111111111001110010100111;
assign LUT_4[43086] = 32'b00000000000000000000000001010011;
assign LUT_4[43087] = 32'b11111111111111111001001101001011;
assign LUT_4[43088] = 32'b00000000000000001000001011101100;
assign LUT_4[43089] = 32'b00000000000000000001010111100100;
assign LUT_4[43090] = 32'b00000000000000000111100110010000;
assign LUT_4[43091] = 32'b00000000000000000000110010001000;
assign LUT_4[43092] = 32'b00000000000000000101001100001000;
assign LUT_4[43093] = 32'b11111111111111111110011000000000;
assign LUT_4[43094] = 32'b00000000000000000100100110101100;
assign LUT_4[43095] = 32'b11111111111111111101110010100100;
assign LUT_4[43096] = 32'b00000000000000000001011000000001;
assign LUT_4[43097] = 32'b11111111111111111010100011111001;
assign LUT_4[43098] = 32'b00000000000000000000110010100101;
assign LUT_4[43099] = 32'b11111111111111111001111110011101;
assign LUT_4[43100] = 32'b11111111111111111110011000011101;
assign LUT_4[43101] = 32'b11111111111111110111100100010101;
assign LUT_4[43102] = 32'b11111111111111111101110011000001;
assign LUT_4[43103] = 32'b11111111111111110110111110111001;
assign LUT_4[43104] = 32'b00000000000000001000110101000101;
assign LUT_4[43105] = 32'b00000000000000000010000000111101;
assign LUT_4[43106] = 32'b00000000000000001000001111101001;
assign LUT_4[43107] = 32'b00000000000000000001011011100001;
assign LUT_4[43108] = 32'b00000000000000000101110101100001;
assign LUT_4[43109] = 32'b11111111111111111111000001011001;
assign LUT_4[43110] = 32'b00000000000000000101010000000101;
assign LUT_4[43111] = 32'b11111111111111111110011011111101;
assign LUT_4[43112] = 32'b00000000000000000010000001011010;
assign LUT_4[43113] = 32'b11111111111111111011001101010010;
assign LUT_4[43114] = 32'b00000000000000000001011011111110;
assign LUT_4[43115] = 32'b11111111111111111010100111110110;
assign LUT_4[43116] = 32'b11111111111111111111000001110110;
assign LUT_4[43117] = 32'b11111111111111111000001101101110;
assign LUT_4[43118] = 32'b11111111111111111110011100011010;
assign LUT_4[43119] = 32'b11111111111111110111101000010010;
assign LUT_4[43120] = 32'b00000000000000000110100110110011;
assign LUT_4[43121] = 32'b11111111111111111111110010101011;
assign LUT_4[43122] = 32'b00000000000000000110000001010111;
assign LUT_4[43123] = 32'b11111111111111111111001101001111;
assign LUT_4[43124] = 32'b00000000000000000011100111001111;
assign LUT_4[43125] = 32'b11111111111111111100110011000111;
assign LUT_4[43126] = 32'b00000000000000000011000001110011;
assign LUT_4[43127] = 32'b11111111111111111100001101101011;
assign LUT_4[43128] = 32'b11111111111111111111110011001000;
assign LUT_4[43129] = 32'b11111111111111111000111111000000;
assign LUT_4[43130] = 32'b11111111111111111111001101101100;
assign LUT_4[43131] = 32'b11111111111111111000011001100100;
assign LUT_4[43132] = 32'b11111111111111111100110011100100;
assign LUT_4[43133] = 32'b11111111111111110101111111011100;
assign LUT_4[43134] = 32'b11111111111111111100001110001000;
assign LUT_4[43135] = 32'b11111111111111110101011010000000;
assign LUT_4[43136] = 32'b00000000000000001011101000110010;
assign LUT_4[43137] = 32'b00000000000000000100110100101010;
assign LUT_4[43138] = 32'b00000000000000001011000011010110;
assign LUT_4[43139] = 32'b00000000000000000100001111001110;
assign LUT_4[43140] = 32'b00000000000000001000101001001110;
assign LUT_4[43141] = 32'b00000000000000000001110101000110;
assign LUT_4[43142] = 32'b00000000000000001000000011110010;
assign LUT_4[43143] = 32'b00000000000000000001001111101010;
assign LUT_4[43144] = 32'b00000000000000000100110101000111;
assign LUT_4[43145] = 32'b11111111111111111110000000111111;
assign LUT_4[43146] = 32'b00000000000000000100001111101011;
assign LUT_4[43147] = 32'b11111111111111111101011011100011;
assign LUT_4[43148] = 32'b00000000000000000001110101100011;
assign LUT_4[43149] = 32'b11111111111111111011000001011011;
assign LUT_4[43150] = 32'b00000000000000000001010000000111;
assign LUT_4[43151] = 32'b11111111111111111010011011111111;
assign LUT_4[43152] = 32'b00000000000000001001011010100000;
assign LUT_4[43153] = 32'b00000000000000000010100110011000;
assign LUT_4[43154] = 32'b00000000000000001000110101000100;
assign LUT_4[43155] = 32'b00000000000000000010000000111100;
assign LUT_4[43156] = 32'b00000000000000000110011010111100;
assign LUT_4[43157] = 32'b11111111111111111111100110110100;
assign LUT_4[43158] = 32'b00000000000000000101110101100000;
assign LUT_4[43159] = 32'b11111111111111111111000001011000;
assign LUT_4[43160] = 32'b00000000000000000010100110110101;
assign LUT_4[43161] = 32'b11111111111111111011110010101101;
assign LUT_4[43162] = 32'b00000000000000000010000001011001;
assign LUT_4[43163] = 32'b11111111111111111011001101010001;
assign LUT_4[43164] = 32'b11111111111111111111100111010001;
assign LUT_4[43165] = 32'b11111111111111111000110011001001;
assign LUT_4[43166] = 32'b11111111111111111111000001110101;
assign LUT_4[43167] = 32'b11111111111111111000001101101101;
assign LUT_4[43168] = 32'b00000000000000001010000011111001;
assign LUT_4[43169] = 32'b00000000000000000011001111110001;
assign LUT_4[43170] = 32'b00000000000000001001011110011101;
assign LUT_4[43171] = 32'b00000000000000000010101010010101;
assign LUT_4[43172] = 32'b00000000000000000111000100010101;
assign LUT_4[43173] = 32'b00000000000000000000010000001101;
assign LUT_4[43174] = 32'b00000000000000000110011110111001;
assign LUT_4[43175] = 32'b11111111111111111111101010110001;
assign LUT_4[43176] = 32'b00000000000000000011010000001110;
assign LUT_4[43177] = 32'b11111111111111111100011100000110;
assign LUT_4[43178] = 32'b00000000000000000010101010110010;
assign LUT_4[43179] = 32'b11111111111111111011110110101010;
assign LUT_4[43180] = 32'b00000000000000000000010000101010;
assign LUT_4[43181] = 32'b11111111111111111001011100100010;
assign LUT_4[43182] = 32'b11111111111111111111101011001110;
assign LUT_4[43183] = 32'b11111111111111111000110111000110;
assign LUT_4[43184] = 32'b00000000000000000111110101100111;
assign LUT_4[43185] = 32'b00000000000000000001000001011111;
assign LUT_4[43186] = 32'b00000000000000000111010000001011;
assign LUT_4[43187] = 32'b00000000000000000000011100000011;
assign LUT_4[43188] = 32'b00000000000000000100110110000011;
assign LUT_4[43189] = 32'b11111111111111111110000001111011;
assign LUT_4[43190] = 32'b00000000000000000100010000100111;
assign LUT_4[43191] = 32'b11111111111111111101011100011111;
assign LUT_4[43192] = 32'b00000000000000000001000001111100;
assign LUT_4[43193] = 32'b11111111111111111010001101110100;
assign LUT_4[43194] = 32'b00000000000000000000011100100000;
assign LUT_4[43195] = 32'b11111111111111111001101000011000;
assign LUT_4[43196] = 32'b11111111111111111110000010011000;
assign LUT_4[43197] = 32'b11111111111111110111001110010000;
assign LUT_4[43198] = 32'b11111111111111111101011100111100;
assign LUT_4[43199] = 32'b11111111111111110110101000110100;
assign LUT_4[43200] = 32'b00000000000000001101000000000110;
assign LUT_4[43201] = 32'b00000000000000000110001011111110;
assign LUT_4[43202] = 32'b00000000000000001100011010101010;
assign LUT_4[43203] = 32'b00000000000000000101100110100010;
assign LUT_4[43204] = 32'b00000000000000001010000000100010;
assign LUT_4[43205] = 32'b00000000000000000011001100011010;
assign LUT_4[43206] = 32'b00000000000000001001011011000110;
assign LUT_4[43207] = 32'b00000000000000000010100110111110;
assign LUT_4[43208] = 32'b00000000000000000110001100011011;
assign LUT_4[43209] = 32'b11111111111111111111011000010011;
assign LUT_4[43210] = 32'b00000000000000000101100110111111;
assign LUT_4[43211] = 32'b11111111111111111110110010110111;
assign LUT_4[43212] = 32'b00000000000000000011001100110111;
assign LUT_4[43213] = 32'b11111111111111111100011000101111;
assign LUT_4[43214] = 32'b00000000000000000010100111011011;
assign LUT_4[43215] = 32'b11111111111111111011110011010011;
assign LUT_4[43216] = 32'b00000000000000001010110001110100;
assign LUT_4[43217] = 32'b00000000000000000011111101101100;
assign LUT_4[43218] = 32'b00000000000000001010001100011000;
assign LUT_4[43219] = 32'b00000000000000000011011000010000;
assign LUT_4[43220] = 32'b00000000000000000111110010010000;
assign LUT_4[43221] = 32'b00000000000000000000111110001000;
assign LUT_4[43222] = 32'b00000000000000000111001100110100;
assign LUT_4[43223] = 32'b00000000000000000000011000101100;
assign LUT_4[43224] = 32'b00000000000000000011111110001001;
assign LUT_4[43225] = 32'b11111111111111111101001010000001;
assign LUT_4[43226] = 32'b00000000000000000011011000101101;
assign LUT_4[43227] = 32'b11111111111111111100100100100101;
assign LUT_4[43228] = 32'b00000000000000000000111110100101;
assign LUT_4[43229] = 32'b11111111111111111010001010011101;
assign LUT_4[43230] = 32'b00000000000000000000011001001001;
assign LUT_4[43231] = 32'b11111111111111111001100101000001;
assign LUT_4[43232] = 32'b00000000000000001011011011001101;
assign LUT_4[43233] = 32'b00000000000000000100100111000101;
assign LUT_4[43234] = 32'b00000000000000001010110101110001;
assign LUT_4[43235] = 32'b00000000000000000100000001101001;
assign LUT_4[43236] = 32'b00000000000000001000011011101001;
assign LUT_4[43237] = 32'b00000000000000000001100111100001;
assign LUT_4[43238] = 32'b00000000000000000111110110001101;
assign LUT_4[43239] = 32'b00000000000000000001000010000101;
assign LUT_4[43240] = 32'b00000000000000000100100111100010;
assign LUT_4[43241] = 32'b11111111111111111101110011011010;
assign LUT_4[43242] = 32'b00000000000000000100000010000110;
assign LUT_4[43243] = 32'b11111111111111111101001101111110;
assign LUT_4[43244] = 32'b00000000000000000001100111111110;
assign LUT_4[43245] = 32'b11111111111111111010110011110110;
assign LUT_4[43246] = 32'b00000000000000000001000010100010;
assign LUT_4[43247] = 32'b11111111111111111010001110011010;
assign LUT_4[43248] = 32'b00000000000000001001001100111011;
assign LUT_4[43249] = 32'b00000000000000000010011000110011;
assign LUT_4[43250] = 32'b00000000000000001000100111011111;
assign LUT_4[43251] = 32'b00000000000000000001110011010111;
assign LUT_4[43252] = 32'b00000000000000000110001101010111;
assign LUT_4[43253] = 32'b11111111111111111111011001001111;
assign LUT_4[43254] = 32'b00000000000000000101100111111011;
assign LUT_4[43255] = 32'b11111111111111111110110011110011;
assign LUT_4[43256] = 32'b00000000000000000010011001010000;
assign LUT_4[43257] = 32'b11111111111111111011100101001000;
assign LUT_4[43258] = 32'b00000000000000000001110011110100;
assign LUT_4[43259] = 32'b11111111111111111010111111101100;
assign LUT_4[43260] = 32'b11111111111111111111011001101100;
assign LUT_4[43261] = 32'b11111111111111111000100101100100;
assign LUT_4[43262] = 32'b11111111111111111110110100010000;
assign LUT_4[43263] = 32'b11111111111111111000000000001000;
assign LUT_4[43264] = 32'b00000000000000001101111110001101;
assign LUT_4[43265] = 32'b00000000000000000111001010000101;
assign LUT_4[43266] = 32'b00000000000000001101011000110001;
assign LUT_4[43267] = 32'b00000000000000000110100100101001;
assign LUT_4[43268] = 32'b00000000000000001010111110101001;
assign LUT_4[43269] = 32'b00000000000000000100001010100001;
assign LUT_4[43270] = 32'b00000000000000001010011001001101;
assign LUT_4[43271] = 32'b00000000000000000011100101000101;
assign LUT_4[43272] = 32'b00000000000000000111001010100010;
assign LUT_4[43273] = 32'b00000000000000000000010110011010;
assign LUT_4[43274] = 32'b00000000000000000110100101000110;
assign LUT_4[43275] = 32'b11111111111111111111110000111110;
assign LUT_4[43276] = 32'b00000000000000000100001010111110;
assign LUT_4[43277] = 32'b11111111111111111101010110110110;
assign LUT_4[43278] = 32'b00000000000000000011100101100010;
assign LUT_4[43279] = 32'b11111111111111111100110001011010;
assign LUT_4[43280] = 32'b00000000000000001011101111111011;
assign LUT_4[43281] = 32'b00000000000000000100111011110011;
assign LUT_4[43282] = 32'b00000000000000001011001010011111;
assign LUT_4[43283] = 32'b00000000000000000100010110010111;
assign LUT_4[43284] = 32'b00000000000000001000110000010111;
assign LUT_4[43285] = 32'b00000000000000000001111100001111;
assign LUT_4[43286] = 32'b00000000000000001000001010111011;
assign LUT_4[43287] = 32'b00000000000000000001010110110011;
assign LUT_4[43288] = 32'b00000000000000000100111100010000;
assign LUT_4[43289] = 32'b11111111111111111110001000001000;
assign LUT_4[43290] = 32'b00000000000000000100010110110100;
assign LUT_4[43291] = 32'b11111111111111111101100010101100;
assign LUT_4[43292] = 32'b00000000000000000001111100101100;
assign LUT_4[43293] = 32'b11111111111111111011001000100100;
assign LUT_4[43294] = 32'b00000000000000000001010111010000;
assign LUT_4[43295] = 32'b11111111111111111010100011001000;
assign LUT_4[43296] = 32'b00000000000000001100011001010100;
assign LUT_4[43297] = 32'b00000000000000000101100101001100;
assign LUT_4[43298] = 32'b00000000000000001011110011111000;
assign LUT_4[43299] = 32'b00000000000000000100111111110000;
assign LUT_4[43300] = 32'b00000000000000001001011001110000;
assign LUT_4[43301] = 32'b00000000000000000010100101101000;
assign LUT_4[43302] = 32'b00000000000000001000110100010100;
assign LUT_4[43303] = 32'b00000000000000000010000000001100;
assign LUT_4[43304] = 32'b00000000000000000101100101101001;
assign LUT_4[43305] = 32'b11111111111111111110110001100001;
assign LUT_4[43306] = 32'b00000000000000000101000000001101;
assign LUT_4[43307] = 32'b11111111111111111110001100000101;
assign LUT_4[43308] = 32'b00000000000000000010100110000101;
assign LUT_4[43309] = 32'b11111111111111111011110001111101;
assign LUT_4[43310] = 32'b00000000000000000010000000101001;
assign LUT_4[43311] = 32'b11111111111111111011001100100001;
assign LUT_4[43312] = 32'b00000000000000001010001011000010;
assign LUT_4[43313] = 32'b00000000000000000011010110111010;
assign LUT_4[43314] = 32'b00000000000000001001100101100110;
assign LUT_4[43315] = 32'b00000000000000000010110001011110;
assign LUT_4[43316] = 32'b00000000000000000111001011011110;
assign LUT_4[43317] = 32'b00000000000000000000010111010110;
assign LUT_4[43318] = 32'b00000000000000000110100110000010;
assign LUT_4[43319] = 32'b11111111111111111111110001111010;
assign LUT_4[43320] = 32'b00000000000000000011010111010111;
assign LUT_4[43321] = 32'b11111111111111111100100011001111;
assign LUT_4[43322] = 32'b00000000000000000010110001111011;
assign LUT_4[43323] = 32'b11111111111111111011111101110011;
assign LUT_4[43324] = 32'b00000000000000000000010111110011;
assign LUT_4[43325] = 32'b11111111111111111001100011101011;
assign LUT_4[43326] = 32'b11111111111111111111110010010111;
assign LUT_4[43327] = 32'b11111111111111111000111110001111;
assign LUT_4[43328] = 32'b00000000000000001111010101100001;
assign LUT_4[43329] = 32'b00000000000000001000100001011001;
assign LUT_4[43330] = 32'b00000000000000001110110000000101;
assign LUT_4[43331] = 32'b00000000000000000111111011111101;
assign LUT_4[43332] = 32'b00000000000000001100010101111101;
assign LUT_4[43333] = 32'b00000000000000000101100001110101;
assign LUT_4[43334] = 32'b00000000000000001011110000100001;
assign LUT_4[43335] = 32'b00000000000000000100111100011001;
assign LUT_4[43336] = 32'b00000000000000001000100001110110;
assign LUT_4[43337] = 32'b00000000000000000001101101101110;
assign LUT_4[43338] = 32'b00000000000000000111111100011010;
assign LUT_4[43339] = 32'b00000000000000000001001000010010;
assign LUT_4[43340] = 32'b00000000000000000101100010010010;
assign LUT_4[43341] = 32'b11111111111111111110101110001010;
assign LUT_4[43342] = 32'b00000000000000000100111100110110;
assign LUT_4[43343] = 32'b11111111111111111110001000101110;
assign LUT_4[43344] = 32'b00000000000000001101000111001111;
assign LUT_4[43345] = 32'b00000000000000000110010011000111;
assign LUT_4[43346] = 32'b00000000000000001100100001110011;
assign LUT_4[43347] = 32'b00000000000000000101101101101011;
assign LUT_4[43348] = 32'b00000000000000001010000111101011;
assign LUT_4[43349] = 32'b00000000000000000011010011100011;
assign LUT_4[43350] = 32'b00000000000000001001100010001111;
assign LUT_4[43351] = 32'b00000000000000000010101110000111;
assign LUT_4[43352] = 32'b00000000000000000110010011100100;
assign LUT_4[43353] = 32'b11111111111111111111011111011100;
assign LUT_4[43354] = 32'b00000000000000000101101110001000;
assign LUT_4[43355] = 32'b11111111111111111110111010000000;
assign LUT_4[43356] = 32'b00000000000000000011010100000000;
assign LUT_4[43357] = 32'b11111111111111111100011111111000;
assign LUT_4[43358] = 32'b00000000000000000010101110100100;
assign LUT_4[43359] = 32'b11111111111111111011111010011100;
assign LUT_4[43360] = 32'b00000000000000001101110000101000;
assign LUT_4[43361] = 32'b00000000000000000110111100100000;
assign LUT_4[43362] = 32'b00000000000000001101001011001100;
assign LUT_4[43363] = 32'b00000000000000000110010111000100;
assign LUT_4[43364] = 32'b00000000000000001010110001000100;
assign LUT_4[43365] = 32'b00000000000000000011111100111100;
assign LUT_4[43366] = 32'b00000000000000001010001011101000;
assign LUT_4[43367] = 32'b00000000000000000011010111100000;
assign LUT_4[43368] = 32'b00000000000000000110111100111101;
assign LUT_4[43369] = 32'b00000000000000000000001000110101;
assign LUT_4[43370] = 32'b00000000000000000110010111100001;
assign LUT_4[43371] = 32'b11111111111111111111100011011001;
assign LUT_4[43372] = 32'b00000000000000000011111101011001;
assign LUT_4[43373] = 32'b11111111111111111101001001010001;
assign LUT_4[43374] = 32'b00000000000000000011010111111101;
assign LUT_4[43375] = 32'b11111111111111111100100011110101;
assign LUT_4[43376] = 32'b00000000000000001011100010010110;
assign LUT_4[43377] = 32'b00000000000000000100101110001110;
assign LUT_4[43378] = 32'b00000000000000001010111100111010;
assign LUT_4[43379] = 32'b00000000000000000100001000110010;
assign LUT_4[43380] = 32'b00000000000000001000100010110010;
assign LUT_4[43381] = 32'b00000000000000000001101110101010;
assign LUT_4[43382] = 32'b00000000000000000111111101010110;
assign LUT_4[43383] = 32'b00000000000000000001001001001110;
assign LUT_4[43384] = 32'b00000000000000000100101110101011;
assign LUT_4[43385] = 32'b11111111111111111101111010100011;
assign LUT_4[43386] = 32'b00000000000000000100001001001111;
assign LUT_4[43387] = 32'b11111111111111111101010101000111;
assign LUT_4[43388] = 32'b00000000000000000001101111000111;
assign LUT_4[43389] = 32'b11111111111111111010111010111111;
assign LUT_4[43390] = 32'b00000000000000000001001001101011;
assign LUT_4[43391] = 32'b11111111111111111010010101100011;
assign LUT_4[43392] = 32'b00000000000000010000100100010101;
assign LUT_4[43393] = 32'b00000000000000001001110000001101;
assign LUT_4[43394] = 32'b00000000000000001111111110111001;
assign LUT_4[43395] = 32'b00000000000000001001001010110001;
assign LUT_4[43396] = 32'b00000000000000001101100100110001;
assign LUT_4[43397] = 32'b00000000000000000110110000101001;
assign LUT_4[43398] = 32'b00000000000000001100111111010101;
assign LUT_4[43399] = 32'b00000000000000000110001011001101;
assign LUT_4[43400] = 32'b00000000000000001001110000101010;
assign LUT_4[43401] = 32'b00000000000000000010111100100010;
assign LUT_4[43402] = 32'b00000000000000001001001011001110;
assign LUT_4[43403] = 32'b00000000000000000010010111000110;
assign LUT_4[43404] = 32'b00000000000000000110110001000110;
assign LUT_4[43405] = 32'b11111111111111111111111100111110;
assign LUT_4[43406] = 32'b00000000000000000110001011101010;
assign LUT_4[43407] = 32'b11111111111111111111010111100010;
assign LUT_4[43408] = 32'b00000000000000001110010110000011;
assign LUT_4[43409] = 32'b00000000000000000111100001111011;
assign LUT_4[43410] = 32'b00000000000000001101110000100111;
assign LUT_4[43411] = 32'b00000000000000000110111100011111;
assign LUT_4[43412] = 32'b00000000000000001011010110011111;
assign LUT_4[43413] = 32'b00000000000000000100100010010111;
assign LUT_4[43414] = 32'b00000000000000001010110001000011;
assign LUT_4[43415] = 32'b00000000000000000011111100111011;
assign LUT_4[43416] = 32'b00000000000000000111100010011000;
assign LUT_4[43417] = 32'b00000000000000000000101110010000;
assign LUT_4[43418] = 32'b00000000000000000110111100111100;
assign LUT_4[43419] = 32'b00000000000000000000001000110100;
assign LUT_4[43420] = 32'b00000000000000000100100010110100;
assign LUT_4[43421] = 32'b11111111111111111101101110101100;
assign LUT_4[43422] = 32'b00000000000000000011111101011000;
assign LUT_4[43423] = 32'b11111111111111111101001001010000;
assign LUT_4[43424] = 32'b00000000000000001110111111011100;
assign LUT_4[43425] = 32'b00000000000000001000001011010100;
assign LUT_4[43426] = 32'b00000000000000001110011010000000;
assign LUT_4[43427] = 32'b00000000000000000111100101111000;
assign LUT_4[43428] = 32'b00000000000000001011111111111000;
assign LUT_4[43429] = 32'b00000000000000000101001011110000;
assign LUT_4[43430] = 32'b00000000000000001011011010011100;
assign LUT_4[43431] = 32'b00000000000000000100100110010100;
assign LUT_4[43432] = 32'b00000000000000001000001011110001;
assign LUT_4[43433] = 32'b00000000000000000001010111101001;
assign LUT_4[43434] = 32'b00000000000000000111100110010101;
assign LUT_4[43435] = 32'b00000000000000000000110010001101;
assign LUT_4[43436] = 32'b00000000000000000101001100001101;
assign LUT_4[43437] = 32'b11111111111111111110011000000101;
assign LUT_4[43438] = 32'b00000000000000000100100110110001;
assign LUT_4[43439] = 32'b11111111111111111101110010101001;
assign LUT_4[43440] = 32'b00000000000000001100110001001010;
assign LUT_4[43441] = 32'b00000000000000000101111101000010;
assign LUT_4[43442] = 32'b00000000000000001100001011101110;
assign LUT_4[43443] = 32'b00000000000000000101010111100110;
assign LUT_4[43444] = 32'b00000000000000001001110001100110;
assign LUT_4[43445] = 32'b00000000000000000010111101011110;
assign LUT_4[43446] = 32'b00000000000000001001001100001010;
assign LUT_4[43447] = 32'b00000000000000000010011000000010;
assign LUT_4[43448] = 32'b00000000000000000101111101011111;
assign LUT_4[43449] = 32'b11111111111111111111001001010111;
assign LUT_4[43450] = 32'b00000000000000000101011000000011;
assign LUT_4[43451] = 32'b11111111111111111110100011111011;
assign LUT_4[43452] = 32'b00000000000000000010111101111011;
assign LUT_4[43453] = 32'b11111111111111111100001001110011;
assign LUT_4[43454] = 32'b00000000000000000010011000011111;
assign LUT_4[43455] = 32'b11111111111111111011100100010111;
assign LUT_4[43456] = 32'b00000000000000010001111011101001;
assign LUT_4[43457] = 32'b00000000000000001011000111100001;
assign LUT_4[43458] = 32'b00000000000000010001010110001101;
assign LUT_4[43459] = 32'b00000000000000001010100010000101;
assign LUT_4[43460] = 32'b00000000000000001110111100000101;
assign LUT_4[43461] = 32'b00000000000000001000000111111101;
assign LUT_4[43462] = 32'b00000000000000001110010110101001;
assign LUT_4[43463] = 32'b00000000000000000111100010100001;
assign LUT_4[43464] = 32'b00000000000000001011000111111110;
assign LUT_4[43465] = 32'b00000000000000000100010011110110;
assign LUT_4[43466] = 32'b00000000000000001010100010100010;
assign LUT_4[43467] = 32'b00000000000000000011101110011010;
assign LUT_4[43468] = 32'b00000000000000001000001000011010;
assign LUT_4[43469] = 32'b00000000000000000001010100010010;
assign LUT_4[43470] = 32'b00000000000000000111100010111110;
assign LUT_4[43471] = 32'b00000000000000000000101110110110;
assign LUT_4[43472] = 32'b00000000000000001111101101010111;
assign LUT_4[43473] = 32'b00000000000000001000111001001111;
assign LUT_4[43474] = 32'b00000000000000001111000111111011;
assign LUT_4[43475] = 32'b00000000000000001000010011110011;
assign LUT_4[43476] = 32'b00000000000000001100101101110011;
assign LUT_4[43477] = 32'b00000000000000000101111001101011;
assign LUT_4[43478] = 32'b00000000000000001100001000010111;
assign LUT_4[43479] = 32'b00000000000000000101010100001111;
assign LUT_4[43480] = 32'b00000000000000001000111001101100;
assign LUT_4[43481] = 32'b00000000000000000010000101100100;
assign LUT_4[43482] = 32'b00000000000000001000010100010000;
assign LUT_4[43483] = 32'b00000000000000000001100000001000;
assign LUT_4[43484] = 32'b00000000000000000101111010001000;
assign LUT_4[43485] = 32'b11111111111111111111000110000000;
assign LUT_4[43486] = 32'b00000000000000000101010100101100;
assign LUT_4[43487] = 32'b11111111111111111110100000100100;
assign LUT_4[43488] = 32'b00000000000000010000010110110000;
assign LUT_4[43489] = 32'b00000000000000001001100010101000;
assign LUT_4[43490] = 32'b00000000000000001111110001010100;
assign LUT_4[43491] = 32'b00000000000000001000111101001100;
assign LUT_4[43492] = 32'b00000000000000001101010111001100;
assign LUT_4[43493] = 32'b00000000000000000110100011000100;
assign LUT_4[43494] = 32'b00000000000000001100110001110000;
assign LUT_4[43495] = 32'b00000000000000000101111101101000;
assign LUT_4[43496] = 32'b00000000000000001001100011000101;
assign LUT_4[43497] = 32'b00000000000000000010101110111101;
assign LUT_4[43498] = 32'b00000000000000001000111101101001;
assign LUT_4[43499] = 32'b00000000000000000010001001100001;
assign LUT_4[43500] = 32'b00000000000000000110100011100001;
assign LUT_4[43501] = 32'b11111111111111111111101111011001;
assign LUT_4[43502] = 32'b00000000000000000101111110000101;
assign LUT_4[43503] = 32'b11111111111111111111001001111101;
assign LUT_4[43504] = 32'b00000000000000001110001000011110;
assign LUT_4[43505] = 32'b00000000000000000111010100010110;
assign LUT_4[43506] = 32'b00000000000000001101100011000010;
assign LUT_4[43507] = 32'b00000000000000000110101110111010;
assign LUT_4[43508] = 32'b00000000000000001011001000111010;
assign LUT_4[43509] = 32'b00000000000000000100010100110010;
assign LUT_4[43510] = 32'b00000000000000001010100011011110;
assign LUT_4[43511] = 32'b00000000000000000011101111010110;
assign LUT_4[43512] = 32'b00000000000000000111010100110011;
assign LUT_4[43513] = 32'b00000000000000000000100000101011;
assign LUT_4[43514] = 32'b00000000000000000110101111010111;
assign LUT_4[43515] = 32'b11111111111111111111111011001111;
assign LUT_4[43516] = 32'b00000000000000000100010101001111;
assign LUT_4[43517] = 32'b11111111111111111101100001000111;
assign LUT_4[43518] = 32'b00000000000000000011101111110011;
assign LUT_4[43519] = 32'b11111111111111111100111011101011;
assign LUT_4[43520] = 32'b00000000000000001000000110110010;
assign LUT_4[43521] = 32'b00000000000000000001010010101010;
assign LUT_4[43522] = 32'b00000000000000000111100001010110;
assign LUT_4[43523] = 32'b00000000000000000000101101001110;
assign LUT_4[43524] = 32'b00000000000000000101000111001110;
assign LUT_4[43525] = 32'b11111111111111111110010011000110;
assign LUT_4[43526] = 32'b00000000000000000100100001110010;
assign LUT_4[43527] = 32'b11111111111111111101101101101010;
assign LUT_4[43528] = 32'b00000000000000000001010011000111;
assign LUT_4[43529] = 32'b11111111111111111010011110111111;
assign LUT_4[43530] = 32'b00000000000000000000101101101011;
assign LUT_4[43531] = 32'b11111111111111111001111001100011;
assign LUT_4[43532] = 32'b11111111111111111110010011100011;
assign LUT_4[43533] = 32'b11111111111111110111011111011011;
assign LUT_4[43534] = 32'b11111111111111111101101110000111;
assign LUT_4[43535] = 32'b11111111111111110110111001111111;
assign LUT_4[43536] = 32'b00000000000000000101111000100000;
assign LUT_4[43537] = 32'b11111111111111111111000100011000;
assign LUT_4[43538] = 32'b00000000000000000101010011000100;
assign LUT_4[43539] = 32'b11111111111111111110011110111100;
assign LUT_4[43540] = 32'b00000000000000000010111000111100;
assign LUT_4[43541] = 32'b11111111111111111100000100110100;
assign LUT_4[43542] = 32'b00000000000000000010010011100000;
assign LUT_4[43543] = 32'b11111111111111111011011111011000;
assign LUT_4[43544] = 32'b11111111111111111111000100110101;
assign LUT_4[43545] = 32'b11111111111111111000010000101101;
assign LUT_4[43546] = 32'b11111111111111111110011111011001;
assign LUT_4[43547] = 32'b11111111111111110111101011010001;
assign LUT_4[43548] = 32'b11111111111111111100000101010001;
assign LUT_4[43549] = 32'b11111111111111110101010001001001;
assign LUT_4[43550] = 32'b11111111111111111011011111110101;
assign LUT_4[43551] = 32'b11111111111111110100101011101101;
assign LUT_4[43552] = 32'b00000000000000000110100001111001;
assign LUT_4[43553] = 32'b11111111111111111111101101110001;
assign LUT_4[43554] = 32'b00000000000000000101111100011101;
assign LUT_4[43555] = 32'b11111111111111111111001000010101;
assign LUT_4[43556] = 32'b00000000000000000011100010010101;
assign LUT_4[43557] = 32'b11111111111111111100101110001101;
assign LUT_4[43558] = 32'b00000000000000000010111100111001;
assign LUT_4[43559] = 32'b11111111111111111100001000110001;
assign LUT_4[43560] = 32'b11111111111111111111101110001110;
assign LUT_4[43561] = 32'b11111111111111111000111010000110;
assign LUT_4[43562] = 32'b11111111111111111111001000110010;
assign LUT_4[43563] = 32'b11111111111111111000010100101010;
assign LUT_4[43564] = 32'b11111111111111111100101110101010;
assign LUT_4[43565] = 32'b11111111111111110101111010100010;
assign LUT_4[43566] = 32'b11111111111111111100001001001110;
assign LUT_4[43567] = 32'b11111111111111110101010101000110;
assign LUT_4[43568] = 32'b00000000000000000100010011100111;
assign LUT_4[43569] = 32'b11111111111111111101011111011111;
assign LUT_4[43570] = 32'b00000000000000000011101110001011;
assign LUT_4[43571] = 32'b11111111111111111100111010000011;
assign LUT_4[43572] = 32'b00000000000000000001010100000011;
assign LUT_4[43573] = 32'b11111111111111111010011111111011;
assign LUT_4[43574] = 32'b00000000000000000000101110100111;
assign LUT_4[43575] = 32'b11111111111111111001111010011111;
assign LUT_4[43576] = 32'b11111111111111111101011111111100;
assign LUT_4[43577] = 32'b11111111111111110110101011110100;
assign LUT_4[43578] = 32'b11111111111111111100111010100000;
assign LUT_4[43579] = 32'b11111111111111110110000110011000;
assign LUT_4[43580] = 32'b11111111111111111010100000011000;
assign LUT_4[43581] = 32'b11111111111111110011101100010000;
assign LUT_4[43582] = 32'b11111111111111111001111010111100;
assign LUT_4[43583] = 32'b11111111111111110011000110110100;
assign LUT_4[43584] = 32'b00000000000000001001011110000110;
assign LUT_4[43585] = 32'b00000000000000000010101001111110;
assign LUT_4[43586] = 32'b00000000000000001000111000101010;
assign LUT_4[43587] = 32'b00000000000000000010000100100010;
assign LUT_4[43588] = 32'b00000000000000000110011110100010;
assign LUT_4[43589] = 32'b11111111111111111111101010011010;
assign LUT_4[43590] = 32'b00000000000000000101111001000110;
assign LUT_4[43591] = 32'b11111111111111111111000100111110;
assign LUT_4[43592] = 32'b00000000000000000010101010011011;
assign LUT_4[43593] = 32'b11111111111111111011110110010011;
assign LUT_4[43594] = 32'b00000000000000000010000100111111;
assign LUT_4[43595] = 32'b11111111111111111011010000110111;
assign LUT_4[43596] = 32'b11111111111111111111101010110111;
assign LUT_4[43597] = 32'b11111111111111111000110110101111;
assign LUT_4[43598] = 32'b11111111111111111111000101011011;
assign LUT_4[43599] = 32'b11111111111111111000010001010011;
assign LUT_4[43600] = 32'b00000000000000000111001111110100;
assign LUT_4[43601] = 32'b00000000000000000000011011101100;
assign LUT_4[43602] = 32'b00000000000000000110101010011000;
assign LUT_4[43603] = 32'b11111111111111111111110110010000;
assign LUT_4[43604] = 32'b00000000000000000100010000010000;
assign LUT_4[43605] = 32'b11111111111111111101011100001000;
assign LUT_4[43606] = 32'b00000000000000000011101010110100;
assign LUT_4[43607] = 32'b11111111111111111100110110101100;
assign LUT_4[43608] = 32'b00000000000000000000011100001001;
assign LUT_4[43609] = 32'b11111111111111111001101000000001;
assign LUT_4[43610] = 32'b11111111111111111111110110101101;
assign LUT_4[43611] = 32'b11111111111111111001000010100101;
assign LUT_4[43612] = 32'b11111111111111111101011100100101;
assign LUT_4[43613] = 32'b11111111111111110110101000011101;
assign LUT_4[43614] = 32'b11111111111111111100110111001001;
assign LUT_4[43615] = 32'b11111111111111110110000011000001;
assign LUT_4[43616] = 32'b00000000000000000111111001001101;
assign LUT_4[43617] = 32'b00000000000000000001000101000101;
assign LUT_4[43618] = 32'b00000000000000000111010011110001;
assign LUT_4[43619] = 32'b00000000000000000000011111101001;
assign LUT_4[43620] = 32'b00000000000000000100111001101001;
assign LUT_4[43621] = 32'b11111111111111111110000101100001;
assign LUT_4[43622] = 32'b00000000000000000100010100001101;
assign LUT_4[43623] = 32'b11111111111111111101100000000101;
assign LUT_4[43624] = 32'b00000000000000000001000101100010;
assign LUT_4[43625] = 32'b11111111111111111010010001011010;
assign LUT_4[43626] = 32'b00000000000000000000100000000110;
assign LUT_4[43627] = 32'b11111111111111111001101011111110;
assign LUT_4[43628] = 32'b11111111111111111110000101111110;
assign LUT_4[43629] = 32'b11111111111111110111010001110110;
assign LUT_4[43630] = 32'b11111111111111111101100000100010;
assign LUT_4[43631] = 32'b11111111111111110110101100011010;
assign LUT_4[43632] = 32'b00000000000000000101101010111011;
assign LUT_4[43633] = 32'b11111111111111111110110110110011;
assign LUT_4[43634] = 32'b00000000000000000101000101011111;
assign LUT_4[43635] = 32'b11111111111111111110010001010111;
assign LUT_4[43636] = 32'b00000000000000000010101011010111;
assign LUT_4[43637] = 32'b11111111111111111011110111001111;
assign LUT_4[43638] = 32'b00000000000000000010000101111011;
assign LUT_4[43639] = 32'b11111111111111111011010001110011;
assign LUT_4[43640] = 32'b11111111111111111110110111010000;
assign LUT_4[43641] = 32'b11111111111111111000000011001000;
assign LUT_4[43642] = 32'b11111111111111111110010001110100;
assign LUT_4[43643] = 32'b11111111111111110111011101101100;
assign LUT_4[43644] = 32'b11111111111111111011110111101100;
assign LUT_4[43645] = 32'b11111111111111110101000011100100;
assign LUT_4[43646] = 32'b11111111111111111011010010010000;
assign LUT_4[43647] = 32'b11111111111111110100011110001000;
assign LUT_4[43648] = 32'b00000000000000001010101100111010;
assign LUT_4[43649] = 32'b00000000000000000011111000110010;
assign LUT_4[43650] = 32'b00000000000000001010000111011110;
assign LUT_4[43651] = 32'b00000000000000000011010011010110;
assign LUT_4[43652] = 32'b00000000000000000111101101010110;
assign LUT_4[43653] = 32'b00000000000000000000111001001110;
assign LUT_4[43654] = 32'b00000000000000000111000111111010;
assign LUT_4[43655] = 32'b00000000000000000000010011110010;
assign LUT_4[43656] = 32'b00000000000000000011111001001111;
assign LUT_4[43657] = 32'b11111111111111111101000101000111;
assign LUT_4[43658] = 32'b00000000000000000011010011110011;
assign LUT_4[43659] = 32'b11111111111111111100011111101011;
assign LUT_4[43660] = 32'b00000000000000000000111001101011;
assign LUT_4[43661] = 32'b11111111111111111010000101100011;
assign LUT_4[43662] = 32'b00000000000000000000010100001111;
assign LUT_4[43663] = 32'b11111111111111111001100000000111;
assign LUT_4[43664] = 32'b00000000000000001000011110101000;
assign LUT_4[43665] = 32'b00000000000000000001101010100000;
assign LUT_4[43666] = 32'b00000000000000000111111001001100;
assign LUT_4[43667] = 32'b00000000000000000001000101000100;
assign LUT_4[43668] = 32'b00000000000000000101011111000100;
assign LUT_4[43669] = 32'b11111111111111111110101010111100;
assign LUT_4[43670] = 32'b00000000000000000100111001101000;
assign LUT_4[43671] = 32'b11111111111111111110000101100000;
assign LUT_4[43672] = 32'b00000000000000000001101010111101;
assign LUT_4[43673] = 32'b11111111111111111010110110110101;
assign LUT_4[43674] = 32'b00000000000000000001000101100001;
assign LUT_4[43675] = 32'b11111111111111111010010001011001;
assign LUT_4[43676] = 32'b11111111111111111110101011011001;
assign LUT_4[43677] = 32'b11111111111111110111110111010001;
assign LUT_4[43678] = 32'b11111111111111111110000101111101;
assign LUT_4[43679] = 32'b11111111111111110111010001110101;
assign LUT_4[43680] = 32'b00000000000000001001001000000001;
assign LUT_4[43681] = 32'b00000000000000000010010011111001;
assign LUT_4[43682] = 32'b00000000000000001000100010100101;
assign LUT_4[43683] = 32'b00000000000000000001101110011101;
assign LUT_4[43684] = 32'b00000000000000000110001000011101;
assign LUT_4[43685] = 32'b11111111111111111111010100010101;
assign LUT_4[43686] = 32'b00000000000000000101100011000001;
assign LUT_4[43687] = 32'b11111111111111111110101110111001;
assign LUT_4[43688] = 32'b00000000000000000010010100010110;
assign LUT_4[43689] = 32'b11111111111111111011100000001110;
assign LUT_4[43690] = 32'b00000000000000000001101110111010;
assign LUT_4[43691] = 32'b11111111111111111010111010110010;
assign LUT_4[43692] = 32'b11111111111111111111010100110010;
assign LUT_4[43693] = 32'b11111111111111111000100000101010;
assign LUT_4[43694] = 32'b11111111111111111110101111010110;
assign LUT_4[43695] = 32'b11111111111111110111111011001110;
assign LUT_4[43696] = 32'b00000000000000000110111001101111;
assign LUT_4[43697] = 32'b00000000000000000000000101100111;
assign LUT_4[43698] = 32'b00000000000000000110010100010011;
assign LUT_4[43699] = 32'b11111111111111111111100000001011;
assign LUT_4[43700] = 32'b00000000000000000011111010001011;
assign LUT_4[43701] = 32'b11111111111111111101000110000011;
assign LUT_4[43702] = 32'b00000000000000000011010100101111;
assign LUT_4[43703] = 32'b11111111111111111100100000100111;
assign LUT_4[43704] = 32'b00000000000000000000000110000100;
assign LUT_4[43705] = 32'b11111111111111111001010001111100;
assign LUT_4[43706] = 32'b11111111111111111111100000101000;
assign LUT_4[43707] = 32'b11111111111111111000101100100000;
assign LUT_4[43708] = 32'b11111111111111111101000110100000;
assign LUT_4[43709] = 32'b11111111111111110110010010011000;
assign LUT_4[43710] = 32'b11111111111111111100100001000100;
assign LUT_4[43711] = 32'b11111111111111110101101100111100;
assign LUT_4[43712] = 32'b00000000000000001100000100001110;
assign LUT_4[43713] = 32'b00000000000000000101010000000110;
assign LUT_4[43714] = 32'b00000000000000001011011110110010;
assign LUT_4[43715] = 32'b00000000000000000100101010101010;
assign LUT_4[43716] = 32'b00000000000000001001000100101010;
assign LUT_4[43717] = 32'b00000000000000000010010000100010;
assign LUT_4[43718] = 32'b00000000000000001000011111001110;
assign LUT_4[43719] = 32'b00000000000000000001101011000110;
assign LUT_4[43720] = 32'b00000000000000000101010000100011;
assign LUT_4[43721] = 32'b11111111111111111110011100011011;
assign LUT_4[43722] = 32'b00000000000000000100101011000111;
assign LUT_4[43723] = 32'b11111111111111111101110110111111;
assign LUT_4[43724] = 32'b00000000000000000010010000111111;
assign LUT_4[43725] = 32'b11111111111111111011011100110111;
assign LUT_4[43726] = 32'b00000000000000000001101011100011;
assign LUT_4[43727] = 32'b11111111111111111010110111011011;
assign LUT_4[43728] = 32'b00000000000000001001110101111100;
assign LUT_4[43729] = 32'b00000000000000000011000001110100;
assign LUT_4[43730] = 32'b00000000000000001001010000100000;
assign LUT_4[43731] = 32'b00000000000000000010011100011000;
assign LUT_4[43732] = 32'b00000000000000000110110110011000;
assign LUT_4[43733] = 32'b00000000000000000000000010010000;
assign LUT_4[43734] = 32'b00000000000000000110010000111100;
assign LUT_4[43735] = 32'b11111111111111111111011100110100;
assign LUT_4[43736] = 32'b00000000000000000011000010010001;
assign LUT_4[43737] = 32'b11111111111111111100001110001001;
assign LUT_4[43738] = 32'b00000000000000000010011100110101;
assign LUT_4[43739] = 32'b11111111111111111011101000101101;
assign LUT_4[43740] = 32'b00000000000000000000000010101101;
assign LUT_4[43741] = 32'b11111111111111111001001110100101;
assign LUT_4[43742] = 32'b11111111111111111111011101010001;
assign LUT_4[43743] = 32'b11111111111111111000101001001001;
assign LUT_4[43744] = 32'b00000000000000001010011111010101;
assign LUT_4[43745] = 32'b00000000000000000011101011001101;
assign LUT_4[43746] = 32'b00000000000000001001111001111001;
assign LUT_4[43747] = 32'b00000000000000000011000101110001;
assign LUT_4[43748] = 32'b00000000000000000111011111110001;
assign LUT_4[43749] = 32'b00000000000000000000101011101001;
assign LUT_4[43750] = 32'b00000000000000000110111010010101;
assign LUT_4[43751] = 32'b00000000000000000000000110001101;
assign LUT_4[43752] = 32'b00000000000000000011101011101010;
assign LUT_4[43753] = 32'b11111111111111111100110111100010;
assign LUT_4[43754] = 32'b00000000000000000011000110001110;
assign LUT_4[43755] = 32'b11111111111111111100010010000110;
assign LUT_4[43756] = 32'b00000000000000000000101100000110;
assign LUT_4[43757] = 32'b11111111111111111001110111111110;
assign LUT_4[43758] = 32'b00000000000000000000000110101010;
assign LUT_4[43759] = 32'b11111111111111111001010010100010;
assign LUT_4[43760] = 32'b00000000000000001000010001000011;
assign LUT_4[43761] = 32'b00000000000000000001011100111011;
assign LUT_4[43762] = 32'b00000000000000000111101011100111;
assign LUT_4[43763] = 32'b00000000000000000000110111011111;
assign LUT_4[43764] = 32'b00000000000000000101010001011111;
assign LUT_4[43765] = 32'b11111111111111111110011101010111;
assign LUT_4[43766] = 32'b00000000000000000100101100000011;
assign LUT_4[43767] = 32'b11111111111111111101110111111011;
assign LUT_4[43768] = 32'b00000000000000000001011101011000;
assign LUT_4[43769] = 32'b11111111111111111010101001010000;
assign LUT_4[43770] = 32'b00000000000000000000110111111100;
assign LUT_4[43771] = 32'b11111111111111111010000011110100;
assign LUT_4[43772] = 32'b11111111111111111110011101110100;
assign LUT_4[43773] = 32'b11111111111111110111101001101100;
assign LUT_4[43774] = 32'b11111111111111111101111000011000;
assign LUT_4[43775] = 32'b11111111111111110111000100010000;
assign LUT_4[43776] = 32'b00000000000000001101000010010101;
assign LUT_4[43777] = 32'b00000000000000000110001110001101;
assign LUT_4[43778] = 32'b00000000000000001100011100111001;
assign LUT_4[43779] = 32'b00000000000000000101101000110001;
assign LUT_4[43780] = 32'b00000000000000001010000010110001;
assign LUT_4[43781] = 32'b00000000000000000011001110101001;
assign LUT_4[43782] = 32'b00000000000000001001011101010101;
assign LUT_4[43783] = 32'b00000000000000000010101001001101;
assign LUT_4[43784] = 32'b00000000000000000110001110101010;
assign LUT_4[43785] = 32'b11111111111111111111011010100010;
assign LUT_4[43786] = 32'b00000000000000000101101001001110;
assign LUT_4[43787] = 32'b11111111111111111110110101000110;
assign LUT_4[43788] = 32'b00000000000000000011001111000110;
assign LUT_4[43789] = 32'b11111111111111111100011010111110;
assign LUT_4[43790] = 32'b00000000000000000010101001101010;
assign LUT_4[43791] = 32'b11111111111111111011110101100010;
assign LUT_4[43792] = 32'b00000000000000001010110100000011;
assign LUT_4[43793] = 32'b00000000000000000011111111111011;
assign LUT_4[43794] = 32'b00000000000000001010001110100111;
assign LUT_4[43795] = 32'b00000000000000000011011010011111;
assign LUT_4[43796] = 32'b00000000000000000111110100011111;
assign LUT_4[43797] = 32'b00000000000000000001000000010111;
assign LUT_4[43798] = 32'b00000000000000000111001111000011;
assign LUT_4[43799] = 32'b00000000000000000000011010111011;
assign LUT_4[43800] = 32'b00000000000000000100000000011000;
assign LUT_4[43801] = 32'b11111111111111111101001100010000;
assign LUT_4[43802] = 32'b00000000000000000011011010111100;
assign LUT_4[43803] = 32'b11111111111111111100100110110100;
assign LUT_4[43804] = 32'b00000000000000000001000000110100;
assign LUT_4[43805] = 32'b11111111111111111010001100101100;
assign LUT_4[43806] = 32'b00000000000000000000011011011000;
assign LUT_4[43807] = 32'b11111111111111111001100111010000;
assign LUT_4[43808] = 32'b00000000000000001011011101011100;
assign LUT_4[43809] = 32'b00000000000000000100101001010100;
assign LUT_4[43810] = 32'b00000000000000001010111000000000;
assign LUT_4[43811] = 32'b00000000000000000100000011111000;
assign LUT_4[43812] = 32'b00000000000000001000011101111000;
assign LUT_4[43813] = 32'b00000000000000000001101001110000;
assign LUT_4[43814] = 32'b00000000000000000111111000011100;
assign LUT_4[43815] = 32'b00000000000000000001000100010100;
assign LUT_4[43816] = 32'b00000000000000000100101001110001;
assign LUT_4[43817] = 32'b11111111111111111101110101101001;
assign LUT_4[43818] = 32'b00000000000000000100000100010101;
assign LUT_4[43819] = 32'b11111111111111111101010000001101;
assign LUT_4[43820] = 32'b00000000000000000001101010001101;
assign LUT_4[43821] = 32'b11111111111111111010110110000101;
assign LUT_4[43822] = 32'b00000000000000000001000100110001;
assign LUT_4[43823] = 32'b11111111111111111010010000101001;
assign LUT_4[43824] = 32'b00000000000000001001001111001010;
assign LUT_4[43825] = 32'b00000000000000000010011011000010;
assign LUT_4[43826] = 32'b00000000000000001000101001101110;
assign LUT_4[43827] = 32'b00000000000000000001110101100110;
assign LUT_4[43828] = 32'b00000000000000000110001111100110;
assign LUT_4[43829] = 32'b11111111111111111111011011011110;
assign LUT_4[43830] = 32'b00000000000000000101101010001010;
assign LUT_4[43831] = 32'b11111111111111111110110110000010;
assign LUT_4[43832] = 32'b00000000000000000010011011011111;
assign LUT_4[43833] = 32'b11111111111111111011100111010111;
assign LUT_4[43834] = 32'b00000000000000000001110110000011;
assign LUT_4[43835] = 32'b11111111111111111011000001111011;
assign LUT_4[43836] = 32'b11111111111111111111011011111011;
assign LUT_4[43837] = 32'b11111111111111111000100111110011;
assign LUT_4[43838] = 32'b11111111111111111110110110011111;
assign LUT_4[43839] = 32'b11111111111111111000000010010111;
assign LUT_4[43840] = 32'b00000000000000001110011001101001;
assign LUT_4[43841] = 32'b00000000000000000111100101100001;
assign LUT_4[43842] = 32'b00000000000000001101110100001101;
assign LUT_4[43843] = 32'b00000000000000000111000000000101;
assign LUT_4[43844] = 32'b00000000000000001011011010000101;
assign LUT_4[43845] = 32'b00000000000000000100100101111101;
assign LUT_4[43846] = 32'b00000000000000001010110100101001;
assign LUT_4[43847] = 32'b00000000000000000100000000100001;
assign LUT_4[43848] = 32'b00000000000000000111100101111110;
assign LUT_4[43849] = 32'b00000000000000000000110001110110;
assign LUT_4[43850] = 32'b00000000000000000111000000100010;
assign LUT_4[43851] = 32'b00000000000000000000001100011010;
assign LUT_4[43852] = 32'b00000000000000000100100110011010;
assign LUT_4[43853] = 32'b11111111111111111101110010010010;
assign LUT_4[43854] = 32'b00000000000000000100000000111110;
assign LUT_4[43855] = 32'b11111111111111111101001100110110;
assign LUT_4[43856] = 32'b00000000000000001100001011010111;
assign LUT_4[43857] = 32'b00000000000000000101010111001111;
assign LUT_4[43858] = 32'b00000000000000001011100101111011;
assign LUT_4[43859] = 32'b00000000000000000100110001110011;
assign LUT_4[43860] = 32'b00000000000000001001001011110011;
assign LUT_4[43861] = 32'b00000000000000000010010111101011;
assign LUT_4[43862] = 32'b00000000000000001000100110010111;
assign LUT_4[43863] = 32'b00000000000000000001110010001111;
assign LUT_4[43864] = 32'b00000000000000000101010111101100;
assign LUT_4[43865] = 32'b11111111111111111110100011100100;
assign LUT_4[43866] = 32'b00000000000000000100110010010000;
assign LUT_4[43867] = 32'b11111111111111111101111110001000;
assign LUT_4[43868] = 32'b00000000000000000010011000001000;
assign LUT_4[43869] = 32'b11111111111111111011100100000000;
assign LUT_4[43870] = 32'b00000000000000000001110010101100;
assign LUT_4[43871] = 32'b11111111111111111010111110100100;
assign LUT_4[43872] = 32'b00000000000000001100110100110000;
assign LUT_4[43873] = 32'b00000000000000000110000000101000;
assign LUT_4[43874] = 32'b00000000000000001100001111010100;
assign LUT_4[43875] = 32'b00000000000000000101011011001100;
assign LUT_4[43876] = 32'b00000000000000001001110101001100;
assign LUT_4[43877] = 32'b00000000000000000011000001000100;
assign LUT_4[43878] = 32'b00000000000000001001001111110000;
assign LUT_4[43879] = 32'b00000000000000000010011011101000;
assign LUT_4[43880] = 32'b00000000000000000110000001000101;
assign LUT_4[43881] = 32'b11111111111111111111001100111101;
assign LUT_4[43882] = 32'b00000000000000000101011011101001;
assign LUT_4[43883] = 32'b11111111111111111110100111100001;
assign LUT_4[43884] = 32'b00000000000000000011000001100001;
assign LUT_4[43885] = 32'b11111111111111111100001101011001;
assign LUT_4[43886] = 32'b00000000000000000010011100000101;
assign LUT_4[43887] = 32'b11111111111111111011100111111101;
assign LUT_4[43888] = 32'b00000000000000001010100110011110;
assign LUT_4[43889] = 32'b00000000000000000011110010010110;
assign LUT_4[43890] = 32'b00000000000000001010000001000010;
assign LUT_4[43891] = 32'b00000000000000000011001100111010;
assign LUT_4[43892] = 32'b00000000000000000111100110111010;
assign LUT_4[43893] = 32'b00000000000000000000110010110010;
assign LUT_4[43894] = 32'b00000000000000000111000001011110;
assign LUT_4[43895] = 32'b00000000000000000000001101010110;
assign LUT_4[43896] = 32'b00000000000000000011110010110011;
assign LUT_4[43897] = 32'b11111111111111111100111110101011;
assign LUT_4[43898] = 32'b00000000000000000011001101010111;
assign LUT_4[43899] = 32'b11111111111111111100011001001111;
assign LUT_4[43900] = 32'b00000000000000000000110011001111;
assign LUT_4[43901] = 32'b11111111111111111001111111000111;
assign LUT_4[43902] = 32'b00000000000000000000001101110011;
assign LUT_4[43903] = 32'b11111111111111111001011001101011;
assign LUT_4[43904] = 32'b00000000000000001111101000011101;
assign LUT_4[43905] = 32'b00000000000000001000110100010101;
assign LUT_4[43906] = 32'b00000000000000001111000011000001;
assign LUT_4[43907] = 32'b00000000000000001000001110111001;
assign LUT_4[43908] = 32'b00000000000000001100101000111001;
assign LUT_4[43909] = 32'b00000000000000000101110100110001;
assign LUT_4[43910] = 32'b00000000000000001100000011011101;
assign LUT_4[43911] = 32'b00000000000000000101001111010101;
assign LUT_4[43912] = 32'b00000000000000001000110100110010;
assign LUT_4[43913] = 32'b00000000000000000010000000101010;
assign LUT_4[43914] = 32'b00000000000000001000001111010110;
assign LUT_4[43915] = 32'b00000000000000000001011011001110;
assign LUT_4[43916] = 32'b00000000000000000101110101001110;
assign LUT_4[43917] = 32'b11111111111111111111000001000110;
assign LUT_4[43918] = 32'b00000000000000000101001111110010;
assign LUT_4[43919] = 32'b11111111111111111110011011101010;
assign LUT_4[43920] = 32'b00000000000000001101011010001011;
assign LUT_4[43921] = 32'b00000000000000000110100110000011;
assign LUT_4[43922] = 32'b00000000000000001100110100101111;
assign LUT_4[43923] = 32'b00000000000000000110000000100111;
assign LUT_4[43924] = 32'b00000000000000001010011010100111;
assign LUT_4[43925] = 32'b00000000000000000011100110011111;
assign LUT_4[43926] = 32'b00000000000000001001110101001011;
assign LUT_4[43927] = 32'b00000000000000000011000001000011;
assign LUT_4[43928] = 32'b00000000000000000110100110100000;
assign LUT_4[43929] = 32'b11111111111111111111110010011000;
assign LUT_4[43930] = 32'b00000000000000000110000001000100;
assign LUT_4[43931] = 32'b11111111111111111111001100111100;
assign LUT_4[43932] = 32'b00000000000000000011100110111100;
assign LUT_4[43933] = 32'b11111111111111111100110010110100;
assign LUT_4[43934] = 32'b00000000000000000011000001100000;
assign LUT_4[43935] = 32'b11111111111111111100001101011000;
assign LUT_4[43936] = 32'b00000000000000001110000011100100;
assign LUT_4[43937] = 32'b00000000000000000111001111011100;
assign LUT_4[43938] = 32'b00000000000000001101011110001000;
assign LUT_4[43939] = 32'b00000000000000000110101010000000;
assign LUT_4[43940] = 32'b00000000000000001011000100000000;
assign LUT_4[43941] = 32'b00000000000000000100001111111000;
assign LUT_4[43942] = 32'b00000000000000001010011110100100;
assign LUT_4[43943] = 32'b00000000000000000011101010011100;
assign LUT_4[43944] = 32'b00000000000000000111001111111001;
assign LUT_4[43945] = 32'b00000000000000000000011011110001;
assign LUT_4[43946] = 32'b00000000000000000110101010011101;
assign LUT_4[43947] = 32'b11111111111111111111110110010101;
assign LUT_4[43948] = 32'b00000000000000000100010000010101;
assign LUT_4[43949] = 32'b11111111111111111101011100001101;
assign LUT_4[43950] = 32'b00000000000000000011101010111001;
assign LUT_4[43951] = 32'b11111111111111111100110110110001;
assign LUT_4[43952] = 32'b00000000000000001011110101010010;
assign LUT_4[43953] = 32'b00000000000000000101000001001010;
assign LUT_4[43954] = 32'b00000000000000001011001111110110;
assign LUT_4[43955] = 32'b00000000000000000100011011101110;
assign LUT_4[43956] = 32'b00000000000000001000110101101110;
assign LUT_4[43957] = 32'b00000000000000000010000001100110;
assign LUT_4[43958] = 32'b00000000000000001000010000010010;
assign LUT_4[43959] = 32'b00000000000000000001011100001010;
assign LUT_4[43960] = 32'b00000000000000000101000001100111;
assign LUT_4[43961] = 32'b11111111111111111110001101011111;
assign LUT_4[43962] = 32'b00000000000000000100011100001011;
assign LUT_4[43963] = 32'b11111111111111111101101000000011;
assign LUT_4[43964] = 32'b00000000000000000010000010000011;
assign LUT_4[43965] = 32'b11111111111111111011001101111011;
assign LUT_4[43966] = 32'b00000000000000000001011100100111;
assign LUT_4[43967] = 32'b11111111111111111010101000011111;
assign LUT_4[43968] = 32'b00000000000000010000111111110001;
assign LUT_4[43969] = 32'b00000000000000001010001011101001;
assign LUT_4[43970] = 32'b00000000000000010000011010010101;
assign LUT_4[43971] = 32'b00000000000000001001100110001101;
assign LUT_4[43972] = 32'b00000000000000001110000000001101;
assign LUT_4[43973] = 32'b00000000000000000111001100000101;
assign LUT_4[43974] = 32'b00000000000000001101011010110001;
assign LUT_4[43975] = 32'b00000000000000000110100110101001;
assign LUT_4[43976] = 32'b00000000000000001010001100000110;
assign LUT_4[43977] = 32'b00000000000000000011010111111110;
assign LUT_4[43978] = 32'b00000000000000001001100110101010;
assign LUT_4[43979] = 32'b00000000000000000010110010100010;
assign LUT_4[43980] = 32'b00000000000000000111001100100010;
assign LUT_4[43981] = 32'b00000000000000000000011000011010;
assign LUT_4[43982] = 32'b00000000000000000110100111000110;
assign LUT_4[43983] = 32'b11111111111111111111110010111110;
assign LUT_4[43984] = 32'b00000000000000001110110001011111;
assign LUT_4[43985] = 32'b00000000000000000111111101010111;
assign LUT_4[43986] = 32'b00000000000000001110001100000011;
assign LUT_4[43987] = 32'b00000000000000000111010111111011;
assign LUT_4[43988] = 32'b00000000000000001011110001111011;
assign LUT_4[43989] = 32'b00000000000000000100111101110011;
assign LUT_4[43990] = 32'b00000000000000001011001100011111;
assign LUT_4[43991] = 32'b00000000000000000100011000010111;
assign LUT_4[43992] = 32'b00000000000000000111111101110100;
assign LUT_4[43993] = 32'b00000000000000000001001001101100;
assign LUT_4[43994] = 32'b00000000000000000111011000011000;
assign LUT_4[43995] = 32'b00000000000000000000100100010000;
assign LUT_4[43996] = 32'b00000000000000000100111110010000;
assign LUT_4[43997] = 32'b11111111111111111110001010001000;
assign LUT_4[43998] = 32'b00000000000000000100011000110100;
assign LUT_4[43999] = 32'b11111111111111111101100100101100;
assign LUT_4[44000] = 32'b00000000000000001111011010111000;
assign LUT_4[44001] = 32'b00000000000000001000100110110000;
assign LUT_4[44002] = 32'b00000000000000001110110101011100;
assign LUT_4[44003] = 32'b00000000000000001000000001010100;
assign LUT_4[44004] = 32'b00000000000000001100011011010100;
assign LUT_4[44005] = 32'b00000000000000000101100111001100;
assign LUT_4[44006] = 32'b00000000000000001011110101111000;
assign LUT_4[44007] = 32'b00000000000000000101000001110000;
assign LUT_4[44008] = 32'b00000000000000001000100111001101;
assign LUT_4[44009] = 32'b00000000000000000001110011000101;
assign LUT_4[44010] = 32'b00000000000000001000000001110001;
assign LUT_4[44011] = 32'b00000000000000000001001101101001;
assign LUT_4[44012] = 32'b00000000000000000101100111101001;
assign LUT_4[44013] = 32'b11111111111111111110110011100001;
assign LUT_4[44014] = 32'b00000000000000000101000010001101;
assign LUT_4[44015] = 32'b11111111111111111110001110000101;
assign LUT_4[44016] = 32'b00000000000000001101001100100110;
assign LUT_4[44017] = 32'b00000000000000000110011000011110;
assign LUT_4[44018] = 32'b00000000000000001100100111001010;
assign LUT_4[44019] = 32'b00000000000000000101110011000010;
assign LUT_4[44020] = 32'b00000000000000001010001101000010;
assign LUT_4[44021] = 32'b00000000000000000011011000111010;
assign LUT_4[44022] = 32'b00000000000000001001100111100110;
assign LUT_4[44023] = 32'b00000000000000000010110011011110;
assign LUT_4[44024] = 32'b00000000000000000110011000111011;
assign LUT_4[44025] = 32'b11111111111111111111100100110011;
assign LUT_4[44026] = 32'b00000000000000000101110011011111;
assign LUT_4[44027] = 32'b11111111111111111110111111010111;
assign LUT_4[44028] = 32'b00000000000000000011011001010111;
assign LUT_4[44029] = 32'b11111111111111111100100101001111;
assign LUT_4[44030] = 32'b00000000000000000010110011111011;
assign LUT_4[44031] = 32'b11111111111111111011111111110011;
assign LUT_4[44032] = 32'b00000000000000001010101101001001;
assign LUT_4[44033] = 32'b00000000000000000011111001000001;
assign LUT_4[44034] = 32'b00000000000000001010000111101101;
assign LUT_4[44035] = 32'b00000000000000000011010011100101;
assign LUT_4[44036] = 32'b00000000000000000111101101100101;
assign LUT_4[44037] = 32'b00000000000000000000111001011101;
assign LUT_4[44038] = 32'b00000000000000000111001000001001;
assign LUT_4[44039] = 32'b00000000000000000000010100000001;
assign LUT_4[44040] = 32'b00000000000000000011111001011110;
assign LUT_4[44041] = 32'b11111111111111111101000101010110;
assign LUT_4[44042] = 32'b00000000000000000011010100000010;
assign LUT_4[44043] = 32'b11111111111111111100011111111010;
assign LUT_4[44044] = 32'b00000000000000000000111001111010;
assign LUT_4[44045] = 32'b11111111111111111010000101110010;
assign LUT_4[44046] = 32'b00000000000000000000010100011110;
assign LUT_4[44047] = 32'b11111111111111111001100000010110;
assign LUT_4[44048] = 32'b00000000000000001000011110110111;
assign LUT_4[44049] = 32'b00000000000000000001101010101111;
assign LUT_4[44050] = 32'b00000000000000000111111001011011;
assign LUT_4[44051] = 32'b00000000000000000001000101010011;
assign LUT_4[44052] = 32'b00000000000000000101011111010011;
assign LUT_4[44053] = 32'b11111111111111111110101011001011;
assign LUT_4[44054] = 32'b00000000000000000100111001110111;
assign LUT_4[44055] = 32'b11111111111111111110000101101111;
assign LUT_4[44056] = 32'b00000000000000000001101011001100;
assign LUT_4[44057] = 32'b11111111111111111010110111000100;
assign LUT_4[44058] = 32'b00000000000000000001000101110000;
assign LUT_4[44059] = 32'b11111111111111111010010001101000;
assign LUT_4[44060] = 32'b11111111111111111110101011101000;
assign LUT_4[44061] = 32'b11111111111111110111110111100000;
assign LUT_4[44062] = 32'b11111111111111111110000110001100;
assign LUT_4[44063] = 32'b11111111111111110111010010000100;
assign LUT_4[44064] = 32'b00000000000000001001001000010000;
assign LUT_4[44065] = 32'b00000000000000000010010100001000;
assign LUT_4[44066] = 32'b00000000000000001000100010110100;
assign LUT_4[44067] = 32'b00000000000000000001101110101100;
assign LUT_4[44068] = 32'b00000000000000000110001000101100;
assign LUT_4[44069] = 32'b11111111111111111111010100100100;
assign LUT_4[44070] = 32'b00000000000000000101100011010000;
assign LUT_4[44071] = 32'b11111111111111111110101111001000;
assign LUT_4[44072] = 32'b00000000000000000010010100100101;
assign LUT_4[44073] = 32'b11111111111111111011100000011101;
assign LUT_4[44074] = 32'b00000000000000000001101111001001;
assign LUT_4[44075] = 32'b11111111111111111010111011000001;
assign LUT_4[44076] = 32'b11111111111111111111010101000001;
assign LUT_4[44077] = 32'b11111111111111111000100000111001;
assign LUT_4[44078] = 32'b11111111111111111110101111100101;
assign LUT_4[44079] = 32'b11111111111111110111111011011101;
assign LUT_4[44080] = 32'b00000000000000000110111001111110;
assign LUT_4[44081] = 32'b00000000000000000000000101110110;
assign LUT_4[44082] = 32'b00000000000000000110010100100010;
assign LUT_4[44083] = 32'b11111111111111111111100000011010;
assign LUT_4[44084] = 32'b00000000000000000011111010011010;
assign LUT_4[44085] = 32'b11111111111111111101000110010010;
assign LUT_4[44086] = 32'b00000000000000000011010100111110;
assign LUT_4[44087] = 32'b11111111111111111100100000110110;
assign LUT_4[44088] = 32'b00000000000000000000000110010011;
assign LUT_4[44089] = 32'b11111111111111111001010010001011;
assign LUT_4[44090] = 32'b11111111111111111111100000110111;
assign LUT_4[44091] = 32'b11111111111111111000101100101111;
assign LUT_4[44092] = 32'b11111111111111111101000110101111;
assign LUT_4[44093] = 32'b11111111111111110110010010100111;
assign LUT_4[44094] = 32'b11111111111111111100100001010011;
assign LUT_4[44095] = 32'b11111111111111110101101101001011;
assign LUT_4[44096] = 32'b00000000000000001100000100011101;
assign LUT_4[44097] = 32'b00000000000000000101010000010101;
assign LUT_4[44098] = 32'b00000000000000001011011111000001;
assign LUT_4[44099] = 32'b00000000000000000100101010111001;
assign LUT_4[44100] = 32'b00000000000000001001000100111001;
assign LUT_4[44101] = 32'b00000000000000000010010000110001;
assign LUT_4[44102] = 32'b00000000000000001000011111011101;
assign LUT_4[44103] = 32'b00000000000000000001101011010101;
assign LUT_4[44104] = 32'b00000000000000000101010000110010;
assign LUT_4[44105] = 32'b11111111111111111110011100101010;
assign LUT_4[44106] = 32'b00000000000000000100101011010110;
assign LUT_4[44107] = 32'b11111111111111111101110111001110;
assign LUT_4[44108] = 32'b00000000000000000010010001001110;
assign LUT_4[44109] = 32'b11111111111111111011011101000110;
assign LUT_4[44110] = 32'b00000000000000000001101011110010;
assign LUT_4[44111] = 32'b11111111111111111010110111101010;
assign LUT_4[44112] = 32'b00000000000000001001110110001011;
assign LUT_4[44113] = 32'b00000000000000000011000010000011;
assign LUT_4[44114] = 32'b00000000000000001001010000101111;
assign LUT_4[44115] = 32'b00000000000000000010011100100111;
assign LUT_4[44116] = 32'b00000000000000000110110110100111;
assign LUT_4[44117] = 32'b00000000000000000000000010011111;
assign LUT_4[44118] = 32'b00000000000000000110010001001011;
assign LUT_4[44119] = 32'b11111111111111111111011101000011;
assign LUT_4[44120] = 32'b00000000000000000011000010100000;
assign LUT_4[44121] = 32'b11111111111111111100001110011000;
assign LUT_4[44122] = 32'b00000000000000000010011101000100;
assign LUT_4[44123] = 32'b11111111111111111011101000111100;
assign LUT_4[44124] = 32'b00000000000000000000000010111100;
assign LUT_4[44125] = 32'b11111111111111111001001110110100;
assign LUT_4[44126] = 32'b11111111111111111111011101100000;
assign LUT_4[44127] = 32'b11111111111111111000101001011000;
assign LUT_4[44128] = 32'b00000000000000001010011111100100;
assign LUT_4[44129] = 32'b00000000000000000011101011011100;
assign LUT_4[44130] = 32'b00000000000000001001111010001000;
assign LUT_4[44131] = 32'b00000000000000000011000110000000;
assign LUT_4[44132] = 32'b00000000000000000111100000000000;
assign LUT_4[44133] = 32'b00000000000000000000101011111000;
assign LUT_4[44134] = 32'b00000000000000000110111010100100;
assign LUT_4[44135] = 32'b00000000000000000000000110011100;
assign LUT_4[44136] = 32'b00000000000000000011101011111001;
assign LUT_4[44137] = 32'b11111111111111111100110111110001;
assign LUT_4[44138] = 32'b00000000000000000011000110011101;
assign LUT_4[44139] = 32'b11111111111111111100010010010101;
assign LUT_4[44140] = 32'b00000000000000000000101100010101;
assign LUT_4[44141] = 32'b11111111111111111001111000001101;
assign LUT_4[44142] = 32'b00000000000000000000000110111001;
assign LUT_4[44143] = 32'b11111111111111111001010010110001;
assign LUT_4[44144] = 32'b00000000000000001000010001010010;
assign LUT_4[44145] = 32'b00000000000000000001011101001010;
assign LUT_4[44146] = 32'b00000000000000000111101011110110;
assign LUT_4[44147] = 32'b00000000000000000000110111101110;
assign LUT_4[44148] = 32'b00000000000000000101010001101110;
assign LUT_4[44149] = 32'b11111111111111111110011101100110;
assign LUT_4[44150] = 32'b00000000000000000100101100010010;
assign LUT_4[44151] = 32'b11111111111111111101111000001010;
assign LUT_4[44152] = 32'b00000000000000000001011101100111;
assign LUT_4[44153] = 32'b11111111111111111010101001011111;
assign LUT_4[44154] = 32'b00000000000000000000111000001011;
assign LUT_4[44155] = 32'b11111111111111111010000100000011;
assign LUT_4[44156] = 32'b11111111111111111110011110000011;
assign LUT_4[44157] = 32'b11111111111111110111101001111011;
assign LUT_4[44158] = 32'b11111111111111111101111000100111;
assign LUT_4[44159] = 32'b11111111111111110111000100011111;
assign LUT_4[44160] = 32'b00000000000000001101010011010001;
assign LUT_4[44161] = 32'b00000000000000000110011111001001;
assign LUT_4[44162] = 32'b00000000000000001100101101110101;
assign LUT_4[44163] = 32'b00000000000000000101111001101101;
assign LUT_4[44164] = 32'b00000000000000001010010011101101;
assign LUT_4[44165] = 32'b00000000000000000011011111100101;
assign LUT_4[44166] = 32'b00000000000000001001101110010001;
assign LUT_4[44167] = 32'b00000000000000000010111010001001;
assign LUT_4[44168] = 32'b00000000000000000110011111100110;
assign LUT_4[44169] = 32'b11111111111111111111101011011110;
assign LUT_4[44170] = 32'b00000000000000000101111010001010;
assign LUT_4[44171] = 32'b11111111111111111111000110000010;
assign LUT_4[44172] = 32'b00000000000000000011100000000010;
assign LUT_4[44173] = 32'b11111111111111111100101011111010;
assign LUT_4[44174] = 32'b00000000000000000010111010100110;
assign LUT_4[44175] = 32'b11111111111111111100000110011110;
assign LUT_4[44176] = 32'b00000000000000001011000100111111;
assign LUT_4[44177] = 32'b00000000000000000100010000110111;
assign LUT_4[44178] = 32'b00000000000000001010011111100011;
assign LUT_4[44179] = 32'b00000000000000000011101011011011;
assign LUT_4[44180] = 32'b00000000000000001000000101011011;
assign LUT_4[44181] = 32'b00000000000000000001010001010011;
assign LUT_4[44182] = 32'b00000000000000000111011111111111;
assign LUT_4[44183] = 32'b00000000000000000000101011110111;
assign LUT_4[44184] = 32'b00000000000000000100010001010100;
assign LUT_4[44185] = 32'b11111111111111111101011101001100;
assign LUT_4[44186] = 32'b00000000000000000011101011111000;
assign LUT_4[44187] = 32'b11111111111111111100110111110000;
assign LUT_4[44188] = 32'b00000000000000000001010001110000;
assign LUT_4[44189] = 32'b11111111111111111010011101101000;
assign LUT_4[44190] = 32'b00000000000000000000101100010100;
assign LUT_4[44191] = 32'b11111111111111111001111000001100;
assign LUT_4[44192] = 32'b00000000000000001011101110011000;
assign LUT_4[44193] = 32'b00000000000000000100111010010000;
assign LUT_4[44194] = 32'b00000000000000001011001000111100;
assign LUT_4[44195] = 32'b00000000000000000100010100110100;
assign LUT_4[44196] = 32'b00000000000000001000101110110100;
assign LUT_4[44197] = 32'b00000000000000000001111010101100;
assign LUT_4[44198] = 32'b00000000000000001000001001011000;
assign LUT_4[44199] = 32'b00000000000000000001010101010000;
assign LUT_4[44200] = 32'b00000000000000000100111010101101;
assign LUT_4[44201] = 32'b11111111111111111110000110100101;
assign LUT_4[44202] = 32'b00000000000000000100010101010001;
assign LUT_4[44203] = 32'b11111111111111111101100001001001;
assign LUT_4[44204] = 32'b00000000000000000001111011001001;
assign LUT_4[44205] = 32'b11111111111111111011000111000001;
assign LUT_4[44206] = 32'b00000000000000000001010101101101;
assign LUT_4[44207] = 32'b11111111111111111010100001100101;
assign LUT_4[44208] = 32'b00000000000000001001100000000110;
assign LUT_4[44209] = 32'b00000000000000000010101011111110;
assign LUT_4[44210] = 32'b00000000000000001000111010101010;
assign LUT_4[44211] = 32'b00000000000000000010000110100010;
assign LUT_4[44212] = 32'b00000000000000000110100000100010;
assign LUT_4[44213] = 32'b11111111111111111111101100011010;
assign LUT_4[44214] = 32'b00000000000000000101111011000110;
assign LUT_4[44215] = 32'b11111111111111111111000110111110;
assign LUT_4[44216] = 32'b00000000000000000010101100011011;
assign LUT_4[44217] = 32'b11111111111111111011111000010011;
assign LUT_4[44218] = 32'b00000000000000000010000110111111;
assign LUT_4[44219] = 32'b11111111111111111011010010110111;
assign LUT_4[44220] = 32'b11111111111111111111101100110111;
assign LUT_4[44221] = 32'b11111111111111111000111000101111;
assign LUT_4[44222] = 32'b11111111111111111111000111011011;
assign LUT_4[44223] = 32'b11111111111111111000010011010011;
assign LUT_4[44224] = 32'b00000000000000001110101010100101;
assign LUT_4[44225] = 32'b00000000000000000111110110011101;
assign LUT_4[44226] = 32'b00000000000000001110000101001001;
assign LUT_4[44227] = 32'b00000000000000000111010001000001;
assign LUT_4[44228] = 32'b00000000000000001011101011000001;
assign LUT_4[44229] = 32'b00000000000000000100110110111001;
assign LUT_4[44230] = 32'b00000000000000001011000101100101;
assign LUT_4[44231] = 32'b00000000000000000100010001011101;
assign LUT_4[44232] = 32'b00000000000000000111110110111010;
assign LUT_4[44233] = 32'b00000000000000000001000010110010;
assign LUT_4[44234] = 32'b00000000000000000111010001011110;
assign LUT_4[44235] = 32'b00000000000000000000011101010110;
assign LUT_4[44236] = 32'b00000000000000000100110111010110;
assign LUT_4[44237] = 32'b11111111111111111110000011001110;
assign LUT_4[44238] = 32'b00000000000000000100010001111010;
assign LUT_4[44239] = 32'b11111111111111111101011101110010;
assign LUT_4[44240] = 32'b00000000000000001100011100010011;
assign LUT_4[44241] = 32'b00000000000000000101101000001011;
assign LUT_4[44242] = 32'b00000000000000001011110110110111;
assign LUT_4[44243] = 32'b00000000000000000101000010101111;
assign LUT_4[44244] = 32'b00000000000000001001011100101111;
assign LUT_4[44245] = 32'b00000000000000000010101000100111;
assign LUT_4[44246] = 32'b00000000000000001000110111010011;
assign LUT_4[44247] = 32'b00000000000000000010000011001011;
assign LUT_4[44248] = 32'b00000000000000000101101000101000;
assign LUT_4[44249] = 32'b11111111111111111110110100100000;
assign LUT_4[44250] = 32'b00000000000000000101000011001100;
assign LUT_4[44251] = 32'b11111111111111111110001111000100;
assign LUT_4[44252] = 32'b00000000000000000010101001000100;
assign LUT_4[44253] = 32'b11111111111111111011110100111100;
assign LUT_4[44254] = 32'b00000000000000000010000011101000;
assign LUT_4[44255] = 32'b11111111111111111011001111100000;
assign LUT_4[44256] = 32'b00000000000000001101000101101100;
assign LUT_4[44257] = 32'b00000000000000000110010001100100;
assign LUT_4[44258] = 32'b00000000000000001100100000010000;
assign LUT_4[44259] = 32'b00000000000000000101101100001000;
assign LUT_4[44260] = 32'b00000000000000001010000110001000;
assign LUT_4[44261] = 32'b00000000000000000011010010000000;
assign LUT_4[44262] = 32'b00000000000000001001100000101100;
assign LUT_4[44263] = 32'b00000000000000000010101100100100;
assign LUT_4[44264] = 32'b00000000000000000110010010000001;
assign LUT_4[44265] = 32'b11111111111111111111011101111001;
assign LUT_4[44266] = 32'b00000000000000000101101100100101;
assign LUT_4[44267] = 32'b11111111111111111110111000011101;
assign LUT_4[44268] = 32'b00000000000000000011010010011101;
assign LUT_4[44269] = 32'b11111111111111111100011110010101;
assign LUT_4[44270] = 32'b00000000000000000010101101000001;
assign LUT_4[44271] = 32'b11111111111111111011111000111001;
assign LUT_4[44272] = 32'b00000000000000001010110111011010;
assign LUT_4[44273] = 32'b00000000000000000100000011010010;
assign LUT_4[44274] = 32'b00000000000000001010010001111110;
assign LUT_4[44275] = 32'b00000000000000000011011101110110;
assign LUT_4[44276] = 32'b00000000000000000111110111110110;
assign LUT_4[44277] = 32'b00000000000000000001000011101110;
assign LUT_4[44278] = 32'b00000000000000000111010010011010;
assign LUT_4[44279] = 32'b00000000000000000000011110010010;
assign LUT_4[44280] = 32'b00000000000000000100000011101111;
assign LUT_4[44281] = 32'b11111111111111111101001111100111;
assign LUT_4[44282] = 32'b00000000000000000011011110010011;
assign LUT_4[44283] = 32'b11111111111111111100101010001011;
assign LUT_4[44284] = 32'b00000000000000000001000100001011;
assign LUT_4[44285] = 32'b11111111111111111010010000000011;
assign LUT_4[44286] = 32'b00000000000000000000011110101111;
assign LUT_4[44287] = 32'b11111111111111111001101010100111;
assign LUT_4[44288] = 32'b00000000000000001111101000101100;
assign LUT_4[44289] = 32'b00000000000000001000110100100100;
assign LUT_4[44290] = 32'b00000000000000001111000011010000;
assign LUT_4[44291] = 32'b00000000000000001000001111001000;
assign LUT_4[44292] = 32'b00000000000000001100101001001000;
assign LUT_4[44293] = 32'b00000000000000000101110101000000;
assign LUT_4[44294] = 32'b00000000000000001100000011101100;
assign LUT_4[44295] = 32'b00000000000000000101001111100100;
assign LUT_4[44296] = 32'b00000000000000001000110101000001;
assign LUT_4[44297] = 32'b00000000000000000010000000111001;
assign LUT_4[44298] = 32'b00000000000000001000001111100101;
assign LUT_4[44299] = 32'b00000000000000000001011011011101;
assign LUT_4[44300] = 32'b00000000000000000101110101011101;
assign LUT_4[44301] = 32'b11111111111111111111000001010101;
assign LUT_4[44302] = 32'b00000000000000000101010000000001;
assign LUT_4[44303] = 32'b11111111111111111110011011111001;
assign LUT_4[44304] = 32'b00000000000000001101011010011010;
assign LUT_4[44305] = 32'b00000000000000000110100110010010;
assign LUT_4[44306] = 32'b00000000000000001100110100111110;
assign LUT_4[44307] = 32'b00000000000000000110000000110110;
assign LUT_4[44308] = 32'b00000000000000001010011010110110;
assign LUT_4[44309] = 32'b00000000000000000011100110101110;
assign LUT_4[44310] = 32'b00000000000000001001110101011010;
assign LUT_4[44311] = 32'b00000000000000000011000001010010;
assign LUT_4[44312] = 32'b00000000000000000110100110101111;
assign LUT_4[44313] = 32'b11111111111111111111110010100111;
assign LUT_4[44314] = 32'b00000000000000000110000001010011;
assign LUT_4[44315] = 32'b11111111111111111111001101001011;
assign LUT_4[44316] = 32'b00000000000000000011100111001011;
assign LUT_4[44317] = 32'b11111111111111111100110011000011;
assign LUT_4[44318] = 32'b00000000000000000011000001101111;
assign LUT_4[44319] = 32'b11111111111111111100001101100111;
assign LUT_4[44320] = 32'b00000000000000001110000011110011;
assign LUT_4[44321] = 32'b00000000000000000111001111101011;
assign LUT_4[44322] = 32'b00000000000000001101011110010111;
assign LUT_4[44323] = 32'b00000000000000000110101010001111;
assign LUT_4[44324] = 32'b00000000000000001011000100001111;
assign LUT_4[44325] = 32'b00000000000000000100010000000111;
assign LUT_4[44326] = 32'b00000000000000001010011110110011;
assign LUT_4[44327] = 32'b00000000000000000011101010101011;
assign LUT_4[44328] = 32'b00000000000000000111010000001000;
assign LUT_4[44329] = 32'b00000000000000000000011100000000;
assign LUT_4[44330] = 32'b00000000000000000110101010101100;
assign LUT_4[44331] = 32'b11111111111111111111110110100100;
assign LUT_4[44332] = 32'b00000000000000000100010000100100;
assign LUT_4[44333] = 32'b11111111111111111101011100011100;
assign LUT_4[44334] = 32'b00000000000000000011101011001000;
assign LUT_4[44335] = 32'b11111111111111111100110111000000;
assign LUT_4[44336] = 32'b00000000000000001011110101100001;
assign LUT_4[44337] = 32'b00000000000000000101000001011001;
assign LUT_4[44338] = 32'b00000000000000001011010000000101;
assign LUT_4[44339] = 32'b00000000000000000100011011111101;
assign LUT_4[44340] = 32'b00000000000000001000110101111101;
assign LUT_4[44341] = 32'b00000000000000000010000001110101;
assign LUT_4[44342] = 32'b00000000000000001000010000100001;
assign LUT_4[44343] = 32'b00000000000000000001011100011001;
assign LUT_4[44344] = 32'b00000000000000000101000001110110;
assign LUT_4[44345] = 32'b11111111111111111110001101101110;
assign LUT_4[44346] = 32'b00000000000000000100011100011010;
assign LUT_4[44347] = 32'b11111111111111111101101000010010;
assign LUT_4[44348] = 32'b00000000000000000010000010010010;
assign LUT_4[44349] = 32'b11111111111111111011001110001010;
assign LUT_4[44350] = 32'b00000000000000000001011100110110;
assign LUT_4[44351] = 32'b11111111111111111010101000101110;
assign LUT_4[44352] = 32'b00000000000000010001000000000000;
assign LUT_4[44353] = 32'b00000000000000001010001011111000;
assign LUT_4[44354] = 32'b00000000000000010000011010100100;
assign LUT_4[44355] = 32'b00000000000000001001100110011100;
assign LUT_4[44356] = 32'b00000000000000001110000000011100;
assign LUT_4[44357] = 32'b00000000000000000111001100010100;
assign LUT_4[44358] = 32'b00000000000000001101011011000000;
assign LUT_4[44359] = 32'b00000000000000000110100110111000;
assign LUT_4[44360] = 32'b00000000000000001010001100010101;
assign LUT_4[44361] = 32'b00000000000000000011011000001101;
assign LUT_4[44362] = 32'b00000000000000001001100110111001;
assign LUT_4[44363] = 32'b00000000000000000010110010110001;
assign LUT_4[44364] = 32'b00000000000000000111001100110001;
assign LUT_4[44365] = 32'b00000000000000000000011000101001;
assign LUT_4[44366] = 32'b00000000000000000110100111010101;
assign LUT_4[44367] = 32'b11111111111111111111110011001101;
assign LUT_4[44368] = 32'b00000000000000001110110001101110;
assign LUT_4[44369] = 32'b00000000000000000111111101100110;
assign LUT_4[44370] = 32'b00000000000000001110001100010010;
assign LUT_4[44371] = 32'b00000000000000000111011000001010;
assign LUT_4[44372] = 32'b00000000000000001011110010001010;
assign LUT_4[44373] = 32'b00000000000000000100111110000010;
assign LUT_4[44374] = 32'b00000000000000001011001100101110;
assign LUT_4[44375] = 32'b00000000000000000100011000100110;
assign LUT_4[44376] = 32'b00000000000000000111111110000011;
assign LUT_4[44377] = 32'b00000000000000000001001001111011;
assign LUT_4[44378] = 32'b00000000000000000111011000100111;
assign LUT_4[44379] = 32'b00000000000000000000100100011111;
assign LUT_4[44380] = 32'b00000000000000000100111110011111;
assign LUT_4[44381] = 32'b11111111111111111110001010010111;
assign LUT_4[44382] = 32'b00000000000000000100011001000011;
assign LUT_4[44383] = 32'b11111111111111111101100100111011;
assign LUT_4[44384] = 32'b00000000000000001111011011000111;
assign LUT_4[44385] = 32'b00000000000000001000100110111111;
assign LUT_4[44386] = 32'b00000000000000001110110101101011;
assign LUT_4[44387] = 32'b00000000000000001000000001100011;
assign LUT_4[44388] = 32'b00000000000000001100011011100011;
assign LUT_4[44389] = 32'b00000000000000000101100111011011;
assign LUT_4[44390] = 32'b00000000000000001011110110000111;
assign LUT_4[44391] = 32'b00000000000000000101000001111111;
assign LUT_4[44392] = 32'b00000000000000001000100111011100;
assign LUT_4[44393] = 32'b00000000000000000001110011010100;
assign LUT_4[44394] = 32'b00000000000000001000000010000000;
assign LUT_4[44395] = 32'b00000000000000000001001101111000;
assign LUT_4[44396] = 32'b00000000000000000101100111111000;
assign LUT_4[44397] = 32'b11111111111111111110110011110000;
assign LUT_4[44398] = 32'b00000000000000000101000010011100;
assign LUT_4[44399] = 32'b11111111111111111110001110010100;
assign LUT_4[44400] = 32'b00000000000000001101001100110101;
assign LUT_4[44401] = 32'b00000000000000000110011000101101;
assign LUT_4[44402] = 32'b00000000000000001100100111011001;
assign LUT_4[44403] = 32'b00000000000000000101110011010001;
assign LUT_4[44404] = 32'b00000000000000001010001101010001;
assign LUT_4[44405] = 32'b00000000000000000011011001001001;
assign LUT_4[44406] = 32'b00000000000000001001100111110101;
assign LUT_4[44407] = 32'b00000000000000000010110011101101;
assign LUT_4[44408] = 32'b00000000000000000110011001001010;
assign LUT_4[44409] = 32'b11111111111111111111100101000010;
assign LUT_4[44410] = 32'b00000000000000000101110011101110;
assign LUT_4[44411] = 32'b11111111111111111110111111100110;
assign LUT_4[44412] = 32'b00000000000000000011011001100110;
assign LUT_4[44413] = 32'b11111111111111111100100101011110;
assign LUT_4[44414] = 32'b00000000000000000010110100001010;
assign LUT_4[44415] = 32'b11111111111111111100000000000010;
assign LUT_4[44416] = 32'b00000000000000010010001110110100;
assign LUT_4[44417] = 32'b00000000000000001011011010101100;
assign LUT_4[44418] = 32'b00000000000000010001101001011000;
assign LUT_4[44419] = 32'b00000000000000001010110101010000;
assign LUT_4[44420] = 32'b00000000000000001111001111010000;
assign LUT_4[44421] = 32'b00000000000000001000011011001000;
assign LUT_4[44422] = 32'b00000000000000001110101001110100;
assign LUT_4[44423] = 32'b00000000000000000111110101101100;
assign LUT_4[44424] = 32'b00000000000000001011011011001001;
assign LUT_4[44425] = 32'b00000000000000000100100111000001;
assign LUT_4[44426] = 32'b00000000000000001010110101101101;
assign LUT_4[44427] = 32'b00000000000000000100000001100101;
assign LUT_4[44428] = 32'b00000000000000001000011011100101;
assign LUT_4[44429] = 32'b00000000000000000001100111011101;
assign LUT_4[44430] = 32'b00000000000000000111110110001001;
assign LUT_4[44431] = 32'b00000000000000000001000010000001;
assign LUT_4[44432] = 32'b00000000000000010000000000100010;
assign LUT_4[44433] = 32'b00000000000000001001001100011010;
assign LUT_4[44434] = 32'b00000000000000001111011011000110;
assign LUT_4[44435] = 32'b00000000000000001000100110111110;
assign LUT_4[44436] = 32'b00000000000000001101000000111110;
assign LUT_4[44437] = 32'b00000000000000000110001100110110;
assign LUT_4[44438] = 32'b00000000000000001100011011100010;
assign LUT_4[44439] = 32'b00000000000000000101100111011010;
assign LUT_4[44440] = 32'b00000000000000001001001100110111;
assign LUT_4[44441] = 32'b00000000000000000010011000101111;
assign LUT_4[44442] = 32'b00000000000000001000100111011011;
assign LUT_4[44443] = 32'b00000000000000000001110011010011;
assign LUT_4[44444] = 32'b00000000000000000110001101010011;
assign LUT_4[44445] = 32'b11111111111111111111011001001011;
assign LUT_4[44446] = 32'b00000000000000000101100111110111;
assign LUT_4[44447] = 32'b11111111111111111110110011101111;
assign LUT_4[44448] = 32'b00000000000000010000101001111011;
assign LUT_4[44449] = 32'b00000000000000001001110101110011;
assign LUT_4[44450] = 32'b00000000000000010000000100011111;
assign LUT_4[44451] = 32'b00000000000000001001010000010111;
assign LUT_4[44452] = 32'b00000000000000001101101010010111;
assign LUT_4[44453] = 32'b00000000000000000110110110001111;
assign LUT_4[44454] = 32'b00000000000000001101000100111011;
assign LUT_4[44455] = 32'b00000000000000000110010000110011;
assign LUT_4[44456] = 32'b00000000000000001001110110010000;
assign LUT_4[44457] = 32'b00000000000000000011000010001000;
assign LUT_4[44458] = 32'b00000000000000001001010000110100;
assign LUT_4[44459] = 32'b00000000000000000010011100101100;
assign LUT_4[44460] = 32'b00000000000000000110110110101100;
assign LUT_4[44461] = 32'b00000000000000000000000010100100;
assign LUT_4[44462] = 32'b00000000000000000110010001010000;
assign LUT_4[44463] = 32'b11111111111111111111011101001000;
assign LUT_4[44464] = 32'b00000000000000001110011011101001;
assign LUT_4[44465] = 32'b00000000000000000111100111100001;
assign LUT_4[44466] = 32'b00000000000000001101110110001101;
assign LUT_4[44467] = 32'b00000000000000000111000010000101;
assign LUT_4[44468] = 32'b00000000000000001011011100000101;
assign LUT_4[44469] = 32'b00000000000000000100100111111101;
assign LUT_4[44470] = 32'b00000000000000001010110110101001;
assign LUT_4[44471] = 32'b00000000000000000100000010100001;
assign LUT_4[44472] = 32'b00000000000000000111100111111110;
assign LUT_4[44473] = 32'b00000000000000000000110011110110;
assign LUT_4[44474] = 32'b00000000000000000111000010100010;
assign LUT_4[44475] = 32'b00000000000000000000001110011010;
assign LUT_4[44476] = 32'b00000000000000000100101000011010;
assign LUT_4[44477] = 32'b11111111111111111101110100010010;
assign LUT_4[44478] = 32'b00000000000000000100000010111110;
assign LUT_4[44479] = 32'b11111111111111111101001110110110;
assign LUT_4[44480] = 32'b00000000000000010011100110001000;
assign LUT_4[44481] = 32'b00000000000000001100110010000000;
assign LUT_4[44482] = 32'b00000000000000010011000000101100;
assign LUT_4[44483] = 32'b00000000000000001100001100100100;
assign LUT_4[44484] = 32'b00000000000000010000100110100100;
assign LUT_4[44485] = 32'b00000000000000001001110010011100;
assign LUT_4[44486] = 32'b00000000000000010000000001001000;
assign LUT_4[44487] = 32'b00000000000000001001001101000000;
assign LUT_4[44488] = 32'b00000000000000001100110010011101;
assign LUT_4[44489] = 32'b00000000000000000101111110010101;
assign LUT_4[44490] = 32'b00000000000000001100001101000001;
assign LUT_4[44491] = 32'b00000000000000000101011000111001;
assign LUT_4[44492] = 32'b00000000000000001001110010111001;
assign LUT_4[44493] = 32'b00000000000000000010111110110001;
assign LUT_4[44494] = 32'b00000000000000001001001101011101;
assign LUT_4[44495] = 32'b00000000000000000010011001010101;
assign LUT_4[44496] = 32'b00000000000000010001010111110110;
assign LUT_4[44497] = 32'b00000000000000001010100011101110;
assign LUT_4[44498] = 32'b00000000000000010000110010011010;
assign LUT_4[44499] = 32'b00000000000000001001111110010010;
assign LUT_4[44500] = 32'b00000000000000001110011000010010;
assign LUT_4[44501] = 32'b00000000000000000111100100001010;
assign LUT_4[44502] = 32'b00000000000000001101110010110110;
assign LUT_4[44503] = 32'b00000000000000000110111110101110;
assign LUT_4[44504] = 32'b00000000000000001010100100001011;
assign LUT_4[44505] = 32'b00000000000000000011110000000011;
assign LUT_4[44506] = 32'b00000000000000001001111110101111;
assign LUT_4[44507] = 32'b00000000000000000011001010100111;
assign LUT_4[44508] = 32'b00000000000000000111100100100111;
assign LUT_4[44509] = 32'b00000000000000000000110000011111;
assign LUT_4[44510] = 32'b00000000000000000110111111001011;
assign LUT_4[44511] = 32'b00000000000000000000001011000011;
assign LUT_4[44512] = 32'b00000000000000010010000001001111;
assign LUT_4[44513] = 32'b00000000000000001011001101000111;
assign LUT_4[44514] = 32'b00000000000000010001011011110011;
assign LUT_4[44515] = 32'b00000000000000001010100111101011;
assign LUT_4[44516] = 32'b00000000000000001111000001101011;
assign LUT_4[44517] = 32'b00000000000000001000001101100011;
assign LUT_4[44518] = 32'b00000000000000001110011100001111;
assign LUT_4[44519] = 32'b00000000000000000111101000000111;
assign LUT_4[44520] = 32'b00000000000000001011001101100100;
assign LUT_4[44521] = 32'b00000000000000000100011001011100;
assign LUT_4[44522] = 32'b00000000000000001010101000001000;
assign LUT_4[44523] = 32'b00000000000000000011110100000000;
assign LUT_4[44524] = 32'b00000000000000001000001110000000;
assign LUT_4[44525] = 32'b00000000000000000001011001111000;
assign LUT_4[44526] = 32'b00000000000000000111101000100100;
assign LUT_4[44527] = 32'b00000000000000000000110100011100;
assign LUT_4[44528] = 32'b00000000000000001111110010111101;
assign LUT_4[44529] = 32'b00000000000000001000111110110101;
assign LUT_4[44530] = 32'b00000000000000001111001101100001;
assign LUT_4[44531] = 32'b00000000000000001000011001011001;
assign LUT_4[44532] = 32'b00000000000000001100110011011001;
assign LUT_4[44533] = 32'b00000000000000000101111111010001;
assign LUT_4[44534] = 32'b00000000000000001100001101111101;
assign LUT_4[44535] = 32'b00000000000000000101011001110101;
assign LUT_4[44536] = 32'b00000000000000001000111111010010;
assign LUT_4[44537] = 32'b00000000000000000010001011001010;
assign LUT_4[44538] = 32'b00000000000000001000011001110110;
assign LUT_4[44539] = 32'b00000000000000000001100101101110;
assign LUT_4[44540] = 32'b00000000000000000101111111101110;
assign LUT_4[44541] = 32'b11111111111111111111001011100110;
assign LUT_4[44542] = 32'b00000000000000000101011010010010;
assign LUT_4[44543] = 32'b11111111111111111110100110001010;
assign LUT_4[44544] = 32'b00000000000000001001110001010001;
assign LUT_4[44545] = 32'b00000000000000000010111101001001;
assign LUT_4[44546] = 32'b00000000000000001001001011110101;
assign LUT_4[44547] = 32'b00000000000000000010010111101101;
assign LUT_4[44548] = 32'b00000000000000000110110001101101;
assign LUT_4[44549] = 32'b11111111111111111111111101100101;
assign LUT_4[44550] = 32'b00000000000000000110001100010001;
assign LUT_4[44551] = 32'b11111111111111111111011000001001;
assign LUT_4[44552] = 32'b00000000000000000010111101100110;
assign LUT_4[44553] = 32'b11111111111111111100001001011110;
assign LUT_4[44554] = 32'b00000000000000000010011000001010;
assign LUT_4[44555] = 32'b11111111111111111011100100000010;
assign LUT_4[44556] = 32'b11111111111111111111111110000010;
assign LUT_4[44557] = 32'b11111111111111111001001001111010;
assign LUT_4[44558] = 32'b11111111111111111111011000100110;
assign LUT_4[44559] = 32'b11111111111111111000100100011110;
assign LUT_4[44560] = 32'b00000000000000000111100010111111;
assign LUT_4[44561] = 32'b00000000000000000000101110110111;
assign LUT_4[44562] = 32'b00000000000000000110111101100011;
assign LUT_4[44563] = 32'b00000000000000000000001001011011;
assign LUT_4[44564] = 32'b00000000000000000100100011011011;
assign LUT_4[44565] = 32'b11111111111111111101101111010011;
assign LUT_4[44566] = 32'b00000000000000000011111101111111;
assign LUT_4[44567] = 32'b11111111111111111101001001110111;
assign LUT_4[44568] = 32'b00000000000000000000101111010100;
assign LUT_4[44569] = 32'b11111111111111111001111011001100;
assign LUT_4[44570] = 32'b00000000000000000000001001111000;
assign LUT_4[44571] = 32'b11111111111111111001010101110000;
assign LUT_4[44572] = 32'b11111111111111111101101111110000;
assign LUT_4[44573] = 32'b11111111111111110110111011101000;
assign LUT_4[44574] = 32'b11111111111111111101001010010100;
assign LUT_4[44575] = 32'b11111111111111110110010110001100;
assign LUT_4[44576] = 32'b00000000000000001000001100011000;
assign LUT_4[44577] = 32'b00000000000000000001011000010000;
assign LUT_4[44578] = 32'b00000000000000000111100110111100;
assign LUT_4[44579] = 32'b00000000000000000000110010110100;
assign LUT_4[44580] = 32'b00000000000000000101001100110100;
assign LUT_4[44581] = 32'b11111111111111111110011000101100;
assign LUT_4[44582] = 32'b00000000000000000100100111011000;
assign LUT_4[44583] = 32'b11111111111111111101110011010000;
assign LUT_4[44584] = 32'b00000000000000000001011000101101;
assign LUT_4[44585] = 32'b11111111111111111010100100100101;
assign LUT_4[44586] = 32'b00000000000000000000110011010001;
assign LUT_4[44587] = 32'b11111111111111111001111111001001;
assign LUT_4[44588] = 32'b11111111111111111110011001001001;
assign LUT_4[44589] = 32'b11111111111111110111100101000001;
assign LUT_4[44590] = 32'b11111111111111111101110011101101;
assign LUT_4[44591] = 32'b11111111111111110110111111100101;
assign LUT_4[44592] = 32'b00000000000000000101111110000110;
assign LUT_4[44593] = 32'b11111111111111111111001001111110;
assign LUT_4[44594] = 32'b00000000000000000101011000101010;
assign LUT_4[44595] = 32'b11111111111111111110100100100010;
assign LUT_4[44596] = 32'b00000000000000000010111110100010;
assign LUT_4[44597] = 32'b11111111111111111100001010011010;
assign LUT_4[44598] = 32'b00000000000000000010011001000110;
assign LUT_4[44599] = 32'b11111111111111111011100100111110;
assign LUT_4[44600] = 32'b11111111111111111111001010011011;
assign LUT_4[44601] = 32'b11111111111111111000010110010011;
assign LUT_4[44602] = 32'b11111111111111111110100100111111;
assign LUT_4[44603] = 32'b11111111111111110111110000110111;
assign LUT_4[44604] = 32'b11111111111111111100001010110111;
assign LUT_4[44605] = 32'b11111111111111110101010110101111;
assign LUT_4[44606] = 32'b11111111111111111011100101011011;
assign LUT_4[44607] = 32'b11111111111111110100110001010011;
assign LUT_4[44608] = 32'b00000000000000001011001000100101;
assign LUT_4[44609] = 32'b00000000000000000100010100011101;
assign LUT_4[44610] = 32'b00000000000000001010100011001001;
assign LUT_4[44611] = 32'b00000000000000000011101111000001;
assign LUT_4[44612] = 32'b00000000000000001000001001000001;
assign LUT_4[44613] = 32'b00000000000000000001010100111001;
assign LUT_4[44614] = 32'b00000000000000000111100011100101;
assign LUT_4[44615] = 32'b00000000000000000000101111011101;
assign LUT_4[44616] = 32'b00000000000000000100010100111010;
assign LUT_4[44617] = 32'b11111111111111111101100000110010;
assign LUT_4[44618] = 32'b00000000000000000011101111011110;
assign LUT_4[44619] = 32'b11111111111111111100111011010110;
assign LUT_4[44620] = 32'b00000000000000000001010101010110;
assign LUT_4[44621] = 32'b11111111111111111010100001001110;
assign LUT_4[44622] = 32'b00000000000000000000101111111010;
assign LUT_4[44623] = 32'b11111111111111111001111011110010;
assign LUT_4[44624] = 32'b00000000000000001000111010010011;
assign LUT_4[44625] = 32'b00000000000000000010000110001011;
assign LUT_4[44626] = 32'b00000000000000001000010100110111;
assign LUT_4[44627] = 32'b00000000000000000001100000101111;
assign LUT_4[44628] = 32'b00000000000000000101111010101111;
assign LUT_4[44629] = 32'b11111111111111111111000110100111;
assign LUT_4[44630] = 32'b00000000000000000101010101010011;
assign LUT_4[44631] = 32'b11111111111111111110100001001011;
assign LUT_4[44632] = 32'b00000000000000000010000110101000;
assign LUT_4[44633] = 32'b11111111111111111011010010100000;
assign LUT_4[44634] = 32'b00000000000000000001100001001100;
assign LUT_4[44635] = 32'b11111111111111111010101101000100;
assign LUT_4[44636] = 32'b11111111111111111111000111000100;
assign LUT_4[44637] = 32'b11111111111111111000010010111100;
assign LUT_4[44638] = 32'b11111111111111111110100001101000;
assign LUT_4[44639] = 32'b11111111111111110111101101100000;
assign LUT_4[44640] = 32'b00000000000000001001100011101100;
assign LUT_4[44641] = 32'b00000000000000000010101111100100;
assign LUT_4[44642] = 32'b00000000000000001000111110010000;
assign LUT_4[44643] = 32'b00000000000000000010001010001000;
assign LUT_4[44644] = 32'b00000000000000000110100100001000;
assign LUT_4[44645] = 32'b11111111111111111111110000000000;
assign LUT_4[44646] = 32'b00000000000000000101111110101100;
assign LUT_4[44647] = 32'b11111111111111111111001010100100;
assign LUT_4[44648] = 32'b00000000000000000010110000000001;
assign LUT_4[44649] = 32'b11111111111111111011111011111001;
assign LUT_4[44650] = 32'b00000000000000000010001010100101;
assign LUT_4[44651] = 32'b11111111111111111011010110011101;
assign LUT_4[44652] = 32'b11111111111111111111110000011101;
assign LUT_4[44653] = 32'b11111111111111111000111100010101;
assign LUT_4[44654] = 32'b11111111111111111111001011000001;
assign LUT_4[44655] = 32'b11111111111111111000010110111001;
assign LUT_4[44656] = 32'b00000000000000000111010101011010;
assign LUT_4[44657] = 32'b00000000000000000000100001010010;
assign LUT_4[44658] = 32'b00000000000000000110101111111110;
assign LUT_4[44659] = 32'b11111111111111111111111011110110;
assign LUT_4[44660] = 32'b00000000000000000100010101110110;
assign LUT_4[44661] = 32'b11111111111111111101100001101110;
assign LUT_4[44662] = 32'b00000000000000000011110000011010;
assign LUT_4[44663] = 32'b11111111111111111100111100010010;
assign LUT_4[44664] = 32'b00000000000000000000100001101111;
assign LUT_4[44665] = 32'b11111111111111111001101101100111;
assign LUT_4[44666] = 32'b11111111111111111111111100010011;
assign LUT_4[44667] = 32'b11111111111111111001001000001011;
assign LUT_4[44668] = 32'b11111111111111111101100010001011;
assign LUT_4[44669] = 32'b11111111111111110110101110000011;
assign LUT_4[44670] = 32'b11111111111111111100111100101111;
assign LUT_4[44671] = 32'b11111111111111110110001000100111;
assign LUT_4[44672] = 32'b00000000000000001100010111011001;
assign LUT_4[44673] = 32'b00000000000000000101100011010001;
assign LUT_4[44674] = 32'b00000000000000001011110001111101;
assign LUT_4[44675] = 32'b00000000000000000100111101110101;
assign LUT_4[44676] = 32'b00000000000000001001010111110101;
assign LUT_4[44677] = 32'b00000000000000000010100011101101;
assign LUT_4[44678] = 32'b00000000000000001000110010011001;
assign LUT_4[44679] = 32'b00000000000000000001111110010001;
assign LUT_4[44680] = 32'b00000000000000000101100011101110;
assign LUT_4[44681] = 32'b11111111111111111110101111100110;
assign LUT_4[44682] = 32'b00000000000000000100111110010010;
assign LUT_4[44683] = 32'b11111111111111111110001010001010;
assign LUT_4[44684] = 32'b00000000000000000010100100001010;
assign LUT_4[44685] = 32'b11111111111111111011110000000010;
assign LUT_4[44686] = 32'b00000000000000000001111110101110;
assign LUT_4[44687] = 32'b11111111111111111011001010100110;
assign LUT_4[44688] = 32'b00000000000000001010001001000111;
assign LUT_4[44689] = 32'b00000000000000000011010100111111;
assign LUT_4[44690] = 32'b00000000000000001001100011101011;
assign LUT_4[44691] = 32'b00000000000000000010101111100011;
assign LUT_4[44692] = 32'b00000000000000000111001001100011;
assign LUT_4[44693] = 32'b00000000000000000000010101011011;
assign LUT_4[44694] = 32'b00000000000000000110100100000111;
assign LUT_4[44695] = 32'b11111111111111111111101111111111;
assign LUT_4[44696] = 32'b00000000000000000011010101011100;
assign LUT_4[44697] = 32'b11111111111111111100100001010100;
assign LUT_4[44698] = 32'b00000000000000000010110000000000;
assign LUT_4[44699] = 32'b11111111111111111011111011111000;
assign LUT_4[44700] = 32'b00000000000000000000010101111000;
assign LUT_4[44701] = 32'b11111111111111111001100001110000;
assign LUT_4[44702] = 32'b11111111111111111111110000011100;
assign LUT_4[44703] = 32'b11111111111111111000111100010100;
assign LUT_4[44704] = 32'b00000000000000001010110010100000;
assign LUT_4[44705] = 32'b00000000000000000011111110011000;
assign LUT_4[44706] = 32'b00000000000000001010001101000100;
assign LUT_4[44707] = 32'b00000000000000000011011000111100;
assign LUT_4[44708] = 32'b00000000000000000111110010111100;
assign LUT_4[44709] = 32'b00000000000000000000111110110100;
assign LUT_4[44710] = 32'b00000000000000000111001101100000;
assign LUT_4[44711] = 32'b00000000000000000000011001011000;
assign LUT_4[44712] = 32'b00000000000000000011111110110101;
assign LUT_4[44713] = 32'b11111111111111111101001010101101;
assign LUT_4[44714] = 32'b00000000000000000011011001011001;
assign LUT_4[44715] = 32'b11111111111111111100100101010001;
assign LUT_4[44716] = 32'b00000000000000000000111111010001;
assign LUT_4[44717] = 32'b11111111111111111010001011001001;
assign LUT_4[44718] = 32'b00000000000000000000011001110101;
assign LUT_4[44719] = 32'b11111111111111111001100101101101;
assign LUT_4[44720] = 32'b00000000000000001000100100001110;
assign LUT_4[44721] = 32'b00000000000000000001110000000110;
assign LUT_4[44722] = 32'b00000000000000000111111110110010;
assign LUT_4[44723] = 32'b00000000000000000001001010101010;
assign LUT_4[44724] = 32'b00000000000000000101100100101010;
assign LUT_4[44725] = 32'b11111111111111111110110000100010;
assign LUT_4[44726] = 32'b00000000000000000100111111001110;
assign LUT_4[44727] = 32'b11111111111111111110001011000110;
assign LUT_4[44728] = 32'b00000000000000000001110000100011;
assign LUT_4[44729] = 32'b11111111111111111010111100011011;
assign LUT_4[44730] = 32'b00000000000000000001001011000111;
assign LUT_4[44731] = 32'b11111111111111111010010110111111;
assign LUT_4[44732] = 32'b11111111111111111110110000111111;
assign LUT_4[44733] = 32'b11111111111111110111111100110111;
assign LUT_4[44734] = 32'b11111111111111111110001011100011;
assign LUT_4[44735] = 32'b11111111111111110111010111011011;
assign LUT_4[44736] = 32'b00000000000000001101101110101101;
assign LUT_4[44737] = 32'b00000000000000000110111010100101;
assign LUT_4[44738] = 32'b00000000000000001101001001010001;
assign LUT_4[44739] = 32'b00000000000000000110010101001001;
assign LUT_4[44740] = 32'b00000000000000001010101111001001;
assign LUT_4[44741] = 32'b00000000000000000011111011000001;
assign LUT_4[44742] = 32'b00000000000000001010001001101101;
assign LUT_4[44743] = 32'b00000000000000000011010101100101;
assign LUT_4[44744] = 32'b00000000000000000110111011000010;
assign LUT_4[44745] = 32'b00000000000000000000000110111010;
assign LUT_4[44746] = 32'b00000000000000000110010101100110;
assign LUT_4[44747] = 32'b11111111111111111111100001011110;
assign LUT_4[44748] = 32'b00000000000000000011111011011110;
assign LUT_4[44749] = 32'b11111111111111111101000111010110;
assign LUT_4[44750] = 32'b00000000000000000011010110000010;
assign LUT_4[44751] = 32'b11111111111111111100100001111010;
assign LUT_4[44752] = 32'b00000000000000001011100000011011;
assign LUT_4[44753] = 32'b00000000000000000100101100010011;
assign LUT_4[44754] = 32'b00000000000000001010111010111111;
assign LUT_4[44755] = 32'b00000000000000000100000110110111;
assign LUT_4[44756] = 32'b00000000000000001000100000110111;
assign LUT_4[44757] = 32'b00000000000000000001101100101111;
assign LUT_4[44758] = 32'b00000000000000000111111011011011;
assign LUT_4[44759] = 32'b00000000000000000001000111010011;
assign LUT_4[44760] = 32'b00000000000000000100101100110000;
assign LUT_4[44761] = 32'b11111111111111111101111000101000;
assign LUT_4[44762] = 32'b00000000000000000100000111010100;
assign LUT_4[44763] = 32'b11111111111111111101010011001100;
assign LUT_4[44764] = 32'b00000000000000000001101101001100;
assign LUT_4[44765] = 32'b11111111111111111010111001000100;
assign LUT_4[44766] = 32'b00000000000000000001000111110000;
assign LUT_4[44767] = 32'b11111111111111111010010011101000;
assign LUT_4[44768] = 32'b00000000000000001100001001110100;
assign LUT_4[44769] = 32'b00000000000000000101010101101100;
assign LUT_4[44770] = 32'b00000000000000001011100100011000;
assign LUT_4[44771] = 32'b00000000000000000100110000010000;
assign LUT_4[44772] = 32'b00000000000000001001001010010000;
assign LUT_4[44773] = 32'b00000000000000000010010110001000;
assign LUT_4[44774] = 32'b00000000000000001000100100110100;
assign LUT_4[44775] = 32'b00000000000000000001110000101100;
assign LUT_4[44776] = 32'b00000000000000000101010110001001;
assign LUT_4[44777] = 32'b11111111111111111110100010000001;
assign LUT_4[44778] = 32'b00000000000000000100110000101101;
assign LUT_4[44779] = 32'b11111111111111111101111100100101;
assign LUT_4[44780] = 32'b00000000000000000010010110100101;
assign LUT_4[44781] = 32'b11111111111111111011100010011101;
assign LUT_4[44782] = 32'b00000000000000000001110001001001;
assign LUT_4[44783] = 32'b11111111111111111010111101000001;
assign LUT_4[44784] = 32'b00000000000000001001111011100010;
assign LUT_4[44785] = 32'b00000000000000000011000111011010;
assign LUT_4[44786] = 32'b00000000000000001001010110000110;
assign LUT_4[44787] = 32'b00000000000000000010100001111110;
assign LUT_4[44788] = 32'b00000000000000000110111011111110;
assign LUT_4[44789] = 32'b00000000000000000000000111110110;
assign LUT_4[44790] = 32'b00000000000000000110010110100010;
assign LUT_4[44791] = 32'b11111111111111111111100010011010;
assign LUT_4[44792] = 32'b00000000000000000011000111110111;
assign LUT_4[44793] = 32'b11111111111111111100010011101111;
assign LUT_4[44794] = 32'b00000000000000000010100010011011;
assign LUT_4[44795] = 32'b11111111111111111011101110010011;
assign LUT_4[44796] = 32'b00000000000000000000001000010011;
assign LUT_4[44797] = 32'b11111111111111111001010100001011;
assign LUT_4[44798] = 32'b11111111111111111111100010110111;
assign LUT_4[44799] = 32'b11111111111111111000101110101111;
assign LUT_4[44800] = 32'b00000000000000001110101100110100;
assign LUT_4[44801] = 32'b00000000000000000111111000101100;
assign LUT_4[44802] = 32'b00000000000000001110000111011000;
assign LUT_4[44803] = 32'b00000000000000000111010011010000;
assign LUT_4[44804] = 32'b00000000000000001011101101010000;
assign LUT_4[44805] = 32'b00000000000000000100111001001000;
assign LUT_4[44806] = 32'b00000000000000001011000111110100;
assign LUT_4[44807] = 32'b00000000000000000100010011101100;
assign LUT_4[44808] = 32'b00000000000000000111111001001001;
assign LUT_4[44809] = 32'b00000000000000000001000101000001;
assign LUT_4[44810] = 32'b00000000000000000111010011101101;
assign LUT_4[44811] = 32'b00000000000000000000011111100101;
assign LUT_4[44812] = 32'b00000000000000000100111001100101;
assign LUT_4[44813] = 32'b11111111111111111110000101011101;
assign LUT_4[44814] = 32'b00000000000000000100010100001001;
assign LUT_4[44815] = 32'b11111111111111111101100000000001;
assign LUT_4[44816] = 32'b00000000000000001100011110100010;
assign LUT_4[44817] = 32'b00000000000000000101101010011010;
assign LUT_4[44818] = 32'b00000000000000001011111001000110;
assign LUT_4[44819] = 32'b00000000000000000101000100111110;
assign LUT_4[44820] = 32'b00000000000000001001011110111110;
assign LUT_4[44821] = 32'b00000000000000000010101010110110;
assign LUT_4[44822] = 32'b00000000000000001000111001100010;
assign LUT_4[44823] = 32'b00000000000000000010000101011010;
assign LUT_4[44824] = 32'b00000000000000000101101010110111;
assign LUT_4[44825] = 32'b11111111111111111110110110101111;
assign LUT_4[44826] = 32'b00000000000000000101000101011011;
assign LUT_4[44827] = 32'b11111111111111111110010001010011;
assign LUT_4[44828] = 32'b00000000000000000010101011010011;
assign LUT_4[44829] = 32'b11111111111111111011110111001011;
assign LUT_4[44830] = 32'b00000000000000000010000101110111;
assign LUT_4[44831] = 32'b11111111111111111011010001101111;
assign LUT_4[44832] = 32'b00000000000000001101000111111011;
assign LUT_4[44833] = 32'b00000000000000000110010011110011;
assign LUT_4[44834] = 32'b00000000000000001100100010011111;
assign LUT_4[44835] = 32'b00000000000000000101101110010111;
assign LUT_4[44836] = 32'b00000000000000001010001000010111;
assign LUT_4[44837] = 32'b00000000000000000011010100001111;
assign LUT_4[44838] = 32'b00000000000000001001100010111011;
assign LUT_4[44839] = 32'b00000000000000000010101110110011;
assign LUT_4[44840] = 32'b00000000000000000110010100010000;
assign LUT_4[44841] = 32'b11111111111111111111100000001000;
assign LUT_4[44842] = 32'b00000000000000000101101110110100;
assign LUT_4[44843] = 32'b11111111111111111110111010101100;
assign LUT_4[44844] = 32'b00000000000000000011010100101100;
assign LUT_4[44845] = 32'b11111111111111111100100000100100;
assign LUT_4[44846] = 32'b00000000000000000010101111010000;
assign LUT_4[44847] = 32'b11111111111111111011111011001000;
assign LUT_4[44848] = 32'b00000000000000001010111001101001;
assign LUT_4[44849] = 32'b00000000000000000100000101100001;
assign LUT_4[44850] = 32'b00000000000000001010010100001101;
assign LUT_4[44851] = 32'b00000000000000000011100000000101;
assign LUT_4[44852] = 32'b00000000000000000111111010000101;
assign LUT_4[44853] = 32'b00000000000000000001000101111101;
assign LUT_4[44854] = 32'b00000000000000000111010100101001;
assign LUT_4[44855] = 32'b00000000000000000000100000100001;
assign LUT_4[44856] = 32'b00000000000000000100000101111110;
assign LUT_4[44857] = 32'b11111111111111111101010001110110;
assign LUT_4[44858] = 32'b00000000000000000011100000100010;
assign LUT_4[44859] = 32'b11111111111111111100101100011010;
assign LUT_4[44860] = 32'b00000000000000000001000110011010;
assign LUT_4[44861] = 32'b11111111111111111010010010010010;
assign LUT_4[44862] = 32'b00000000000000000000100000111110;
assign LUT_4[44863] = 32'b11111111111111111001101100110110;
assign LUT_4[44864] = 32'b00000000000000010000000100001000;
assign LUT_4[44865] = 32'b00000000000000001001010000000000;
assign LUT_4[44866] = 32'b00000000000000001111011110101100;
assign LUT_4[44867] = 32'b00000000000000001000101010100100;
assign LUT_4[44868] = 32'b00000000000000001101000100100100;
assign LUT_4[44869] = 32'b00000000000000000110010000011100;
assign LUT_4[44870] = 32'b00000000000000001100011111001000;
assign LUT_4[44871] = 32'b00000000000000000101101011000000;
assign LUT_4[44872] = 32'b00000000000000001001010000011101;
assign LUT_4[44873] = 32'b00000000000000000010011100010101;
assign LUT_4[44874] = 32'b00000000000000001000101011000001;
assign LUT_4[44875] = 32'b00000000000000000001110110111001;
assign LUT_4[44876] = 32'b00000000000000000110010000111001;
assign LUT_4[44877] = 32'b11111111111111111111011100110001;
assign LUT_4[44878] = 32'b00000000000000000101101011011101;
assign LUT_4[44879] = 32'b11111111111111111110110111010101;
assign LUT_4[44880] = 32'b00000000000000001101110101110110;
assign LUT_4[44881] = 32'b00000000000000000111000001101110;
assign LUT_4[44882] = 32'b00000000000000001101010000011010;
assign LUT_4[44883] = 32'b00000000000000000110011100010010;
assign LUT_4[44884] = 32'b00000000000000001010110110010010;
assign LUT_4[44885] = 32'b00000000000000000100000010001010;
assign LUT_4[44886] = 32'b00000000000000001010010000110110;
assign LUT_4[44887] = 32'b00000000000000000011011100101110;
assign LUT_4[44888] = 32'b00000000000000000111000010001011;
assign LUT_4[44889] = 32'b00000000000000000000001110000011;
assign LUT_4[44890] = 32'b00000000000000000110011100101111;
assign LUT_4[44891] = 32'b11111111111111111111101000100111;
assign LUT_4[44892] = 32'b00000000000000000100000010100111;
assign LUT_4[44893] = 32'b11111111111111111101001110011111;
assign LUT_4[44894] = 32'b00000000000000000011011101001011;
assign LUT_4[44895] = 32'b11111111111111111100101001000011;
assign LUT_4[44896] = 32'b00000000000000001110011111001111;
assign LUT_4[44897] = 32'b00000000000000000111101011000111;
assign LUT_4[44898] = 32'b00000000000000001101111001110011;
assign LUT_4[44899] = 32'b00000000000000000111000101101011;
assign LUT_4[44900] = 32'b00000000000000001011011111101011;
assign LUT_4[44901] = 32'b00000000000000000100101011100011;
assign LUT_4[44902] = 32'b00000000000000001010111010001111;
assign LUT_4[44903] = 32'b00000000000000000100000110000111;
assign LUT_4[44904] = 32'b00000000000000000111101011100100;
assign LUT_4[44905] = 32'b00000000000000000000110111011100;
assign LUT_4[44906] = 32'b00000000000000000111000110001000;
assign LUT_4[44907] = 32'b00000000000000000000010010000000;
assign LUT_4[44908] = 32'b00000000000000000100101100000000;
assign LUT_4[44909] = 32'b11111111111111111101110111111000;
assign LUT_4[44910] = 32'b00000000000000000100000110100100;
assign LUT_4[44911] = 32'b11111111111111111101010010011100;
assign LUT_4[44912] = 32'b00000000000000001100010000111101;
assign LUT_4[44913] = 32'b00000000000000000101011100110101;
assign LUT_4[44914] = 32'b00000000000000001011101011100001;
assign LUT_4[44915] = 32'b00000000000000000100110111011001;
assign LUT_4[44916] = 32'b00000000000000001001010001011001;
assign LUT_4[44917] = 32'b00000000000000000010011101010001;
assign LUT_4[44918] = 32'b00000000000000001000101011111101;
assign LUT_4[44919] = 32'b00000000000000000001110111110101;
assign LUT_4[44920] = 32'b00000000000000000101011101010010;
assign LUT_4[44921] = 32'b11111111111111111110101001001010;
assign LUT_4[44922] = 32'b00000000000000000100110111110110;
assign LUT_4[44923] = 32'b11111111111111111110000011101110;
assign LUT_4[44924] = 32'b00000000000000000010011101101110;
assign LUT_4[44925] = 32'b11111111111111111011101001100110;
assign LUT_4[44926] = 32'b00000000000000000001111000010010;
assign LUT_4[44927] = 32'b11111111111111111011000100001010;
assign LUT_4[44928] = 32'b00000000000000010001010010111100;
assign LUT_4[44929] = 32'b00000000000000001010011110110100;
assign LUT_4[44930] = 32'b00000000000000010000101101100000;
assign LUT_4[44931] = 32'b00000000000000001001111001011000;
assign LUT_4[44932] = 32'b00000000000000001110010011011000;
assign LUT_4[44933] = 32'b00000000000000000111011111010000;
assign LUT_4[44934] = 32'b00000000000000001101101101111100;
assign LUT_4[44935] = 32'b00000000000000000110111001110100;
assign LUT_4[44936] = 32'b00000000000000001010011111010001;
assign LUT_4[44937] = 32'b00000000000000000011101011001001;
assign LUT_4[44938] = 32'b00000000000000001001111001110101;
assign LUT_4[44939] = 32'b00000000000000000011000101101101;
assign LUT_4[44940] = 32'b00000000000000000111011111101101;
assign LUT_4[44941] = 32'b00000000000000000000101011100101;
assign LUT_4[44942] = 32'b00000000000000000110111010010001;
assign LUT_4[44943] = 32'b00000000000000000000000110001001;
assign LUT_4[44944] = 32'b00000000000000001111000100101010;
assign LUT_4[44945] = 32'b00000000000000001000010000100010;
assign LUT_4[44946] = 32'b00000000000000001110011111001110;
assign LUT_4[44947] = 32'b00000000000000000111101011000110;
assign LUT_4[44948] = 32'b00000000000000001100000101000110;
assign LUT_4[44949] = 32'b00000000000000000101010000111110;
assign LUT_4[44950] = 32'b00000000000000001011011111101010;
assign LUT_4[44951] = 32'b00000000000000000100101011100010;
assign LUT_4[44952] = 32'b00000000000000001000010000111111;
assign LUT_4[44953] = 32'b00000000000000000001011100110111;
assign LUT_4[44954] = 32'b00000000000000000111101011100011;
assign LUT_4[44955] = 32'b00000000000000000000110111011011;
assign LUT_4[44956] = 32'b00000000000000000101010001011011;
assign LUT_4[44957] = 32'b11111111111111111110011101010011;
assign LUT_4[44958] = 32'b00000000000000000100101011111111;
assign LUT_4[44959] = 32'b11111111111111111101110111110111;
assign LUT_4[44960] = 32'b00000000000000001111101110000011;
assign LUT_4[44961] = 32'b00000000000000001000111001111011;
assign LUT_4[44962] = 32'b00000000000000001111001000100111;
assign LUT_4[44963] = 32'b00000000000000001000010100011111;
assign LUT_4[44964] = 32'b00000000000000001100101110011111;
assign LUT_4[44965] = 32'b00000000000000000101111010010111;
assign LUT_4[44966] = 32'b00000000000000001100001001000011;
assign LUT_4[44967] = 32'b00000000000000000101010100111011;
assign LUT_4[44968] = 32'b00000000000000001000111010011000;
assign LUT_4[44969] = 32'b00000000000000000010000110010000;
assign LUT_4[44970] = 32'b00000000000000001000010100111100;
assign LUT_4[44971] = 32'b00000000000000000001100000110100;
assign LUT_4[44972] = 32'b00000000000000000101111010110100;
assign LUT_4[44973] = 32'b11111111111111111111000110101100;
assign LUT_4[44974] = 32'b00000000000000000101010101011000;
assign LUT_4[44975] = 32'b11111111111111111110100001010000;
assign LUT_4[44976] = 32'b00000000000000001101011111110001;
assign LUT_4[44977] = 32'b00000000000000000110101011101001;
assign LUT_4[44978] = 32'b00000000000000001100111010010101;
assign LUT_4[44979] = 32'b00000000000000000110000110001101;
assign LUT_4[44980] = 32'b00000000000000001010100000001101;
assign LUT_4[44981] = 32'b00000000000000000011101100000101;
assign LUT_4[44982] = 32'b00000000000000001001111010110001;
assign LUT_4[44983] = 32'b00000000000000000011000110101001;
assign LUT_4[44984] = 32'b00000000000000000110101100000110;
assign LUT_4[44985] = 32'b11111111111111111111110111111110;
assign LUT_4[44986] = 32'b00000000000000000110000110101010;
assign LUT_4[44987] = 32'b11111111111111111111010010100010;
assign LUT_4[44988] = 32'b00000000000000000011101100100010;
assign LUT_4[44989] = 32'b11111111111111111100111000011010;
assign LUT_4[44990] = 32'b00000000000000000011000111000110;
assign LUT_4[44991] = 32'b11111111111111111100010010111110;
assign LUT_4[44992] = 32'b00000000000000010010101010010000;
assign LUT_4[44993] = 32'b00000000000000001011110110001000;
assign LUT_4[44994] = 32'b00000000000000010010000100110100;
assign LUT_4[44995] = 32'b00000000000000001011010000101100;
assign LUT_4[44996] = 32'b00000000000000001111101010101100;
assign LUT_4[44997] = 32'b00000000000000001000110110100100;
assign LUT_4[44998] = 32'b00000000000000001111000101010000;
assign LUT_4[44999] = 32'b00000000000000001000010001001000;
assign LUT_4[45000] = 32'b00000000000000001011110110100101;
assign LUT_4[45001] = 32'b00000000000000000101000010011101;
assign LUT_4[45002] = 32'b00000000000000001011010001001001;
assign LUT_4[45003] = 32'b00000000000000000100011101000001;
assign LUT_4[45004] = 32'b00000000000000001000110111000001;
assign LUT_4[45005] = 32'b00000000000000000010000010111001;
assign LUT_4[45006] = 32'b00000000000000001000010001100101;
assign LUT_4[45007] = 32'b00000000000000000001011101011101;
assign LUT_4[45008] = 32'b00000000000000010000011011111110;
assign LUT_4[45009] = 32'b00000000000000001001100111110110;
assign LUT_4[45010] = 32'b00000000000000001111110110100010;
assign LUT_4[45011] = 32'b00000000000000001001000010011010;
assign LUT_4[45012] = 32'b00000000000000001101011100011010;
assign LUT_4[45013] = 32'b00000000000000000110101000010010;
assign LUT_4[45014] = 32'b00000000000000001100110110111110;
assign LUT_4[45015] = 32'b00000000000000000110000010110110;
assign LUT_4[45016] = 32'b00000000000000001001101000010011;
assign LUT_4[45017] = 32'b00000000000000000010110100001011;
assign LUT_4[45018] = 32'b00000000000000001001000010110111;
assign LUT_4[45019] = 32'b00000000000000000010001110101111;
assign LUT_4[45020] = 32'b00000000000000000110101000101111;
assign LUT_4[45021] = 32'b11111111111111111111110100100111;
assign LUT_4[45022] = 32'b00000000000000000110000011010011;
assign LUT_4[45023] = 32'b11111111111111111111001111001011;
assign LUT_4[45024] = 32'b00000000000000010001000101010111;
assign LUT_4[45025] = 32'b00000000000000001010010001001111;
assign LUT_4[45026] = 32'b00000000000000010000011111111011;
assign LUT_4[45027] = 32'b00000000000000001001101011110011;
assign LUT_4[45028] = 32'b00000000000000001110000101110011;
assign LUT_4[45029] = 32'b00000000000000000111010001101011;
assign LUT_4[45030] = 32'b00000000000000001101100000010111;
assign LUT_4[45031] = 32'b00000000000000000110101100001111;
assign LUT_4[45032] = 32'b00000000000000001010010001101100;
assign LUT_4[45033] = 32'b00000000000000000011011101100100;
assign LUT_4[45034] = 32'b00000000000000001001101100010000;
assign LUT_4[45035] = 32'b00000000000000000010111000001000;
assign LUT_4[45036] = 32'b00000000000000000111010010001000;
assign LUT_4[45037] = 32'b00000000000000000000011110000000;
assign LUT_4[45038] = 32'b00000000000000000110101100101100;
assign LUT_4[45039] = 32'b11111111111111111111111000100100;
assign LUT_4[45040] = 32'b00000000000000001110110111000101;
assign LUT_4[45041] = 32'b00000000000000001000000010111101;
assign LUT_4[45042] = 32'b00000000000000001110010001101001;
assign LUT_4[45043] = 32'b00000000000000000111011101100001;
assign LUT_4[45044] = 32'b00000000000000001011110111100001;
assign LUT_4[45045] = 32'b00000000000000000101000011011001;
assign LUT_4[45046] = 32'b00000000000000001011010010000101;
assign LUT_4[45047] = 32'b00000000000000000100011101111101;
assign LUT_4[45048] = 32'b00000000000000001000000011011010;
assign LUT_4[45049] = 32'b00000000000000000001001111010010;
assign LUT_4[45050] = 32'b00000000000000000111011101111110;
assign LUT_4[45051] = 32'b00000000000000000000101001110110;
assign LUT_4[45052] = 32'b00000000000000000101000011110110;
assign LUT_4[45053] = 32'b11111111111111111110001111101110;
assign LUT_4[45054] = 32'b00000000000000000100011110011010;
assign LUT_4[45055] = 32'b11111111111111111101101010010010;
assign LUT_4[45056] = 32'b00000000000000001001110011010001;
assign LUT_4[45057] = 32'b00000000000000000010111111001001;
assign LUT_4[45058] = 32'b00000000000000001001001101110101;
assign LUT_4[45059] = 32'b00000000000000000010011001101101;
assign LUT_4[45060] = 32'b00000000000000000110110011101101;
assign LUT_4[45061] = 32'b11111111111111111111111111100101;
assign LUT_4[45062] = 32'b00000000000000000110001110010001;
assign LUT_4[45063] = 32'b11111111111111111111011010001001;
assign LUT_4[45064] = 32'b00000000000000000010111111100110;
assign LUT_4[45065] = 32'b11111111111111111100001011011110;
assign LUT_4[45066] = 32'b00000000000000000010011010001010;
assign LUT_4[45067] = 32'b11111111111111111011100110000010;
assign LUT_4[45068] = 32'b00000000000000000000000000000010;
assign LUT_4[45069] = 32'b11111111111111111001001011111010;
assign LUT_4[45070] = 32'b11111111111111111111011010100110;
assign LUT_4[45071] = 32'b11111111111111111000100110011110;
assign LUT_4[45072] = 32'b00000000000000000111100100111111;
assign LUT_4[45073] = 32'b00000000000000000000110000110111;
assign LUT_4[45074] = 32'b00000000000000000110111111100011;
assign LUT_4[45075] = 32'b00000000000000000000001011011011;
assign LUT_4[45076] = 32'b00000000000000000100100101011011;
assign LUT_4[45077] = 32'b11111111111111111101110001010011;
assign LUT_4[45078] = 32'b00000000000000000011111111111111;
assign LUT_4[45079] = 32'b11111111111111111101001011110111;
assign LUT_4[45080] = 32'b00000000000000000000110001010100;
assign LUT_4[45081] = 32'b11111111111111111001111101001100;
assign LUT_4[45082] = 32'b00000000000000000000001011111000;
assign LUT_4[45083] = 32'b11111111111111111001010111110000;
assign LUT_4[45084] = 32'b11111111111111111101110001110000;
assign LUT_4[45085] = 32'b11111111111111110110111101101000;
assign LUT_4[45086] = 32'b11111111111111111101001100010100;
assign LUT_4[45087] = 32'b11111111111111110110011000001100;
assign LUT_4[45088] = 32'b00000000000000001000001110011000;
assign LUT_4[45089] = 32'b00000000000000000001011010010000;
assign LUT_4[45090] = 32'b00000000000000000111101000111100;
assign LUT_4[45091] = 32'b00000000000000000000110100110100;
assign LUT_4[45092] = 32'b00000000000000000101001110110100;
assign LUT_4[45093] = 32'b11111111111111111110011010101100;
assign LUT_4[45094] = 32'b00000000000000000100101001011000;
assign LUT_4[45095] = 32'b11111111111111111101110101010000;
assign LUT_4[45096] = 32'b00000000000000000001011010101101;
assign LUT_4[45097] = 32'b11111111111111111010100110100101;
assign LUT_4[45098] = 32'b00000000000000000000110101010001;
assign LUT_4[45099] = 32'b11111111111111111010000001001001;
assign LUT_4[45100] = 32'b11111111111111111110011011001001;
assign LUT_4[45101] = 32'b11111111111111110111100111000001;
assign LUT_4[45102] = 32'b11111111111111111101110101101101;
assign LUT_4[45103] = 32'b11111111111111110111000001100101;
assign LUT_4[45104] = 32'b00000000000000000110000000000110;
assign LUT_4[45105] = 32'b11111111111111111111001011111110;
assign LUT_4[45106] = 32'b00000000000000000101011010101010;
assign LUT_4[45107] = 32'b11111111111111111110100110100010;
assign LUT_4[45108] = 32'b00000000000000000011000000100010;
assign LUT_4[45109] = 32'b11111111111111111100001100011010;
assign LUT_4[45110] = 32'b00000000000000000010011011000110;
assign LUT_4[45111] = 32'b11111111111111111011100110111110;
assign LUT_4[45112] = 32'b11111111111111111111001100011011;
assign LUT_4[45113] = 32'b11111111111111111000011000010011;
assign LUT_4[45114] = 32'b11111111111111111110100110111111;
assign LUT_4[45115] = 32'b11111111111111110111110010110111;
assign LUT_4[45116] = 32'b11111111111111111100001100110111;
assign LUT_4[45117] = 32'b11111111111111110101011000101111;
assign LUT_4[45118] = 32'b11111111111111111011100111011011;
assign LUT_4[45119] = 32'b11111111111111110100110011010011;
assign LUT_4[45120] = 32'b00000000000000001011001010100101;
assign LUT_4[45121] = 32'b00000000000000000100010110011101;
assign LUT_4[45122] = 32'b00000000000000001010100101001001;
assign LUT_4[45123] = 32'b00000000000000000011110001000001;
assign LUT_4[45124] = 32'b00000000000000001000001011000001;
assign LUT_4[45125] = 32'b00000000000000000001010110111001;
assign LUT_4[45126] = 32'b00000000000000000111100101100101;
assign LUT_4[45127] = 32'b00000000000000000000110001011101;
assign LUT_4[45128] = 32'b00000000000000000100010110111010;
assign LUT_4[45129] = 32'b11111111111111111101100010110010;
assign LUT_4[45130] = 32'b00000000000000000011110001011110;
assign LUT_4[45131] = 32'b11111111111111111100111101010110;
assign LUT_4[45132] = 32'b00000000000000000001010111010110;
assign LUT_4[45133] = 32'b11111111111111111010100011001110;
assign LUT_4[45134] = 32'b00000000000000000000110001111010;
assign LUT_4[45135] = 32'b11111111111111111001111101110010;
assign LUT_4[45136] = 32'b00000000000000001000111100010011;
assign LUT_4[45137] = 32'b00000000000000000010001000001011;
assign LUT_4[45138] = 32'b00000000000000001000010110110111;
assign LUT_4[45139] = 32'b00000000000000000001100010101111;
assign LUT_4[45140] = 32'b00000000000000000101111100101111;
assign LUT_4[45141] = 32'b11111111111111111111001000100111;
assign LUT_4[45142] = 32'b00000000000000000101010111010011;
assign LUT_4[45143] = 32'b11111111111111111110100011001011;
assign LUT_4[45144] = 32'b00000000000000000010001000101000;
assign LUT_4[45145] = 32'b11111111111111111011010100100000;
assign LUT_4[45146] = 32'b00000000000000000001100011001100;
assign LUT_4[45147] = 32'b11111111111111111010101111000100;
assign LUT_4[45148] = 32'b11111111111111111111001001000100;
assign LUT_4[45149] = 32'b11111111111111111000010100111100;
assign LUT_4[45150] = 32'b11111111111111111110100011101000;
assign LUT_4[45151] = 32'b11111111111111110111101111100000;
assign LUT_4[45152] = 32'b00000000000000001001100101101100;
assign LUT_4[45153] = 32'b00000000000000000010110001100100;
assign LUT_4[45154] = 32'b00000000000000001001000000010000;
assign LUT_4[45155] = 32'b00000000000000000010001100001000;
assign LUT_4[45156] = 32'b00000000000000000110100110001000;
assign LUT_4[45157] = 32'b11111111111111111111110010000000;
assign LUT_4[45158] = 32'b00000000000000000110000000101100;
assign LUT_4[45159] = 32'b11111111111111111111001100100100;
assign LUT_4[45160] = 32'b00000000000000000010110010000001;
assign LUT_4[45161] = 32'b11111111111111111011111101111001;
assign LUT_4[45162] = 32'b00000000000000000010001100100101;
assign LUT_4[45163] = 32'b11111111111111111011011000011101;
assign LUT_4[45164] = 32'b11111111111111111111110010011101;
assign LUT_4[45165] = 32'b11111111111111111000111110010101;
assign LUT_4[45166] = 32'b11111111111111111111001101000001;
assign LUT_4[45167] = 32'b11111111111111111000011000111001;
assign LUT_4[45168] = 32'b00000000000000000111010111011010;
assign LUT_4[45169] = 32'b00000000000000000000100011010010;
assign LUT_4[45170] = 32'b00000000000000000110110001111110;
assign LUT_4[45171] = 32'b11111111111111111111111101110110;
assign LUT_4[45172] = 32'b00000000000000000100010111110110;
assign LUT_4[45173] = 32'b11111111111111111101100011101110;
assign LUT_4[45174] = 32'b00000000000000000011110010011010;
assign LUT_4[45175] = 32'b11111111111111111100111110010010;
assign LUT_4[45176] = 32'b00000000000000000000100011101111;
assign LUT_4[45177] = 32'b11111111111111111001101111100111;
assign LUT_4[45178] = 32'b11111111111111111111111110010011;
assign LUT_4[45179] = 32'b11111111111111111001001010001011;
assign LUT_4[45180] = 32'b11111111111111111101100100001011;
assign LUT_4[45181] = 32'b11111111111111110110110000000011;
assign LUT_4[45182] = 32'b11111111111111111100111110101111;
assign LUT_4[45183] = 32'b11111111111111110110001010100111;
assign LUT_4[45184] = 32'b00000000000000001100011001011001;
assign LUT_4[45185] = 32'b00000000000000000101100101010001;
assign LUT_4[45186] = 32'b00000000000000001011110011111101;
assign LUT_4[45187] = 32'b00000000000000000100111111110101;
assign LUT_4[45188] = 32'b00000000000000001001011001110101;
assign LUT_4[45189] = 32'b00000000000000000010100101101101;
assign LUT_4[45190] = 32'b00000000000000001000110100011001;
assign LUT_4[45191] = 32'b00000000000000000010000000010001;
assign LUT_4[45192] = 32'b00000000000000000101100101101110;
assign LUT_4[45193] = 32'b11111111111111111110110001100110;
assign LUT_4[45194] = 32'b00000000000000000101000000010010;
assign LUT_4[45195] = 32'b11111111111111111110001100001010;
assign LUT_4[45196] = 32'b00000000000000000010100110001010;
assign LUT_4[45197] = 32'b11111111111111111011110010000010;
assign LUT_4[45198] = 32'b00000000000000000010000000101110;
assign LUT_4[45199] = 32'b11111111111111111011001100100110;
assign LUT_4[45200] = 32'b00000000000000001010001011000111;
assign LUT_4[45201] = 32'b00000000000000000011010110111111;
assign LUT_4[45202] = 32'b00000000000000001001100101101011;
assign LUT_4[45203] = 32'b00000000000000000010110001100011;
assign LUT_4[45204] = 32'b00000000000000000111001011100011;
assign LUT_4[45205] = 32'b00000000000000000000010111011011;
assign LUT_4[45206] = 32'b00000000000000000110100110000111;
assign LUT_4[45207] = 32'b11111111111111111111110001111111;
assign LUT_4[45208] = 32'b00000000000000000011010111011100;
assign LUT_4[45209] = 32'b11111111111111111100100011010100;
assign LUT_4[45210] = 32'b00000000000000000010110010000000;
assign LUT_4[45211] = 32'b11111111111111111011111101111000;
assign LUT_4[45212] = 32'b00000000000000000000010111111000;
assign LUT_4[45213] = 32'b11111111111111111001100011110000;
assign LUT_4[45214] = 32'b11111111111111111111110010011100;
assign LUT_4[45215] = 32'b11111111111111111000111110010100;
assign LUT_4[45216] = 32'b00000000000000001010110100100000;
assign LUT_4[45217] = 32'b00000000000000000100000000011000;
assign LUT_4[45218] = 32'b00000000000000001010001111000100;
assign LUT_4[45219] = 32'b00000000000000000011011010111100;
assign LUT_4[45220] = 32'b00000000000000000111110100111100;
assign LUT_4[45221] = 32'b00000000000000000001000000110100;
assign LUT_4[45222] = 32'b00000000000000000111001111100000;
assign LUT_4[45223] = 32'b00000000000000000000011011011000;
assign LUT_4[45224] = 32'b00000000000000000100000000110101;
assign LUT_4[45225] = 32'b11111111111111111101001100101101;
assign LUT_4[45226] = 32'b00000000000000000011011011011001;
assign LUT_4[45227] = 32'b11111111111111111100100111010001;
assign LUT_4[45228] = 32'b00000000000000000001000001010001;
assign LUT_4[45229] = 32'b11111111111111111010001101001001;
assign LUT_4[45230] = 32'b00000000000000000000011011110101;
assign LUT_4[45231] = 32'b11111111111111111001100111101101;
assign LUT_4[45232] = 32'b00000000000000001000100110001110;
assign LUT_4[45233] = 32'b00000000000000000001110010000110;
assign LUT_4[45234] = 32'b00000000000000001000000000110010;
assign LUT_4[45235] = 32'b00000000000000000001001100101010;
assign LUT_4[45236] = 32'b00000000000000000101100110101010;
assign LUT_4[45237] = 32'b11111111111111111110110010100010;
assign LUT_4[45238] = 32'b00000000000000000101000001001110;
assign LUT_4[45239] = 32'b11111111111111111110001101000110;
assign LUT_4[45240] = 32'b00000000000000000001110010100011;
assign LUT_4[45241] = 32'b11111111111111111010111110011011;
assign LUT_4[45242] = 32'b00000000000000000001001101000111;
assign LUT_4[45243] = 32'b11111111111111111010011000111111;
assign LUT_4[45244] = 32'b11111111111111111110110010111111;
assign LUT_4[45245] = 32'b11111111111111110111111110110111;
assign LUT_4[45246] = 32'b11111111111111111110001101100011;
assign LUT_4[45247] = 32'b11111111111111110111011001011011;
assign LUT_4[45248] = 32'b00000000000000001101110000101101;
assign LUT_4[45249] = 32'b00000000000000000110111100100101;
assign LUT_4[45250] = 32'b00000000000000001101001011010001;
assign LUT_4[45251] = 32'b00000000000000000110010111001001;
assign LUT_4[45252] = 32'b00000000000000001010110001001001;
assign LUT_4[45253] = 32'b00000000000000000011111101000001;
assign LUT_4[45254] = 32'b00000000000000001010001011101101;
assign LUT_4[45255] = 32'b00000000000000000011010111100101;
assign LUT_4[45256] = 32'b00000000000000000110111101000010;
assign LUT_4[45257] = 32'b00000000000000000000001000111010;
assign LUT_4[45258] = 32'b00000000000000000110010111100110;
assign LUT_4[45259] = 32'b11111111111111111111100011011110;
assign LUT_4[45260] = 32'b00000000000000000011111101011110;
assign LUT_4[45261] = 32'b11111111111111111101001001010110;
assign LUT_4[45262] = 32'b00000000000000000011011000000010;
assign LUT_4[45263] = 32'b11111111111111111100100011111010;
assign LUT_4[45264] = 32'b00000000000000001011100010011011;
assign LUT_4[45265] = 32'b00000000000000000100101110010011;
assign LUT_4[45266] = 32'b00000000000000001010111100111111;
assign LUT_4[45267] = 32'b00000000000000000100001000110111;
assign LUT_4[45268] = 32'b00000000000000001000100010110111;
assign LUT_4[45269] = 32'b00000000000000000001101110101111;
assign LUT_4[45270] = 32'b00000000000000000111111101011011;
assign LUT_4[45271] = 32'b00000000000000000001001001010011;
assign LUT_4[45272] = 32'b00000000000000000100101110110000;
assign LUT_4[45273] = 32'b11111111111111111101111010101000;
assign LUT_4[45274] = 32'b00000000000000000100001001010100;
assign LUT_4[45275] = 32'b11111111111111111101010101001100;
assign LUT_4[45276] = 32'b00000000000000000001101111001100;
assign LUT_4[45277] = 32'b11111111111111111010111011000100;
assign LUT_4[45278] = 32'b00000000000000000001001001110000;
assign LUT_4[45279] = 32'b11111111111111111010010101101000;
assign LUT_4[45280] = 32'b00000000000000001100001011110100;
assign LUT_4[45281] = 32'b00000000000000000101010111101100;
assign LUT_4[45282] = 32'b00000000000000001011100110011000;
assign LUT_4[45283] = 32'b00000000000000000100110010010000;
assign LUT_4[45284] = 32'b00000000000000001001001100010000;
assign LUT_4[45285] = 32'b00000000000000000010011000001000;
assign LUT_4[45286] = 32'b00000000000000001000100110110100;
assign LUT_4[45287] = 32'b00000000000000000001110010101100;
assign LUT_4[45288] = 32'b00000000000000000101011000001001;
assign LUT_4[45289] = 32'b11111111111111111110100100000001;
assign LUT_4[45290] = 32'b00000000000000000100110010101101;
assign LUT_4[45291] = 32'b11111111111111111101111110100101;
assign LUT_4[45292] = 32'b00000000000000000010011000100101;
assign LUT_4[45293] = 32'b11111111111111111011100100011101;
assign LUT_4[45294] = 32'b00000000000000000001110011001001;
assign LUT_4[45295] = 32'b11111111111111111010111111000001;
assign LUT_4[45296] = 32'b00000000000000001001111101100010;
assign LUT_4[45297] = 32'b00000000000000000011001001011010;
assign LUT_4[45298] = 32'b00000000000000001001011000000110;
assign LUT_4[45299] = 32'b00000000000000000010100011111110;
assign LUT_4[45300] = 32'b00000000000000000110111101111110;
assign LUT_4[45301] = 32'b00000000000000000000001001110110;
assign LUT_4[45302] = 32'b00000000000000000110011000100010;
assign LUT_4[45303] = 32'b11111111111111111111100100011010;
assign LUT_4[45304] = 32'b00000000000000000011001001110111;
assign LUT_4[45305] = 32'b11111111111111111100010101101111;
assign LUT_4[45306] = 32'b00000000000000000010100100011011;
assign LUT_4[45307] = 32'b11111111111111111011110000010011;
assign LUT_4[45308] = 32'b00000000000000000000001010010011;
assign LUT_4[45309] = 32'b11111111111111111001010110001011;
assign LUT_4[45310] = 32'b11111111111111111111100100110111;
assign LUT_4[45311] = 32'b11111111111111111000110000101111;
assign LUT_4[45312] = 32'b00000000000000001110101110110100;
assign LUT_4[45313] = 32'b00000000000000000111111010101100;
assign LUT_4[45314] = 32'b00000000000000001110001001011000;
assign LUT_4[45315] = 32'b00000000000000000111010101010000;
assign LUT_4[45316] = 32'b00000000000000001011101111010000;
assign LUT_4[45317] = 32'b00000000000000000100111011001000;
assign LUT_4[45318] = 32'b00000000000000001011001001110100;
assign LUT_4[45319] = 32'b00000000000000000100010101101100;
assign LUT_4[45320] = 32'b00000000000000000111111011001001;
assign LUT_4[45321] = 32'b00000000000000000001000111000001;
assign LUT_4[45322] = 32'b00000000000000000111010101101101;
assign LUT_4[45323] = 32'b00000000000000000000100001100101;
assign LUT_4[45324] = 32'b00000000000000000100111011100101;
assign LUT_4[45325] = 32'b11111111111111111110000111011101;
assign LUT_4[45326] = 32'b00000000000000000100010110001001;
assign LUT_4[45327] = 32'b11111111111111111101100010000001;
assign LUT_4[45328] = 32'b00000000000000001100100000100010;
assign LUT_4[45329] = 32'b00000000000000000101101100011010;
assign LUT_4[45330] = 32'b00000000000000001011111011000110;
assign LUT_4[45331] = 32'b00000000000000000101000110111110;
assign LUT_4[45332] = 32'b00000000000000001001100000111110;
assign LUT_4[45333] = 32'b00000000000000000010101100110110;
assign LUT_4[45334] = 32'b00000000000000001000111011100010;
assign LUT_4[45335] = 32'b00000000000000000010000111011010;
assign LUT_4[45336] = 32'b00000000000000000101101100110111;
assign LUT_4[45337] = 32'b11111111111111111110111000101111;
assign LUT_4[45338] = 32'b00000000000000000101000111011011;
assign LUT_4[45339] = 32'b11111111111111111110010011010011;
assign LUT_4[45340] = 32'b00000000000000000010101101010011;
assign LUT_4[45341] = 32'b11111111111111111011111001001011;
assign LUT_4[45342] = 32'b00000000000000000010000111110111;
assign LUT_4[45343] = 32'b11111111111111111011010011101111;
assign LUT_4[45344] = 32'b00000000000000001101001001111011;
assign LUT_4[45345] = 32'b00000000000000000110010101110011;
assign LUT_4[45346] = 32'b00000000000000001100100100011111;
assign LUT_4[45347] = 32'b00000000000000000101110000010111;
assign LUT_4[45348] = 32'b00000000000000001010001010010111;
assign LUT_4[45349] = 32'b00000000000000000011010110001111;
assign LUT_4[45350] = 32'b00000000000000001001100100111011;
assign LUT_4[45351] = 32'b00000000000000000010110000110011;
assign LUT_4[45352] = 32'b00000000000000000110010110010000;
assign LUT_4[45353] = 32'b11111111111111111111100010001000;
assign LUT_4[45354] = 32'b00000000000000000101110000110100;
assign LUT_4[45355] = 32'b11111111111111111110111100101100;
assign LUT_4[45356] = 32'b00000000000000000011010110101100;
assign LUT_4[45357] = 32'b11111111111111111100100010100100;
assign LUT_4[45358] = 32'b00000000000000000010110001010000;
assign LUT_4[45359] = 32'b11111111111111111011111101001000;
assign LUT_4[45360] = 32'b00000000000000001010111011101001;
assign LUT_4[45361] = 32'b00000000000000000100000111100001;
assign LUT_4[45362] = 32'b00000000000000001010010110001101;
assign LUT_4[45363] = 32'b00000000000000000011100010000101;
assign LUT_4[45364] = 32'b00000000000000000111111100000101;
assign LUT_4[45365] = 32'b00000000000000000001000111111101;
assign LUT_4[45366] = 32'b00000000000000000111010110101001;
assign LUT_4[45367] = 32'b00000000000000000000100010100001;
assign LUT_4[45368] = 32'b00000000000000000100000111111110;
assign LUT_4[45369] = 32'b11111111111111111101010011110110;
assign LUT_4[45370] = 32'b00000000000000000011100010100010;
assign LUT_4[45371] = 32'b11111111111111111100101110011010;
assign LUT_4[45372] = 32'b00000000000000000001001000011010;
assign LUT_4[45373] = 32'b11111111111111111010010100010010;
assign LUT_4[45374] = 32'b00000000000000000000100010111110;
assign LUT_4[45375] = 32'b11111111111111111001101110110110;
assign LUT_4[45376] = 32'b00000000000000010000000110001000;
assign LUT_4[45377] = 32'b00000000000000001001010010000000;
assign LUT_4[45378] = 32'b00000000000000001111100000101100;
assign LUT_4[45379] = 32'b00000000000000001000101100100100;
assign LUT_4[45380] = 32'b00000000000000001101000110100100;
assign LUT_4[45381] = 32'b00000000000000000110010010011100;
assign LUT_4[45382] = 32'b00000000000000001100100001001000;
assign LUT_4[45383] = 32'b00000000000000000101101101000000;
assign LUT_4[45384] = 32'b00000000000000001001010010011101;
assign LUT_4[45385] = 32'b00000000000000000010011110010101;
assign LUT_4[45386] = 32'b00000000000000001000101101000001;
assign LUT_4[45387] = 32'b00000000000000000001111000111001;
assign LUT_4[45388] = 32'b00000000000000000110010010111001;
assign LUT_4[45389] = 32'b11111111111111111111011110110001;
assign LUT_4[45390] = 32'b00000000000000000101101101011101;
assign LUT_4[45391] = 32'b11111111111111111110111001010101;
assign LUT_4[45392] = 32'b00000000000000001101110111110110;
assign LUT_4[45393] = 32'b00000000000000000111000011101110;
assign LUT_4[45394] = 32'b00000000000000001101010010011010;
assign LUT_4[45395] = 32'b00000000000000000110011110010010;
assign LUT_4[45396] = 32'b00000000000000001010111000010010;
assign LUT_4[45397] = 32'b00000000000000000100000100001010;
assign LUT_4[45398] = 32'b00000000000000001010010010110110;
assign LUT_4[45399] = 32'b00000000000000000011011110101110;
assign LUT_4[45400] = 32'b00000000000000000111000100001011;
assign LUT_4[45401] = 32'b00000000000000000000010000000011;
assign LUT_4[45402] = 32'b00000000000000000110011110101111;
assign LUT_4[45403] = 32'b11111111111111111111101010100111;
assign LUT_4[45404] = 32'b00000000000000000100000100100111;
assign LUT_4[45405] = 32'b11111111111111111101010000011111;
assign LUT_4[45406] = 32'b00000000000000000011011111001011;
assign LUT_4[45407] = 32'b11111111111111111100101011000011;
assign LUT_4[45408] = 32'b00000000000000001110100001001111;
assign LUT_4[45409] = 32'b00000000000000000111101101000111;
assign LUT_4[45410] = 32'b00000000000000001101111011110011;
assign LUT_4[45411] = 32'b00000000000000000111000111101011;
assign LUT_4[45412] = 32'b00000000000000001011100001101011;
assign LUT_4[45413] = 32'b00000000000000000100101101100011;
assign LUT_4[45414] = 32'b00000000000000001010111100001111;
assign LUT_4[45415] = 32'b00000000000000000100001000000111;
assign LUT_4[45416] = 32'b00000000000000000111101101100100;
assign LUT_4[45417] = 32'b00000000000000000000111001011100;
assign LUT_4[45418] = 32'b00000000000000000111001000001000;
assign LUT_4[45419] = 32'b00000000000000000000010100000000;
assign LUT_4[45420] = 32'b00000000000000000100101110000000;
assign LUT_4[45421] = 32'b11111111111111111101111001111000;
assign LUT_4[45422] = 32'b00000000000000000100001000100100;
assign LUT_4[45423] = 32'b11111111111111111101010100011100;
assign LUT_4[45424] = 32'b00000000000000001100010010111101;
assign LUT_4[45425] = 32'b00000000000000000101011110110101;
assign LUT_4[45426] = 32'b00000000000000001011101101100001;
assign LUT_4[45427] = 32'b00000000000000000100111001011001;
assign LUT_4[45428] = 32'b00000000000000001001010011011001;
assign LUT_4[45429] = 32'b00000000000000000010011111010001;
assign LUT_4[45430] = 32'b00000000000000001000101101111101;
assign LUT_4[45431] = 32'b00000000000000000001111001110101;
assign LUT_4[45432] = 32'b00000000000000000101011111010010;
assign LUT_4[45433] = 32'b11111111111111111110101011001010;
assign LUT_4[45434] = 32'b00000000000000000100111001110110;
assign LUT_4[45435] = 32'b11111111111111111110000101101110;
assign LUT_4[45436] = 32'b00000000000000000010011111101110;
assign LUT_4[45437] = 32'b11111111111111111011101011100110;
assign LUT_4[45438] = 32'b00000000000000000001111010010010;
assign LUT_4[45439] = 32'b11111111111111111011000110001010;
assign LUT_4[45440] = 32'b00000000000000010001010100111100;
assign LUT_4[45441] = 32'b00000000000000001010100000110100;
assign LUT_4[45442] = 32'b00000000000000010000101111100000;
assign LUT_4[45443] = 32'b00000000000000001001111011011000;
assign LUT_4[45444] = 32'b00000000000000001110010101011000;
assign LUT_4[45445] = 32'b00000000000000000111100001010000;
assign LUT_4[45446] = 32'b00000000000000001101101111111100;
assign LUT_4[45447] = 32'b00000000000000000110111011110100;
assign LUT_4[45448] = 32'b00000000000000001010100001010001;
assign LUT_4[45449] = 32'b00000000000000000011101101001001;
assign LUT_4[45450] = 32'b00000000000000001001111011110101;
assign LUT_4[45451] = 32'b00000000000000000011000111101101;
assign LUT_4[45452] = 32'b00000000000000000111100001101101;
assign LUT_4[45453] = 32'b00000000000000000000101101100101;
assign LUT_4[45454] = 32'b00000000000000000110111100010001;
assign LUT_4[45455] = 32'b00000000000000000000001000001001;
assign LUT_4[45456] = 32'b00000000000000001111000110101010;
assign LUT_4[45457] = 32'b00000000000000001000010010100010;
assign LUT_4[45458] = 32'b00000000000000001110100001001110;
assign LUT_4[45459] = 32'b00000000000000000111101101000110;
assign LUT_4[45460] = 32'b00000000000000001100000111000110;
assign LUT_4[45461] = 32'b00000000000000000101010010111110;
assign LUT_4[45462] = 32'b00000000000000001011100001101010;
assign LUT_4[45463] = 32'b00000000000000000100101101100010;
assign LUT_4[45464] = 32'b00000000000000001000010010111111;
assign LUT_4[45465] = 32'b00000000000000000001011110110111;
assign LUT_4[45466] = 32'b00000000000000000111101101100011;
assign LUT_4[45467] = 32'b00000000000000000000111001011011;
assign LUT_4[45468] = 32'b00000000000000000101010011011011;
assign LUT_4[45469] = 32'b11111111111111111110011111010011;
assign LUT_4[45470] = 32'b00000000000000000100101101111111;
assign LUT_4[45471] = 32'b11111111111111111101111001110111;
assign LUT_4[45472] = 32'b00000000000000001111110000000011;
assign LUT_4[45473] = 32'b00000000000000001000111011111011;
assign LUT_4[45474] = 32'b00000000000000001111001010100111;
assign LUT_4[45475] = 32'b00000000000000001000010110011111;
assign LUT_4[45476] = 32'b00000000000000001100110000011111;
assign LUT_4[45477] = 32'b00000000000000000101111100010111;
assign LUT_4[45478] = 32'b00000000000000001100001011000011;
assign LUT_4[45479] = 32'b00000000000000000101010110111011;
assign LUT_4[45480] = 32'b00000000000000001000111100011000;
assign LUT_4[45481] = 32'b00000000000000000010001000010000;
assign LUT_4[45482] = 32'b00000000000000001000010110111100;
assign LUT_4[45483] = 32'b00000000000000000001100010110100;
assign LUT_4[45484] = 32'b00000000000000000101111100110100;
assign LUT_4[45485] = 32'b11111111111111111111001000101100;
assign LUT_4[45486] = 32'b00000000000000000101010111011000;
assign LUT_4[45487] = 32'b11111111111111111110100011010000;
assign LUT_4[45488] = 32'b00000000000000001101100001110001;
assign LUT_4[45489] = 32'b00000000000000000110101101101001;
assign LUT_4[45490] = 32'b00000000000000001100111100010101;
assign LUT_4[45491] = 32'b00000000000000000110001000001101;
assign LUT_4[45492] = 32'b00000000000000001010100010001101;
assign LUT_4[45493] = 32'b00000000000000000011101110000101;
assign LUT_4[45494] = 32'b00000000000000001001111100110001;
assign LUT_4[45495] = 32'b00000000000000000011001000101001;
assign LUT_4[45496] = 32'b00000000000000000110101110000110;
assign LUT_4[45497] = 32'b11111111111111111111111001111110;
assign LUT_4[45498] = 32'b00000000000000000110001000101010;
assign LUT_4[45499] = 32'b11111111111111111111010100100010;
assign LUT_4[45500] = 32'b00000000000000000011101110100010;
assign LUT_4[45501] = 32'b11111111111111111100111010011010;
assign LUT_4[45502] = 32'b00000000000000000011001001000110;
assign LUT_4[45503] = 32'b11111111111111111100010100111110;
assign LUT_4[45504] = 32'b00000000000000010010101100010000;
assign LUT_4[45505] = 32'b00000000000000001011111000001000;
assign LUT_4[45506] = 32'b00000000000000010010000110110100;
assign LUT_4[45507] = 32'b00000000000000001011010010101100;
assign LUT_4[45508] = 32'b00000000000000001111101100101100;
assign LUT_4[45509] = 32'b00000000000000001000111000100100;
assign LUT_4[45510] = 32'b00000000000000001111000111010000;
assign LUT_4[45511] = 32'b00000000000000001000010011001000;
assign LUT_4[45512] = 32'b00000000000000001011111000100101;
assign LUT_4[45513] = 32'b00000000000000000101000100011101;
assign LUT_4[45514] = 32'b00000000000000001011010011001001;
assign LUT_4[45515] = 32'b00000000000000000100011111000001;
assign LUT_4[45516] = 32'b00000000000000001000111001000001;
assign LUT_4[45517] = 32'b00000000000000000010000100111001;
assign LUT_4[45518] = 32'b00000000000000001000010011100101;
assign LUT_4[45519] = 32'b00000000000000000001011111011101;
assign LUT_4[45520] = 32'b00000000000000010000011101111110;
assign LUT_4[45521] = 32'b00000000000000001001101001110110;
assign LUT_4[45522] = 32'b00000000000000001111111000100010;
assign LUT_4[45523] = 32'b00000000000000001001000100011010;
assign LUT_4[45524] = 32'b00000000000000001101011110011010;
assign LUT_4[45525] = 32'b00000000000000000110101010010010;
assign LUT_4[45526] = 32'b00000000000000001100111000111110;
assign LUT_4[45527] = 32'b00000000000000000110000100110110;
assign LUT_4[45528] = 32'b00000000000000001001101010010011;
assign LUT_4[45529] = 32'b00000000000000000010110110001011;
assign LUT_4[45530] = 32'b00000000000000001001000100110111;
assign LUT_4[45531] = 32'b00000000000000000010010000101111;
assign LUT_4[45532] = 32'b00000000000000000110101010101111;
assign LUT_4[45533] = 32'b11111111111111111111110110100111;
assign LUT_4[45534] = 32'b00000000000000000110000101010011;
assign LUT_4[45535] = 32'b11111111111111111111010001001011;
assign LUT_4[45536] = 32'b00000000000000010001000111010111;
assign LUT_4[45537] = 32'b00000000000000001010010011001111;
assign LUT_4[45538] = 32'b00000000000000010000100001111011;
assign LUT_4[45539] = 32'b00000000000000001001101101110011;
assign LUT_4[45540] = 32'b00000000000000001110000111110011;
assign LUT_4[45541] = 32'b00000000000000000111010011101011;
assign LUT_4[45542] = 32'b00000000000000001101100010010111;
assign LUT_4[45543] = 32'b00000000000000000110101110001111;
assign LUT_4[45544] = 32'b00000000000000001010010011101100;
assign LUT_4[45545] = 32'b00000000000000000011011111100100;
assign LUT_4[45546] = 32'b00000000000000001001101110010000;
assign LUT_4[45547] = 32'b00000000000000000010111010001000;
assign LUT_4[45548] = 32'b00000000000000000111010100001000;
assign LUT_4[45549] = 32'b00000000000000000000100000000000;
assign LUT_4[45550] = 32'b00000000000000000110101110101100;
assign LUT_4[45551] = 32'b11111111111111111111111010100100;
assign LUT_4[45552] = 32'b00000000000000001110111001000101;
assign LUT_4[45553] = 32'b00000000000000001000000100111101;
assign LUT_4[45554] = 32'b00000000000000001110010011101001;
assign LUT_4[45555] = 32'b00000000000000000111011111100001;
assign LUT_4[45556] = 32'b00000000000000001011111001100001;
assign LUT_4[45557] = 32'b00000000000000000101000101011001;
assign LUT_4[45558] = 32'b00000000000000001011010100000101;
assign LUT_4[45559] = 32'b00000000000000000100011111111101;
assign LUT_4[45560] = 32'b00000000000000001000000101011010;
assign LUT_4[45561] = 32'b00000000000000000001010001010010;
assign LUT_4[45562] = 32'b00000000000000000111011111111110;
assign LUT_4[45563] = 32'b00000000000000000000101011110110;
assign LUT_4[45564] = 32'b00000000000000000101000101110110;
assign LUT_4[45565] = 32'b11111111111111111110010001101110;
assign LUT_4[45566] = 32'b00000000000000000100100000011010;
assign LUT_4[45567] = 32'b11111111111111111101101100010010;
assign LUT_4[45568] = 32'b00000000000000001000110111011001;
assign LUT_4[45569] = 32'b00000000000000000010000011010001;
assign LUT_4[45570] = 32'b00000000000000001000010001111101;
assign LUT_4[45571] = 32'b00000000000000000001011101110101;
assign LUT_4[45572] = 32'b00000000000000000101110111110101;
assign LUT_4[45573] = 32'b11111111111111111111000011101101;
assign LUT_4[45574] = 32'b00000000000000000101010010011001;
assign LUT_4[45575] = 32'b11111111111111111110011110010001;
assign LUT_4[45576] = 32'b00000000000000000010000011101110;
assign LUT_4[45577] = 32'b11111111111111111011001111100110;
assign LUT_4[45578] = 32'b00000000000000000001011110010010;
assign LUT_4[45579] = 32'b11111111111111111010101010001010;
assign LUT_4[45580] = 32'b11111111111111111111000100001010;
assign LUT_4[45581] = 32'b11111111111111111000010000000010;
assign LUT_4[45582] = 32'b11111111111111111110011110101110;
assign LUT_4[45583] = 32'b11111111111111110111101010100110;
assign LUT_4[45584] = 32'b00000000000000000110101001000111;
assign LUT_4[45585] = 32'b11111111111111111111110100111111;
assign LUT_4[45586] = 32'b00000000000000000110000011101011;
assign LUT_4[45587] = 32'b11111111111111111111001111100011;
assign LUT_4[45588] = 32'b00000000000000000011101001100011;
assign LUT_4[45589] = 32'b11111111111111111100110101011011;
assign LUT_4[45590] = 32'b00000000000000000011000100000111;
assign LUT_4[45591] = 32'b11111111111111111100001111111111;
assign LUT_4[45592] = 32'b11111111111111111111110101011100;
assign LUT_4[45593] = 32'b11111111111111111001000001010100;
assign LUT_4[45594] = 32'b11111111111111111111010000000000;
assign LUT_4[45595] = 32'b11111111111111111000011011111000;
assign LUT_4[45596] = 32'b11111111111111111100110101111000;
assign LUT_4[45597] = 32'b11111111111111110110000001110000;
assign LUT_4[45598] = 32'b11111111111111111100010000011100;
assign LUT_4[45599] = 32'b11111111111111110101011100010100;
assign LUT_4[45600] = 32'b00000000000000000111010010100000;
assign LUT_4[45601] = 32'b00000000000000000000011110011000;
assign LUT_4[45602] = 32'b00000000000000000110101101000100;
assign LUT_4[45603] = 32'b11111111111111111111111000111100;
assign LUT_4[45604] = 32'b00000000000000000100010010111100;
assign LUT_4[45605] = 32'b11111111111111111101011110110100;
assign LUT_4[45606] = 32'b00000000000000000011101101100000;
assign LUT_4[45607] = 32'b11111111111111111100111001011000;
assign LUT_4[45608] = 32'b00000000000000000000011110110101;
assign LUT_4[45609] = 32'b11111111111111111001101010101101;
assign LUT_4[45610] = 32'b11111111111111111111111001011001;
assign LUT_4[45611] = 32'b11111111111111111001000101010001;
assign LUT_4[45612] = 32'b11111111111111111101011111010001;
assign LUT_4[45613] = 32'b11111111111111110110101011001001;
assign LUT_4[45614] = 32'b11111111111111111100111001110101;
assign LUT_4[45615] = 32'b11111111111111110110000101101101;
assign LUT_4[45616] = 32'b00000000000000000101000100001110;
assign LUT_4[45617] = 32'b11111111111111111110010000000110;
assign LUT_4[45618] = 32'b00000000000000000100011110110010;
assign LUT_4[45619] = 32'b11111111111111111101101010101010;
assign LUT_4[45620] = 32'b00000000000000000010000100101010;
assign LUT_4[45621] = 32'b11111111111111111011010000100010;
assign LUT_4[45622] = 32'b00000000000000000001011111001110;
assign LUT_4[45623] = 32'b11111111111111111010101011000110;
assign LUT_4[45624] = 32'b11111111111111111110010000100011;
assign LUT_4[45625] = 32'b11111111111111110111011100011011;
assign LUT_4[45626] = 32'b11111111111111111101101011000111;
assign LUT_4[45627] = 32'b11111111111111110110110110111111;
assign LUT_4[45628] = 32'b11111111111111111011010000111111;
assign LUT_4[45629] = 32'b11111111111111110100011100110111;
assign LUT_4[45630] = 32'b11111111111111111010101011100011;
assign LUT_4[45631] = 32'b11111111111111110011110111011011;
assign LUT_4[45632] = 32'b00000000000000001010001110101101;
assign LUT_4[45633] = 32'b00000000000000000011011010100101;
assign LUT_4[45634] = 32'b00000000000000001001101001010001;
assign LUT_4[45635] = 32'b00000000000000000010110101001001;
assign LUT_4[45636] = 32'b00000000000000000111001111001001;
assign LUT_4[45637] = 32'b00000000000000000000011011000001;
assign LUT_4[45638] = 32'b00000000000000000110101001101101;
assign LUT_4[45639] = 32'b11111111111111111111110101100101;
assign LUT_4[45640] = 32'b00000000000000000011011011000010;
assign LUT_4[45641] = 32'b11111111111111111100100110111010;
assign LUT_4[45642] = 32'b00000000000000000010110101100110;
assign LUT_4[45643] = 32'b11111111111111111100000001011110;
assign LUT_4[45644] = 32'b00000000000000000000011011011110;
assign LUT_4[45645] = 32'b11111111111111111001100111010110;
assign LUT_4[45646] = 32'b11111111111111111111110110000010;
assign LUT_4[45647] = 32'b11111111111111111001000001111010;
assign LUT_4[45648] = 32'b00000000000000001000000000011011;
assign LUT_4[45649] = 32'b00000000000000000001001100010011;
assign LUT_4[45650] = 32'b00000000000000000111011010111111;
assign LUT_4[45651] = 32'b00000000000000000000100110110111;
assign LUT_4[45652] = 32'b00000000000000000101000000110111;
assign LUT_4[45653] = 32'b11111111111111111110001100101111;
assign LUT_4[45654] = 32'b00000000000000000100011011011011;
assign LUT_4[45655] = 32'b11111111111111111101100111010011;
assign LUT_4[45656] = 32'b00000000000000000001001100110000;
assign LUT_4[45657] = 32'b11111111111111111010011000101000;
assign LUT_4[45658] = 32'b00000000000000000000100111010100;
assign LUT_4[45659] = 32'b11111111111111111001110011001100;
assign LUT_4[45660] = 32'b11111111111111111110001101001100;
assign LUT_4[45661] = 32'b11111111111111110111011001000100;
assign LUT_4[45662] = 32'b11111111111111111101100111110000;
assign LUT_4[45663] = 32'b11111111111111110110110011101000;
assign LUT_4[45664] = 32'b00000000000000001000101001110100;
assign LUT_4[45665] = 32'b00000000000000000001110101101100;
assign LUT_4[45666] = 32'b00000000000000001000000100011000;
assign LUT_4[45667] = 32'b00000000000000000001010000010000;
assign LUT_4[45668] = 32'b00000000000000000101101010010000;
assign LUT_4[45669] = 32'b11111111111111111110110110001000;
assign LUT_4[45670] = 32'b00000000000000000101000100110100;
assign LUT_4[45671] = 32'b11111111111111111110010000101100;
assign LUT_4[45672] = 32'b00000000000000000001110110001001;
assign LUT_4[45673] = 32'b11111111111111111011000010000001;
assign LUT_4[45674] = 32'b00000000000000000001010000101101;
assign LUT_4[45675] = 32'b11111111111111111010011100100101;
assign LUT_4[45676] = 32'b11111111111111111110110110100101;
assign LUT_4[45677] = 32'b11111111111111111000000010011101;
assign LUT_4[45678] = 32'b11111111111111111110010001001001;
assign LUT_4[45679] = 32'b11111111111111110111011101000001;
assign LUT_4[45680] = 32'b00000000000000000110011011100010;
assign LUT_4[45681] = 32'b11111111111111111111100111011010;
assign LUT_4[45682] = 32'b00000000000000000101110110000110;
assign LUT_4[45683] = 32'b11111111111111111111000001111110;
assign LUT_4[45684] = 32'b00000000000000000011011011111110;
assign LUT_4[45685] = 32'b11111111111111111100100111110110;
assign LUT_4[45686] = 32'b00000000000000000010110110100010;
assign LUT_4[45687] = 32'b11111111111111111100000010011010;
assign LUT_4[45688] = 32'b11111111111111111111100111110111;
assign LUT_4[45689] = 32'b11111111111111111000110011101111;
assign LUT_4[45690] = 32'b11111111111111111111000010011011;
assign LUT_4[45691] = 32'b11111111111111111000001110010011;
assign LUT_4[45692] = 32'b11111111111111111100101000010011;
assign LUT_4[45693] = 32'b11111111111111110101110100001011;
assign LUT_4[45694] = 32'b11111111111111111100000010110111;
assign LUT_4[45695] = 32'b11111111111111110101001110101111;
assign LUT_4[45696] = 32'b00000000000000001011011101100001;
assign LUT_4[45697] = 32'b00000000000000000100101001011001;
assign LUT_4[45698] = 32'b00000000000000001010111000000101;
assign LUT_4[45699] = 32'b00000000000000000100000011111101;
assign LUT_4[45700] = 32'b00000000000000001000011101111101;
assign LUT_4[45701] = 32'b00000000000000000001101001110101;
assign LUT_4[45702] = 32'b00000000000000000111111000100001;
assign LUT_4[45703] = 32'b00000000000000000001000100011001;
assign LUT_4[45704] = 32'b00000000000000000100101001110110;
assign LUT_4[45705] = 32'b11111111111111111101110101101110;
assign LUT_4[45706] = 32'b00000000000000000100000100011010;
assign LUT_4[45707] = 32'b11111111111111111101010000010010;
assign LUT_4[45708] = 32'b00000000000000000001101010010010;
assign LUT_4[45709] = 32'b11111111111111111010110110001010;
assign LUT_4[45710] = 32'b00000000000000000001000100110110;
assign LUT_4[45711] = 32'b11111111111111111010010000101110;
assign LUT_4[45712] = 32'b00000000000000001001001111001111;
assign LUT_4[45713] = 32'b00000000000000000010011011000111;
assign LUT_4[45714] = 32'b00000000000000001000101001110011;
assign LUT_4[45715] = 32'b00000000000000000001110101101011;
assign LUT_4[45716] = 32'b00000000000000000110001111101011;
assign LUT_4[45717] = 32'b11111111111111111111011011100011;
assign LUT_4[45718] = 32'b00000000000000000101101010001111;
assign LUT_4[45719] = 32'b11111111111111111110110110000111;
assign LUT_4[45720] = 32'b00000000000000000010011011100100;
assign LUT_4[45721] = 32'b11111111111111111011100111011100;
assign LUT_4[45722] = 32'b00000000000000000001110110001000;
assign LUT_4[45723] = 32'b11111111111111111011000010000000;
assign LUT_4[45724] = 32'b11111111111111111111011100000000;
assign LUT_4[45725] = 32'b11111111111111111000100111111000;
assign LUT_4[45726] = 32'b11111111111111111110110110100100;
assign LUT_4[45727] = 32'b11111111111111111000000010011100;
assign LUT_4[45728] = 32'b00000000000000001001111000101000;
assign LUT_4[45729] = 32'b00000000000000000011000100100000;
assign LUT_4[45730] = 32'b00000000000000001001010011001100;
assign LUT_4[45731] = 32'b00000000000000000010011111000100;
assign LUT_4[45732] = 32'b00000000000000000110111001000100;
assign LUT_4[45733] = 32'b00000000000000000000000100111100;
assign LUT_4[45734] = 32'b00000000000000000110010011101000;
assign LUT_4[45735] = 32'b11111111111111111111011111100000;
assign LUT_4[45736] = 32'b00000000000000000011000100111101;
assign LUT_4[45737] = 32'b11111111111111111100010000110101;
assign LUT_4[45738] = 32'b00000000000000000010011111100001;
assign LUT_4[45739] = 32'b11111111111111111011101011011001;
assign LUT_4[45740] = 32'b00000000000000000000000101011001;
assign LUT_4[45741] = 32'b11111111111111111001010001010001;
assign LUT_4[45742] = 32'b11111111111111111111011111111101;
assign LUT_4[45743] = 32'b11111111111111111000101011110101;
assign LUT_4[45744] = 32'b00000000000000000111101010010110;
assign LUT_4[45745] = 32'b00000000000000000000110110001110;
assign LUT_4[45746] = 32'b00000000000000000111000100111010;
assign LUT_4[45747] = 32'b00000000000000000000010000110010;
assign LUT_4[45748] = 32'b00000000000000000100101010110010;
assign LUT_4[45749] = 32'b11111111111111111101110110101010;
assign LUT_4[45750] = 32'b00000000000000000100000101010110;
assign LUT_4[45751] = 32'b11111111111111111101010001001110;
assign LUT_4[45752] = 32'b00000000000000000000110110101011;
assign LUT_4[45753] = 32'b11111111111111111010000010100011;
assign LUT_4[45754] = 32'b00000000000000000000010001001111;
assign LUT_4[45755] = 32'b11111111111111111001011101000111;
assign LUT_4[45756] = 32'b11111111111111111101110111000111;
assign LUT_4[45757] = 32'b11111111111111110111000010111111;
assign LUT_4[45758] = 32'b11111111111111111101010001101011;
assign LUT_4[45759] = 32'b11111111111111110110011101100011;
assign LUT_4[45760] = 32'b00000000000000001100110100110101;
assign LUT_4[45761] = 32'b00000000000000000110000000101101;
assign LUT_4[45762] = 32'b00000000000000001100001111011001;
assign LUT_4[45763] = 32'b00000000000000000101011011010001;
assign LUT_4[45764] = 32'b00000000000000001001110101010001;
assign LUT_4[45765] = 32'b00000000000000000011000001001001;
assign LUT_4[45766] = 32'b00000000000000001001001111110101;
assign LUT_4[45767] = 32'b00000000000000000010011011101101;
assign LUT_4[45768] = 32'b00000000000000000110000001001010;
assign LUT_4[45769] = 32'b11111111111111111111001101000010;
assign LUT_4[45770] = 32'b00000000000000000101011011101110;
assign LUT_4[45771] = 32'b11111111111111111110100111100110;
assign LUT_4[45772] = 32'b00000000000000000011000001100110;
assign LUT_4[45773] = 32'b11111111111111111100001101011110;
assign LUT_4[45774] = 32'b00000000000000000010011100001010;
assign LUT_4[45775] = 32'b11111111111111111011101000000010;
assign LUT_4[45776] = 32'b00000000000000001010100110100011;
assign LUT_4[45777] = 32'b00000000000000000011110010011011;
assign LUT_4[45778] = 32'b00000000000000001010000001000111;
assign LUT_4[45779] = 32'b00000000000000000011001100111111;
assign LUT_4[45780] = 32'b00000000000000000111100110111111;
assign LUT_4[45781] = 32'b00000000000000000000110010110111;
assign LUT_4[45782] = 32'b00000000000000000111000001100011;
assign LUT_4[45783] = 32'b00000000000000000000001101011011;
assign LUT_4[45784] = 32'b00000000000000000011110010111000;
assign LUT_4[45785] = 32'b11111111111111111100111110110000;
assign LUT_4[45786] = 32'b00000000000000000011001101011100;
assign LUT_4[45787] = 32'b11111111111111111100011001010100;
assign LUT_4[45788] = 32'b00000000000000000000110011010100;
assign LUT_4[45789] = 32'b11111111111111111001111111001100;
assign LUT_4[45790] = 32'b00000000000000000000001101111000;
assign LUT_4[45791] = 32'b11111111111111111001011001110000;
assign LUT_4[45792] = 32'b00000000000000001011001111111100;
assign LUT_4[45793] = 32'b00000000000000000100011011110100;
assign LUT_4[45794] = 32'b00000000000000001010101010100000;
assign LUT_4[45795] = 32'b00000000000000000011110110011000;
assign LUT_4[45796] = 32'b00000000000000001000010000011000;
assign LUT_4[45797] = 32'b00000000000000000001011100010000;
assign LUT_4[45798] = 32'b00000000000000000111101010111100;
assign LUT_4[45799] = 32'b00000000000000000000110110110100;
assign LUT_4[45800] = 32'b00000000000000000100011100010001;
assign LUT_4[45801] = 32'b11111111111111111101101000001001;
assign LUT_4[45802] = 32'b00000000000000000011110110110101;
assign LUT_4[45803] = 32'b11111111111111111101000010101101;
assign LUT_4[45804] = 32'b00000000000000000001011100101101;
assign LUT_4[45805] = 32'b11111111111111111010101000100101;
assign LUT_4[45806] = 32'b00000000000000000000110111010001;
assign LUT_4[45807] = 32'b11111111111111111010000011001001;
assign LUT_4[45808] = 32'b00000000000000001001000001101010;
assign LUT_4[45809] = 32'b00000000000000000010001101100010;
assign LUT_4[45810] = 32'b00000000000000001000011100001110;
assign LUT_4[45811] = 32'b00000000000000000001101000000110;
assign LUT_4[45812] = 32'b00000000000000000110000010000110;
assign LUT_4[45813] = 32'b11111111111111111111001101111110;
assign LUT_4[45814] = 32'b00000000000000000101011100101010;
assign LUT_4[45815] = 32'b11111111111111111110101000100010;
assign LUT_4[45816] = 32'b00000000000000000010001101111111;
assign LUT_4[45817] = 32'b11111111111111111011011001110111;
assign LUT_4[45818] = 32'b00000000000000000001101000100011;
assign LUT_4[45819] = 32'b11111111111111111010110100011011;
assign LUT_4[45820] = 32'b11111111111111111111001110011011;
assign LUT_4[45821] = 32'b11111111111111111000011010010011;
assign LUT_4[45822] = 32'b11111111111111111110101000111111;
assign LUT_4[45823] = 32'b11111111111111110111110100110111;
assign LUT_4[45824] = 32'b00000000000000001101110010111100;
assign LUT_4[45825] = 32'b00000000000000000110111110110100;
assign LUT_4[45826] = 32'b00000000000000001101001101100000;
assign LUT_4[45827] = 32'b00000000000000000110011001011000;
assign LUT_4[45828] = 32'b00000000000000001010110011011000;
assign LUT_4[45829] = 32'b00000000000000000011111111010000;
assign LUT_4[45830] = 32'b00000000000000001010001101111100;
assign LUT_4[45831] = 32'b00000000000000000011011001110100;
assign LUT_4[45832] = 32'b00000000000000000110111111010001;
assign LUT_4[45833] = 32'b00000000000000000000001011001001;
assign LUT_4[45834] = 32'b00000000000000000110011001110101;
assign LUT_4[45835] = 32'b11111111111111111111100101101101;
assign LUT_4[45836] = 32'b00000000000000000011111111101101;
assign LUT_4[45837] = 32'b11111111111111111101001011100101;
assign LUT_4[45838] = 32'b00000000000000000011011010010001;
assign LUT_4[45839] = 32'b11111111111111111100100110001001;
assign LUT_4[45840] = 32'b00000000000000001011100100101010;
assign LUT_4[45841] = 32'b00000000000000000100110000100010;
assign LUT_4[45842] = 32'b00000000000000001010111111001110;
assign LUT_4[45843] = 32'b00000000000000000100001011000110;
assign LUT_4[45844] = 32'b00000000000000001000100101000110;
assign LUT_4[45845] = 32'b00000000000000000001110000111110;
assign LUT_4[45846] = 32'b00000000000000000111111111101010;
assign LUT_4[45847] = 32'b00000000000000000001001011100010;
assign LUT_4[45848] = 32'b00000000000000000100110000111111;
assign LUT_4[45849] = 32'b11111111111111111101111100110111;
assign LUT_4[45850] = 32'b00000000000000000100001011100011;
assign LUT_4[45851] = 32'b11111111111111111101010111011011;
assign LUT_4[45852] = 32'b00000000000000000001110001011011;
assign LUT_4[45853] = 32'b11111111111111111010111101010011;
assign LUT_4[45854] = 32'b00000000000000000001001011111111;
assign LUT_4[45855] = 32'b11111111111111111010010111110111;
assign LUT_4[45856] = 32'b00000000000000001100001110000011;
assign LUT_4[45857] = 32'b00000000000000000101011001111011;
assign LUT_4[45858] = 32'b00000000000000001011101000100111;
assign LUT_4[45859] = 32'b00000000000000000100110100011111;
assign LUT_4[45860] = 32'b00000000000000001001001110011111;
assign LUT_4[45861] = 32'b00000000000000000010011010010111;
assign LUT_4[45862] = 32'b00000000000000001000101001000011;
assign LUT_4[45863] = 32'b00000000000000000001110100111011;
assign LUT_4[45864] = 32'b00000000000000000101011010011000;
assign LUT_4[45865] = 32'b11111111111111111110100110010000;
assign LUT_4[45866] = 32'b00000000000000000100110100111100;
assign LUT_4[45867] = 32'b11111111111111111110000000110100;
assign LUT_4[45868] = 32'b00000000000000000010011010110100;
assign LUT_4[45869] = 32'b11111111111111111011100110101100;
assign LUT_4[45870] = 32'b00000000000000000001110101011000;
assign LUT_4[45871] = 32'b11111111111111111011000001010000;
assign LUT_4[45872] = 32'b00000000000000001001111111110001;
assign LUT_4[45873] = 32'b00000000000000000011001011101001;
assign LUT_4[45874] = 32'b00000000000000001001011010010101;
assign LUT_4[45875] = 32'b00000000000000000010100110001101;
assign LUT_4[45876] = 32'b00000000000000000111000000001101;
assign LUT_4[45877] = 32'b00000000000000000000001100000101;
assign LUT_4[45878] = 32'b00000000000000000110011010110001;
assign LUT_4[45879] = 32'b11111111111111111111100110101001;
assign LUT_4[45880] = 32'b00000000000000000011001100000110;
assign LUT_4[45881] = 32'b11111111111111111100010111111110;
assign LUT_4[45882] = 32'b00000000000000000010100110101010;
assign LUT_4[45883] = 32'b11111111111111111011110010100010;
assign LUT_4[45884] = 32'b00000000000000000000001100100010;
assign LUT_4[45885] = 32'b11111111111111111001011000011010;
assign LUT_4[45886] = 32'b11111111111111111111100111000110;
assign LUT_4[45887] = 32'b11111111111111111000110010111110;
assign LUT_4[45888] = 32'b00000000000000001111001010010000;
assign LUT_4[45889] = 32'b00000000000000001000010110001000;
assign LUT_4[45890] = 32'b00000000000000001110100100110100;
assign LUT_4[45891] = 32'b00000000000000000111110000101100;
assign LUT_4[45892] = 32'b00000000000000001100001010101100;
assign LUT_4[45893] = 32'b00000000000000000101010110100100;
assign LUT_4[45894] = 32'b00000000000000001011100101010000;
assign LUT_4[45895] = 32'b00000000000000000100110001001000;
assign LUT_4[45896] = 32'b00000000000000001000010110100101;
assign LUT_4[45897] = 32'b00000000000000000001100010011101;
assign LUT_4[45898] = 32'b00000000000000000111110001001001;
assign LUT_4[45899] = 32'b00000000000000000000111101000001;
assign LUT_4[45900] = 32'b00000000000000000101010111000001;
assign LUT_4[45901] = 32'b11111111111111111110100010111001;
assign LUT_4[45902] = 32'b00000000000000000100110001100101;
assign LUT_4[45903] = 32'b11111111111111111101111101011101;
assign LUT_4[45904] = 32'b00000000000000001100111011111110;
assign LUT_4[45905] = 32'b00000000000000000110000111110110;
assign LUT_4[45906] = 32'b00000000000000001100010110100010;
assign LUT_4[45907] = 32'b00000000000000000101100010011010;
assign LUT_4[45908] = 32'b00000000000000001001111100011010;
assign LUT_4[45909] = 32'b00000000000000000011001000010010;
assign LUT_4[45910] = 32'b00000000000000001001010110111110;
assign LUT_4[45911] = 32'b00000000000000000010100010110110;
assign LUT_4[45912] = 32'b00000000000000000110001000010011;
assign LUT_4[45913] = 32'b11111111111111111111010100001011;
assign LUT_4[45914] = 32'b00000000000000000101100010110111;
assign LUT_4[45915] = 32'b11111111111111111110101110101111;
assign LUT_4[45916] = 32'b00000000000000000011001000101111;
assign LUT_4[45917] = 32'b11111111111111111100010100100111;
assign LUT_4[45918] = 32'b00000000000000000010100011010011;
assign LUT_4[45919] = 32'b11111111111111111011101111001011;
assign LUT_4[45920] = 32'b00000000000000001101100101010111;
assign LUT_4[45921] = 32'b00000000000000000110110001001111;
assign LUT_4[45922] = 32'b00000000000000001100111111111011;
assign LUT_4[45923] = 32'b00000000000000000110001011110011;
assign LUT_4[45924] = 32'b00000000000000001010100101110011;
assign LUT_4[45925] = 32'b00000000000000000011110001101011;
assign LUT_4[45926] = 32'b00000000000000001010000000010111;
assign LUT_4[45927] = 32'b00000000000000000011001100001111;
assign LUT_4[45928] = 32'b00000000000000000110110001101100;
assign LUT_4[45929] = 32'b11111111111111111111111101100100;
assign LUT_4[45930] = 32'b00000000000000000110001100010000;
assign LUT_4[45931] = 32'b11111111111111111111011000001000;
assign LUT_4[45932] = 32'b00000000000000000011110010001000;
assign LUT_4[45933] = 32'b11111111111111111100111110000000;
assign LUT_4[45934] = 32'b00000000000000000011001100101100;
assign LUT_4[45935] = 32'b11111111111111111100011000100100;
assign LUT_4[45936] = 32'b00000000000000001011010111000101;
assign LUT_4[45937] = 32'b00000000000000000100100010111101;
assign LUT_4[45938] = 32'b00000000000000001010110001101001;
assign LUT_4[45939] = 32'b00000000000000000011111101100001;
assign LUT_4[45940] = 32'b00000000000000001000010111100001;
assign LUT_4[45941] = 32'b00000000000000000001100011011001;
assign LUT_4[45942] = 32'b00000000000000000111110010000101;
assign LUT_4[45943] = 32'b00000000000000000000111101111101;
assign LUT_4[45944] = 32'b00000000000000000100100011011010;
assign LUT_4[45945] = 32'b11111111111111111101101111010010;
assign LUT_4[45946] = 32'b00000000000000000011111101111110;
assign LUT_4[45947] = 32'b11111111111111111101001001110110;
assign LUT_4[45948] = 32'b00000000000000000001100011110110;
assign LUT_4[45949] = 32'b11111111111111111010101111101110;
assign LUT_4[45950] = 32'b00000000000000000000111110011010;
assign LUT_4[45951] = 32'b11111111111111111010001010010010;
assign LUT_4[45952] = 32'b00000000000000010000011001000100;
assign LUT_4[45953] = 32'b00000000000000001001100100111100;
assign LUT_4[45954] = 32'b00000000000000001111110011101000;
assign LUT_4[45955] = 32'b00000000000000001000111111100000;
assign LUT_4[45956] = 32'b00000000000000001101011001100000;
assign LUT_4[45957] = 32'b00000000000000000110100101011000;
assign LUT_4[45958] = 32'b00000000000000001100110100000100;
assign LUT_4[45959] = 32'b00000000000000000101111111111100;
assign LUT_4[45960] = 32'b00000000000000001001100101011001;
assign LUT_4[45961] = 32'b00000000000000000010110001010001;
assign LUT_4[45962] = 32'b00000000000000001000111111111101;
assign LUT_4[45963] = 32'b00000000000000000010001011110101;
assign LUT_4[45964] = 32'b00000000000000000110100101110101;
assign LUT_4[45965] = 32'b11111111111111111111110001101101;
assign LUT_4[45966] = 32'b00000000000000000110000000011001;
assign LUT_4[45967] = 32'b11111111111111111111001100010001;
assign LUT_4[45968] = 32'b00000000000000001110001010110010;
assign LUT_4[45969] = 32'b00000000000000000111010110101010;
assign LUT_4[45970] = 32'b00000000000000001101100101010110;
assign LUT_4[45971] = 32'b00000000000000000110110001001110;
assign LUT_4[45972] = 32'b00000000000000001011001011001110;
assign LUT_4[45973] = 32'b00000000000000000100010111000110;
assign LUT_4[45974] = 32'b00000000000000001010100101110010;
assign LUT_4[45975] = 32'b00000000000000000011110001101010;
assign LUT_4[45976] = 32'b00000000000000000111010111000111;
assign LUT_4[45977] = 32'b00000000000000000000100010111111;
assign LUT_4[45978] = 32'b00000000000000000110110001101011;
assign LUT_4[45979] = 32'b11111111111111111111111101100011;
assign LUT_4[45980] = 32'b00000000000000000100010111100011;
assign LUT_4[45981] = 32'b11111111111111111101100011011011;
assign LUT_4[45982] = 32'b00000000000000000011110010000111;
assign LUT_4[45983] = 32'b11111111111111111100111101111111;
assign LUT_4[45984] = 32'b00000000000000001110110100001011;
assign LUT_4[45985] = 32'b00000000000000001000000000000011;
assign LUT_4[45986] = 32'b00000000000000001110001110101111;
assign LUT_4[45987] = 32'b00000000000000000111011010100111;
assign LUT_4[45988] = 32'b00000000000000001011110100100111;
assign LUT_4[45989] = 32'b00000000000000000101000000011111;
assign LUT_4[45990] = 32'b00000000000000001011001111001011;
assign LUT_4[45991] = 32'b00000000000000000100011011000011;
assign LUT_4[45992] = 32'b00000000000000001000000000100000;
assign LUT_4[45993] = 32'b00000000000000000001001100011000;
assign LUT_4[45994] = 32'b00000000000000000111011011000100;
assign LUT_4[45995] = 32'b00000000000000000000100110111100;
assign LUT_4[45996] = 32'b00000000000000000101000000111100;
assign LUT_4[45997] = 32'b11111111111111111110001100110100;
assign LUT_4[45998] = 32'b00000000000000000100011011100000;
assign LUT_4[45999] = 32'b11111111111111111101100111011000;
assign LUT_4[46000] = 32'b00000000000000001100100101111001;
assign LUT_4[46001] = 32'b00000000000000000101110001110001;
assign LUT_4[46002] = 32'b00000000000000001100000000011101;
assign LUT_4[46003] = 32'b00000000000000000101001100010101;
assign LUT_4[46004] = 32'b00000000000000001001100110010101;
assign LUT_4[46005] = 32'b00000000000000000010110010001101;
assign LUT_4[46006] = 32'b00000000000000001001000000111001;
assign LUT_4[46007] = 32'b00000000000000000010001100110001;
assign LUT_4[46008] = 32'b00000000000000000101110010001110;
assign LUT_4[46009] = 32'b11111111111111111110111110000110;
assign LUT_4[46010] = 32'b00000000000000000101001100110010;
assign LUT_4[46011] = 32'b11111111111111111110011000101010;
assign LUT_4[46012] = 32'b00000000000000000010110010101010;
assign LUT_4[46013] = 32'b11111111111111111011111110100010;
assign LUT_4[46014] = 32'b00000000000000000010001101001110;
assign LUT_4[46015] = 32'b11111111111111111011011001000110;
assign LUT_4[46016] = 32'b00000000000000010001110000011000;
assign LUT_4[46017] = 32'b00000000000000001010111100010000;
assign LUT_4[46018] = 32'b00000000000000010001001010111100;
assign LUT_4[46019] = 32'b00000000000000001010010110110100;
assign LUT_4[46020] = 32'b00000000000000001110110000110100;
assign LUT_4[46021] = 32'b00000000000000000111111100101100;
assign LUT_4[46022] = 32'b00000000000000001110001011011000;
assign LUT_4[46023] = 32'b00000000000000000111010111010000;
assign LUT_4[46024] = 32'b00000000000000001010111100101101;
assign LUT_4[46025] = 32'b00000000000000000100001000100101;
assign LUT_4[46026] = 32'b00000000000000001010010111010001;
assign LUT_4[46027] = 32'b00000000000000000011100011001001;
assign LUT_4[46028] = 32'b00000000000000000111111101001001;
assign LUT_4[46029] = 32'b00000000000000000001001001000001;
assign LUT_4[46030] = 32'b00000000000000000111010111101101;
assign LUT_4[46031] = 32'b00000000000000000000100011100101;
assign LUT_4[46032] = 32'b00000000000000001111100010000110;
assign LUT_4[46033] = 32'b00000000000000001000101101111110;
assign LUT_4[46034] = 32'b00000000000000001110111100101010;
assign LUT_4[46035] = 32'b00000000000000001000001000100010;
assign LUT_4[46036] = 32'b00000000000000001100100010100010;
assign LUT_4[46037] = 32'b00000000000000000101101110011010;
assign LUT_4[46038] = 32'b00000000000000001011111101000110;
assign LUT_4[46039] = 32'b00000000000000000101001000111110;
assign LUT_4[46040] = 32'b00000000000000001000101110011011;
assign LUT_4[46041] = 32'b00000000000000000001111010010011;
assign LUT_4[46042] = 32'b00000000000000001000001000111111;
assign LUT_4[46043] = 32'b00000000000000000001010100110111;
assign LUT_4[46044] = 32'b00000000000000000101101110110111;
assign LUT_4[46045] = 32'b11111111111111111110111010101111;
assign LUT_4[46046] = 32'b00000000000000000101001001011011;
assign LUT_4[46047] = 32'b11111111111111111110010101010011;
assign LUT_4[46048] = 32'b00000000000000010000001011011111;
assign LUT_4[46049] = 32'b00000000000000001001010111010111;
assign LUT_4[46050] = 32'b00000000000000001111100110000011;
assign LUT_4[46051] = 32'b00000000000000001000110001111011;
assign LUT_4[46052] = 32'b00000000000000001101001011111011;
assign LUT_4[46053] = 32'b00000000000000000110010111110011;
assign LUT_4[46054] = 32'b00000000000000001100100110011111;
assign LUT_4[46055] = 32'b00000000000000000101110010010111;
assign LUT_4[46056] = 32'b00000000000000001001010111110100;
assign LUT_4[46057] = 32'b00000000000000000010100011101100;
assign LUT_4[46058] = 32'b00000000000000001000110010011000;
assign LUT_4[46059] = 32'b00000000000000000001111110010000;
assign LUT_4[46060] = 32'b00000000000000000110011000010000;
assign LUT_4[46061] = 32'b11111111111111111111100100001000;
assign LUT_4[46062] = 32'b00000000000000000101110010110100;
assign LUT_4[46063] = 32'b11111111111111111110111110101100;
assign LUT_4[46064] = 32'b00000000000000001101111101001101;
assign LUT_4[46065] = 32'b00000000000000000111001001000101;
assign LUT_4[46066] = 32'b00000000000000001101010111110001;
assign LUT_4[46067] = 32'b00000000000000000110100011101001;
assign LUT_4[46068] = 32'b00000000000000001010111101101001;
assign LUT_4[46069] = 32'b00000000000000000100001001100001;
assign LUT_4[46070] = 32'b00000000000000001010011000001101;
assign LUT_4[46071] = 32'b00000000000000000011100100000101;
assign LUT_4[46072] = 32'b00000000000000000111001001100010;
assign LUT_4[46073] = 32'b00000000000000000000010101011010;
assign LUT_4[46074] = 32'b00000000000000000110100100000110;
assign LUT_4[46075] = 32'b11111111111111111111101111111110;
assign LUT_4[46076] = 32'b00000000000000000100001001111110;
assign LUT_4[46077] = 32'b11111111111111111101010101110110;
assign LUT_4[46078] = 32'b00000000000000000011100100100010;
assign LUT_4[46079] = 32'b11111111111111111100110000011010;
assign LUT_4[46080] = 32'b00000000000000001011011101110000;
assign LUT_4[46081] = 32'b00000000000000000100101001101000;
assign LUT_4[46082] = 32'b00000000000000001010111000010100;
assign LUT_4[46083] = 32'b00000000000000000100000100001100;
assign LUT_4[46084] = 32'b00000000000000001000011110001100;
assign LUT_4[46085] = 32'b00000000000000000001101010000100;
assign LUT_4[46086] = 32'b00000000000000000111111000110000;
assign LUT_4[46087] = 32'b00000000000000000001000100101000;
assign LUT_4[46088] = 32'b00000000000000000100101010000101;
assign LUT_4[46089] = 32'b11111111111111111101110101111101;
assign LUT_4[46090] = 32'b00000000000000000100000100101001;
assign LUT_4[46091] = 32'b11111111111111111101010000100001;
assign LUT_4[46092] = 32'b00000000000000000001101010100001;
assign LUT_4[46093] = 32'b11111111111111111010110110011001;
assign LUT_4[46094] = 32'b00000000000000000001000101000101;
assign LUT_4[46095] = 32'b11111111111111111010010000111101;
assign LUT_4[46096] = 32'b00000000000000001001001111011110;
assign LUT_4[46097] = 32'b00000000000000000010011011010110;
assign LUT_4[46098] = 32'b00000000000000001000101010000010;
assign LUT_4[46099] = 32'b00000000000000000001110101111010;
assign LUT_4[46100] = 32'b00000000000000000110001111111010;
assign LUT_4[46101] = 32'b11111111111111111111011011110010;
assign LUT_4[46102] = 32'b00000000000000000101101010011110;
assign LUT_4[46103] = 32'b11111111111111111110110110010110;
assign LUT_4[46104] = 32'b00000000000000000010011011110011;
assign LUT_4[46105] = 32'b11111111111111111011100111101011;
assign LUT_4[46106] = 32'b00000000000000000001110110010111;
assign LUT_4[46107] = 32'b11111111111111111011000010001111;
assign LUT_4[46108] = 32'b11111111111111111111011100001111;
assign LUT_4[46109] = 32'b11111111111111111000101000000111;
assign LUT_4[46110] = 32'b11111111111111111110110110110011;
assign LUT_4[46111] = 32'b11111111111111111000000010101011;
assign LUT_4[46112] = 32'b00000000000000001001111000110111;
assign LUT_4[46113] = 32'b00000000000000000011000100101111;
assign LUT_4[46114] = 32'b00000000000000001001010011011011;
assign LUT_4[46115] = 32'b00000000000000000010011111010011;
assign LUT_4[46116] = 32'b00000000000000000110111001010011;
assign LUT_4[46117] = 32'b00000000000000000000000101001011;
assign LUT_4[46118] = 32'b00000000000000000110010011110111;
assign LUT_4[46119] = 32'b11111111111111111111011111101111;
assign LUT_4[46120] = 32'b00000000000000000011000101001100;
assign LUT_4[46121] = 32'b11111111111111111100010001000100;
assign LUT_4[46122] = 32'b00000000000000000010011111110000;
assign LUT_4[46123] = 32'b11111111111111111011101011101000;
assign LUT_4[46124] = 32'b00000000000000000000000101101000;
assign LUT_4[46125] = 32'b11111111111111111001010001100000;
assign LUT_4[46126] = 32'b11111111111111111111100000001100;
assign LUT_4[46127] = 32'b11111111111111111000101100000100;
assign LUT_4[46128] = 32'b00000000000000000111101010100101;
assign LUT_4[46129] = 32'b00000000000000000000110110011101;
assign LUT_4[46130] = 32'b00000000000000000111000101001001;
assign LUT_4[46131] = 32'b00000000000000000000010001000001;
assign LUT_4[46132] = 32'b00000000000000000100101011000001;
assign LUT_4[46133] = 32'b11111111111111111101110110111001;
assign LUT_4[46134] = 32'b00000000000000000100000101100101;
assign LUT_4[46135] = 32'b11111111111111111101010001011101;
assign LUT_4[46136] = 32'b00000000000000000000110110111010;
assign LUT_4[46137] = 32'b11111111111111111010000010110010;
assign LUT_4[46138] = 32'b00000000000000000000010001011110;
assign LUT_4[46139] = 32'b11111111111111111001011101010110;
assign LUT_4[46140] = 32'b11111111111111111101110111010110;
assign LUT_4[46141] = 32'b11111111111111110111000011001110;
assign LUT_4[46142] = 32'b11111111111111111101010001111010;
assign LUT_4[46143] = 32'b11111111111111110110011101110010;
assign LUT_4[46144] = 32'b00000000000000001100110101000100;
assign LUT_4[46145] = 32'b00000000000000000110000000111100;
assign LUT_4[46146] = 32'b00000000000000001100001111101000;
assign LUT_4[46147] = 32'b00000000000000000101011011100000;
assign LUT_4[46148] = 32'b00000000000000001001110101100000;
assign LUT_4[46149] = 32'b00000000000000000011000001011000;
assign LUT_4[46150] = 32'b00000000000000001001010000000100;
assign LUT_4[46151] = 32'b00000000000000000010011011111100;
assign LUT_4[46152] = 32'b00000000000000000110000001011001;
assign LUT_4[46153] = 32'b11111111111111111111001101010001;
assign LUT_4[46154] = 32'b00000000000000000101011011111101;
assign LUT_4[46155] = 32'b11111111111111111110100111110101;
assign LUT_4[46156] = 32'b00000000000000000011000001110101;
assign LUT_4[46157] = 32'b11111111111111111100001101101101;
assign LUT_4[46158] = 32'b00000000000000000010011100011001;
assign LUT_4[46159] = 32'b11111111111111111011101000010001;
assign LUT_4[46160] = 32'b00000000000000001010100110110010;
assign LUT_4[46161] = 32'b00000000000000000011110010101010;
assign LUT_4[46162] = 32'b00000000000000001010000001010110;
assign LUT_4[46163] = 32'b00000000000000000011001101001110;
assign LUT_4[46164] = 32'b00000000000000000111100111001110;
assign LUT_4[46165] = 32'b00000000000000000000110011000110;
assign LUT_4[46166] = 32'b00000000000000000111000001110010;
assign LUT_4[46167] = 32'b00000000000000000000001101101010;
assign LUT_4[46168] = 32'b00000000000000000011110011000111;
assign LUT_4[46169] = 32'b11111111111111111100111110111111;
assign LUT_4[46170] = 32'b00000000000000000011001101101011;
assign LUT_4[46171] = 32'b11111111111111111100011001100011;
assign LUT_4[46172] = 32'b00000000000000000000110011100011;
assign LUT_4[46173] = 32'b11111111111111111001111111011011;
assign LUT_4[46174] = 32'b00000000000000000000001110000111;
assign LUT_4[46175] = 32'b11111111111111111001011001111111;
assign LUT_4[46176] = 32'b00000000000000001011010000001011;
assign LUT_4[46177] = 32'b00000000000000000100011100000011;
assign LUT_4[46178] = 32'b00000000000000001010101010101111;
assign LUT_4[46179] = 32'b00000000000000000011110110100111;
assign LUT_4[46180] = 32'b00000000000000001000010000100111;
assign LUT_4[46181] = 32'b00000000000000000001011100011111;
assign LUT_4[46182] = 32'b00000000000000000111101011001011;
assign LUT_4[46183] = 32'b00000000000000000000110111000011;
assign LUT_4[46184] = 32'b00000000000000000100011100100000;
assign LUT_4[46185] = 32'b11111111111111111101101000011000;
assign LUT_4[46186] = 32'b00000000000000000011110111000100;
assign LUT_4[46187] = 32'b11111111111111111101000010111100;
assign LUT_4[46188] = 32'b00000000000000000001011100111100;
assign LUT_4[46189] = 32'b11111111111111111010101000110100;
assign LUT_4[46190] = 32'b00000000000000000000110111100000;
assign LUT_4[46191] = 32'b11111111111111111010000011011000;
assign LUT_4[46192] = 32'b00000000000000001001000001111001;
assign LUT_4[46193] = 32'b00000000000000000010001101110001;
assign LUT_4[46194] = 32'b00000000000000001000011100011101;
assign LUT_4[46195] = 32'b00000000000000000001101000010101;
assign LUT_4[46196] = 32'b00000000000000000110000010010101;
assign LUT_4[46197] = 32'b11111111111111111111001110001101;
assign LUT_4[46198] = 32'b00000000000000000101011100111001;
assign LUT_4[46199] = 32'b11111111111111111110101000110001;
assign LUT_4[46200] = 32'b00000000000000000010001110001110;
assign LUT_4[46201] = 32'b11111111111111111011011010000110;
assign LUT_4[46202] = 32'b00000000000000000001101000110010;
assign LUT_4[46203] = 32'b11111111111111111010110100101010;
assign LUT_4[46204] = 32'b11111111111111111111001110101010;
assign LUT_4[46205] = 32'b11111111111111111000011010100010;
assign LUT_4[46206] = 32'b11111111111111111110101001001110;
assign LUT_4[46207] = 32'b11111111111111110111110101000110;
assign LUT_4[46208] = 32'b00000000000000001110000011111000;
assign LUT_4[46209] = 32'b00000000000000000111001111110000;
assign LUT_4[46210] = 32'b00000000000000001101011110011100;
assign LUT_4[46211] = 32'b00000000000000000110101010010100;
assign LUT_4[46212] = 32'b00000000000000001011000100010100;
assign LUT_4[46213] = 32'b00000000000000000100010000001100;
assign LUT_4[46214] = 32'b00000000000000001010011110111000;
assign LUT_4[46215] = 32'b00000000000000000011101010110000;
assign LUT_4[46216] = 32'b00000000000000000111010000001101;
assign LUT_4[46217] = 32'b00000000000000000000011100000101;
assign LUT_4[46218] = 32'b00000000000000000110101010110001;
assign LUT_4[46219] = 32'b11111111111111111111110110101001;
assign LUT_4[46220] = 32'b00000000000000000100010000101001;
assign LUT_4[46221] = 32'b11111111111111111101011100100001;
assign LUT_4[46222] = 32'b00000000000000000011101011001101;
assign LUT_4[46223] = 32'b11111111111111111100110111000101;
assign LUT_4[46224] = 32'b00000000000000001011110101100110;
assign LUT_4[46225] = 32'b00000000000000000101000001011110;
assign LUT_4[46226] = 32'b00000000000000001011010000001010;
assign LUT_4[46227] = 32'b00000000000000000100011100000010;
assign LUT_4[46228] = 32'b00000000000000001000110110000010;
assign LUT_4[46229] = 32'b00000000000000000010000001111010;
assign LUT_4[46230] = 32'b00000000000000001000010000100110;
assign LUT_4[46231] = 32'b00000000000000000001011100011110;
assign LUT_4[46232] = 32'b00000000000000000101000001111011;
assign LUT_4[46233] = 32'b11111111111111111110001101110011;
assign LUT_4[46234] = 32'b00000000000000000100011100011111;
assign LUT_4[46235] = 32'b11111111111111111101101000010111;
assign LUT_4[46236] = 32'b00000000000000000010000010010111;
assign LUT_4[46237] = 32'b11111111111111111011001110001111;
assign LUT_4[46238] = 32'b00000000000000000001011100111011;
assign LUT_4[46239] = 32'b11111111111111111010101000110011;
assign LUT_4[46240] = 32'b00000000000000001100011110111111;
assign LUT_4[46241] = 32'b00000000000000000101101010110111;
assign LUT_4[46242] = 32'b00000000000000001011111001100011;
assign LUT_4[46243] = 32'b00000000000000000101000101011011;
assign LUT_4[46244] = 32'b00000000000000001001011111011011;
assign LUT_4[46245] = 32'b00000000000000000010101011010011;
assign LUT_4[46246] = 32'b00000000000000001000111001111111;
assign LUT_4[46247] = 32'b00000000000000000010000101110111;
assign LUT_4[46248] = 32'b00000000000000000101101011010100;
assign LUT_4[46249] = 32'b11111111111111111110110111001100;
assign LUT_4[46250] = 32'b00000000000000000101000101111000;
assign LUT_4[46251] = 32'b11111111111111111110010001110000;
assign LUT_4[46252] = 32'b00000000000000000010101011110000;
assign LUT_4[46253] = 32'b11111111111111111011110111101000;
assign LUT_4[46254] = 32'b00000000000000000010000110010100;
assign LUT_4[46255] = 32'b11111111111111111011010010001100;
assign LUT_4[46256] = 32'b00000000000000001010010000101101;
assign LUT_4[46257] = 32'b00000000000000000011011100100101;
assign LUT_4[46258] = 32'b00000000000000001001101011010001;
assign LUT_4[46259] = 32'b00000000000000000010110111001001;
assign LUT_4[46260] = 32'b00000000000000000111010001001001;
assign LUT_4[46261] = 32'b00000000000000000000011101000001;
assign LUT_4[46262] = 32'b00000000000000000110101011101101;
assign LUT_4[46263] = 32'b11111111111111111111110111100101;
assign LUT_4[46264] = 32'b00000000000000000011011101000010;
assign LUT_4[46265] = 32'b11111111111111111100101000111010;
assign LUT_4[46266] = 32'b00000000000000000010110111100110;
assign LUT_4[46267] = 32'b11111111111111111100000011011110;
assign LUT_4[46268] = 32'b00000000000000000000011101011110;
assign LUT_4[46269] = 32'b11111111111111111001101001010110;
assign LUT_4[46270] = 32'b11111111111111111111111000000010;
assign LUT_4[46271] = 32'b11111111111111111001000011111010;
assign LUT_4[46272] = 32'b00000000000000001111011011001100;
assign LUT_4[46273] = 32'b00000000000000001000100111000100;
assign LUT_4[46274] = 32'b00000000000000001110110101110000;
assign LUT_4[46275] = 32'b00000000000000001000000001101000;
assign LUT_4[46276] = 32'b00000000000000001100011011101000;
assign LUT_4[46277] = 32'b00000000000000000101100111100000;
assign LUT_4[46278] = 32'b00000000000000001011110110001100;
assign LUT_4[46279] = 32'b00000000000000000101000010000100;
assign LUT_4[46280] = 32'b00000000000000001000100111100001;
assign LUT_4[46281] = 32'b00000000000000000001110011011001;
assign LUT_4[46282] = 32'b00000000000000001000000010000101;
assign LUT_4[46283] = 32'b00000000000000000001001101111101;
assign LUT_4[46284] = 32'b00000000000000000101100111111101;
assign LUT_4[46285] = 32'b11111111111111111110110011110101;
assign LUT_4[46286] = 32'b00000000000000000101000010100001;
assign LUT_4[46287] = 32'b11111111111111111110001110011001;
assign LUT_4[46288] = 32'b00000000000000001101001100111010;
assign LUT_4[46289] = 32'b00000000000000000110011000110010;
assign LUT_4[46290] = 32'b00000000000000001100100111011110;
assign LUT_4[46291] = 32'b00000000000000000101110011010110;
assign LUT_4[46292] = 32'b00000000000000001010001101010110;
assign LUT_4[46293] = 32'b00000000000000000011011001001110;
assign LUT_4[46294] = 32'b00000000000000001001100111111010;
assign LUT_4[46295] = 32'b00000000000000000010110011110010;
assign LUT_4[46296] = 32'b00000000000000000110011001001111;
assign LUT_4[46297] = 32'b11111111111111111111100101000111;
assign LUT_4[46298] = 32'b00000000000000000101110011110011;
assign LUT_4[46299] = 32'b11111111111111111110111111101011;
assign LUT_4[46300] = 32'b00000000000000000011011001101011;
assign LUT_4[46301] = 32'b11111111111111111100100101100011;
assign LUT_4[46302] = 32'b00000000000000000010110100001111;
assign LUT_4[46303] = 32'b11111111111111111100000000000111;
assign LUT_4[46304] = 32'b00000000000000001101110110010011;
assign LUT_4[46305] = 32'b00000000000000000111000010001011;
assign LUT_4[46306] = 32'b00000000000000001101010000110111;
assign LUT_4[46307] = 32'b00000000000000000110011100101111;
assign LUT_4[46308] = 32'b00000000000000001010110110101111;
assign LUT_4[46309] = 32'b00000000000000000100000010100111;
assign LUT_4[46310] = 32'b00000000000000001010010001010011;
assign LUT_4[46311] = 32'b00000000000000000011011101001011;
assign LUT_4[46312] = 32'b00000000000000000111000010101000;
assign LUT_4[46313] = 32'b00000000000000000000001110100000;
assign LUT_4[46314] = 32'b00000000000000000110011101001100;
assign LUT_4[46315] = 32'b11111111111111111111101001000100;
assign LUT_4[46316] = 32'b00000000000000000100000011000100;
assign LUT_4[46317] = 32'b11111111111111111101001110111100;
assign LUT_4[46318] = 32'b00000000000000000011011101101000;
assign LUT_4[46319] = 32'b11111111111111111100101001100000;
assign LUT_4[46320] = 32'b00000000000000001011101000000001;
assign LUT_4[46321] = 32'b00000000000000000100110011111001;
assign LUT_4[46322] = 32'b00000000000000001011000010100101;
assign LUT_4[46323] = 32'b00000000000000000100001110011101;
assign LUT_4[46324] = 32'b00000000000000001000101000011101;
assign LUT_4[46325] = 32'b00000000000000000001110100010101;
assign LUT_4[46326] = 32'b00000000000000001000000011000001;
assign LUT_4[46327] = 32'b00000000000000000001001110111001;
assign LUT_4[46328] = 32'b00000000000000000100110100010110;
assign LUT_4[46329] = 32'b11111111111111111110000000001110;
assign LUT_4[46330] = 32'b00000000000000000100001110111010;
assign LUT_4[46331] = 32'b11111111111111111101011010110010;
assign LUT_4[46332] = 32'b00000000000000000001110100110010;
assign LUT_4[46333] = 32'b11111111111111111011000000101010;
assign LUT_4[46334] = 32'b00000000000000000001001111010110;
assign LUT_4[46335] = 32'b11111111111111111010011011001110;
assign LUT_4[46336] = 32'b00000000000000010000011001010011;
assign LUT_4[46337] = 32'b00000000000000001001100101001011;
assign LUT_4[46338] = 32'b00000000000000001111110011110111;
assign LUT_4[46339] = 32'b00000000000000001000111111101111;
assign LUT_4[46340] = 32'b00000000000000001101011001101111;
assign LUT_4[46341] = 32'b00000000000000000110100101100111;
assign LUT_4[46342] = 32'b00000000000000001100110100010011;
assign LUT_4[46343] = 32'b00000000000000000110000000001011;
assign LUT_4[46344] = 32'b00000000000000001001100101101000;
assign LUT_4[46345] = 32'b00000000000000000010110001100000;
assign LUT_4[46346] = 32'b00000000000000001001000000001100;
assign LUT_4[46347] = 32'b00000000000000000010001100000100;
assign LUT_4[46348] = 32'b00000000000000000110100110000100;
assign LUT_4[46349] = 32'b11111111111111111111110001111100;
assign LUT_4[46350] = 32'b00000000000000000110000000101000;
assign LUT_4[46351] = 32'b11111111111111111111001100100000;
assign LUT_4[46352] = 32'b00000000000000001110001011000001;
assign LUT_4[46353] = 32'b00000000000000000111010110111001;
assign LUT_4[46354] = 32'b00000000000000001101100101100101;
assign LUT_4[46355] = 32'b00000000000000000110110001011101;
assign LUT_4[46356] = 32'b00000000000000001011001011011101;
assign LUT_4[46357] = 32'b00000000000000000100010111010101;
assign LUT_4[46358] = 32'b00000000000000001010100110000001;
assign LUT_4[46359] = 32'b00000000000000000011110001111001;
assign LUT_4[46360] = 32'b00000000000000000111010111010110;
assign LUT_4[46361] = 32'b00000000000000000000100011001110;
assign LUT_4[46362] = 32'b00000000000000000110110001111010;
assign LUT_4[46363] = 32'b11111111111111111111111101110010;
assign LUT_4[46364] = 32'b00000000000000000100010111110010;
assign LUT_4[46365] = 32'b11111111111111111101100011101010;
assign LUT_4[46366] = 32'b00000000000000000011110010010110;
assign LUT_4[46367] = 32'b11111111111111111100111110001110;
assign LUT_4[46368] = 32'b00000000000000001110110100011010;
assign LUT_4[46369] = 32'b00000000000000001000000000010010;
assign LUT_4[46370] = 32'b00000000000000001110001110111110;
assign LUT_4[46371] = 32'b00000000000000000111011010110110;
assign LUT_4[46372] = 32'b00000000000000001011110100110110;
assign LUT_4[46373] = 32'b00000000000000000101000000101110;
assign LUT_4[46374] = 32'b00000000000000001011001111011010;
assign LUT_4[46375] = 32'b00000000000000000100011011010010;
assign LUT_4[46376] = 32'b00000000000000001000000000101111;
assign LUT_4[46377] = 32'b00000000000000000001001100100111;
assign LUT_4[46378] = 32'b00000000000000000111011011010011;
assign LUT_4[46379] = 32'b00000000000000000000100111001011;
assign LUT_4[46380] = 32'b00000000000000000101000001001011;
assign LUT_4[46381] = 32'b11111111111111111110001101000011;
assign LUT_4[46382] = 32'b00000000000000000100011011101111;
assign LUT_4[46383] = 32'b11111111111111111101100111100111;
assign LUT_4[46384] = 32'b00000000000000001100100110001000;
assign LUT_4[46385] = 32'b00000000000000000101110010000000;
assign LUT_4[46386] = 32'b00000000000000001100000000101100;
assign LUT_4[46387] = 32'b00000000000000000101001100100100;
assign LUT_4[46388] = 32'b00000000000000001001100110100100;
assign LUT_4[46389] = 32'b00000000000000000010110010011100;
assign LUT_4[46390] = 32'b00000000000000001001000001001000;
assign LUT_4[46391] = 32'b00000000000000000010001101000000;
assign LUT_4[46392] = 32'b00000000000000000101110010011101;
assign LUT_4[46393] = 32'b11111111111111111110111110010101;
assign LUT_4[46394] = 32'b00000000000000000101001101000001;
assign LUT_4[46395] = 32'b11111111111111111110011000111001;
assign LUT_4[46396] = 32'b00000000000000000010110010111001;
assign LUT_4[46397] = 32'b11111111111111111011111110110001;
assign LUT_4[46398] = 32'b00000000000000000010001101011101;
assign LUT_4[46399] = 32'b11111111111111111011011001010101;
assign LUT_4[46400] = 32'b00000000000000010001110000100111;
assign LUT_4[46401] = 32'b00000000000000001010111100011111;
assign LUT_4[46402] = 32'b00000000000000010001001011001011;
assign LUT_4[46403] = 32'b00000000000000001010010111000011;
assign LUT_4[46404] = 32'b00000000000000001110110001000011;
assign LUT_4[46405] = 32'b00000000000000000111111100111011;
assign LUT_4[46406] = 32'b00000000000000001110001011100111;
assign LUT_4[46407] = 32'b00000000000000000111010111011111;
assign LUT_4[46408] = 32'b00000000000000001010111100111100;
assign LUT_4[46409] = 32'b00000000000000000100001000110100;
assign LUT_4[46410] = 32'b00000000000000001010010111100000;
assign LUT_4[46411] = 32'b00000000000000000011100011011000;
assign LUT_4[46412] = 32'b00000000000000000111111101011000;
assign LUT_4[46413] = 32'b00000000000000000001001001010000;
assign LUT_4[46414] = 32'b00000000000000000111010111111100;
assign LUT_4[46415] = 32'b00000000000000000000100011110100;
assign LUT_4[46416] = 32'b00000000000000001111100010010101;
assign LUT_4[46417] = 32'b00000000000000001000101110001101;
assign LUT_4[46418] = 32'b00000000000000001110111100111001;
assign LUT_4[46419] = 32'b00000000000000001000001000110001;
assign LUT_4[46420] = 32'b00000000000000001100100010110001;
assign LUT_4[46421] = 32'b00000000000000000101101110101001;
assign LUT_4[46422] = 32'b00000000000000001011111101010101;
assign LUT_4[46423] = 32'b00000000000000000101001001001101;
assign LUT_4[46424] = 32'b00000000000000001000101110101010;
assign LUT_4[46425] = 32'b00000000000000000001111010100010;
assign LUT_4[46426] = 32'b00000000000000001000001001001110;
assign LUT_4[46427] = 32'b00000000000000000001010101000110;
assign LUT_4[46428] = 32'b00000000000000000101101111000110;
assign LUT_4[46429] = 32'b11111111111111111110111010111110;
assign LUT_4[46430] = 32'b00000000000000000101001001101010;
assign LUT_4[46431] = 32'b11111111111111111110010101100010;
assign LUT_4[46432] = 32'b00000000000000010000001011101110;
assign LUT_4[46433] = 32'b00000000000000001001010111100110;
assign LUT_4[46434] = 32'b00000000000000001111100110010010;
assign LUT_4[46435] = 32'b00000000000000001000110010001010;
assign LUT_4[46436] = 32'b00000000000000001101001100001010;
assign LUT_4[46437] = 32'b00000000000000000110011000000010;
assign LUT_4[46438] = 32'b00000000000000001100100110101110;
assign LUT_4[46439] = 32'b00000000000000000101110010100110;
assign LUT_4[46440] = 32'b00000000000000001001011000000011;
assign LUT_4[46441] = 32'b00000000000000000010100011111011;
assign LUT_4[46442] = 32'b00000000000000001000110010100111;
assign LUT_4[46443] = 32'b00000000000000000001111110011111;
assign LUT_4[46444] = 32'b00000000000000000110011000011111;
assign LUT_4[46445] = 32'b11111111111111111111100100010111;
assign LUT_4[46446] = 32'b00000000000000000101110011000011;
assign LUT_4[46447] = 32'b11111111111111111110111110111011;
assign LUT_4[46448] = 32'b00000000000000001101111101011100;
assign LUT_4[46449] = 32'b00000000000000000111001001010100;
assign LUT_4[46450] = 32'b00000000000000001101011000000000;
assign LUT_4[46451] = 32'b00000000000000000110100011111000;
assign LUT_4[46452] = 32'b00000000000000001010111101111000;
assign LUT_4[46453] = 32'b00000000000000000100001001110000;
assign LUT_4[46454] = 32'b00000000000000001010011000011100;
assign LUT_4[46455] = 32'b00000000000000000011100100010100;
assign LUT_4[46456] = 32'b00000000000000000111001001110001;
assign LUT_4[46457] = 32'b00000000000000000000010101101001;
assign LUT_4[46458] = 32'b00000000000000000110100100010101;
assign LUT_4[46459] = 32'b11111111111111111111110000001101;
assign LUT_4[46460] = 32'b00000000000000000100001010001101;
assign LUT_4[46461] = 32'b11111111111111111101010110000101;
assign LUT_4[46462] = 32'b00000000000000000011100100110001;
assign LUT_4[46463] = 32'b11111111111111111100110000101001;
assign LUT_4[46464] = 32'b00000000000000010010111111011011;
assign LUT_4[46465] = 32'b00000000000000001100001011010011;
assign LUT_4[46466] = 32'b00000000000000010010011001111111;
assign LUT_4[46467] = 32'b00000000000000001011100101110111;
assign LUT_4[46468] = 32'b00000000000000001111111111110111;
assign LUT_4[46469] = 32'b00000000000000001001001011101111;
assign LUT_4[46470] = 32'b00000000000000001111011010011011;
assign LUT_4[46471] = 32'b00000000000000001000100110010011;
assign LUT_4[46472] = 32'b00000000000000001100001011110000;
assign LUT_4[46473] = 32'b00000000000000000101010111101000;
assign LUT_4[46474] = 32'b00000000000000001011100110010100;
assign LUT_4[46475] = 32'b00000000000000000100110010001100;
assign LUT_4[46476] = 32'b00000000000000001001001100001100;
assign LUT_4[46477] = 32'b00000000000000000010011000000100;
assign LUT_4[46478] = 32'b00000000000000001000100110110000;
assign LUT_4[46479] = 32'b00000000000000000001110010101000;
assign LUT_4[46480] = 32'b00000000000000010000110001001001;
assign LUT_4[46481] = 32'b00000000000000001001111101000001;
assign LUT_4[46482] = 32'b00000000000000010000001011101101;
assign LUT_4[46483] = 32'b00000000000000001001010111100101;
assign LUT_4[46484] = 32'b00000000000000001101110001100101;
assign LUT_4[46485] = 32'b00000000000000000110111101011101;
assign LUT_4[46486] = 32'b00000000000000001101001100001001;
assign LUT_4[46487] = 32'b00000000000000000110011000000001;
assign LUT_4[46488] = 32'b00000000000000001001111101011110;
assign LUT_4[46489] = 32'b00000000000000000011001001010110;
assign LUT_4[46490] = 32'b00000000000000001001011000000010;
assign LUT_4[46491] = 32'b00000000000000000010100011111010;
assign LUT_4[46492] = 32'b00000000000000000110111101111010;
assign LUT_4[46493] = 32'b00000000000000000000001001110010;
assign LUT_4[46494] = 32'b00000000000000000110011000011110;
assign LUT_4[46495] = 32'b11111111111111111111100100010110;
assign LUT_4[46496] = 32'b00000000000000010001011010100010;
assign LUT_4[46497] = 32'b00000000000000001010100110011010;
assign LUT_4[46498] = 32'b00000000000000010000110101000110;
assign LUT_4[46499] = 32'b00000000000000001010000000111110;
assign LUT_4[46500] = 32'b00000000000000001110011010111110;
assign LUT_4[46501] = 32'b00000000000000000111100110110110;
assign LUT_4[46502] = 32'b00000000000000001101110101100010;
assign LUT_4[46503] = 32'b00000000000000000111000001011010;
assign LUT_4[46504] = 32'b00000000000000001010100110110111;
assign LUT_4[46505] = 32'b00000000000000000011110010101111;
assign LUT_4[46506] = 32'b00000000000000001010000001011011;
assign LUT_4[46507] = 32'b00000000000000000011001101010011;
assign LUT_4[46508] = 32'b00000000000000000111100111010011;
assign LUT_4[46509] = 32'b00000000000000000000110011001011;
assign LUT_4[46510] = 32'b00000000000000000111000001110111;
assign LUT_4[46511] = 32'b00000000000000000000001101101111;
assign LUT_4[46512] = 32'b00000000000000001111001100010000;
assign LUT_4[46513] = 32'b00000000000000001000011000001000;
assign LUT_4[46514] = 32'b00000000000000001110100110110100;
assign LUT_4[46515] = 32'b00000000000000000111110010101100;
assign LUT_4[46516] = 32'b00000000000000001100001100101100;
assign LUT_4[46517] = 32'b00000000000000000101011000100100;
assign LUT_4[46518] = 32'b00000000000000001011100111010000;
assign LUT_4[46519] = 32'b00000000000000000100110011001000;
assign LUT_4[46520] = 32'b00000000000000001000011000100101;
assign LUT_4[46521] = 32'b00000000000000000001100100011101;
assign LUT_4[46522] = 32'b00000000000000000111110011001001;
assign LUT_4[46523] = 32'b00000000000000000000111111000001;
assign LUT_4[46524] = 32'b00000000000000000101011001000001;
assign LUT_4[46525] = 32'b11111111111111111110100100111001;
assign LUT_4[46526] = 32'b00000000000000000100110011100101;
assign LUT_4[46527] = 32'b11111111111111111101111111011101;
assign LUT_4[46528] = 32'b00000000000000010100010110101111;
assign LUT_4[46529] = 32'b00000000000000001101100010100111;
assign LUT_4[46530] = 32'b00000000000000010011110001010011;
assign LUT_4[46531] = 32'b00000000000000001100111101001011;
assign LUT_4[46532] = 32'b00000000000000010001010111001011;
assign LUT_4[46533] = 32'b00000000000000001010100011000011;
assign LUT_4[46534] = 32'b00000000000000010000110001101111;
assign LUT_4[46535] = 32'b00000000000000001001111101100111;
assign LUT_4[46536] = 32'b00000000000000001101100011000100;
assign LUT_4[46537] = 32'b00000000000000000110101110111100;
assign LUT_4[46538] = 32'b00000000000000001100111101101000;
assign LUT_4[46539] = 32'b00000000000000000110001001100000;
assign LUT_4[46540] = 32'b00000000000000001010100011100000;
assign LUT_4[46541] = 32'b00000000000000000011101111011000;
assign LUT_4[46542] = 32'b00000000000000001001111110000100;
assign LUT_4[46543] = 32'b00000000000000000011001001111100;
assign LUT_4[46544] = 32'b00000000000000010010001000011101;
assign LUT_4[46545] = 32'b00000000000000001011010100010101;
assign LUT_4[46546] = 32'b00000000000000010001100011000001;
assign LUT_4[46547] = 32'b00000000000000001010101110111001;
assign LUT_4[46548] = 32'b00000000000000001111001000111001;
assign LUT_4[46549] = 32'b00000000000000001000010100110001;
assign LUT_4[46550] = 32'b00000000000000001110100011011101;
assign LUT_4[46551] = 32'b00000000000000000111101111010101;
assign LUT_4[46552] = 32'b00000000000000001011010100110010;
assign LUT_4[46553] = 32'b00000000000000000100100000101010;
assign LUT_4[46554] = 32'b00000000000000001010101111010110;
assign LUT_4[46555] = 32'b00000000000000000011111011001110;
assign LUT_4[46556] = 32'b00000000000000001000010101001110;
assign LUT_4[46557] = 32'b00000000000000000001100001000110;
assign LUT_4[46558] = 32'b00000000000000000111101111110010;
assign LUT_4[46559] = 32'b00000000000000000000111011101010;
assign LUT_4[46560] = 32'b00000000000000010010110001110110;
assign LUT_4[46561] = 32'b00000000000000001011111101101110;
assign LUT_4[46562] = 32'b00000000000000010010001100011010;
assign LUT_4[46563] = 32'b00000000000000001011011000010010;
assign LUT_4[46564] = 32'b00000000000000001111110010010010;
assign LUT_4[46565] = 32'b00000000000000001000111110001010;
assign LUT_4[46566] = 32'b00000000000000001111001100110110;
assign LUT_4[46567] = 32'b00000000000000001000011000101110;
assign LUT_4[46568] = 32'b00000000000000001011111110001011;
assign LUT_4[46569] = 32'b00000000000000000101001010000011;
assign LUT_4[46570] = 32'b00000000000000001011011000101111;
assign LUT_4[46571] = 32'b00000000000000000100100100100111;
assign LUT_4[46572] = 32'b00000000000000001000111110100111;
assign LUT_4[46573] = 32'b00000000000000000010001010011111;
assign LUT_4[46574] = 32'b00000000000000001000011001001011;
assign LUT_4[46575] = 32'b00000000000000000001100101000011;
assign LUT_4[46576] = 32'b00000000000000010000100011100100;
assign LUT_4[46577] = 32'b00000000000000001001101111011100;
assign LUT_4[46578] = 32'b00000000000000001111111110001000;
assign LUT_4[46579] = 32'b00000000000000001001001010000000;
assign LUT_4[46580] = 32'b00000000000000001101100100000000;
assign LUT_4[46581] = 32'b00000000000000000110101111111000;
assign LUT_4[46582] = 32'b00000000000000001100111110100100;
assign LUT_4[46583] = 32'b00000000000000000110001010011100;
assign LUT_4[46584] = 32'b00000000000000001001101111111001;
assign LUT_4[46585] = 32'b00000000000000000010111011110001;
assign LUT_4[46586] = 32'b00000000000000001001001010011101;
assign LUT_4[46587] = 32'b00000000000000000010010110010101;
assign LUT_4[46588] = 32'b00000000000000000110110000010101;
assign LUT_4[46589] = 32'b11111111111111111111111100001101;
assign LUT_4[46590] = 32'b00000000000000000110001010111001;
assign LUT_4[46591] = 32'b11111111111111111111010110110001;
assign LUT_4[46592] = 32'b00000000000000001010100001111000;
assign LUT_4[46593] = 32'b00000000000000000011101101110000;
assign LUT_4[46594] = 32'b00000000000000001001111100011100;
assign LUT_4[46595] = 32'b00000000000000000011001000010100;
assign LUT_4[46596] = 32'b00000000000000000111100010010100;
assign LUT_4[46597] = 32'b00000000000000000000101110001100;
assign LUT_4[46598] = 32'b00000000000000000110111100111000;
assign LUT_4[46599] = 32'b00000000000000000000001000110000;
assign LUT_4[46600] = 32'b00000000000000000011101110001101;
assign LUT_4[46601] = 32'b11111111111111111100111010000101;
assign LUT_4[46602] = 32'b00000000000000000011001000110001;
assign LUT_4[46603] = 32'b11111111111111111100010100101001;
assign LUT_4[46604] = 32'b00000000000000000000101110101001;
assign LUT_4[46605] = 32'b11111111111111111001111010100001;
assign LUT_4[46606] = 32'b00000000000000000000001001001101;
assign LUT_4[46607] = 32'b11111111111111111001010101000101;
assign LUT_4[46608] = 32'b00000000000000001000010011100110;
assign LUT_4[46609] = 32'b00000000000000000001011111011110;
assign LUT_4[46610] = 32'b00000000000000000111101110001010;
assign LUT_4[46611] = 32'b00000000000000000000111010000010;
assign LUT_4[46612] = 32'b00000000000000000101010100000010;
assign LUT_4[46613] = 32'b11111111111111111110011111111010;
assign LUT_4[46614] = 32'b00000000000000000100101110100110;
assign LUT_4[46615] = 32'b11111111111111111101111010011110;
assign LUT_4[46616] = 32'b00000000000000000001011111111011;
assign LUT_4[46617] = 32'b11111111111111111010101011110011;
assign LUT_4[46618] = 32'b00000000000000000000111010011111;
assign LUT_4[46619] = 32'b11111111111111111010000110010111;
assign LUT_4[46620] = 32'b11111111111111111110100000010111;
assign LUT_4[46621] = 32'b11111111111111110111101100001111;
assign LUT_4[46622] = 32'b11111111111111111101111010111011;
assign LUT_4[46623] = 32'b11111111111111110111000110110011;
assign LUT_4[46624] = 32'b00000000000000001000111100111111;
assign LUT_4[46625] = 32'b00000000000000000010001000110111;
assign LUT_4[46626] = 32'b00000000000000001000010111100011;
assign LUT_4[46627] = 32'b00000000000000000001100011011011;
assign LUT_4[46628] = 32'b00000000000000000101111101011011;
assign LUT_4[46629] = 32'b11111111111111111111001001010011;
assign LUT_4[46630] = 32'b00000000000000000101010111111111;
assign LUT_4[46631] = 32'b11111111111111111110100011110111;
assign LUT_4[46632] = 32'b00000000000000000010001001010100;
assign LUT_4[46633] = 32'b11111111111111111011010101001100;
assign LUT_4[46634] = 32'b00000000000000000001100011111000;
assign LUT_4[46635] = 32'b11111111111111111010101111110000;
assign LUT_4[46636] = 32'b11111111111111111111001001110000;
assign LUT_4[46637] = 32'b11111111111111111000010101101000;
assign LUT_4[46638] = 32'b11111111111111111110100100010100;
assign LUT_4[46639] = 32'b11111111111111110111110000001100;
assign LUT_4[46640] = 32'b00000000000000000110101110101101;
assign LUT_4[46641] = 32'b11111111111111111111111010100101;
assign LUT_4[46642] = 32'b00000000000000000110001001010001;
assign LUT_4[46643] = 32'b11111111111111111111010101001001;
assign LUT_4[46644] = 32'b00000000000000000011101111001001;
assign LUT_4[46645] = 32'b11111111111111111100111011000001;
assign LUT_4[46646] = 32'b00000000000000000011001001101101;
assign LUT_4[46647] = 32'b11111111111111111100010101100101;
assign LUT_4[46648] = 32'b11111111111111111111111011000010;
assign LUT_4[46649] = 32'b11111111111111111001000110111010;
assign LUT_4[46650] = 32'b11111111111111111111010101100110;
assign LUT_4[46651] = 32'b11111111111111111000100001011110;
assign LUT_4[46652] = 32'b11111111111111111100111011011110;
assign LUT_4[46653] = 32'b11111111111111110110000111010110;
assign LUT_4[46654] = 32'b11111111111111111100010110000010;
assign LUT_4[46655] = 32'b11111111111111110101100001111010;
assign LUT_4[46656] = 32'b00000000000000001011111001001100;
assign LUT_4[46657] = 32'b00000000000000000101000101000100;
assign LUT_4[46658] = 32'b00000000000000001011010011110000;
assign LUT_4[46659] = 32'b00000000000000000100011111101000;
assign LUT_4[46660] = 32'b00000000000000001000111001101000;
assign LUT_4[46661] = 32'b00000000000000000010000101100000;
assign LUT_4[46662] = 32'b00000000000000001000010100001100;
assign LUT_4[46663] = 32'b00000000000000000001100000000100;
assign LUT_4[46664] = 32'b00000000000000000101000101100001;
assign LUT_4[46665] = 32'b11111111111111111110010001011001;
assign LUT_4[46666] = 32'b00000000000000000100100000000101;
assign LUT_4[46667] = 32'b11111111111111111101101011111101;
assign LUT_4[46668] = 32'b00000000000000000010000101111101;
assign LUT_4[46669] = 32'b11111111111111111011010001110101;
assign LUT_4[46670] = 32'b00000000000000000001100000100001;
assign LUT_4[46671] = 32'b11111111111111111010101100011001;
assign LUT_4[46672] = 32'b00000000000000001001101010111010;
assign LUT_4[46673] = 32'b00000000000000000010110110110010;
assign LUT_4[46674] = 32'b00000000000000001001000101011110;
assign LUT_4[46675] = 32'b00000000000000000010010001010110;
assign LUT_4[46676] = 32'b00000000000000000110101011010110;
assign LUT_4[46677] = 32'b11111111111111111111110111001110;
assign LUT_4[46678] = 32'b00000000000000000110000101111010;
assign LUT_4[46679] = 32'b11111111111111111111010001110010;
assign LUT_4[46680] = 32'b00000000000000000010110111001111;
assign LUT_4[46681] = 32'b11111111111111111100000011000111;
assign LUT_4[46682] = 32'b00000000000000000010010001110011;
assign LUT_4[46683] = 32'b11111111111111111011011101101011;
assign LUT_4[46684] = 32'b11111111111111111111110111101011;
assign LUT_4[46685] = 32'b11111111111111111001000011100011;
assign LUT_4[46686] = 32'b11111111111111111111010010001111;
assign LUT_4[46687] = 32'b11111111111111111000011110000111;
assign LUT_4[46688] = 32'b00000000000000001010010100010011;
assign LUT_4[46689] = 32'b00000000000000000011100000001011;
assign LUT_4[46690] = 32'b00000000000000001001101110110111;
assign LUT_4[46691] = 32'b00000000000000000010111010101111;
assign LUT_4[46692] = 32'b00000000000000000111010100101111;
assign LUT_4[46693] = 32'b00000000000000000000100000100111;
assign LUT_4[46694] = 32'b00000000000000000110101111010011;
assign LUT_4[46695] = 32'b11111111111111111111111011001011;
assign LUT_4[46696] = 32'b00000000000000000011100000101000;
assign LUT_4[46697] = 32'b11111111111111111100101100100000;
assign LUT_4[46698] = 32'b00000000000000000010111011001100;
assign LUT_4[46699] = 32'b11111111111111111100000111000100;
assign LUT_4[46700] = 32'b00000000000000000000100001000100;
assign LUT_4[46701] = 32'b11111111111111111001101100111100;
assign LUT_4[46702] = 32'b11111111111111111111111011101000;
assign LUT_4[46703] = 32'b11111111111111111001000111100000;
assign LUT_4[46704] = 32'b00000000000000001000000110000001;
assign LUT_4[46705] = 32'b00000000000000000001010001111001;
assign LUT_4[46706] = 32'b00000000000000000111100000100101;
assign LUT_4[46707] = 32'b00000000000000000000101100011101;
assign LUT_4[46708] = 32'b00000000000000000101000110011101;
assign LUT_4[46709] = 32'b11111111111111111110010010010101;
assign LUT_4[46710] = 32'b00000000000000000100100001000001;
assign LUT_4[46711] = 32'b11111111111111111101101100111001;
assign LUT_4[46712] = 32'b00000000000000000001010010010110;
assign LUT_4[46713] = 32'b11111111111111111010011110001110;
assign LUT_4[46714] = 32'b00000000000000000000101100111010;
assign LUT_4[46715] = 32'b11111111111111111001111000110010;
assign LUT_4[46716] = 32'b11111111111111111110010010110010;
assign LUT_4[46717] = 32'b11111111111111110111011110101010;
assign LUT_4[46718] = 32'b11111111111111111101101101010110;
assign LUT_4[46719] = 32'b11111111111111110110111001001110;
assign LUT_4[46720] = 32'b00000000000000001101001000000000;
assign LUT_4[46721] = 32'b00000000000000000110010011111000;
assign LUT_4[46722] = 32'b00000000000000001100100010100100;
assign LUT_4[46723] = 32'b00000000000000000101101110011100;
assign LUT_4[46724] = 32'b00000000000000001010001000011100;
assign LUT_4[46725] = 32'b00000000000000000011010100010100;
assign LUT_4[46726] = 32'b00000000000000001001100011000000;
assign LUT_4[46727] = 32'b00000000000000000010101110111000;
assign LUT_4[46728] = 32'b00000000000000000110010100010101;
assign LUT_4[46729] = 32'b11111111111111111111100000001101;
assign LUT_4[46730] = 32'b00000000000000000101101110111001;
assign LUT_4[46731] = 32'b11111111111111111110111010110001;
assign LUT_4[46732] = 32'b00000000000000000011010100110001;
assign LUT_4[46733] = 32'b11111111111111111100100000101001;
assign LUT_4[46734] = 32'b00000000000000000010101111010101;
assign LUT_4[46735] = 32'b11111111111111111011111011001101;
assign LUT_4[46736] = 32'b00000000000000001010111001101110;
assign LUT_4[46737] = 32'b00000000000000000100000101100110;
assign LUT_4[46738] = 32'b00000000000000001010010100010010;
assign LUT_4[46739] = 32'b00000000000000000011100000001010;
assign LUT_4[46740] = 32'b00000000000000000111111010001010;
assign LUT_4[46741] = 32'b00000000000000000001000110000010;
assign LUT_4[46742] = 32'b00000000000000000111010100101110;
assign LUT_4[46743] = 32'b00000000000000000000100000100110;
assign LUT_4[46744] = 32'b00000000000000000100000110000011;
assign LUT_4[46745] = 32'b11111111111111111101010001111011;
assign LUT_4[46746] = 32'b00000000000000000011100000100111;
assign LUT_4[46747] = 32'b11111111111111111100101100011111;
assign LUT_4[46748] = 32'b00000000000000000001000110011111;
assign LUT_4[46749] = 32'b11111111111111111010010010010111;
assign LUT_4[46750] = 32'b00000000000000000000100001000011;
assign LUT_4[46751] = 32'b11111111111111111001101100111011;
assign LUT_4[46752] = 32'b00000000000000001011100011000111;
assign LUT_4[46753] = 32'b00000000000000000100101110111111;
assign LUT_4[46754] = 32'b00000000000000001010111101101011;
assign LUT_4[46755] = 32'b00000000000000000100001001100011;
assign LUT_4[46756] = 32'b00000000000000001000100011100011;
assign LUT_4[46757] = 32'b00000000000000000001101111011011;
assign LUT_4[46758] = 32'b00000000000000000111111110000111;
assign LUT_4[46759] = 32'b00000000000000000001001001111111;
assign LUT_4[46760] = 32'b00000000000000000100101111011100;
assign LUT_4[46761] = 32'b11111111111111111101111011010100;
assign LUT_4[46762] = 32'b00000000000000000100001010000000;
assign LUT_4[46763] = 32'b11111111111111111101010101111000;
assign LUT_4[46764] = 32'b00000000000000000001101111111000;
assign LUT_4[46765] = 32'b11111111111111111010111011110000;
assign LUT_4[46766] = 32'b00000000000000000001001010011100;
assign LUT_4[46767] = 32'b11111111111111111010010110010100;
assign LUT_4[46768] = 32'b00000000000000001001010100110101;
assign LUT_4[46769] = 32'b00000000000000000010100000101101;
assign LUT_4[46770] = 32'b00000000000000001000101111011001;
assign LUT_4[46771] = 32'b00000000000000000001111011010001;
assign LUT_4[46772] = 32'b00000000000000000110010101010001;
assign LUT_4[46773] = 32'b11111111111111111111100001001001;
assign LUT_4[46774] = 32'b00000000000000000101101111110101;
assign LUT_4[46775] = 32'b11111111111111111110111011101101;
assign LUT_4[46776] = 32'b00000000000000000010100001001010;
assign LUT_4[46777] = 32'b11111111111111111011101101000010;
assign LUT_4[46778] = 32'b00000000000000000001111011101110;
assign LUT_4[46779] = 32'b11111111111111111011000111100110;
assign LUT_4[46780] = 32'b11111111111111111111100001100110;
assign LUT_4[46781] = 32'b11111111111111111000101101011110;
assign LUT_4[46782] = 32'b11111111111111111110111100001010;
assign LUT_4[46783] = 32'b11111111111111111000001000000010;
assign LUT_4[46784] = 32'b00000000000000001110011111010100;
assign LUT_4[46785] = 32'b00000000000000000111101011001100;
assign LUT_4[46786] = 32'b00000000000000001101111001111000;
assign LUT_4[46787] = 32'b00000000000000000111000101110000;
assign LUT_4[46788] = 32'b00000000000000001011011111110000;
assign LUT_4[46789] = 32'b00000000000000000100101011101000;
assign LUT_4[46790] = 32'b00000000000000001010111010010100;
assign LUT_4[46791] = 32'b00000000000000000100000110001100;
assign LUT_4[46792] = 32'b00000000000000000111101011101001;
assign LUT_4[46793] = 32'b00000000000000000000110111100001;
assign LUT_4[46794] = 32'b00000000000000000111000110001101;
assign LUT_4[46795] = 32'b00000000000000000000010010000101;
assign LUT_4[46796] = 32'b00000000000000000100101100000101;
assign LUT_4[46797] = 32'b11111111111111111101110111111101;
assign LUT_4[46798] = 32'b00000000000000000100000110101001;
assign LUT_4[46799] = 32'b11111111111111111101010010100001;
assign LUT_4[46800] = 32'b00000000000000001100010001000010;
assign LUT_4[46801] = 32'b00000000000000000101011100111010;
assign LUT_4[46802] = 32'b00000000000000001011101011100110;
assign LUT_4[46803] = 32'b00000000000000000100110111011110;
assign LUT_4[46804] = 32'b00000000000000001001010001011110;
assign LUT_4[46805] = 32'b00000000000000000010011101010110;
assign LUT_4[46806] = 32'b00000000000000001000101100000010;
assign LUT_4[46807] = 32'b00000000000000000001110111111010;
assign LUT_4[46808] = 32'b00000000000000000101011101010111;
assign LUT_4[46809] = 32'b11111111111111111110101001001111;
assign LUT_4[46810] = 32'b00000000000000000100110111111011;
assign LUT_4[46811] = 32'b11111111111111111110000011110011;
assign LUT_4[46812] = 32'b00000000000000000010011101110011;
assign LUT_4[46813] = 32'b11111111111111111011101001101011;
assign LUT_4[46814] = 32'b00000000000000000001111000010111;
assign LUT_4[46815] = 32'b11111111111111111011000100001111;
assign LUT_4[46816] = 32'b00000000000000001100111010011011;
assign LUT_4[46817] = 32'b00000000000000000110000110010011;
assign LUT_4[46818] = 32'b00000000000000001100010100111111;
assign LUT_4[46819] = 32'b00000000000000000101100000110111;
assign LUT_4[46820] = 32'b00000000000000001001111010110111;
assign LUT_4[46821] = 32'b00000000000000000011000110101111;
assign LUT_4[46822] = 32'b00000000000000001001010101011011;
assign LUT_4[46823] = 32'b00000000000000000010100001010011;
assign LUT_4[46824] = 32'b00000000000000000110000110110000;
assign LUT_4[46825] = 32'b11111111111111111111010010101000;
assign LUT_4[46826] = 32'b00000000000000000101100001010100;
assign LUT_4[46827] = 32'b11111111111111111110101101001100;
assign LUT_4[46828] = 32'b00000000000000000011000111001100;
assign LUT_4[46829] = 32'b11111111111111111100010011000100;
assign LUT_4[46830] = 32'b00000000000000000010100001110000;
assign LUT_4[46831] = 32'b11111111111111111011101101101000;
assign LUT_4[46832] = 32'b00000000000000001010101100001001;
assign LUT_4[46833] = 32'b00000000000000000011111000000001;
assign LUT_4[46834] = 32'b00000000000000001010000110101101;
assign LUT_4[46835] = 32'b00000000000000000011010010100101;
assign LUT_4[46836] = 32'b00000000000000000111101100100101;
assign LUT_4[46837] = 32'b00000000000000000000111000011101;
assign LUT_4[46838] = 32'b00000000000000000111000111001001;
assign LUT_4[46839] = 32'b00000000000000000000010011000001;
assign LUT_4[46840] = 32'b00000000000000000011111000011110;
assign LUT_4[46841] = 32'b11111111111111111101000100010110;
assign LUT_4[46842] = 32'b00000000000000000011010011000010;
assign LUT_4[46843] = 32'b11111111111111111100011110111010;
assign LUT_4[46844] = 32'b00000000000000000000111000111010;
assign LUT_4[46845] = 32'b11111111111111111010000100110010;
assign LUT_4[46846] = 32'b00000000000000000000010011011110;
assign LUT_4[46847] = 32'b11111111111111111001011111010110;
assign LUT_4[46848] = 32'b00000000000000001111011101011011;
assign LUT_4[46849] = 32'b00000000000000001000101001010011;
assign LUT_4[46850] = 32'b00000000000000001110110111111111;
assign LUT_4[46851] = 32'b00000000000000001000000011110111;
assign LUT_4[46852] = 32'b00000000000000001100011101110111;
assign LUT_4[46853] = 32'b00000000000000000101101001101111;
assign LUT_4[46854] = 32'b00000000000000001011111000011011;
assign LUT_4[46855] = 32'b00000000000000000101000100010011;
assign LUT_4[46856] = 32'b00000000000000001000101001110000;
assign LUT_4[46857] = 32'b00000000000000000001110101101000;
assign LUT_4[46858] = 32'b00000000000000001000000100010100;
assign LUT_4[46859] = 32'b00000000000000000001010000001100;
assign LUT_4[46860] = 32'b00000000000000000101101010001100;
assign LUT_4[46861] = 32'b11111111111111111110110110000100;
assign LUT_4[46862] = 32'b00000000000000000101000100110000;
assign LUT_4[46863] = 32'b11111111111111111110010000101000;
assign LUT_4[46864] = 32'b00000000000000001101001111001001;
assign LUT_4[46865] = 32'b00000000000000000110011011000001;
assign LUT_4[46866] = 32'b00000000000000001100101001101101;
assign LUT_4[46867] = 32'b00000000000000000101110101100101;
assign LUT_4[46868] = 32'b00000000000000001010001111100101;
assign LUT_4[46869] = 32'b00000000000000000011011011011101;
assign LUT_4[46870] = 32'b00000000000000001001101010001001;
assign LUT_4[46871] = 32'b00000000000000000010110110000001;
assign LUT_4[46872] = 32'b00000000000000000110011011011110;
assign LUT_4[46873] = 32'b11111111111111111111100111010110;
assign LUT_4[46874] = 32'b00000000000000000101110110000010;
assign LUT_4[46875] = 32'b11111111111111111111000001111010;
assign LUT_4[46876] = 32'b00000000000000000011011011111010;
assign LUT_4[46877] = 32'b11111111111111111100100111110010;
assign LUT_4[46878] = 32'b00000000000000000010110110011110;
assign LUT_4[46879] = 32'b11111111111111111100000010010110;
assign LUT_4[46880] = 32'b00000000000000001101111000100010;
assign LUT_4[46881] = 32'b00000000000000000111000100011010;
assign LUT_4[46882] = 32'b00000000000000001101010011000110;
assign LUT_4[46883] = 32'b00000000000000000110011110111110;
assign LUT_4[46884] = 32'b00000000000000001010111000111110;
assign LUT_4[46885] = 32'b00000000000000000100000100110110;
assign LUT_4[46886] = 32'b00000000000000001010010011100010;
assign LUT_4[46887] = 32'b00000000000000000011011111011010;
assign LUT_4[46888] = 32'b00000000000000000111000100110111;
assign LUT_4[46889] = 32'b00000000000000000000010000101111;
assign LUT_4[46890] = 32'b00000000000000000110011111011011;
assign LUT_4[46891] = 32'b11111111111111111111101011010011;
assign LUT_4[46892] = 32'b00000000000000000100000101010011;
assign LUT_4[46893] = 32'b11111111111111111101010001001011;
assign LUT_4[46894] = 32'b00000000000000000011011111110111;
assign LUT_4[46895] = 32'b11111111111111111100101011101111;
assign LUT_4[46896] = 32'b00000000000000001011101010010000;
assign LUT_4[46897] = 32'b00000000000000000100110110001000;
assign LUT_4[46898] = 32'b00000000000000001011000100110100;
assign LUT_4[46899] = 32'b00000000000000000100010000101100;
assign LUT_4[46900] = 32'b00000000000000001000101010101100;
assign LUT_4[46901] = 32'b00000000000000000001110110100100;
assign LUT_4[46902] = 32'b00000000000000001000000101010000;
assign LUT_4[46903] = 32'b00000000000000000001010001001000;
assign LUT_4[46904] = 32'b00000000000000000100110110100101;
assign LUT_4[46905] = 32'b11111111111111111110000010011101;
assign LUT_4[46906] = 32'b00000000000000000100010001001001;
assign LUT_4[46907] = 32'b11111111111111111101011101000001;
assign LUT_4[46908] = 32'b00000000000000000001110111000001;
assign LUT_4[46909] = 32'b11111111111111111011000010111001;
assign LUT_4[46910] = 32'b00000000000000000001010001100101;
assign LUT_4[46911] = 32'b11111111111111111010011101011101;
assign LUT_4[46912] = 32'b00000000000000010000110100101111;
assign LUT_4[46913] = 32'b00000000000000001010000000100111;
assign LUT_4[46914] = 32'b00000000000000010000001111010011;
assign LUT_4[46915] = 32'b00000000000000001001011011001011;
assign LUT_4[46916] = 32'b00000000000000001101110101001011;
assign LUT_4[46917] = 32'b00000000000000000111000001000011;
assign LUT_4[46918] = 32'b00000000000000001101001111101111;
assign LUT_4[46919] = 32'b00000000000000000110011011100111;
assign LUT_4[46920] = 32'b00000000000000001010000001000100;
assign LUT_4[46921] = 32'b00000000000000000011001100111100;
assign LUT_4[46922] = 32'b00000000000000001001011011101000;
assign LUT_4[46923] = 32'b00000000000000000010100111100000;
assign LUT_4[46924] = 32'b00000000000000000111000001100000;
assign LUT_4[46925] = 32'b00000000000000000000001101011000;
assign LUT_4[46926] = 32'b00000000000000000110011100000100;
assign LUT_4[46927] = 32'b11111111111111111111100111111100;
assign LUT_4[46928] = 32'b00000000000000001110100110011101;
assign LUT_4[46929] = 32'b00000000000000000111110010010101;
assign LUT_4[46930] = 32'b00000000000000001110000001000001;
assign LUT_4[46931] = 32'b00000000000000000111001100111001;
assign LUT_4[46932] = 32'b00000000000000001011100110111001;
assign LUT_4[46933] = 32'b00000000000000000100110010110001;
assign LUT_4[46934] = 32'b00000000000000001011000001011101;
assign LUT_4[46935] = 32'b00000000000000000100001101010101;
assign LUT_4[46936] = 32'b00000000000000000111110010110010;
assign LUT_4[46937] = 32'b00000000000000000000111110101010;
assign LUT_4[46938] = 32'b00000000000000000111001101010110;
assign LUT_4[46939] = 32'b00000000000000000000011001001110;
assign LUT_4[46940] = 32'b00000000000000000100110011001110;
assign LUT_4[46941] = 32'b11111111111111111101111111000110;
assign LUT_4[46942] = 32'b00000000000000000100001101110010;
assign LUT_4[46943] = 32'b11111111111111111101011001101010;
assign LUT_4[46944] = 32'b00000000000000001111001111110110;
assign LUT_4[46945] = 32'b00000000000000001000011011101110;
assign LUT_4[46946] = 32'b00000000000000001110101010011010;
assign LUT_4[46947] = 32'b00000000000000000111110110010010;
assign LUT_4[46948] = 32'b00000000000000001100010000010010;
assign LUT_4[46949] = 32'b00000000000000000101011100001010;
assign LUT_4[46950] = 32'b00000000000000001011101010110110;
assign LUT_4[46951] = 32'b00000000000000000100110110101110;
assign LUT_4[46952] = 32'b00000000000000001000011100001011;
assign LUT_4[46953] = 32'b00000000000000000001101000000011;
assign LUT_4[46954] = 32'b00000000000000000111110110101111;
assign LUT_4[46955] = 32'b00000000000000000001000010100111;
assign LUT_4[46956] = 32'b00000000000000000101011100100111;
assign LUT_4[46957] = 32'b11111111111111111110101000011111;
assign LUT_4[46958] = 32'b00000000000000000100110111001011;
assign LUT_4[46959] = 32'b11111111111111111110000011000011;
assign LUT_4[46960] = 32'b00000000000000001101000001100100;
assign LUT_4[46961] = 32'b00000000000000000110001101011100;
assign LUT_4[46962] = 32'b00000000000000001100011100001000;
assign LUT_4[46963] = 32'b00000000000000000101101000000000;
assign LUT_4[46964] = 32'b00000000000000001010000010000000;
assign LUT_4[46965] = 32'b00000000000000000011001101111000;
assign LUT_4[46966] = 32'b00000000000000001001011100100100;
assign LUT_4[46967] = 32'b00000000000000000010101000011100;
assign LUT_4[46968] = 32'b00000000000000000110001101111001;
assign LUT_4[46969] = 32'b11111111111111111111011001110001;
assign LUT_4[46970] = 32'b00000000000000000101101000011101;
assign LUT_4[46971] = 32'b11111111111111111110110100010101;
assign LUT_4[46972] = 32'b00000000000000000011001110010101;
assign LUT_4[46973] = 32'b11111111111111111100011010001101;
assign LUT_4[46974] = 32'b00000000000000000010101000111001;
assign LUT_4[46975] = 32'b11111111111111111011110100110001;
assign LUT_4[46976] = 32'b00000000000000010010000011100011;
assign LUT_4[46977] = 32'b00000000000000001011001111011011;
assign LUT_4[46978] = 32'b00000000000000010001011110000111;
assign LUT_4[46979] = 32'b00000000000000001010101001111111;
assign LUT_4[46980] = 32'b00000000000000001111000011111111;
assign LUT_4[46981] = 32'b00000000000000001000001111110111;
assign LUT_4[46982] = 32'b00000000000000001110011110100011;
assign LUT_4[46983] = 32'b00000000000000000111101010011011;
assign LUT_4[46984] = 32'b00000000000000001011001111111000;
assign LUT_4[46985] = 32'b00000000000000000100011011110000;
assign LUT_4[46986] = 32'b00000000000000001010101010011100;
assign LUT_4[46987] = 32'b00000000000000000011110110010100;
assign LUT_4[46988] = 32'b00000000000000001000010000010100;
assign LUT_4[46989] = 32'b00000000000000000001011100001100;
assign LUT_4[46990] = 32'b00000000000000000111101010111000;
assign LUT_4[46991] = 32'b00000000000000000000110110110000;
assign LUT_4[46992] = 32'b00000000000000001111110101010001;
assign LUT_4[46993] = 32'b00000000000000001001000001001001;
assign LUT_4[46994] = 32'b00000000000000001111001111110101;
assign LUT_4[46995] = 32'b00000000000000001000011011101101;
assign LUT_4[46996] = 32'b00000000000000001100110101101101;
assign LUT_4[46997] = 32'b00000000000000000110000001100101;
assign LUT_4[46998] = 32'b00000000000000001100010000010001;
assign LUT_4[46999] = 32'b00000000000000000101011100001001;
assign LUT_4[47000] = 32'b00000000000000001001000001100110;
assign LUT_4[47001] = 32'b00000000000000000010001101011110;
assign LUT_4[47002] = 32'b00000000000000001000011100001010;
assign LUT_4[47003] = 32'b00000000000000000001101000000010;
assign LUT_4[47004] = 32'b00000000000000000110000010000010;
assign LUT_4[47005] = 32'b11111111111111111111001101111010;
assign LUT_4[47006] = 32'b00000000000000000101011100100110;
assign LUT_4[47007] = 32'b11111111111111111110101000011110;
assign LUT_4[47008] = 32'b00000000000000010000011110101010;
assign LUT_4[47009] = 32'b00000000000000001001101010100010;
assign LUT_4[47010] = 32'b00000000000000001111111001001110;
assign LUT_4[47011] = 32'b00000000000000001001000101000110;
assign LUT_4[47012] = 32'b00000000000000001101011111000110;
assign LUT_4[47013] = 32'b00000000000000000110101010111110;
assign LUT_4[47014] = 32'b00000000000000001100111001101010;
assign LUT_4[47015] = 32'b00000000000000000110000101100010;
assign LUT_4[47016] = 32'b00000000000000001001101010111111;
assign LUT_4[47017] = 32'b00000000000000000010110110110111;
assign LUT_4[47018] = 32'b00000000000000001001000101100011;
assign LUT_4[47019] = 32'b00000000000000000010010001011011;
assign LUT_4[47020] = 32'b00000000000000000110101011011011;
assign LUT_4[47021] = 32'b11111111111111111111110111010011;
assign LUT_4[47022] = 32'b00000000000000000110000101111111;
assign LUT_4[47023] = 32'b11111111111111111111010001110111;
assign LUT_4[47024] = 32'b00000000000000001110010000011000;
assign LUT_4[47025] = 32'b00000000000000000111011100010000;
assign LUT_4[47026] = 32'b00000000000000001101101010111100;
assign LUT_4[47027] = 32'b00000000000000000110110110110100;
assign LUT_4[47028] = 32'b00000000000000001011010000110100;
assign LUT_4[47029] = 32'b00000000000000000100011100101100;
assign LUT_4[47030] = 32'b00000000000000001010101011011000;
assign LUT_4[47031] = 32'b00000000000000000011110111010000;
assign LUT_4[47032] = 32'b00000000000000000111011100101101;
assign LUT_4[47033] = 32'b00000000000000000000101000100101;
assign LUT_4[47034] = 32'b00000000000000000110110111010001;
assign LUT_4[47035] = 32'b00000000000000000000000011001001;
assign LUT_4[47036] = 32'b00000000000000000100011101001001;
assign LUT_4[47037] = 32'b11111111111111111101101001000001;
assign LUT_4[47038] = 32'b00000000000000000011110111101101;
assign LUT_4[47039] = 32'b11111111111111111101000011100101;
assign LUT_4[47040] = 32'b00000000000000010011011010110111;
assign LUT_4[47041] = 32'b00000000000000001100100110101111;
assign LUT_4[47042] = 32'b00000000000000010010110101011011;
assign LUT_4[47043] = 32'b00000000000000001100000001010011;
assign LUT_4[47044] = 32'b00000000000000010000011011010011;
assign LUT_4[47045] = 32'b00000000000000001001100111001011;
assign LUT_4[47046] = 32'b00000000000000001111110101110111;
assign LUT_4[47047] = 32'b00000000000000001001000001101111;
assign LUT_4[47048] = 32'b00000000000000001100100111001100;
assign LUT_4[47049] = 32'b00000000000000000101110011000100;
assign LUT_4[47050] = 32'b00000000000000001100000001110000;
assign LUT_4[47051] = 32'b00000000000000000101001101101000;
assign LUT_4[47052] = 32'b00000000000000001001100111101000;
assign LUT_4[47053] = 32'b00000000000000000010110011100000;
assign LUT_4[47054] = 32'b00000000000000001001000010001100;
assign LUT_4[47055] = 32'b00000000000000000010001110000100;
assign LUT_4[47056] = 32'b00000000000000010001001100100101;
assign LUT_4[47057] = 32'b00000000000000001010011000011101;
assign LUT_4[47058] = 32'b00000000000000010000100111001001;
assign LUT_4[47059] = 32'b00000000000000001001110011000001;
assign LUT_4[47060] = 32'b00000000000000001110001101000001;
assign LUT_4[47061] = 32'b00000000000000000111011000111001;
assign LUT_4[47062] = 32'b00000000000000001101100111100101;
assign LUT_4[47063] = 32'b00000000000000000110110011011101;
assign LUT_4[47064] = 32'b00000000000000001010011000111010;
assign LUT_4[47065] = 32'b00000000000000000011100100110010;
assign LUT_4[47066] = 32'b00000000000000001001110011011110;
assign LUT_4[47067] = 32'b00000000000000000010111111010110;
assign LUT_4[47068] = 32'b00000000000000000111011001010110;
assign LUT_4[47069] = 32'b00000000000000000000100101001110;
assign LUT_4[47070] = 32'b00000000000000000110110011111010;
assign LUT_4[47071] = 32'b11111111111111111111111111110010;
assign LUT_4[47072] = 32'b00000000000000010001110101111110;
assign LUT_4[47073] = 32'b00000000000000001011000001110110;
assign LUT_4[47074] = 32'b00000000000000010001010000100010;
assign LUT_4[47075] = 32'b00000000000000001010011100011010;
assign LUT_4[47076] = 32'b00000000000000001110110110011010;
assign LUT_4[47077] = 32'b00000000000000001000000010010010;
assign LUT_4[47078] = 32'b00000000000000001110010000111110;
assign LUT_4[47079] = 32'b00000000000000000111011100110110;
assign LUT_4[47080] = 32'b00000000000000001011000010010011;
assign LUT_4[47081] = 32'b00000000000000000100001110001011;
assign LUT_4[47082] = 32'b00000000000000001010011100110111;
assign LUT_4[47083] = 32'b00000000000000000011101000101111;
assign LUT_4[47084] = 32'b00000000000000001000000010101111;
assign LUT_4[47085] = 32'b00000000000000000001001110100111;
assign LUT_4[47086] = 32'b00000000000000000111011101010011;
assign LUT_4[47087] = 32'b00000000000000000000101001001011;
assign LUT_4[47088] = 32'b00000000000000001111100111101100;
assign LUT_4[47089] = 32'b00000000000000001000110011100100;
assign LUT_4[47090] = 32'b00000000000000001111000010010000;
assign LUT_4[47091] = 32'b00000000000000001000001110001000;
assign LUT_4[47092] = 32'b00000000000000001100101000001000;
assign LUT_4[47093] = 32'b00000000000000000101110100000000;
assign LUT_4[47094] = 32'b00000000000000001100000010101100;
assign LUT_4[47095] = 32'b00000000000000000101001110100100;
assign LUT_4[47096] = 32'b00000000000000001000110100000001;
assign LUT_4[47097] = 32'b00000000000000000001111111111001;
assign LUT_4[47098] = 32'b00000000000000001000001110100101;
assign LUT_4[47099] = 32'b00000000000000000001011010011101;
assign LUT_4[47100] = 32'b00000000000000000101110100011101;
assign LUT_4[47101] = 32'b11111111111111111111000000010101;
assign LUT_4[47102] = 32'b00000000000000000101001111000001;
assign LUT_4[47103] = 32'b11111111111111111110011010111001;
assign LUT_4[47104] = 32'b00000000000000000101010010011011;
assign LUT_4[47105] = 32'b11111111111111111110011110010011;
assign LUT_4[47106] = 32'b00000000000000000100101100111111;
assign LUT_4[47107] = 32'b11111111111111111101111000110111;
assign LUT_4[47108] = 32'b00000000000000000010010010110111;
assign LUT_4[47109] = 32'b11111111111111111011011110101111;
assign LUT_4[47110] = 32'b00000000000000000001101101011011;
assign LUT_4[47111] = 32'b11111111111111111010111001010011;
assign LUT_4[47112] = 32'b11111111111111111110011110110000;
assign LUT_4[47113] = 32'b11111111111111110111101010101000;
assign LUT_4[47114] = 32'b11111111111111111101111001010100;
assign LUT_4[47115] = 32'b11111111111111110111000101001100;
assign LUT_4[47116] = 32'b11111111111111111011011111001100;
assign LUT_4[47117] = 32'b11111111111111110100101011000100;
assign LUT_4[47118] = 32'b11111111111111111010111001110000;
assign LUT_4[47119] = 32'b11111111111111110100000101101000;
assign LUT_4[47120] = 32'b00000000000000000011000100001001;
assign LUT_4[47121] = 32'b11111111111111111100010000000001;
assign LUT_4[47122] = 32'b00000000000000000010011110101101;
assign LUT_4[47123] = 32'b11111111111111111011101010100101;
assign LUT_4[47124] = 32'b00000000000000000000000100100101;
assign LUT_4[47125] = 32'b11111111111111111001010000011101;
assign LUT_4[47126] = 32'b11111111111111111111011111001001;
assign LUT_4[47127] = 32'b11111111111111111000101011000001;
assign LUT_4[47128] = 32'b11111111111111111100010000011110;
assign LUT_4[47129] = 32'b11111111111111110101011100010110;
assign LUT_4[47130] = 32'b11111111111111111011101011000010;
assign LUT_4[47131] = 32'b11111111111111110100110110111010;
assign LUT_4[47132] = 32'b11111111111111111001010000111010;
assign LUT_4[47133] = 32'b11111111111111110010011100110010;
assign LUT_4[47134] = 32'b11111111111111111000101011011110;
assign LUT_4[47135] = 32'b11111111111111110001110111010110;
assign LUT_4[47136] = 32'b00000000000000000011101101100010;
assign LUT_4[47137] = 32'b11111111111111111100111001011010;
assign LUT_4[47138] = 32'b00000000000000000011001000000110;
assign LUT_4[47139] = 32'b11111111111111111100010011111110;
assign LUT_4[47140] = 32'b00000000000000000000101101111110;
assign LUT_4[47141] = 32'b11111111111111111001111001110110;
assign LUT_4[47142] = 32'b00000000000000000000001000100010;
assign LUT_4[47143] = 32'b11111111111111111001010100011010;
assign LUT_4[47144] = 32'b11111111111111111100111001110111;
assign LUT_4[47145] = 32'b11111111111111110110000101101111;
assign LUT_4[47146] = 32'b11111111111111111100010100011011;
assign LUT_4[47147] = 32'b11111111111111110101100000010011;
assign LUT_4[47148] = 32'b11111111111111111001111010010011;
assign LUT_4[47149] = 32'b11111111111111110011000110001011;
assign LUT_4[47150] = 32'b11111111111111111001010100110111;
assign LUT_4[47151] = 32'b11111111111111110010100000101111;
assign LUT_4[47152] = 32'b00000000000000000001011111010000;
assign LUT_4[47153] = 32'b11111111111111111010101011001000;
assign LUT_4[47154] = 32'b00000000000000000000111001110100;
assign LUT_4[47155] = 32'b11111111111111111010000101101100;
assign LUT_4[47156] = 32'b11111111111111111110011111101100;
assign LUT_4[47157] = 32'b11111111111111110111101011100100;
assign LUT_4[47158] = 32'b11111111111111111101111010010000;
assign LUT_4[47159] = 32'b11111111111111110111000110001000;
assign LUT_4[47160] = 32'b11111111111111111010101011100101;
assign LUT_4[47161] = 32'b11111111111111110011110111011101;
assign LUT_4[47162] = 32'b11111111111111111010000110001001;
assign LUT_4[47163] = 32'b11111111111111110011010010000001;
assign LUT_4[47164] = 32'b11111111111111110111101100000001;
assign LUT_4[47165] = 32'b11111111111111110000110111111001;
assign LUT_4[47166] = 32'b11111111111111110111000110100101;
assign LUT_4[47167] = 32'b11111111111111110000010010011101;
assign LUT_4[47168] = 32'b00000000000000000110101001101111;
assign LUT_4[47169] = 32'b11111111111111111111110101100111;
assign LUT_4[47170] = 32'b00000000000000000110000100010011;
assign LUT_4[47171] = 32'b11111111111111111111010000001011;
assign LUT_4[47172] = 32'b00000000000000000011101010001011;
assign LUT_4[47173] = 32'b11111111111111111100110110000011;
assign LUT_4[47174] = 32'b00000000000000000011000100101111;
assign LUT_4[47175] = 32'b11111111111111111100010000100111;
assign LUT_4[47176] = 32'b11111111111111111111110110000100;
assign LUT_4[47177] = 32'b11111111111111111001000001111100;
assign LUT_4[47178] = 32'b11111111111111111111010000101000;
assign LUT_4[47179] = 32'b11111111111111111000011100100000;
assign LUT_4[47180] = 32'b11111111111111111100110110100000;
assign LUT_4[47181] = 32'b11111111111111110110000010011000;
assign LUT_4[47182] = 32'b11111111111111111100010001000100;
assign LUT_4[47183] = 32'b11111111111111110101011100111100;
assign LUT_4[47184] = 32'b00000000000000000100011011011101;
assign LUT_4[47185] = 32'b11111111111111111101100111010101;
assign LUT_4[47186] = 32'b00000000000000000011110110000001;
assign LUT_4[47187] = 32'b11111111111111111101000001111001;
assign LUT_4[47188] = 32'b00000000000000000001011011111001;
assign LUT_4[47189] = 32'b11111111111111111010100111110001;
assign LUT_4[47190] = 32'b00000000000000000000110110011101;
assign LUT_4[47191] = 32'b11111111111111111010000010010101;
assign LUT_4[47192] = 32'b11111111111111111101100111110010;
assign LUT_4[47193] = 32'b11111111111111110110110011101010;
assign LUT_4[47194] = 32'b11111111111111111101000010010110;
assign LUT_4[47195] = 32'b11111111111111110110001110001110;
assign LUT_4[47196] = 32'b11111111111111111010101000001110;
assign LUT_4[47197] = 32'b11111111111111110011110100000110;
assign LUT_4[47198] = 32'b11111111111111111010000010110010;
assign LUT_4[47199] = 32'b11111111111111110011001110101010;
assign LUT_4[47200] = 32'b00000000000000000101000100110110;
assign LUT_4[47201] = 32'b11111111111111111110010000101110;
assign LUT_4[47202] = 32'b00000000000000000100011111011010;
assign LUT_4[47203] = 32'b11111111111111111101101011010010;
assign LUT_4[47204] = 32'b00000000000000000010000101010010;
assign LUT_4[47205] = 32'b11111111111111111011010001001010;
assign LUT_4[47206] = 32'b00000000000000000001011111110110;
assign LUT_4[47207] = 32'b11111111111111111010101011101110;
assign LUT_4[47208] = 32'b11111111111111111110010001001011;
assign LUT_4[47209] = 32'b11111111111111110111011101000011;
assign LUT_4[47210] = 32'b11111111111111111101101011101111;
assign LUT_4[47211] = 32'b11111111111111110110110111100111;
assign LUT_4[47212] = 32'b11111111111111111011010001100111;
assign LUT_4[47213] = 32'b11111111111111110100011101011111;
assign LUT_4[47214] = 32'b11111111111111111010101100001011;
assign LUT_4[47215] = 32'b11111111111111110011111000000011;
assign LUT_4[47216] = 32'b00000000000000000010110110100100;
assign LUT_4[47217] = 32'b11111111111111111100000010011100;
assign LUT_4[47218] = 32'b00000000000000000010010001001000;
assign LUT_4[47219] = 32'b11111111111111111011011101000000;
assign LUT_4[47220] = 32'b11111111111111111111110111000000;
assign LUT_4[47221] = 32'b11111111111111111001000010111000;
assign LUT_4[47222] = 32'b11111111111111111111010001100100;
assign LUT_4[47223] = 32'b11111111111111111000011101011100;
assign LUT_4[47224] = 32'b11111111111111111100000010111001;
assign LUT_4[47225] = 32'b11111111111111110101001110110001;
assign LUT_4[47226] = 32'b11111111111111111011011101011101;
assign LUT_4[47227] = 32'b11111111111111110100101001010101;
assign LUT_4[47228] = 32'b11111111111111111001000011010101;
assign LUT_4[47229] = 32'b11111111111111110010001111001101;
assign LUT_4[47230] = 32'b11111111111111111000011101111001;
assign LUT_4[47231] = 32'b11111111111111110001101001110001;
assign LUT_4[47232] = 32'b00000000000000000111111000100011;
assign LUT_4[47233] = 32'b00000000000000000001000100011011;
assign LUT_4[47234] = 32'b00000000000000000111010011000111;
assign LUT_4[47235] = 32'b00000000000000000000011110111111;
assign LUT_4[47236] = 32'b00000000000000000100111000111111;
assign LUT_4[47237] = 32'b11111111111111111110000100110111;
assign LUT_4[47238] = 32'b00000000000000000100010011100011;
assign LUT_4[47239] = 32'b11111111111111111101011111011011;
assign LUT_4[47240] = 32'b00000000000000000001000100111000;
assign LUT_4[47241] = 32'b11111111111111111010010000110000;
assign LUT_4[47242] = 32'b00000000000000000000011111011100;
assign LUT_4[47243] = 32'b11111111111111111001101011010100;
assign LUT_4[47244] = 32'b11111111111111111110000101010100;
assign LUT_4[47245] = 32'b11111111111111110111010001001100;
assign LUT_4[47246] = 32'b11111111111111111101011111111000;
assign LUT_4[47247] = 32'b11111111111111110110101011110000;
assign LUT_4[47248] = 32'b00000000000000000101101010010001;
assign LUT_4[47249] = 32'b11111111111111111110110110001001;
assign LUT_4[47250] = 32'b00000000000000000101000100110101;
assign LUT_4[47251] = 32'b11111111111111111110010000101101;
assign LUT_4[47252] = 32'b00000000000000000010101010101101;
assign LUT_4[47253] = 32'b11111111111111111011110110100101;
assign LUT_4[47254] = 32'b00000000000000000010000101010001;
assign LUT_4[47255] = 32'b11111111111111111011010001001001;
assign LUT_4[47256] = 32'b11111111111111111110110110100110;
assign LUT_4[47257] = 32'b11111111111111111000000010011110;
assign LUT_4[47258] = 32'b11111111111111111110010001001010;
assign LUT_4[47259] = 32'b11111111111111110111011101000010;
assign LUT_4[47260] = 32'b11111111111111111011110111000010;
assign LUT_4[47261] = 32'b11111111111111110101000010111010;
assign LUT_4[47262] = 32'b11111111111111111011010001100110;
assign LUT_4[47263] = 32'b11111111111111110100011101011110;
assign LUT_4[47264] = 32'b00000000000000000110010011101010;
assign LUT_4[47265] = 32'b11111111111111111111011111100010;
assign LUT_4[47266] = 32'b00000000000000000101101110001110;
assign LUT_4[47267] = 32'b11111111111111111110111010000110;
assign LUT_4[47268] = 32'b00000000000000000011010100000110;
assign LUT_4[47269] = 32'b11111111111111111100011111111110;
assign LUT_4[47270] = 32'b00000000000000000010101110101010;
assign LUT_4[47271] = 32'b11111111111111111011111010100010;
assign LUT_4[47272] = 32'b11111111111111111111011111111111;
assign LUT_4[47273] = 32'b11111111111111111000101011110111;
assign LUT_4[47274] = 32'b11111111111111111110111010100011;
assign LUT_4[47275] = 32'b11111111111111111000000110011011;
assign LUT_4[47276] = 32'b11111111111111111100100000011011;
assign LUT_4[47277] = 32'b11111111111111110101101100010011;
assign LUT_4[47278] = 32'b11111111111111111011111010111111;
assign LUT_4[47279] = 32'b11111111111111110101000110110111;
assign LUT_4[47280] = 32'b00000000000000000100000101011000;
assign LUT_4[47281] = 32'b11111111111111111101010001010000;
assign LUT_4[47282] = 32'b00000000000000000011011111111100;
assign LUT_4[47283] = 32'b11111111111111111100101011110100;
assign LUT_4[47284] = 32'b00000000000000000001000101110100;
assign LUT_4[47285] = 32'b11111111111111111010010001101100;
assign LUT_4[47286] = 32'b00000000000000000000100000011000;
assign LUT_4[47287] = 32'b11111111111111111001101100010000;
assign LUT_4[47288] = 32'b11111111111111111101010001101101;
assign LUT_4[47289] = 32'b11111111111111110110011101100101;
assign LUT_4[47290] = 32'b11111111111111111100101100010001;
assign LUT_4[47291] = 32'b11111111111111110101111000001001;
assign LUT_4[47292] = 32'b11111111111111111010010010001001;
assign LUT_4[47293] = 32'b11111111111111110011011110000001;
assign LUT_4[47294] = 32'b11111111111111111001101100101101;
assign LUT_4[47295] = 32'b11111111111111110010111000100101;
assign LUT_4[47296] = 32'b00000000000000001001001111110111;
assign LUT_4[47297] = 32'b00000000000000000010011011101111;
assign LUT_4[47298] = 32'b00000000000000001000101010011011;
assign LUT_4[47299] = 32'b00000000000000000001110110010011;
assign LUT_4[47300] = 32'b00000000000000000110010000010011;
assign LUT_4[47301] = 32'b11111111111111111111011100001011;
assign LUT_4[47302] = 32'b00000000000000000101101010110111;
assign LUT_4[47303] = 32'b11111111111111111110110110101111;
assign LUT_4[47304] = 32'b00000000000000000010011100001100;
assign LUT_4[47305] = 32'b11111111111111111011101000000100;
assign LUT_4[47306] = 32'b00000000000000000001110110110000;
assign LUT_4[47307] = 32'b11111111111111111011000010101000;
assign LUT_4[47308] = 32'b11111111111111111111011100101000;
assign LUT_4[47309] = 32'b11111111111111111000101000100000;
assign LUT_4[47310] = 32'b11111111111111111110110111001100;
assign LUT_4[47311] = 32'b11111111111111111000000011000100;
assign LUT_4[47312] = 32'b00000000000000000111000001100101;
assign LUT_4[47313] = 32'b00000000000000000000001101011101;
assign LUT_4[47314] = 32'b00000000000000000110011100001001;
assign LUT_4[47315] = 32'b11111111111111111111101000000001;
assign LUT_4[47316] = 32'b00000000000000000100000010000001;
assign LUT_4[47317] = 32'b11111111111111111101001101111001;
assign LUT_4[47318] = 32'b00000000000000000011011100100101;
assign LUT_4[47319] = 32'b11111111111111111100101000011101;
assign LUT_4[47320] = 32'b00000000000000000000001101111010;
assign LUT_4[47321] = 32'b11111111111111111001011001110010;
assign LUT_4[47322] = 32'b11111111111111111111101000011110;
assign LUT_4[47323] = 32'b11111111111111111000110100010110;
assign LUT_4[47324] = 32'b11111111111111111101001110010110;
assign LUT_4[47325] = 32'b11111111111111110110011010001110;
assign LUT_4[47326] = 32'b11111111111111111100101000111010;
assign LUT_4[47327] = 32'b11111111111111110101110100110010;
assign LUT_4[47328] = 32'b00000000000000000111101010111110;
assign LUT_4[47329] = 32'b00000000000000000000110110110110;
assign LUT_4[47330] = 32'b00000000000000000111000101100010;
assign LUT_4[47331] = 32'b00000000000000000000010001011010;
assign LUT_4[47332] = 32'b00000000000000000100101011011010;
assign LUT_4[47333] = 32'b11111111111111111101110111010010;
assign LUT_4[47334] = 32'b00000000000000000100000101111110;
assign LUT_4[47335] = 32'b11111111111111111101010001110110;
assign LUT_4[47336] = 32'b00000000000000000000110111010011;
assign LUT_4[47337] = 32'b11111111111111111010000011001011;
assign LUT_4[47338] = 32'b00000000000000000000010001110111;
assign LUT_4[47339] = 32'b11111111111111111001011101101111;
assign LUT_4[47340] = 32'b11111111111111111101110111101111;
assign LUT_4[47341] = 32'b11111111111111110111000011100111;
assign LUT_4[47342] = 32'b11111111111111111101010010010011;
assign LUT_4[47343] = 32'b11111111111111110110011110001011;
assign LUT_4[47344] = 32'b00000000000000000101011100101100;
assign LUT_4[47345] = 32'b11111111111111111110101000100100;
assign LUT_4[47346] = 32'b00000000000000000100110111010000;
assign LUT_4[47347] = 32'b11111111111111111110000011001000;
assign LUT_4[47348] = 32'b00000000000000000010011101001000;
assign LUT_4[47349] = 32'b11111111111111111011101001000000;
assign LUT_4[47350] = 32'b00000000000000000001110111101100;
assign LUT_4[47351] = 32'b11111111111111111011000011100100;
assign LUT_4[47352] = 32'b11111111111111111110101001000001;
assign LUT_4[47353] = 32'b11111111111111110111110100111001;
assign LUT_4[47354] = 32'b11111111111111111110000011100101;
assign LUT_4[47355] = 32'b11111111111111110111001111011101;
assign LUT_4[47356] = 32'b11111111111111111011101001011101;
assign LUT_4[47357] = 32'b11111111111111110100110101010101;
assign LUT_4[47358] = 32'b11111111111111111011000100000001;
assign LUT_4[47359] = 32'b11111111111111110100001111111001;
assign LUT_4[47360] = 32'b00000000000000001010001101111110;
assign LUT_4[47361] = 32'b00000000000000000011011001110110;
assign LUT_4[47362] = 32'b00000000000000001001101000100010;
assign LUT_4[47363] = 32'b00000000000000000010110100011010;
assign LUT_4[47364] = 32'b00000000000000000111001110011010;
assign LUT_4[47365] = 32'b00000000000000000000011010010010;
assign LUT_4[47366] = 32'b00000000000000000110101000111110;
assign LUT_4[47367] = 32'b11111111111111111111110100110110;
assign LUT_4[47368] = 32'b00000000000000000011011010010011;
assign LUT_4[47369] = 32'b11111111111111111100100110001011;
assign LUT_4[47370] = 32'b00000000000000000010110100110111;
assign LUT_4[47371] = 32'b11111111111111111100000000101111;
assign LUT_4[47372] = 32'b00000000000000000000011010101111;
assign LUT_4[47373] = 32'b11111111111111111001100110100111;
assign LUT_4[47374] = 32'b11111111111111111111110101010011;
assign LUT_4[47375] = 32'b11111111111111111001000001001011;
assign LUT_4[47376] = 32'b00000000000000000111111111101100;
assign LUT_4[47377] = 32'b00000000000000000001001011100100;
assign LUT_4[47378] = 32'b00000000000000000111011010010000;
assign LUT_4[47379] = 32'b00000000000000000000100110001000;
assign LUT_4[47380] = 32'b00000000000000000101000000001000;
assign LUT_4[47381] = 32'b11111111111111111110001100000000;
assign LUT_4[47382] = 32'b00000000000000000100011010101100;
assign LUT_4[47383] = 32'b11111111111111111101100110100100;
assign LUT_4[47384] = 32'b00000000000000000001001100000001;
assign LUT_4[47385] = 32'b11111111111111111010010111111001;
assign LUT_4[47386] = 32'b00000000000000000000100110100101;
assign LUT_4[47387] = 32'b11111111111111111001110010011101;
assign LUT_4[47388] = 32'b11111111111111111110001100011101;
assign LUT_4[47389] = 32'b11111111111111110111011000010101;
assign LUT_4[47390] = 32'b11111111111111111101100111000001;
assign LUT_4[47391] = 32'b11111111111111110110110010111001;
assign LUT_4[47392] = 32'b00000000000000001000101001000101;
assign LUT_4[47393] = 32'b00000000000000000001110100111101;
assign LUT_4[47394] = 32'b00000000000000001000000011101001;
assign LUT_4[47395] = 32'b00000000000000000001001111100001;
assign LUT_4[47396] = 32'b00000000000000000101101001100001;
assign LUT_4[47397] = 32'b11111111111111111110110101011001;
assign LUT_4[47398] = 32'b00000000000000000101000100000101;
assign LUT_4[47399] = 32'b11111111111111111110001111111101;
assign LUT_4[47400] = 32'b00000000000000000001110101011010;
assign LUT_4[47401] = 32'b11111111111111111011000001010010;
assign LUT_4[47402] = 32'b00000000000000000001001111111110;
assign LUT_4[47403] = 32'b11111111111111111010011011110110;
assign LUT_4[47404] = 32'b11111111111111111110110101110110;
assign LUT_4[47405] = 32'b11111111111111111000000001101110;
assign LUT_4[47406] = 32'b11111111111111111110010000011010;
assign LUT_4[47407] = 32'b11111111111111110111011100010010;
assign LUT_4[47408] = 32'b00000000000000000110011010110011;
assign LUT_4[47409] = 32'b11111111111111111111100110101011;
assign LUT_4[47410] = 32'b00000000000000000101110101010111;
assign LUT_4[47411] = 32'b11111111111111111111000001001111;
assign LUT_4[47412] = 32'b00000000000000000011011011001111;
assign LUT_4[47413] = 32'b11111111111111111100100111000111;
assign LUT_4[47414] = 32'b00000000000000000010110101110011;
assign LUT_4[47415] = 32'b11111111111111111100000001101011;
assign LUT_4[47416] = 32'b11111111111111111111100111001000;
assign LUT_4[47417] = 32'b11111111111111111000110011000000;
assign LUT_4[47418] = 32'b11111111111111111111000001101100;
assign LUT_4[47419] = 32'b11111111111111111000001101100100;
assign LUT_4[47420] = 32'b11111111111111111100100111100100;
assign LUT_4[47421] = 32'b11111111111111110101110011011100;
assign LUT_4[47422] = 32'b11111111111111111100000010001000;
assign LUT_4[47423] = 32'b11111111111111110101001110000000;
assign LUT_4[47424] = 32'b00000000000000001011100101010010;
assign LUT_4[47425] = 32'b00000000000000000100110001001010;
assign LUT_4[47426] = 32'b00000000000000001010111111110110;
assign LUT_4[47427] = 32'b00000000000000000100001011101110;
assign LUT_4[47428] = 32'b00000000000000001000100101101110;
assign LUT_4[47429] = 32'b00000000000000000001110001100110;
assign LUT_4[47430] = 32'b00000000000000001000000000010010;
assign LUT_4[47431] = 32'b00000000000000000001001100001010;
assign LUT_4[47432] = 32'b00000000000000000100110001100111;
assign LUT_4[47433] = 32'b11111111111111111101111101011111;
assign LUT_4[47434] = 32'b00000000000000000100001100001011;
assign LUT_4[47435] = 32'b11111111111111111101011000000011;
assign LUT_4[47436] = 32'b00000000000000000001110010000011;
assign LUT_4[47437] = 32'b11111111111111111010111101111011;
assign LUT_4[47438] = 32'b00000000000000000001001100100111;
assign LUT_4[47439] = 32'b11111111111111111010011000011111;
assign LUT_4[47440] = 32'b00000000000000001001010111000000;
assign LUT_4[47441] = 32'b00000000000000000010100010111000;
assign LUT_4[47442] = 32'b00000000000000001000110001100100;
assign LUT_4[47443] = 32'b00000000000000000001111101011100;
assign LUT_4[47444] = 32'b00000000000000000110010111011100;
assign LUT_4[47445] = 32'b11111111111111111111100011010100;
assign LUT_4[47446] = 32'b00000000000000000101110010000000;
assign LUT_4[47447] = 32'b11111111111111111110111101111000;
assign LUT_4[47448] = 32'b00000000000000000010100011010101;
assign LUT_4[47449] = 32'b11111111111111111011101111001101;
assign LUT_4[47450] = 32'b00000000000000000001111101111001;
assign LUT_4[47451] = 32'b11111111111111111011001001110001;
assign LUT_4[47452] = 32'b11111111111111111111100011110001;
assign LUT_4[47453] = 32'b11111111111111111000101111101001;
assign LUT_4[47454] = 32'b11111111111111111110111110010101;
assign LUT_4[47455] = 32'b11111111111111111000001010001101;
assign LUT_4[47456] = 32'b00000000000000001010000000011001;
assign LUT_4[47457] = 32'b00000000000000000011001100010001;
assign LUT_4[47458] = 32'b00000000000000001001011010111101;
assign LUT_4[47459] = 32'b00000000000000000010100110110101;
assign LUT_4[47460] = 32'b00000000000000000111000000110101;
assign LUT_4[47461] = 32'b00000000000000000000001100101101;
assign LUT_4[47462] = 32'b00000000000000000110011011011001;
assign LUT_4[47463] = 32'b11111111111111111111100111010001;
assign LUT_4[47464] = 32'b00000000000000000011001100101110;
assign LUT_4[47465] = 32'b11111111111111111100011000100110;
assign LUT_4[47466] = 32'b00000000000000000010100111010010;
assign LUT_4[47467] = 32'b11111111111111111011110011001010;
assign LUT_4[47468] = 32'b00000000000000000000001101001010;
assign LUT_4[47469] = 32'b11111111111111111001011001000010;
assign LUT_4[47470] = 32'b11111111111111111111100111101110;
assign LUT_4[47471] = 32'b11111111111111111000110011100110;
assign LUT_4[47472] = 32'b00000000000000000111110010000111;
assign LUT_4[47473] = 32'b00000000000000000000111101111111;
assign LUT_4[47474] = 32'b00000000000000000111001100101011;
assign LUT_4[47475] = 32'b00000000000000000000011000100011;
assign LUT_4[47476] = 32'b00000000000000000100110010100011;
assign LUT_4[47477] = 32'b11111111111111111101111110011011;
assign LUT_4[47478] = 32'b00000000000000000100001101000111;
assign LUT_4[47479] = 32'b11111111111111111101011000111111;
assign LUT_4[47480] = 32'b00000000000000000000111110011100;
assign LUT_4[47481] = 32'b11111111111111111010001010010100;
assign LUT_4[47482] = 32'b00000000000000000000011001000000;
assign LUT_4[47483] = 32'b11111111111111111001100100111000;
assign LUT_4[47484] = 32'b11111111111111111101111110111000;
assign LUT_4[47485] = 32'b11111111111111110111001010110000;
assign LUT_4[47486] = 32'b11111111111111111101011001011100;
assign LUT_4[47487] = 32'b11111111111111110110100101010100;
assign LUT_4[47488] = 32'b00000000000000001100110100000110;
assign LUT_4[47489] = 32'b00000000000000000101111111111110;
assign LUT_4[47490] = 32'b00000000000000001100001110101010;
assign LUT_4[47491] = 32'b00000000000000000101011010100010;
assign LUT_4[47492] = 32'b00000000000000001001110100100010;
assign LUT_4[47493] = 32'b00000000000000000011000000011010;
assign LUT_4[47494] = 32'b00000000000000001001001111000110;
assign LUT_4[47495] = 32'b00000000000000000010011010111110;
assign LUT_4[47496] = 32'b00000000000000000110000000011011;
assign LUT_4[47497] = 32'b11111111111111111111001100010011;
assign LUT_4[47498] = 32'b00000000000000000101011010111111;
assign LUT_4[47499] = 32'b11111111111111111110100110110111;
assign LUT_4[47500] = 32'b00000000000000000011000000110111;
assign LUT_4[47501] = 32'b11111111111111111100001100101111;
assign LUT_4[47502] = 32'b00000000000000000010011011011011;
assign LUT_4[47503] = 32'b11111111111111111011100111010011;
assign LUT_4[47504] = 32'b00000000000000001010100101110100;
assign LUT_4[47505] = 32'b00000000000000000011110001101100;
assign LUT_4[47506] = 32'b00000000000000001010000000011000;
assign LUT_4[47507] = 32'b00000000000000000011001100010000;
assign LUT_4[47508] = 32'b00000000000000000111100110010000;
assign LUT_4[47509] = 32'b00000000000000000000110010001000;
assign LUT_4[47510] = 32'b00000000000000000111000000110100;
assign LUT_4[47511] = 32'b00000000000000000000001100101100;
assign LUT_4[47512] = 32'b00000000000000000011110010001001;
assign LUT_4[47513] = 32'b11111111111111111100111110000001;
assign LUT_4[47514] = 32'b00000000000000000011001100101101;
assign LUT_4[47515] = 32'b11111111111111111100011000100101;
assign LUT_4[47516] = 32'b00000000000000000000110010100101;
assign LUT_4[47517] = 32'b11111111111111111001111110011101;
assign LUT_4[47518] = 32'b00000000000000000000001101001001;
assign LUT_4[47519] = 32'b11111111111111111001011001000001;
assign LUT_4[47520] = 32'b00000000000000001011001111001101;
assign LUT_4[47521] = 32'b00000000000000000100011011000101;
assign LUT_4[47522] = 32'b00000000000000001010101001110001;
assign LUT_4[47523] = 32'b00000000000000000011110101101001;
assign LUT_4[47524] = 32'b00000000000000001000001111101001;
assign LUT_4[47525] = 32'b00000000000000000001011011100001;
assign LUT_4[47526] = 32'b00000000000000000111101010001101;
assign LUT_4[47527] = 32'b00000000000000000000110110000101;
assign LUT_4[47528] = 32'b00000000000000000100011011100010;
assign LUT_4[47529] = 32'b11111111111111111101100111011010;
assign LUT_4[47530] = 32'b00000000000000000011110110000110;
assign LUT_4[47531] = 32'b11111111111111111101000001111110;
assign LUT_4[47532] = 32'b00000000000000000001011011111110;
assign LUT_4[47533] = 32'b11111111111111111010100111110110;
assign LUT_4[47534] = 32'b00000000000000000000110110100010;
assign LUT_4[47535] = 32'b11111111111111111010000010011010;
assign LUT_4[47536] = 32'b00000000000000001001000000111011;
assign LUT_4[47537] = 32'b00000000000000000010001100110011;
assign LUT_4[47538] = 32'b00000000000000001000011011011111;
assign LUT_4[47539] = 32'b00000000000000000001100111010111;
assign LUT_4[47540] = 32'b00000000000000000110000001010111;
assign LUT_4[47541] = 32'b11111111111111111111001101001111;
assign LUT_4[47542] = 32'b00000000000000000101011011111011;
assign LUT_4[47543] = 32'b11111111111111111110100111110011;
assign LUT_4[47544] = 32'b00000000000000000010001101010000;
assign LUT_4[47545] = 32'b11111111111111111011011001001000;
assign LUT_4[47546] = 32'b00000000000000000001100111110100;
assign LUT_4[47547] = 32'b11111111111111111010110011101100;
assign LUT_4[47548] = 32'b11111111111111111111001101101100;
assign LUT_4[47549] = 32'b11111111111111111000011001100100;
assign LUT_4[47550] = 32'b11111111111111111110101000010000;
assign LUT_4[47551] = 32'b11111111111111110111110100001000;
assign LUT_4[47552] = 32'b00000000000000001110001011011010;
assign LUT_4[47553] = 32'b00000000000000000111010111010010;
assign LUT_4[47554] = 32'b00000000000000001101100101111110;
assign LUT_4[47555] = 32'b00000000000000000110110001110110;
assign LUT_4[47556] = 32'b00000000000000001011001011110110;
assign LUT_4[47557] = 32'b00000000000000000100010111101110;
assign LUT_4[47558] = 32'b00000000000000001010100110011010;
assign LUT_4[47559] = 32'b00000000000000000011110010010010;
assign LUT_4[47560] = 32'b00000000000000000111010111101111;
assign LUT_4[47561] = 32'b00000000000000000000100011100111;
assign LUT_4[47562] = 32'b00000000000000000110110010010011;
assign LUT_4[47563] = 32'b11111111111111111111111110001011;
assign LUT_4[47564] = 32'b00000000000000000100011000001011;
assign LUT_4[47565] = 32'b11111111111111111101100100000011;
assign LUT_4[47566] = 32'b00000000000000000011110010101111;
assign LUT_4[47567] = 32'b11111111111111111100111110100111;
assign LUT_4[47568] = 32'b00000000000000001011111101001000;
assign LUT_4[47569] = 32'b00000000000000000101001001000000;
assign LUT_4[47570] = 32'b00000000000000001011010111101100;
assign LUT_4[47571] = 32'b00000000000000000100100011100100;
assign LUT_4[47572] = 32'b00000000000000001000111101100100;
assign LUT_4[47573] = 32'b00000000000000000010001001011100;
assign LUT_4[47574] = 32'b00000000000000001000011000001000;
assign LUT_4[47575] = 32'b00000000000000000001100100000000;
assign LUT_4[47576] = 32'b00000000000000000101001001011101;
assign LUT_4[47577] = 32'b11111111111111111110010101010101;
assign LUT_4[47578] = 32'b00000000000000000100100100000001;
assign LUT_4[47579] = 32'b11111111111111111101101111111001;
assign LUT_4[47580] = 32'b00000000000000000010001001111001;
assign LUT_4[47581] = 32'b11111111111111111011010101110001;
assign LUT_4[47582] = 32'b00000000000000000001100100011101;
assign LUT_4[47583] = 32'b11111111111111111010110000010101;
assign LUT_4[47584] = 32'b00000000000000001100100110100001;
assign LUT_4[47585] = 32'b00000000000000000101110010011001;
assign LUT_4[47586] = 32'b00000000000000001100000001000101;
assign LUT_4[47587] = 32'b00000000000000000101001100111101;
assign LUT_4[47588] = 32'b00000000000000001001100110111101;
assign LUT_4[47589] = 32'b00000000000000000010110010110101;
assign LUT_4[47590] = 32'b00000000000000001001000001100001;
assign LUT_4[47591] = 32'b00000000000000000010001101011001;
assign LUT_4[47592] = 32'b00000000000000000101110010110110;
assign LUT_4[47593] = 32'b11111111111111111110111110101110;
assign LUT_4[47594] = 32'b00000000000000000101001101011010;
assign LUT_4[47595] = 32'b11111111111111111110011001010010;
assign LUT_4[47596] = 32'b00000000000000000010110011010010;
assign LUT_4[47597] = 32'b11111111111111111011111111001010;
assign LUT_4[47598] = 32'b00000000000000000010001101110110;
assign LUT_4[47599] = 32'b11111111111111111011011001101110;
assign LUT_4[47600] = 32'b00000000000000001010011000001111;
assign LUT_4[47601] = 32'b00000000000000000011100100000111;
assign LUT_4[47602] = 32'b00000000000000001001110010110011;
assign LUT_4[47603] = 32'b00000000000000000010111110101011;
assign LUT_4[47604] = 32'b00000000000000000111011000101011;
assign LUT_4[47605] = 32'b00000000000000000000100100100011;
assign LUT_4[47606] = 32'b00000000000000000110110011001111;
assign LUT_4[47607] = 32'b11111111111111111111111111000111;
assign LUT_4[47608] = 32'b00000000000000000011100100100100;
assign LUT_4[47609] = 32'b11111111111111111100110000011100;
assign LUT_4[47610] = 32'b00000000000000000010111111001000;
assign LUT_4[47611] = 32'b11111111111111111100001011000000;
assign LUT_4[47612] = 32'b00000000000000000000100101000000;
assign LUT_4[47613] = 32'b11111111111111111001110000111000;
assign LUT_4[47614] = 32'b11111111111111111111111111100100;
assign LUT_4[47615] = 32'b11111111111111111001001011011100;
assign LUT_4[47616] = 32'b00000000000000000100010110100011;
assign LUT_4[47617] = 32'b11111111111111111101100010011011;
assign LUT_4[47618] = 32'b00000000000000000011110001000111;
assign LUT_4[47619] = 32'b11111111111111111100111100111111;
assign LUT_4[47620] = 32'b00000000000000000001010110111111;
assign LUT_4[47621] = 32'b11111111111111111010100010110111;
assign LUT_4[47622] = 32'b00000000000000000000110001100011;
assign LUT_4[47623] = 32'b11111111111111111001111101011011;
assign LUT_4[47624] = 32'b11111111111111111101100010111000;
assign LUT_4[47625] = 32'b11111111111111110110101110110000;
assign LUT_4[47626] = 32'b11111111111111111100111101011100;
assign LUT_4[47627] = 32'b11111111111111110110001001010100;
assign LUT_4[47628] = 32'b11111111111111111010100011010100;
assign LUT_4[47629] = 32'b11111111111111110011101111001100;
assign LUT_4[47630] = 32'b11111111111111111001111101111000;
assign LUT_4[47631] = 32'b11111111111111110011001001110000;
assign LUT_4[47632] = 32'b00000000000000000010001000010001;
assign LUT_4[47633] = 32'b11111111111111111011010100001001;
assign LUT_4[47634] = 32'b00000000000000000001100010110101;
assign LUT_4[47635] = 32'b11111111111111111010101110101101;
assign LUT_4[47636] = 32'b11111111111111111111001000101101;
assign LUT_4[47637] = 32'b11111111111111111000010100100101;
assign LUT_4[47638] = 32'b11111111111111111110100011010001;
assign LUT_4[47639] = 32'b11111111111111110111101111001001;
assign LUT_4[47640] = 32'b11111111111111111011010100100110;
assign LUT_4[47641] = 32'b11111111111111110100100000011110;
assign LUT_4[47642] = 32'b11111111111111111010101111001010;
assign LUT_4[47643] = 32'b11111111111111110011111011000010;
assign LUT_4[47644] = 32'b11111111111111111000010101000010;
assign LUT_4[47645] = 32'b11111111111111110001100000111010;
assign LUT_4[47646] = 32'b11111111111111110111101111100110;
assign LUT_4[47647] = 32'b11111111111111110000111011011110;
assign LUT_4[47648] = 32'b00000000000000000010110001101010;
assign LUT_4[47649] = 32'b11111111111111111011111101100010;
assign LUT_4[47650] = 32'b00000000000000000010001100001110;
assign LUT_4[47651] = 32'b11111111111111111011011000000110;
assign LUT_4[47652] = 32'b11111111111111111111110010000110;
assign LUT_4[47653] = 32'b11111111111111111000111101111110;
assign LUT_4[47654] = 32'b11111111111111111111001100101010;
assign LUT_4[47655] = 32'b11111111111111111000011000100010;
assign LUT_4[47656] = 32'b11111111111111111011111101111111;
assign LUT_4[47657] = 32'b11111111111111110101001001110111;
assign LUT_4[47658] = 32'b11111111111111111011011000100011;
assign LUT_4[47659] = 32'b11111111111111110100100100011011;
assign LUT_4[47660] = 32'b11111111111111111000111110011011;
assign LUT_4[47661] = 32'b11111111111111110010001010010011;
assign LUT_4[47662] = 32'b11111111111111111000011000111111;
assign LUT_4[47663] = 32'b11111111111111110001100100110111;
assign LUT_4[47664] = 32'b00000000000000000000100011011000;
assign LUT_4[47665] = 32'b11111111111111111001101111010000;
assign LUT_4[47666] = 32'b11111111111111111111111101111100;
assign LUT_4[47667] = 32'b11111111111111111001001001110100;
assign LUT_4[47668] = 32'b11111111111111111101100011110100;
assign LUT_4[47669] = 32'b11111111111111110110101111101100;
assign LUT_4[47670] = 32'b11111111111111111100111110011000;
assign LUT_4[47671] = 32'b11111111111111110110001010010000;
assign LUT_4[47672] = 32'b11111111111111111001101111101101;
assign LUT_4[47673] = 32'b11111111111111110010111011100101;
assign LUT_4[47674] = 32'b11111111111111111001001010010001;
assign LUT_4[47675] = 32'b11111111111111110010010110001001;
assign LUT_4[47676] = 32'b11111111111111110110110000001001;
assign LUT_4[47677] = 32'b11111111111111101111111100000001;
assign LUT_4[47678] = 32'b11111111111111110110001010101101;
assign LUT_4[47679] = 32'b11111111111111101111010110100101;
assign LUT_4[47680] = 32'b00000000000000000101101101110111;
assign LUT_4[47681] = 32'b11111111111111111110111001101111;
assign LUT_4[47682] = 32'b00000000000000000101001000011011;
assign LUT_4[47683] = 32'b11111111111111111110010100010011;
assign LUT_4[47684] = 32'b00000000000000000010101110010011;
assign LUT_4[47685] = 32'b11111111111111111011111010001011;
assign LUT_4[47686] = 32'b00000000000000000010001000110111;
assign LUT_4[47687] = 32'b11111111111111111011010100101111;
assign LUT_4[47688] = 32'b11111111111111111110111010001100;
assign LUT_4[47689] = 32'b11111111111111111000000110000100;
assign LUT_4[47690] = 32'b11111111111111111110010100110000;
assign LUT_4[47691] = 32'b11111111111111110111100000101000;
assign LUT_4[47692] = 32'b11111111111111111011111010101000;
assign LUT_4[47693] = 32'b11111111111111110101000110100000;
assign LUT_4[47694] = 32'b11111111111111111011010101001100;
assign LUT_4[47695] = 32'b11111111111111110100100001000100;
assign LUT_4[47696] = 32'b00000000000000000011011111100101;
assign LUT_4[47697] = 32'b11111111111111111100101011011101;
assign LUT_4[47698] = 32'b00000000000000000010111010001001;
assign LUT_4[47699] = 32'b11111111111111111100000110000001;
assign LUT_4[47700] = 32'b00000000000000000000100000000001;
assign LUT_4[47701] = 32'b11111111111111111001101011111001;
assign LUT_4[47702] = 32'b11111111111111111111111010100101;
assign LUT_4[47703] = 32'b11111111111111111001000110011101;
assign LUT_4[47704] = 32'b11111111111111111100101011111010;
assign LUT_4[47705] = 32'b11111111111111110101110111110010;
assign LUT_4[47706] = 32'b11111111111111111100000110011110;
assign LUT_4[47707] = 32'b11111111111111110101010010010110;
assign LUT_4[47708] = 32'b11111111111111111001101100010110;
assign LUT_4[47709] = 32'b11111111111111110010111000001110;
assign LUT_4[47710] = 32'b11111111111111111001000110111010;
assign LUT_4[47711] = 32'b11111111111111110010010010110010;
assign LUT_4[47712] = 32'b00000000000000000100001000111110;
assign LUT_4[47713] = 32'b11111111111111111101010100110110;
assign LUT_4[47714] = 32'b00000000000000000011100011100010;
assign LUT_4[47715] = 32'b11111111111111111100101111011010;
assign LUT_4[47716] = 32'b00000000000000000001001001011010;
assign LUT_4[47717] = 32'b11111111111111111010010101010010;
assign LUT_4[47718] = 32'b00000000000000000000100011111110;
assign LUT_4[47719] = 32'b11111111111111111001101111110110;
assign LUT_4[47720] = 32'b11111111111111111101010101010011;
assign LUT_4[47721] = 32'b11111111111111110110100001001011;
assign LUT_4[47722] = 32'b11111111111111111100101111110111;
assign LUT_4[47723] = 32'b11111111111111110101111011101111;
assign LUT_4[47724] = 32'b11111111111111111010010101101111;
assign LUT_4[47725] = 32'b11111111111111110011100001100111;
assign LUT_4[47726] = 32'b11111111111111111001110000010011;
assign LUT_4[47727] = 32'b11111111111111110010111100001011;
assign LUT_4[47728] = 32'b00000000000000000001111010101100;
assign LUT_4[47729] = 32'b11111111111111111011000110100100;
assign LUT_4[47730] = 32'b00000000000000000001010101010000;
assign LUT_4[47731] = 32'b11111111111111111010100001001000;
assign LUT_4[47732] = 32'b11111111111111111110111011001000;
assign LUT_4[47733] = 32'b11111111111111111000000111000000;
assign LUT_4[47734] = 32'b11111111111111111110010101101100;
assign LUT_4[47735] = 32'b11111111111111110111100001100100;
assign LUT_4[47736] = 32'b11111111111111111011000111000001;
assign LUT_4[47737] = 32'b11111111111111110100010010111001;
assign LUT_4[47738] = 32'b11111111111111111010100001100101;
assign LUT_4[47739] = 32'b11111111111111110011101101011101;
assign LUT_4[47740] = 32'b11111111111111111000000111011101;
assign LUT_4[47741] = 32'b11111111111111110001010011010101;
assign LUT_4[47742] = 32'b11111111111111110111100010000001;
assign LUT_4[47743] = 32'b11111111111111110000101101111001;
assign LUT_4[47744] = 32'b00000000000000000110111100101011;
assign LUT_4[47745] = 32'b00000000000000000000001000100011;
assign LUT_4[47746] = 32'b00000000000000000110010111001111;
assign LUT_4[47747] = 32'b11111111111111111111100011000111;
assign LUT_4[47748] = 32'b00000000000000000011111101000111;
assign LUT_4[47749] = 32'b11111111111111111101001000111111;
assign LUT_4[47750] = 32'b00000000000000000011010111101011;
assign LUT_4[47751] = 32'b11111111111111111100100011100011;
assign LUT_4[47752] = 32'b00000000000000000000001001000000;
assign LUT_4[47753] = 32'b11111111111111111001010100111000;
assign LUT_4[47754] = 32'b11111111111111111111100011100100;
assign LUT_4[47755] = 32'b11111111111111111000101111011100;
assign LUT_4[47756] = 32'b11111111111111111101001001011100;
assign LUT_4[47757] = 32'b11111111111111110110010101010100;
assign LUT_4[47758] = 32'b11111111111111111100100100000000;
assign LUT_4[47759] = 32'b11111111111111110101101111111000;
assign LUT_4[47760] = 32'b00000000000000000100101110011001;
assign LUT_4[47761] = 32'b11111111111111111101111010010001;
assign LUT_4[47762] = 32'b00000000000000000100001000111101;
assign LUT_4[47763] = 32'b11111111111111111101010100110101;
assign LUT_4[47764] = 32'b00000000000000000001101110110101;
assign LUT_4[47765] = 32'b11111111111111111010111010101101;
assign LUT_4[47766] = 32'b00000000000000000001001001011001;
assign LUT_4[47767] = 32'b11111111111111111010010101010001;
assign LUT_4[47768] = 32'b11111111111111111101111010101110;
assign LUT_4[47769] = 32'b11111111111111110111000110100110;
assign LUT_4[47770] = 32'b11111111111111111101010101010010;
assign LUT_4[47771] = 32'b11111111111111110110100001001010;
assign LUT_4[47772] = 32'b11111111111111111010111011001010;
assign LUT_4[47773] = 32'b11111111111111110100000111000010;
assign LUT_4[47774] = 32'b11111111111111111010010101101110;
assign LUT_4[47775] = 32'b11111111111111110011100001100110;
assign LUT_4[47776] = 32'b00000000000000000101010111110010;
assign LUT_4[47777] = 32'b11111111111111111110100011101010;
assign LUT_4[47778] = 32'b00000000000000000100110010010110;
assign LUT_4[47779] = 32'b11111111111111111101111110001110;
assign LUT_4[47780] = 32'b00000000000000000010011000001110;
assign LUT_4[47781] = 32'b11111111111111111011100100000110;
assign LUT_4[47782] = 32'b00000000000000000001110010110010;
assign LUT_4[47783] = 32'b11111111111111111010111110101010;
assign LUT_4[47784] = 32'b11111111111111111110100100000111;
assign LUT_4[47785] = 32'b11111111111111110111101111111111;
assign LUT_4[47786] = 32'b11111111111111111101111110101011;
assign LUT_4[47787] = 32'b11111111111111110111001010100011;
assign LUT_4[47788] = 32'b11111111111111111011100100100011;
assign LUT_4[47789] = 32'b11111111111111110100110000011011;
assign LUT_4[47790] = 32'b11111111111111111010111111000111;
assign LUT_4[47791] = 32'b11111111111111110100001010111111;
assign LUT_4[47792] = 32'b00000000000000000011001001100000;
assign LUT_4[47793] = 32'b11111111111111111100010101011000;
assign LUT_4[47794] = 32'b00000000000000000010100100000100;
assign LUT_4[47795] = 32'b11111111111111111011101111111100;
assign LUT_4[47796] = 32'b00000000000000000000001001111100;
assign LUT_4[47797] = 32'b11111111111111111001010101110100;
assign LUT_4[47798] = 32'b11111111111111111111100100100000;
assign LUT_4[47799] = 32'b11111111111111111000110000011000;
assign LUT_4[47800] = 32'b11111111111111111100010101110101;
assign LUT_4[47801] = 32'b11111111111111110101100001101101;
assign LUT_4[47802] = 32'b11111111111111111011110000011001;
assign LUT_4[47803] = 32'b11111111111111110100111100010001;
assign LUT_4[47804] = 32'b11111111111111111001010110010001;
assign LUT_4[47805] = 32'b11111111111111110010100010001001;
assign LUT_4[47806] = 32'b11111111111111111000110000110101;
assign LUT_4[47807] = 32'b11111111111111110001111100101101;
assign LUT_4[47808] = 32'b00000000000000001000010011111111;
assign LUT_4[47809] = 32'b00000000000000000001011111110111;
assign LUT_4[47810] = 32'b00000000000000000111101110100011;
assign LUT_4[47811] = 32'b00000000000000000000111010011011;
assign LUT_4[47812] = 32'b00000000000000000101010100011011;
assign LUT_4[47813] = 32'b11111111111111111110100000010011;
assign LUT_4[47814] = 32'b00000000000000000100101110111111;
assign LUT_4[47815] = 32'b11111111111111111101111010110111;
assign LUT_4[47816] = 32'b00000000000000000001100000010100;
assign LUT_4[47817] = 32'b11111111111111111010101100001100;
assign LUT_4[47818] = 32'b00000000000000000000111010111000;
assign LUT_4[47819] = 32'b11111111111111111010000110110000;
assign LUT_4[47820] = 32'b11111111111111111110100000110000;
assign LUT_4[47821] = 32'b11111111111111110111101100101000;
assign LUT_4[47822] = 32'b11111111111111111101111011010100;
assign LUT_4[47823] = 32'b11111111111111110111000111001100;
assign LUT_4[47824] = 32'b00000000000000000110000101101101;
assign LUT_4[47825] = 32'b11111111111111111111010001100101;
assign LUT_4[47826] = 32'b00000000000000000101100000010001;
assign LUT_4[47827] = 32'b11111111111111111110101100001001;
assign LUT_4[47828] = 32'b00000000000000000011000110001001;
assign LUT_4[47829] = 32'b11111111111111111100010010000001;
assign LUT_4[47830] = 32'b00000000000000000010100000101101;
assign LUT_4[47831] = 32'b11111111111111111011101100100101;
assign LUT_4[47832] = 32'b11111111111111111111010010000010;
assign LUT_4[47833] = 32'b11111111111111111000011101111010;
assign LUT_4[47834] = 32'b11111111111111111110101100100110;
assign LUT_4[47835] = 32'b11111111111111110111111000011110;
assign LUT_4[47836] = 32'b11111111111111111100010010011110;
assign LUT_4[47837] = 32'b11111111111111110101011110010110;
assign LUT_4[47838] = 32'b11111111111111111011101101000010;
assign LUT_4[47839] = 32'b11111111111111110100111000111010;
assign LUT_4[47840] = 32'b00000000000000000110101111000110;
assign LUT_4[47841] = 32'b11111111111111111111111010111110;
assign LUT_4[47842] = 32'b00000000000000000110001001101010;
assign LUT_4[47843] = 32'b11111111111111111111010101100010;
assign LUT_4[47844] = 32'b00000000000000000011101111100010;
assign LUT_4[47845] = 32'b11111111111111111100111011011010;
assign LUT_4[47846] = 32'b00000000000000000011001010000110;
assign LUT_4[47847] = 32'b11111111111111111100010101111110;
assign LUT_4[47848] = 32'b11111111111111111111111011011011;
assign LUT_4[47849] = 32'b11111111111111111001000111010011;
assign LUT_4[47850] = 32'b11111111111111111111010101111111;
assign LUT_4[47851] = 32'b11111111111111111000100001110111;
assign LUT_4[47852] = 32'b11111111111111111100111011110111;
assign LUT_4[47853] = 32'b11111111111111110110000111101111;
assign LUT_4[47854] = 32'b11111111111111111100010110011011;
assign LUT_4[47855] = 32'b11111111111111110101100010010011;
assign LUT_4[47856] = 32'b00000000000000000100100000110100;
assign LUT_4[47857] = 32'b11111111111111111101101100101100;
assign LUT_4[47858] = 32'b00000000000000000011111011011000;
assign LUT_4[47859] = 32'b11111111111111111101000111010000;
assign LUT_4[47860] = 32'b00000000000000000001100001010000;
assign LUT_4[47861] = 32'b11111111111111111010101101001000;
assign LUT_4[47862] = 32'b00000000000000000000111011110100;
assign LUT_4[47863] = 32'b11111111111111111010000111101100;
assign LUT_4[47864] = 32'b11111111111111111101101101001001;
assign LUT_4[47865] = 32'b11111111111111110110111001000001;
assign LUT_4[47866] = 32'b11111111111111111101000111101101;
assign LUT_4[47867] = 32'b11111111111111110110010011100101;
assign LUT_4[47868] = 32'b11111111111111111010101101100101;
assign LUT_4[47869] = 32'b11111111111111110011111001011101;
assign LUT_4[47870] = 32'b11111111111111111010001000001001;
assign LUT_4[47871] = 32'b11111111111111110011010100000001;
assign LUT_4[47872] = 32'b00000000000000001001010010000110;
assign LUT_4[47873] = 32'b00000000000000000010011101111110;
assign LUT_4[47874] = 32'b00000000000000001000101100101010;
assign LUT_4[47875] = 32'b00000000000000000001111000100010;
assign LUT_4[47876] = 32'b00000000000000000110010010100010;
assign LUT_4[47877] = 32'b11111111111111111111011110011010;
assign LUT_4[47878] = 32'b00000000000000000101101101000110;
assign LUT_4[47879] = 32'b11111111111111111110111000111110;
assign LUT_4[47880] = 32'b00000000000000000010011110011011;
assign LUT_4[47881] = 32'b11111111111111111011101010010011;
assign LUT_4[47882] = 32'b00000000000000000001111000111111;
assign LUT_4[47883] = 32'b11111111111111111011000100110111;
assign LUT_4[47884] = 32'b11111111111111111111011110110111;
assign LUT_4[47885] = 32'b11111111111111111000101010101111;
assign LUT_4[47886] = 32'b11111111111111111110111001011011;
assign LUT_4[47887] = 32'b11111111111111111000000101010011;
assign LUT_4[47888] = 32'b00000000000000000111000011110100;
assign LUT_4[47889] = 32'b00000000000000000000001111101100;
assign LUT_4[47890] = 32'b00000000000000000110011110011000;
assign LUT_4[47891] = 32'b11111111111111111111101010010000;
assign LUT_4[47892] = 32'b00000000000000000100000100010000;
assign LUT_4[47893] = 32'b11111111111111111101010000001000;
assign LUT_4[47894] = 32'b00000000000000000011011110110100;
assign LUT_4[47895] = 32'b11111111111111111100101010101100;
assign LUT_4[47896] = 32'b00000000000000000000010000001001;
assign LUT_4[47897] = 32'b11111111111111111001011100000001;
assign LUT_4[47898] = 32'b11111111111111111111101010101101;
assign LUT_4[47899] = 32'b11111111111111111000110110100101;
assign LUT_4[47900] = 32'b11111111111111111101010000100101;
assign LUT_4[47901] = 32'b11111111111111110110011100011101;
assign LUT_4[47902] = 32'b11111111111111111100101011001001;
assign LUT_4[47903] = 32'b11111111111111110101110111000001;
assign LUT_4[47904] = 32'b00000000000000000111101101001101;
assign LUT_4[47905] = 32'b00000000000000000000111001000101;
assign LUT_4[47906] = 32'b00000000000000000111000111110001;
assign LUT_4[47907] = 32'b00000000000000000000010011101001;
assign LUT_4[47908] = 32'b00000000000000000100101101101001;
assign LUT_4[47909] = 32'b11111111111111111101111001100001;
assign LUT_4[47910] = 32'b00000000000000000100001000001101;
assign LUT_4[47911] = 32'b11111111111111111101010100000101;
assign LUT_4[47912] = 32'b00000000000000000000111001100010;
assign LUT_4[47913] = 32'b11111111111111111010000101011010;
assign LUT_4[47914] = 32'b00000000000000000000010100000110;
assign LUT_4[47915] = 32'b11111111111111111001011111111110;
assign LUT_4[47916] = 32'b11111111111111111101111001111110;
assign LUT_4[47917] = 32'b11111111111111110111000101110110;
assign LUT_4[47918] = 32'b11111111111111111101010100100010;
assign LUT_4[47919] = 32'b11111111111111110110100000011010;
assign LUT_4[47920] = 32'b00000000000000000101011110111011;
assign LUT_4[47921] = 32'b11111111111111111110101010110011;
assign LUT_4[47922] = 32'b00000000000000000100111001011111;
assign LUT_4[47923] = 32'b11111111111111111110000101010111;
assign LUT_4[47924] = 32'b00000000000000000010011111010111;
assign LUT_4[47925] = 32'b11111111111111111011101011001111;
assign LUT_4[47926] = 32'b00000000000000000001111001111011;
assign LUT_4[47927] = 32'b11111111111111111011000101110011;
assign LUT_4[47928] = 32'b11111111111111111110101011010000;
assign LUT_4[47929] = 32'b11111111111111110111110111001000;
assign LUT_4[47930] = 32'b11111111111111111110000101110100;
assign LUT_4[47931] = 32'b11111111111111110111010001101100;
assign LUT_4[47932] = 32'b11111111111111111011101011101100;
assign LUT_4[47933] = 32'b11111111111111110100110111100100;
assign LUT_4[47934] = 32'b11111111111111111011000110010000;
assign LUT_4[47935] = 32'b11111111111111110100010010001000;
assign LUT_4[47936] = 32'b00000000000000001010101001011010;
assign LUT_4[47937] = 32'b00000000000000000011110101010010;
assign LUT_4[47938] = 32'b00000000000000001010000011111110;
assign LUT_4[47939] = 32'b00000000000000000011001111110110;
assign LUT_4[47940] = 32'b00000000000000000111101001110110;
assign LUT_4[47941] = 32'b00000000000000000000110101101110;
assign LUT_4[47942] = 32'b00000000000000000111000100011010;
assign LUT_4[47943] = 32'b00000000000000000000010000010010;
assign LUT_4[47944] = 32'b00000000000000000011110101101111;
assign LUT_4[47945] = 32'b11111111111111111101000001100111;
assign LUT_4[47946] = 32'b00000000000000000011010000010011;
assign LUT_4[47947] = 32'b11111111111111111100011100001011;
assign LUT_4[47948] = 32'b00000000000000000000110110001011;
assign LUT_4[47949] = 32'b11111111111111111010000010000011;
assign LUT_4[47950] = 32'b00000000000000000000010000101111;
assign LUT_4[47951] = 32'b11111111111111111001011100100111;
assign LUT_4[47952] = 32'b00000000000000001000011011001000;
assign LUT_4[47953] = 32'b00000000000000000001100111000000;
assign LUT_4[47954] = 32'b00000000000000000111110101101100;
assign LUT_4[47955] = 32'b00000000000000000001000001100100;
assign LUT_4[47956] = 32'b00000000000000000101011011100100;
assign LUT_4[47957] = 32'b11111111111111111110100111011100;
assign LUT_4[47958] = 32'b00000000000000000100110110001000;
assign LUT_4[47959] = 32'b11111111111111111110000010000000;
assign LUT_4[47960] = 32'b00000000000000000001100111011101;
assign LUT_4[47961] = 32'b11111111111111111010110011010101;
assign LUT_4[47962] = 32'b00000000000000000001000010000001;
assign LUT_4[47963] = 32'b11111111111111111010001101111001;
assign LUT_4[47964] = 32'b11111111111111111110100111111001;
assign LUT_4[47965] = 32'b11111111111111110111110011110001;
assign LUT_4[47966] = 32'b11111111111111111110000010011101;
assign LUT_4[47967] = 32'b11111111111111110111001110010101;
assign LUT_4[47968] = 32'b00000000000000001001000100100001;
assign LUT_4[47969] = 32'b00000000000000000010010000011001;
assign LUT_4[47970] = 32'b00000000000000001000011111000101;
assign LUT_4[47971] = 32'b00000000000000000001101010111101;
assign LUT_4[47972] = 32'b00000000000000000110000100111101;
assign LUT_4[47973] = 32'b11111111111111111111010000110101;
assign LUT_4[47974] = 32'b00000000000000000101011111100001;
assign LUT_4[47975] = 32'b11111111111111111110101011011001;
assign LUT_4[47976] = 32'b00000000000000000010010000110110;
assign LUT_4[47977] = 32'b11111111111111111011011100101110;
assign LUT_4[47978] = 32'b00000000000000000001101011011010;
assign LUT_4[47979] = 32'b11111111111111111010110111010010;
assign LUT_4[47980] = 32'b11111111111111111111010001010010;
assign LUT_4[47981] = 32'b11111111111111111000011101001010;
assign LUT_4[47982] = 32'b11111111111111111110101011110110;
assign LUT_4[47983] = 32'b11111111111111110111110111101110;
assign LUT_4[47984] = 32'b00000000000000000110110110001111;
assign LUT_4[47985] = 32'b00000000000000000000000010000111;
assign LUT_4[47986] = 32'b00000000000000000110010000110011;
assign LUT_4[47987] = 32'b11111111111111111111011100101011;
assign LUT_4[47988] = 32'b00000000000000000011110110101011;
assign LUT_4[47989] = 32'b11111111111111111101000010100011;
assign LUT_4[47990] = 32'b00000000000000000011010001001111;
assign LUT_4[47991] = 32'b11111111111111111100011101000111;
assign LUT_4[47992] = 32'b00000000000000000000000010100100;
assign LUT_4[47993] = 32'b11111111111111111001001110011100;
assign LUT_4[47994] = 32'b11111111111111111111011101001000;
assign LUT_4[47995] = 32'b11111111111111111000101001000000;
assign LUT_4[47996] = 32'b11111111111111111101000011000000;
assign LUT_4[47997] = 32'b11111111111111110110001110111000;
assign LUT_4[47998] = 32'b11111111111111111100011101100100;
assign LUT_4[47999] = 32'b11111111111111110101101001011100;
assign LUT_4[48000] = 32'b00000000000000001011111000001110;
assign LUT_4[48001] = 32'b00000000000000000101000100000110;
assign LUT_4[48002] = 32'b00000000000000001011010010110010;
assign LUT_4[48003] = 32'b00000000000000000100011110101010;
assign LUT_4[48004] = 32'b00000000000000001000111000101010;
assign LUT_4[48005] = 32'b00000000000000000010000100100010;
assign LUT_4[48006] = 32'b00000000000000001000010011001110;
assign LUT_4[48007] = 32'b00000000000000000001011111000110;
assign LUT_4[48008] = 32'b00000000000000000101000100100011;
assign LUT_4[48009] = 32'b11111111111111111110010000011011;
assign LUT_4[48010] = 32'b00000000000000000100011111000111;
assign LUT_4[48011] = 32'b11111111111111111101101010111111;
assign LUT_4[48012] = 32'b00000000000000000010000100111111;
assign LUT_4[48013] = 32'b11111111111111111011010000110111;
assign LUT_4[48014] = 32'b00000000000000000001011111100011;
assign LUT_4[48015] = 32'b11111111111111111010101011011011;
assign LUT_4[48016] = 32'b00000000000000001001101001111100;
assign LUT_4[48017] = 32'b00000000000000000010110101110100;
assign LUT_4[48018] = 32'b00000000000000001001000100100000;
assign LUT_4[48019] = 32'b00000000000000000010010000011000;
assign LUT_4[48020] = 32'b00000000000000000110101010011000;
assign LUT_4[48021] = 32'b11111111111111111111110110010000;
assign LUT_4[48022] = 32'b00000000000000000110000100111100;
assign LUT_4[48023] = 32'b11111111111111111111010000110100;
assign LUT_4[48024] = 32'b00000000000000000010110110010001;
assign LUT_4[48025] = 32'b11111111111111111100000010001001;
assign LUT_4[48026] = 32'b00000000000000000010010000110101;
assign LUT_4[48027] = 32'b11111111111111111011011100101101;
assign LUT_4[48028] = 32'b11111111111111111111110110101101;
assign LUT_4[48029] = 32'b11111111111111111001000010100101;
assign LUT_4[48030] = 32'b11111111111111111111010001010001;
assign LUT_4[48031] = 32'b11111111111111111000011101001001;
assign LUT_4[48032] = 32'b00000000000000001010010011010101;
assign LUT_4[48033] = 32'b00000000000000000011011111001101;
assign LUT_4[48034] = 32'b00000000000000001001101101111001;
assign LUT_4[48035] = 32'b00000000000000000010111001110001;
assign LUT_4[48036] = 32'b00000000000000000111010011110001;
assign LUT_4[48037] = 32'b00000000000000000000011111101001;
assign LUT_4[48038] = 32'b00000000000000000110101110010101;
assign LUT_4[48039] = 32'b11111111111111111111111010001101;
assign LUT_4[48040] = 32'b00000000000000000011011111101010;
assign LUT_4[48041] = 32'b11111111111111111100101011100010;
assign LUT_4[48042] = 32'b00000000000000000010111010001110;
assign LUT_4[48043] = 32'b11111111111111111100000110000110;
assign LUT_4[48044] = 32'b00000000000000000000100000000110;
assign LUT_4[48045] = 32'b11111111111111111001101011111110;
assign LUT_4[48046] = 32'b11111111111111111111111010101010;
assign LUT_4[48047] = 32'b11111111111111111001000110100010;
assign LUT_4[48048] = 32'b00000000000000001000000101000011;
assign LUT_4[48049] = 32'b00000000000000000001010000111011;
assign LUT_4[48050] = 32'b00000000000000000111011111100111;
assign LUT_4[48051] = 32'b00000000000000000000101011011111;
assign LUT_4[48052] = 32'b00000000000000000101000101011111;
assign LUT_4[48053] = 32'b11111111111111111110010001010111;
assign LUT_4[48054] = 32'b00000000000000000100100000000011;
assign LUT_4[48055] = 32'b11111111111111111101101011111011;
assign LUT_4[48056] = 32'b00000000000000000001010001011000;
assign LUT_4[48057] = 32'b11111111111111111010011101010000;
assign LUT_4[48058] = 32'b00000000000000000000101011111100;
assign LUT_4[48059] = 32'b11111111111111111001110111110100;
assign LUT_4[48060] = 32'b11111111111111111110010001110100;
assign LUT_4[48061] = 32'b11111111111111110111011101101100;
assign LUT_4[48062] = 32'b11111111111111111101101100011000;
assign LUT_4[48063] = 32'b11111111111111110110111000010000;
assign LUT_4[48064] = 32'b00000000000000001101001111100010;
assign LUT_4[48065] = 32'b00000000000000000110011011011010;
assign LUT_4[48066] = 32'b00000000000000001100101010000110;
assign LUT_4[48067] = 32'b00000000000000000101110101111110;
assign LUT_4[48068] = 32'b00000000000000001010001111111110;
assign LUT_4[48069] = 32'b00000000000000000011011011110110;
assign LUT_4[48070] = 32'b00000000000000001001101010100010;
assign LUT_4[48071] = 32'b00000000000000000010110110011010;
assign LUT_4[48072] = 32'b00000000000000000110011011110111;
assign LUT_4[48073] = 32'b11111111111111111111100111101111;
assign LUT_4[48074] = 32'b00000000000000000101110110011011;
assign LUT_4[48075] = 32'b11111111111111111111000010010011;
assign LUT_4[48076] = 32'b00000000000000000011011100010011;
assign LUT_4[48077] = 32'b11111111111111111100101000001011;
assign LUT_4[48078] = 32'b00000000000000000010110110110111;
assign LUT_4[48079] = 32'b11111111111111111100000010101111;
assign LUT_4[48080] = 32'b00000000000000001011000001010000;
assign LUT_4[48081] = 32'b00000000000000000100001101001000;
assign LUT_4[48082] = 32'b00000000000000001010011011110100;
assign LUT_4[48083] = 32'b00000000000000000011100111101100;
assign LUT_4[48084] = 32'b00000000000000001000000001101100;
assign LUT_4[48085] = 32'b00000000000000000001001101100100;
assign LUT_4[48086] = 32'b00000000000000000111011100010000;
assign LUT_4[48087] = 32'b00000000000000000000101000001000;
assign LUT_4[48088] = 32'b00000000000000000100001101100101;
assign LUT_4[48089] = 32'b11111111111111111101011001011101;
assign LUT_4[48090] = 32'b00000000000000000011101000001001;
assign LUT_4[48091] = 32'b11111111111111111100110100000001;
assign LUT_4[48092] = 32'b00000000000000000001001110000001;
assign LUT_4[48093] = 32'b11111111111111111010011001111001;
assign LUT_4[48094] = 32'b00000000000000000000101000100101;
assign LUT_4[48095] = 32'b11111111111111111001110100011101;
assign LUT_4[48096] = 32'b00000000000000001011101010101001;
assign LUT_4[48097] = 32'b00000000000000000100110110100001;
assign LUT_4[48098] = 32'b00000000000000001011000101001101;
assign LUT_4[48099] = 32'b00000000000000000100010001000101;
assign LUT_4[48100] = 32'b00000000000000001000101011000101;
assign LUT_4[48101] = 32'b00000000000000000001110110111101;
assign LUT_4[48102] = 32'b00000000000000001000000101101001;
assign LUT_4[48103] = 32'b00000000000000000001010001100001;
assign LUT_4[48104] = 32'b00000000000000000100110110111110;
assign LUT_4[48105] = 32'b11111111111111111110000010110110;
assign LUT_4[48106] = 32'b00000000000000000100010001100010;
assign LUT_4[48107] = 32'b11111111111111111101011101011010;
assign LUT_4[48108] = 32'b00000000000000000001110111011010;
assign LUT_4[48109] = 32'b11111111111111111011000011010010;
assign LUT_4[48110] = 32'b00000000000000000001010001111110;
assign LUT_4[48111] = 32'b11111111111111111010011101110110;
assign LUT_4[48112] = 32'b00000000000000001001011100010111;
assign LUT_4[48113] = 32'b00000000000000000010101000001111;
assign LUT_4[48114] = 32'b00000000000000001000110110111011;
assign LUT_4[48115] = 32'b00000000000000000010000010110011;
assign LUT_4[48116] = 32'b00000000000000000110011100110011;
assign LUT_4[48117] = 32'b11111111111111111111101000101011;
assign LUT_4[48118] = 32'b00000000000000000101110111010111;
assign LUT_4[48119] = 32'b11111111111111111111000011001111;
assign LUT_4[48120] = 32'b00000000000000000010101000101100;
assign LUT_4[48121] = 32'b11111111111111111011110100100100;
assign LUT_4[48122] = 32'b00000000000000000010000011010000;
assign LUT_4[48123] = 32'b11111111111111111011001111001000;
assign LUT_4[48124] = 32'b11111111111111111111101001001000;
assign LUT_4[48125] = 32'b11111111111111111000110101000000;
assign LUT_4[48126] = 32'b11111111111111111111000011101100;
assign LUT_4[48127] = 32'b11111111111111111000001111100100;
assign LUT_4[48128] = 32'b00000000000000000110111100111010;
assign LUT_4[48129] = 32'b00000000000000000000001000110010;
assign LUT_4[48130] = 32'b00000000000000000110010111011110;
assign LUT_4[48131] = 32'b11111111111111111111100011010110;
assign LUT_4[48132] = 32'b00000000000000000011111101010110;
assign LUT_4[48133] = 32'b11111111111111111101001001001110;
assign LUT_4[48134] = 32'b00000000000000000011010111111010;
assign LUT_4[48135] = 32'b11111111111111111100100011110010;
assign LUT_4[48136] = 32'b00000000000000000000001001001111;
assign LUT_4[48137] = 32'b11111111111111111001010101000111;
assign LUT_4[48138] = 32'b11111111111111111111100011110011;
assign LUT_4[48139] = 32'b11111111111111111000101111101011;
assign LUT_4[48140] = 32'b11111111111111111101001001101011;
assign LUT_4[48141] = 32'b11111111111111110110010101100011;
assign LUT_4[48142] = 32'b11111111111111111100100100001111;
assign LUT_4[48143] = 32'b11111111111111110101110000000111;
assign LUT_4[48144] = 32'b00000000000000000100101110101000;
assign LUT_4[48145] = 32'b11111111111111111101111010100000;
assign LUT_4[48146] = 32'b00000000000000000100001001001100;
assign LUT_4[48147] = 32'b11111111111111111101010101000100;
assign LUT_4[48148] = 32'b00000000000000000001101111000100;
assign LUT_4[48149] = 32'b11111111111111111010111010111100;
assign LUT_4[48150] = 32'b00000000000000000001001001101000;
assign LUT_4[48151] = 32'b11111111111111111010010101100000;
assign LUT_4[48152] = 32'b11111111111111111101111010111101;
assign LUT_4[48153] = 32'b11111111111111110111000110110101;
assign LUT_4[48154] = 32'b11111111111111111101010101100001;
assign LUT_4[48155] = 32'b11111111111111110110100001011001;
assign LUT_4[48156] = 32'b11111111111111111010111011011001;
assign LUT_4[48157] = 32'b11111111111111110100000111010001;
assign LUT_4[48158] = 32'b11111111111111111010010101111101;
assign LUT_4[48159] = 32'b11111111111111110011100001110101;
assign LUT_4[48160] = 32'b00000000000000000101011000000001;
assign LUT_4[48161] = 32'b11111111111111111110100011111001;
assign LUT_4[48162] = 32'b00000000000000000100110010100101;
assign LUT_4[48163] = 32'b11111111111111111101111110011101;
assign LUT_4[48164] = 32'b00000000000000000010011000011101;
assign LUT_4[48165] = 32'b11111111111111111011100100010101;
assign LUT_4[48166] = 32'b00000000000000000001110011000001;
assign LUT_4[48167] = 32'b11111111111111111010111110111001;
assign LUT_4[48168] = 32'b11111111111111111110100100010110;
assign LUT_4[48169] = 32'b11111111111111110111110000001110;
assign LUT_4[48170] = 32'b11111111111111111101111110111010;
assign LUT_4[48171] = 32'b11111111111111110111001010110010;
assign LUT_4[48172] = 32'b11111111111111111011100100110010;
assign LUT_4[48173] = 32'b11111111111111110100110000101010;
assign LUT_4[48174] = 32'b11111111111111111010111111010110;
assign LUT_4[48175] = 32'b11111111111111110100001011001110;
assign LUT_4[48176] = 32'b00000000000000000011001001101111;
assign LUT_4[48177] = 32'b11111111111111111100010101100111;
assign LUT_4[48178] = 32'b00000000000000000010100100010011;
assign LUT_4[48179] = 32'b11111111111111111011110000001011;
assign LUT_4[48180] = 32'b00000000000000000000001010001011;
assign LUT_4[48181] = 32'b11111111111111111001010110000011;
assign LUT_4[48182] = 32'b11111111111111111111100100101111;
assign LUT_4[48183] = 32'b11111111111111111000110000100111;
assign LUT_4[48184] = 32'b11111111111111111100010110000100;
assign LUT_4[48185] = 32'b11111111111111110101100001111100;
assign LUT_4[48186] = 32'b11111111111111111011110000101000;
assign LUT_4[48187] = 32'b11111111111111110100111100100000;
assign LUT_4[48188] = 32'b11111111111111111001010110100000;
assign LUT_4[48189] = 32'b11111111111111110010100010011000;
assign LUT_4[48190] = 32'b11111111111111111000110001000100;
assign LUT_4[48191] = 32'b11111111111111110001111100111100;
assign LUT_4[48192] = 32'b00000000000000001000010100001110;
assign LUT_4[48193] = 32'b00000000000000000001100000000110;
assign LUT_4[48194] = 32'b00000000000000000111101110110010;
assign LUT_4[48195] = 32'b00000000000000000000111010101010;
assign LUT_4[48196] = 32'b00000000000000000101010100101010;
assign LUT_4[48197] = 32'b11111111111111111110100000100010;
assign LUT_4[48198] = 32'b00000000000000000100101111001110;
assign LUT_4[48199] = 32'b11111111111111111101111011000110;
assign LUT_4[48200] = 32'b00000000000000000001100000100011;
assign LUT_4[48201] = 32'b11111111111111111010101100011011;
assign LUT_4[48202] = 32'b00000000000000000000111011000111;
assign LUT_4[48203] = 32'b11111111111111111010000110111111;
assign LUT_4[48204] = 32'b11111111111111111110100000111111;
assign LUT_4[48205] = 32'b11111111111111110111101100110111;
assign LUT_4[48206] = 32'b11111111111111111101111011100011;
assign LUT_4[48207] = 32'b11111111111111110111000111011011;
assign LUT_4[48208] = 32'b00000000000000000110000101111100;
assign LUT_4[48209] = 32'b11111111111111111111010001110100;
assign LUT_4[48210] = 32'b00000000000000000101100000100000;
assign LUT_4[48211] = 32'b11111111111111111110101100011000;
assign LUT_4[48212] = 32'b00000000000000000011000110011000;
assign LUT_4[48213] = 32'b11111111111111111100010010010000;
assign LUT_4[48214] = 32'b00000000000000000010100000111100;
assign LUT_4[48215] = 32'b11111111111111111011101100110100;
assign LUT_4[48216] = 32'b11111111111111111111010010010001;
assign LUT_4[48217] = 32'b11111111111111111000011110001001;
assign LUT_4[48218] = 32'b11111111111111111110101100110101;
assign LUT_4[48219] = 32'b11111111111111110111111000101101;
assign LUT_4[48220] = 32'b11111111111111111100010010101101;
assign LUT_4[48221] = 32'b11111111111111110101011110100101;
assign LUT_4[48222] = 32'b11111111111111111011101101010001;
assign LUT_4[48223] = 32'b11111111111111110100111001001001;
assign LUT_4[48224] = 32'b00000000000000000110101111010101;
assign LUT_4[48225] = 32'b11111111111111111111111011001101;
assign LUT_4[48226] = 32'b00000000000000000110001001111001;
assign LUT_4[48227] = 32'b11111111111111111111010101110001;
assign LUT_4[48228] = 32'b00000000000000000011101111110001;
assign LUT_4[48229] = 32'b11111111111111111100111011101001;
assign LUT_4[48230] = 32'b00000000000000000011001010010101;
assign LUT_4[48231] = 32'b11111111111111111100010110001101;
assign LUT_4[48232] = 32'b11111111111111111111111011101010;
assign LUT_4[48233] = 32'b11111111111111111001000111100010;
assign LUT_4[48234] = 32'b11111111111111111111010110001110;
assign LUT_4[48235] = 32'b11111111111111111000100010000110;
assign LUT_4[48236] = 32'b11111111111111111100111100000110;
assign LUT_4[48237] = 32'b11111111111111110110000111111110;
assign LUT_4[48238] = 32'b11111111111111111100010110101010;
assign LUT_4[48239] = 32'b11111111111111110101100010100010;
assign LUT_4[48240] = 32'b00000000000000000100100001000011;
assign LUT_4[48241] = 32'b11111111111111111101101100111011;
assign LUT_4[48242] = 32'b00000000000000000011111011100111;
assign LUT_4[48243] = 32'b11111111111111111101000111011111;
assign LUT_4[48244] = 32'b00000000000000000001100001011111;
assign LUT_4[48245] = 32'b11111111111111111010101101010111;
assign LUT_4[48246] = 32'b00000000000000000000111100000011;
assign LUT_4[48247] = 32'b11111111111111111010000111111011;
assign LUT_4[48248] = 32'b11111111111111111101101101011000;
assign LUT_4[48249] = 32'b11111111111111110110111001010000;
assign LUT_4[48250] = 32'b11111111111111111101000111111100;
assign LUT_4[48251] = 32'b11111111111111110110010011110100;
assign LUT_4[48252] = 32'b11111111111111111010101101110100;
assign LUT_4[48253] = 32'b11111111111111110011111001101100;
assign LUT_4[48254] = 32'b11111111111111111010001000011000;
assign LUT_4[48255] = 32'b11111111111111110011010100010000;
assign LUT_4[48256] = 32'b00000000000000001001100011000010;
assign LUT_4[48257] = 32'b00000000000000000010101110111010;
assign LUT_4[48258] = 32'b00000000000000001000111101100110;
assign LUT_4[48259] = 32'b00000000000000000010001001011110;
assign LUT_4[48260] = 32'b00000000000000000110100011011110;
assign LUT_4[48261] = 32'b11111111111111111111101111010110;
assign LUT_4[48262] = 32'b00000000000000000101111110000010;
assign LUT_4[48263] = 32'b11111111111111111111001001111010;
assign LUT_4[48264] = 32'b00000000000000000010101111010111;
assign LUT_4[48265] = 32'b11111111111111111011111011001111;
assign LUT_4[48266] = 32'b00000000000000000010001001111011;
assign LUT_4[48267] = 32'b11111111111111111011010101110011;
assign LUT_4[48268] = 32'b11111111111111111111101111110011;
assign LUT_4[48269] = 32'b11111111111111111000111011101011;
assign LUT_4[48270] = 32'b11111111111111111111001010010111;
assign LUT_4[48271] = 32'b11111111111111111000010110001111;
assign LUT_4[48272] = 32'b00000000000000000111010100110000;
assign LUT_4[48273] = 32'b00000000000000000000100000101000;
assign LUT_4[48274] = 32'b00000000000000000110101111010100;
assign LUT_4[48275] = 32'b11111111111111111111111011001100;
assign LUT_4[48276] = 32'b00000000000000000100010101001100;
assign LUT_4[48277] = 32'b11111111111111111101100001000100;
assign LUT_4[48278] = 32'b00000000000000000011101111110000;
assign LUT_4[48279] = 32'b11111111111111111100111011101000;
assign LUT_4[48280] = 32'b00000000000000000000100001000101;
assign LUT_4[48281] = 32'b11111111111111111001101100111101;
assign LUT_4[48282] = 32'b11111111111111111111111011101001;
assign LUT_4[48283] = 32'b11111111111111111001000111100001;
assign LUT_4[48284] = 32'b11111111111111111101100001100001;
assign LUT_4[48285] = 32'b11111111111111110110101101011001;
assign LUT_4[48286] = 32'b11111111111111111100111100000101;
assign LUT_4[48287] = 32'b11111111111111110110000111111101;
assign LUT_4[48288] = 32'b00000000000000000111111110001001;
assign LUT_4[48289] = 32'b00000000000000000001001010000001;
assign LUT_4[48290] = 32'b00000000000000000111011000101101;
assign LUT_4[48291] = 32'b00000000000000000000100100100101;
assign LUT_4[48292] = 32'b00000000000000000100111110100101;
assign LUT_4[48293] = 32'b11111111111111111110001010011101;
assign LUT_4[48294] = 32'b00000000000000000100011001001001;
assign LUT_4[48295] = 32'b11111111111111111101100101000001;
assign LUT_4[48296] = 32'b00000000000000000001001010011110;
assign LUT_4[48297] = 32'b11111111111111111010010110010110;
assign LUT_4[48298] = 32'b00000000000000000000100101000010;
assign LUT_4[48299] = 32'b11111111111111111001110000111010;
assign LUT_4[48300] = 32'b11111111111111111110001010111010;
assign LUT_4[48301] = 32'b11111111111111110111010110110010;
assign LUT_4[48302] = 32'b11111111111111111101100101011110;
assign LUT_4[48303] = 32'b11111111111111110110110001010110;
assign LUT_4[48304] = 32'b00000000000000000101101111110111;
assign LUT_4[48305] = 32'b11111111111111111110111011101111;
assign LUT_4[48306] = 32'b00000000000000000101001010011011;
assign LUT_4[48307] = 32'b11111111111111111110010110010011;
assign LUT_4[48308] = 32'b00000000000000000010110000010011;
assign LUT_4[48309] = 32'b11111111111111111011111100001011;
assign LUT_4[48310] = 32'b00000000000000000010001010110111;
assign LUT_4[48311] = 32'b11111111111111111011010110101111;
assign LUT_4[48312] = 32'b11111111111111111110111100001100;
assign LUT_4[48313] = 32'b11111111111111111000001000000100;
assign LUT_4[48314] = 32'b11111111111111111110010110110000;
assign LUT_4[48315] = 32'b11111111111111110111100010101000;
assign LUT_4[48316] = 32'b11111111111111111011111100101000;
assign LUT_4[48317] = 32'b11111111111111110101001000100000;
assign LUT_4[48318] = 32'b11111111111111111011010111001100;
assign LUT_4[48319] = 32'b11111111111111110100100011000100;
assign LUT_4[48320] = 32'b00000000000000001010111010010110;
assign LUT_4[48321] = 32'b00000000000000000100000110001110;
assign LUT_4[48322] = 32'b00000000000000001010010100111010;
assign LUT_4[48323] = 32'b00000000000000000011100000110010;
assign LUT_4[48324] = 32'b00000000000000000111111010110010;
assign LUT_4[48325] = 32'b00000000000000000001000110101010;
assign LUT_4[48326] = 32'b00000000000000000111010101010110;
assign LUT_4[48327] = 32'b00000000000000000000100001001110;
assign LUT_4[48328] = 32'b00000000000000000100000110101011;
assign LUT_4[48329] = 32'b11111111111111111101010010100011;
assign LUT_4[48330] = 32'b00000000000000000011100001001111;
assign LUT_4[48331] = 32'b11111111111111111100101101000111;
assign LUT_4[48332] = 32'b00000000000000000001000111000111;
assign LUT_4[48333] = 32'b11111111111111111010010010111111;
assign LUT_4[48334] = 32'b00000000000000000000100001101011;
assign LUT_4[48335] = 32'b11111111111111111001101101100011;
assign LUT_4[48336] = 32'b00000000000000001000101100000100;
assign LUT_4[48337] = 32'b00000000000000000001110111111100;
assign LUT_4[48338] = 32'b00000000000000001000000110101000;
assign LUT_4[48339] = 32'b00000000000000000001010010100000;
assign LUT_4[48340] = 32'b00000000000000000101101100100000;
assign LUT_4[48341] = 32'b11111111111111111110111000011000;
assign LUT_4[48342] = 32'b00000000000000000101000111000100;
assign LUT_4[48343] = 32'b11111111111111111110010010111100;
assign LUT_4[48344] = 32'b00000000000000000001111000011001;
assign LUT_4[48345] = 32'b11111111111111111011000100010001;
assign LUT_4[48346] = 32'b00000000000000000001010010111101;
assign LUT_4[48347] = 32'b11111111111111111010011110110101;
assign LUT_4[48348] = 32'b11111111111111111110111000110101;
assign LUT_4[48349] = 32'b11111111111111111000000100101101;
assign LUT_4[48350] = 32'b11111111111111111110010011011001;
assign LUT_4[48351] = 32'b11111111111111110111011111010001;
assign LUT_4[48352] = 32'b00000000000000001001010101011101;
assign LUT_4[48353] = 32'b00000000000000000010100001010101;
assign LUT_4[48354] = 32'b00000000000000001000110000000001;
assign LUT_4[48355] = 32'b00000000000000000001111011111001;
assign LUT_4[48356] = 32'b00000000000000000110010101111001;
assign LUT_4[48357] = 32'b11111111111111111111100001110001;
assign LUT_4[48358] = 32'b00000000000000000101110000011101;
assign LUT_4[48359] = 32'b11111111111111111110111100010101;
assign LUT_4[48360] = 32'b00000000000000000010100001110010;
assign LUT_4[48361] = 32'b11111111111111111011101101101010;
assign LUT_4[48362] = 32'b00000000000000000001111100010110;
assign LUT_4[48363] = 32'b11111111111111111011001000001110;
assign LUT_4[48364] = 32'b11111111111111111111100010001110;
assign LUT_4[48365] = 32'b11111111111111111000101110000110;
assign LUT_4[48366] = 32'b11111111111111111110111100110010;
assign LUT_4[48367] = 32'b11111111111111111000001000101010;
assign LUT_4[48368] = 32'b00000000000000000111000111001011;
assign LUT_4[48369] = 32'b00000000000000000000010011000011;
assign LUT_4[48370] = 32'b00000000000000000110100001101111;
assign LUT_4[48371] = 32'b11111111111111111111101101100111;
assign LUT_4[48372] = 32'b00000000000000000100000111100111;
assign LUT_4[48373] = 32'b11111111111111111101010011011111;
assign LUT_4[48374] = 32'b00000000000000000011100010001011;
assign LUT_4[48375] = 32'b11111111111111111100101110000011;
assign LUT_4[48376] = 32'b00000000000000000000010011100000;
assign LUT_4[48377] = 32'b11111111111111111001011111011000;
assign LUT_4[48378] = 32'b11111111111111111111101110000100;
assign LUT_4[48379] = 32'b11111111111111111000111001111100;
assign LUT_4[48380] = 32'b11111111111111111101010011111100;
assign LUT_4[48381] = 32'b11111111111111110110011111110100;
assign LUT_4[48382] = 32'b11111111111111111100101110100000;
assign LUT_4[48383] = 32'b11111111111111110101111010011000;
assign LUT_4[48384] = 32'b00000000000000001011111000011101;
assign LUT_4[48385] = 32'b00000000000000000101000100010101;
assign LUT_4[48386] = 32'b00000000000000001011010011000001;
assign LUT_4[48387] = 32'b00000000000000000100011110111001;
assign LUT_4[48388] = 32'b00000000000000001000111000111001;
assign LUT_4[48389] = 32'b00000000000000000010000100110001;
assign LUT_4[48390] = 32'b00000000000000001000010011011101;
assign LUT_4[48391] = 32'b00000000000000000001011111010101;
assign LUT_4[48392] = 32'b00000000000000000101000100110010;
assign LUT_4[48393] = 32'b11111111111111111110010000101010;
assign LUT_4[48394] = 32'b00000000000000000100011111010110;
assign LUT_4[48395] = 32'b11111111111111111101101011001110;
assign LUT_4[48396] = 32'b00000000000000000010000101001110;
assign LUT_4[48397] = 32'b11111111111111111011010001000110;
assign LUT_4[48398] = 32'b00000000000000000001011111110010;
assign LUT_4[48399] = 32'b11111111111111111010101011101010;
assign LUT_4[48400] = 32'b00000000000000001001101010001011;
assign LUT_4[48401] = 32'b00000000000000000010110110000011;
assign LUT_4[48402] = 32'b00000000000000001001000100101111;
assign LUT_4[48403] = 32'b00000000000000000010010000100111;
assign LUT_4[48404] = 32'b00000000000000000110101010100111;
assign LUT_4[48405] = 32'b11111111111111111111110110011111;
assign LUT_4[48406] = 32'b00000000000000000110000101001011;
assign LUT_4[48407] = 32'b11111111111111111111010001000011;
assign LUT_4[48408] = 32'b00000000000000000010110110100000;
assign LUT_4[48409] = 32'b11111111111111111100000010011000;
assign LUT_4[48410] = 32'b00000000000000000010010001000100;
assign LUT_4[48411] = 32'b11111111111111111011011100111100;
assign LUT_4[48412] = 32'b11111111111111111111110110111100;
assign LUT_4[48413] = 32'b11111111111111111001000010110100;
assign LUT_4[48414] = 32'b11111111111111111111010001100000;
assign LUT_4[48415] = 32'b11111111111111111000011101011000;
assign LUT_4[48416] = 32'b00000000000000001010010011100100;
assign LUT_4[48417] = 32'b00000000000000000011011111011100;
assign LUT_4[48418] = 32'b00000000000000001001101110001000;
assign LUT_4[48419] = 32'b00000000000000000010111010000000;
assign LUT_4[48420] = 32'b00000000000000000111010100000000;
assign LUT_4[48421] = 32'b00000000000000000000011111111000;
assign LUT_4[48422] = 32'b00000000000000000110101110100100;
assign LUT_4[48423] = 32'b11111111111111111111111010011100;
assign LUT_4[48424] = 32'b00000000000000000011011111111001;
assign LUT_4[48425] = 32'b11111111111111111100101011110001;
assign LUT_4[48426] = 32'b00000000000000000010111010011101;
assign LUT_4[48427] = 32'b11111111111111111100000110010101;
assign LUT_4[48428] = 32'b00000000000000000000100000010101;
assign LUT_4[48429] = 32'b11111111111111111001101100001101;
assign LUT_4[48430] = 32'b11111111111111111111111010111001;
assign LUT_4[48431] = 32'b11111111111111111001000110110001;
assign LUT_4[48432] = 32'b00000000000000001000000101010010;
assign LUT_4[48433] = 32'b00000000000000000001010001001010;
assign LUT_4[48434] = 32'b00000000000000000111011111110110;
assign LUT_4[48435] = 32'b00000000000000000000101011101110;
assign LUT_4[48436] = 32'b00000000000000000101000101101110;
assign LUT_4[48437] = 32'b11111111111111111110010001100110;
assign LUT_4[48438] = 32'b00000000000000000100100000010010;
assign LUT_4[48439] = 32'b11111111111111111101101100001010;
assign LUT_4[48440] = 32'b00000000000000000001010001100111;
assign LUT_4[48441] = 32'b11111111111111111010011101011111;
assign LUT_4[48442] = 32'b00000000000000000000101100001011;
assign LUT_4[48443] = 32'b11111111111111111001111000000011;
assign LUT_4[48444] = 32'b11111111111111111110010010000011;
assign LUT_4[48445] = 32'b11111111111111110111011101111011;
assign LUT_4[48446] = 32'b11111111111111111101101100100111;
assign LUT_4[48447] = 32'b11111111111111110110111000011111;
assign LUT_4[48448] = 32'b00000000000000001101001111110001;
assign LUT_4[48449] = 32'b00000000000000000110011011101001;
assign LUT_4[48450] = 32'b00000000000000001100101010010101;
assign LUT_4[48451] = 32'b00000000000000000101110110001101;
assign LUT_4[48452] = 32'b00000000000000001010010000001101;
assign LUT_4[48453] = 32'b00000000000000000011011100000101;
assign LUT_4[48454] = 32'b00000000000000001001101010110001;
assign LUT_4[48455] = 32'b00000000000000000010110110101001;
assign LUT_4[48456] = 32'b00000000000000000110011100000110;
assign LUT_4[48457] = 32'b11111111111111111111100111111110;
assign LUT_4[48458] = 32'b00000000000000000101110110101010;
assign LUT_4[48459] = 32'b11111111111111111111000010100010;
assign LUT_4[48460] = 32'b00000000000000000011011100100010;
assign LUT_4[48461] = 32'b11111111111111111100101000011010;
assign LUT_4[48462] = 32'b00000000000000000010110111000110;
assign LUT_4[48463] = 32'b11111111111111111100000010111110;
assign LUT_4[48464] = 32'b00000000000000001011000001011111;
assign LUT_4[48465] = 32'b00000000000000000100001101010111;
assign LUT_4[48466] = 32'b00000000000000001010011100000011;
assign LUT_4[48467] = 32'b00000000000000000011100111111011;
assign LUT_4[48468] = 32'b00000000000000001000000001111011;
assign LUT_4[48469] = 32'b00000000000000000001001101110011;
assign LUT_4[48470] = 32'b00000000000000000111011100011111;
assign LUT_4[48471] = 32'b00000000000000000000101000010111;
assign LUT_4[48472] = 32'b00000000000000000100001101110100;
assign LUT_4[48473] = 32'b11111111111111111101011001101100;
assign LUT_4[48474] = 32'b00000000000000000011101000011000;
assign LUT_4[48475] = 32'b11111111111111111100110100010000;
assign LUT_4[48476] = 32'b00000000000000000001001110010000;
assign LUT_4[48477] = 32'b11111111111111111010011010001000;
assign LUT_4[48478] = 32'b00000000000000000000101000110100;
assign LUT_4[48479] = 32'b11111111111111111001110100101100;
assign LUT_4[48480] = 32'b00000000000000001011101010111000;
assign LUT_4[48481] = 32'b00000000000000000100110110110000;
assign LUT_4[48482] = 32'b00000000000000001011000101011100;
assign LUT_4[48483] = 32'b00000000000000000100010001010100;
assign LUT_4[48484] = 32'b00000000000000001000101011010100;
assign LUT_4[48485] = 32'b00000000000000000001110111001100;
assign LUT_4[48486] = 32'b00000000000000001000000101111000;
assign LUT_4[48487] = 32'b00000000000000000001010001110000;
assign LUT_4[48488] = 32'b00000000000000000100110111001101;
assign LUT_4[48489] = 32'b11111111111111111110000011000101;
assign LUT_4[48490] = 32'b00000000000000000100010001110001;
assign LUT_4[48491] = 32'b11111111111111111101011101101001;
assign LUT_4[48492] = 32'b00000000000000000001110111101001;
assign LUT_4[48493] = 32'b11111111111111111011000011100001;
assign LUT_4[48494] = 32'b00000000000000000001010010001101;
assign LUT_4[48495] = 32'b11111111111111111010011110000101;
assign LUT_4[48496] = 32'b00000000000000001001011100100110;
assign LUT_4[48497] = 32'b00000000000000000010101000011110;
assign LUT_4[48498] = 32'b00000000000000001000110111001010;
assign LUT_4[48499] = 32'b00000000000000000010000011000010;
assign LUT_4[48500] = 32'b00000000000000000110011101000010;
assign LUT_4[48501] = 32'b11111111111111111111101000111010;
assign LUT_4[48502] = 32'b00000000000000000101110111100110;
assign LUT_4[48503] = 32'b11111111111111111111000011011110;
assign LUT_4[48504] = 32'b00000000000000000010101000111011;
assign LUT_4[48505] = 32'b11111111111111111011110100110011;
assign LUT_4[48506] = 32'b00000000000000000010000011011111;
assign LUT_4[48507] = 32'b11111111111111111011001111010111;
assign LUT_4[48508] = 32'b11111111111111111111101001010111;
assign LUT_4[48509] = 32'b11111111111111111000110101001111;
assign LUT_4[48510] = 32'b11111111111111111111000011111011;
assign LUT_4[48511] = 32'b11111111111111111000001111110011;
assign LUT_4[48512] = 32'b00000000000000001110011110100101;
assign LUT_4[48513] = 32'b00000000000000000111101010011101;
assign LUT_4[48514] = 32'b00000000000000001101111001001001;
assign LUT_4[48515] = 32'b00000000000000000111000101000001;
assign LUT_4[48516] = 32'b00000000000000001011011111000001;
assign LUT_4[48517] = 32'b00000000000000000100101010111001;
assign LUT_4[48518] = 32'b00000000000000001010111001100101;
assign LUT_4[48519] = 32'b00000000000000000100000101011101;
assign LUT_4[48520] = 32'b00000000000000000111101010111010;
assign LUT_4[48521] = 32'b00000000000000000000110110110010;
assign LUT_4[48522] = 32'b00000000000000000111000101011110;
assign LUT_4[48523] = 32'b00000000000000000000010001010110;
assign LUT_4[48524] = 32'b00000000000000000100101011010110;
assign LUT_4[48525] = 32'b11111111111111111101110111001110;
assign LUT_4[48526] = 32'b00000000000000000100000101111010;
assign LUT_4[48527] = 32'b11111111111111111101010001110010;
assign LUT_4[48528] = 32'b00000000000000001100010000010011;
assign LUT_4[48529] = 32'b00000000000000000101011100001011;
assign LUT_4[48530] = 32'b00000000000000001011101010110111;
assign LUT_4[48531] = 32'b00000000000000000100110110101111;
assign LUT_4[48532] = 32'b00000000000000001001010000101111;
assign LUT_4[48533] = 32'b00000000000000000010011100100111;
assign LUT_4[48534] = 32'b00000000000000001000101011010011;
assign LUT_4[48535] = 32'b00000000000000000001110111001011;
assign LUT_4[48536] = 32'b00000000000000000101011100101000;
assign LUT_4[48537] = 32'b11111111111111111110101000100000;
assign LUT_4[48538] = 32'b00000000000000000100110111001100;
assign LUT_4[48539] = 32'b11111111111111111110000011000100;
assign LUT_4[48540] = 32'b00000000000000000010011101000100;
assign LUT_4[48541] = 32'b11111111111111111011101000111100;
assign LUT_4[48542] = 32'b00000000000000000001110111101000;
assign LUT_4[48543] = 32'b11111111111111111011000011100000;
assign LUT_4[48544] = 32'b00000000000000001100111001101100;
assign LUT_4[48545] = 32'b00000000000000000110000101100100;
assign LUT_4[48546] = 32'b00000000000000001100010100010000;
assign LUT_4[48547] = 32'b00000000000000000101100000001000;
assign LUT_4[48548] = 32'b00000000000000001001111010001000;
assign LUT_4[48549] = 32'b00000000000000000011000110000000;
assign LUT_4[48550] = 32'b00000000000000001001010100101100;
assign LUT_4[48551] = 32'b00000000000000000010100000100100;
assign LUT_4[48552] = 32'b00000000000000000110000110000001;
assign LUT_4[48553] = 32'b11111111111111111111010001111001;
assign LUT_4[48554] = 32'b00000000000000000101100000100101;
assign LUT_4[48555] = 32'b11111111111111111110101100011101;
assign LUT_4[48556] = 32'b00000000000000000011000110011101;
assign LUT_4[48557] = 32'b11111111111111111100010010010101;
assign LUT_4[48558] = 32'b00000000000000000010100001000001;
assign LUT_4[48559] = 32'b11111111111111111011101100111001;
assign LUT_4[48560] = 32'b00000000000000001010101011011010;
assign LUT_4[48561] = 32'b00000000000000000011110111010010;
assign LUT_4[48562] = 32'b00000000000000001010000101111110;
assign LUT_4[48563] = 32'b00000000000000000011010001110110;
assign LUT_4[48564] = 32'b00000000000000000111101011110110;
assign LUT_4[48565] = 32'b00000000000000000000110111101110;
assign LUT_4[48566] = 32'b00000000000000000111000110011010;
assign LUT_4[48567] = 32'b00000000000000000000010010010010;
assign LUT_4[48568] = 32'b00000000000000000011110111101111;
assign LUT_4[48569] = 32'b11111111111111111101000011100111;
assign LUT_4[48570] = 32'b00000000000000000011010010010011;
assign LUT_4[48571] = 32'b11111111111111111100011110001011;
assign LUT_4[48572] = 32'b00000000000000000000111000001011;
assign LUT_4[48573] = 32'b11111111111111111010000100000011;
assign LUT_4[48574] = 32'b00000000000000000000010010101111;
assign LUT_4[48575] = 32'b11111111111111111001011110100111;
assign LUT_4[48576] = 32'b00000000000000001111110101111001;
assign LUT_4[48577] = 32'b00000000000000001001000001110001;
assign LUT_4[48578] = 32'b00000000000000001111010000011101;
assign LUT_4[48579] = 32'b00000000000000001000011100010101;
assign LUT_4[48580] = 32'b00000000000000001100110110010101;
assign LUT_4[48581] = 32'b00000000000000000110000010001101;
assign LUT_4[48582] = 32'b00000000000000001100010000111001;
assign LUT_4[48583] = 32'b00000000000000000101011100110001;
assign LUT_4[48584] = 32'b00000000000000001001000010001110;
assign LUT_4[48585] = 32'b00000000000000000010001110000110;
assign LUT_4[48586] = 32'b00000000000000001000011100110010;
assign LUT_4[48587] = 32'b00000000000000000001101000101010;
assign LUT_4[48588] = 32'b00000000000000000110000010101010;
assign LUT_4[48589] = 32'b11111111111111111111001110100010;
assign LUT_4[48590] = 32'b00000000000000000101011101001110;
assign LUT_4[48591] = 32'b11111111111111111110101001000110;
assign LUT_4[48592] = 32'b00000000000000001101100111100111;
assign LUT_4[48593] = 32'b00000000000000000110110011011111;
assign LUT_4[48594] = 32'b00000000000000001101000010001011;
assign LUT_4[48595] = 32'b00000000000000000110001110000011;
assign LUT_4[48596] = 32'b00000000000000001010101000000011;
assign LUT_4[48597] = 32'b00000000000000000011110011111011;
assign LUT_4[48598] = 32'b00000000000000001010000010100111;
assign LUT_4[48599] = 32'b00000000000000000011001110011111;
assign LUT_4[48600] = 32'b00000000000000000110110011111100;
assign LUT_4[48601] = 32'b11111111111111111111111111110100;
assign LUT_4[48602] = 32'b00000000000000000110001110100000;
assign LUT_4[48603] = 32'b11111111111111111111011010011000;
assign LUT_4[48604] = 32'b00000000000000000011110100011000;
assign LUT_4[48605] = 32'b11111111111111111101000000010000;
assign LUT_4[48606] = 32'b00000000000000000011001110111100;
assign LUT_4[48607] = 32'b11111111111111111100011010110100;
assign LUT_4[48608] = 32'b00000000000000001110010001000000;
assign LUT_4[48609] = 32'b00000000000000000111011100111000;
assign LUT_4[48610] = 32'b00000000000000001101101011100100;
assign LUT_4[48611] = 32'b00000000000000000110110111011100;
assign LUT_4[48612] = 32'b00000000000000001011010001011100;
assign LUT_4[48613] = 32'b00000000000000000100011101010100;
assign LUT_4[48614] = 32'b00000000000000001010101100000000;
assign LUT_4[48615] = 32'b00000000000000000011110111111000;
assign LUT_4[48616] = 32'b00000000000000000111011101010101;
assign LUT_4[48617] = 32'b00000000000000000000101001001101;
assign LUT_4[48618] = 32'b00000000000000000110110111111001;
assign LUT_4[48619] = 32'b00000000000000000000000011110001;
assign LUT_4[48620] = 32'b00000000000000000100011101110001;
assign LUT_4[48621] = 32'b11111111111111111101101001101001;
assign LUT_4[48622] = 32'b00000000000000000011111000010101;
assign LUT_4[48623] = 32'b11111111111111111101000100001101;
assign LUT_4[48624] = 32'b00000000000000001100000010101110;
assign LUT_4[48625] = 32'b00000000000000000101001110100110;
assign LUT_4[48626] = 32'b00000000000000001011011101010010;
assign LUT_4[48627] = 32'b00000000000000000100101001001010;
assign LUT_4[48628] = 32'b00000000000000001001000011001010;
assign LUT_4[48629] = 32'b00000000000000000010001111000010;
assign LUT_4[48630] = 32'b00000000000000001000011101101110;
assign LUT_4[48631] = 32'b00000000000000000001101001100110;
assign LUT_4[48632] = 32'b00000000000000000101001111000011;
assign LUT_4[48633] = 32'b11111111111111111110011010111011;
assign LUT_4[48634] = 32'b00000000000000000100101001100111;
assign LUT_4[48635] = 32'b11111111111111111101110101011111;
assign LUT_4[48636] = 32'b00000000000000000010001111011111;
assign LUT_4[48637] = 32'b11111111111111111011011011010111;
assign LUT_4[48638] = 32'b00000000000000000001101010000011;
assign LUT_4[48639] = 32'b11111111111111111010110101111011;
assign LUT_4[48640] = 32'b00000000000000000110000001000010;
assign LUT_4[48641] = 32'b11111111111111111111001100111010;
assign LUT_4[48642] = 32'b00000000000000000101011011100110;
assign LUT_4[48643] = 32'b11111111111111111110100111011110;
assign LUT_4[48644] = 32'b00000000000000000011000001011110;
assign LUT_4[48645] = 32'b11111111111111111100001101010110;
assign LUT_4[48646] = 32'b00000000000000000010011100000010;
assign LUT_4[48647] = 32'b11111111111111111011100111111010;
assign LUT_4[48648] = 32'b11111111111111111111001101010111;
assign LUT_4[48649] = 32'b11111111111111111000011001001111;
assign LUT_4[48650] = 32'b11111111111111111110100111111011;
assign LUT_4[48651] = 32'b11111111111111110111110011110011;
assign LUT_4[48652] = 32'b11111111111111111100001101110011;
assign LUT_4[48653] = 32'b11111111111111110101011001101011;
assign LUT_4[48654] = 32'b11111111111111111011101000010111;
assign LUT_4[48655] = 32'b11111111111111110100110100001111;
assign LUT_4[48656] = 32'b00000000000000000011110010110000;
assign LUT_4[48657] = 32'b11111111111111111100111110101000;
assign LUT_4[48658] = 32'b00000000000000000011001101010100;
assign LUT_4[48659] = 32'b11111111111111111100011001001100;
assign LUT_4[48660] = 32'b00000000000000000000110011001100;
assign LUT_4[48661] = 32'b11111111111111111001111111000100;
assign LUT_4[48662] = 32'b00000000000000000000001101110000;
assign LUT_4[48663] = 32'b11111111111111111001011001101000;
assign LUT_4[48664] = 32'b11111111111111111100111111000101;
assign LUT_4[48665] = 32'b11111111111111110110001010111101;
assign LUT_4[48666] = 32'b11111111111111111100011001101001;
assign LUT_4[48667] = 32'b11111111111111110101100101100001;
assign LUT_4[48668] = 32'b11111111111111111001111111100001;
assign LUT_4[48669] = 32'b11111111111111110011001011011001;
assign LUT_4[48670] = 32'b11111111111111111001011010000101;
assign LUT_4[48671] = 32'b11111111111111110010100101111101;
assign LUT_4[48672] = 32'b00000000000000000100011100001001;
assign LUT_4[48673] = 32'b11111111111111111101101000000001;
assign LUT_4[48674] = 32'b00000000000000000011110110101101;
assign LUT_4[48675] = 32'b11111111111111111101000010100101;
assign LUT_4[48676] = 32'b00000000000000000001011100100101;
assign LUT_4[48677] = 32'b11111111111111111010101000011101;
assign LUT_4[48678] = 32'b00000000000000000000110111001001;
assign LUT_4[48679] = 32'b11111111111111111010000011000001;
assign LUT_4[48680] = 32'b11111111111111111101101000011110;
assign LUT_4[48681] = 32'b11111111111111110110110100010110;
assign LUT_4[48682] = 32'b11111111111111111101000011000010;
assign LUT_4[48683] = 32'b11111111111111110110001110111010;
assign LUT_4[48684] = 32'b11111111111111111010101000111010;
assign LUT_4[48685] = 32'b11111111111111110011110100110010;
assign LUT_4[48686] = 32'b11111111111111111010000011011110;
assign LUT_4[48687] = 32'b11111111111111110011001111010110;
assign LUT_4[48688] = 32'b00000000000000000010001101110111;
assign LUT_4[48689] = 32'b11111111111111111011011001101111;
assign LUT_4[48690] = 32'b00000000000000000001101000011011;
assign LUT_4[48691] = 32'b11111111111111111010110100010011;
assign LUT_4[48692] = 32'b11111111111111111111001110010011;
assign LUT_4[48693] = 32'b11111111111111111000011010001011;
assign LUT_4[48694] = 32'b11111111111111111110101000110111;
assign LUT_4[48695] = 32'b11111111111111110111110100101111;
assign LUT_4[48696] = 32'b11111111111111111011011010001100;
assign LUT_4[48697] = 32'b11111111111111110100100110000100;
assign LUT_4[48698] = 32'b11111111111111111010110100110000;
assign LUT_4[48699] = 32'b11111111111111110100000000101000;
assign LUT_4[48700] = 32'b11111111111111111000011010101000;
assign LUT_4[48701] = 32'b11111111111111110001100110100000;
assign LUT_4[48702] = 32'b11111111111111110111110101001100;
assign LUT_4[48703] = 32'b11111111111111110001000001000100;
assign LUT_4[48704] = 32'b00000000000000000111011000010110;
assign LUT_4[48705] = 32'b00000000000000000000100100001110;
assign LUT_4[48706] = 32'b00000000000000000110110010111010;
assign LUT_4[48707] = 32'b11111111111111111111111110110010;
assign LUT_4[48708] = 32'b00000000000000000100011000110010;
assign LUT_4[48709] = 32'b11111111111111111101100100101010;
assign LUT_4[48710] = 32'b00000000000000000011110011010110;
assign LUT_4[48711] = 32'b11111111111111111100111111001110;
assign LUT_4[48712] = 32'b00000000000000000000100100101011;
assign LUT_4[48713] = 32'b11111111111111111001110000100011;
assign LUT_4[48714] = 32'b11111111111111111111111111001111;
assign LUT_4[48715] = 32'b11111111111111111001001011000111;
assign LUT_4[48716] = 32'b11111111111111111101100101000111;
assign LUT_4[48717] = 32'b11111111111111110110110000111111;
assign LUT_4[48718] = 32'b11111111111111111100111111101011;
assign LUT_4[48719] = 32'b11111111111111110110001011100011;
assign LUT_4[48720] = 32'b00000000000000000101001010000100;
assign LUT_4[48721] = 32'b11111111111111111110010101111100;
assign LUT_4[48722] = 32'b00000000000000000100100100101000;
assign LUT_4[48723] = 32'b11111111111111111101110000100000;
assign LUT_4[48724] = 32'b00000000000000000010001010100000;
assign LUT_4[48725] = 32'b11111111111111111011010110011000;
assign LUT_4[48726] = 32'b00000000000000000001100101000100;
assign LUT_4[48727] = 32'b11111111111111111010110000111100;
assign LUT_4[48728] = 32'b11111111111111111110010110011001;
assign LUT_4[48729] = 32'b11111111111111110111100010010001;
assign LUT_4[48730] = 32'b11111111111111111101110000111101;
assign LUT_4[48731] = 32'b11111111111111110110111100110101;
assign LUT_4[48732] = 32'b11111111111111111011010110110101;
assign LUT_4[48733] = 32'b11111111111111110100100010101101;
assign LUT_4[48734] = 32'b11111111111111111010110001011001;
assign LUT_4[48735] = 32'b11111111111111110011111101010001;
assign LUT_4[48736] = 32'b00000000000000000101110011011101;
assign LUT_4[48737] = 32'b11111111111111111110111111010101;
assign LUT_4[48738] = 32'b00000000000000000101001110000001;
assign LUT_4[48739] = 32'b11111111111111111110011001111001;
assign LUT_4[48740] = 32'b00000000000000000010110011111001;
assign LUT_4[48741] = 32'b11111111111111111011111111110001;
assign LUT_4[48742] = 32'b00000000000000000010001110011101;
assign LUT_4[48743] = 32'b11111111111111111011011010010101;
assign LUT_4[48744] = 32'b11111111111111111110111111110010;
assign LUT_4[48745] = 32'b11111111111111111000001011101010;
assign LUT_4[48746] = 32'b11111111111111111110011010010110;
assign LUT_4[48747] = 32'b11111111111111110111100110001110;
assign LUT_4[48748] = 32'b11111111111111111100000000001110;
assign LUT_4[48749] = 32'b11111111111111110101001100000110;
assign LUT_4[48750] = 32'b11111111111111111011011010110010;
assign LUT_4[48751] = 32'b11111111111111110100100110101010;
assign LUT_4[48752] = 32'b00000000000000000011100101001011;
assign LUT_4[48753] = 32'b11111111111111111100110001000011;
assign LUT_4[48754] = 32'b00000000000000000010111111101111;
assign LUT_4[48755] = 32'b11111111111111111100001011100111;
assign LUT_4[48756] = 32'b00000000000000000000100101100111;
assign LUT_4[48757] = 32'b11111111111111111001110001011111;
assign LUT_4[48758] = 32'b00000000000000000000000000001011;
assign LUT_4[48759] = 32'b11111111111111111001001100000011;
assign LUT_4[48760] = 32'b11111111111111111100110001100000;
assign LUT_4[48761] = 32'b11111111111111110101111101011000;
assign LUT_4[48762] = 32'b11111111111111111100001100000100;
assign LUT_4[48763] = 32'b11111111111111110101010111111100;
assign LUT_4[48764] = 32'b11111111111111111001110001111100;
assign LUT_4[48765] = 32'b11111111111111110010111101110100;
assign LUT_4[48766] = 32'b11111111111111111001001100100000;
assign LUT_4[48767] = 32'b11111111111111110010011000011000;
assign LUT_4[48768] = 32'b00000000000000001000100111001010;
assign LUT_4[48769] = 32'b00000000000000000001110011000010;
assign LUT_4[48770] = 32'b00000000000000001000000001101110;
assign LUT_4[48771] = 32'b00000000000000000001001101100110;
assign LUT_4[48772] = 32'b00000000000000000101100111100110;
assign LUT_4[48773] = 32'b11111111111111111110110011011110;
assign LUT_4[48774] = 32'b00000000000000000101000010001010;
assign LUT_4[48775] = 32'b11111111111111111110001110000010;
assign LUT_4[48776] = 32'b00000000000000000001110011011111;
assign LUT_4[48777] = 32'b11111111111111111010111111010111;
assign LUT_4[48778] = 32'b00000000000000000001001110000011;
assign LUT_4[48779] = 32'b11111111111111111010011001111011;
assign LUT_4[48780] = 32'b11111111111111111110110011111011;
assign LUT_4[48781] = 32'b11111111111111110111111111110011;
assign LUT_4[48782] = 32'b11111111111111111110001110011111;
assign LUT_4[48783] = 32'b11111111111111110111011010010111;
assign LUT_4[48784] = 32'b00000000000000000110011000111000;
assign LUT_4[48785] = 32'b11111111111111111111100100110000;
assign LUT_4[48786] = 32'b00000000000000000101110011011100;
assign LUT_4[48787] = 32'b11111111111111111110111111010100;
assign LUT_4[48788] = 32'b00000000000000000011011001010100;
assign LUT_4[48789] = 32'b11111111111111111100100101001100;
assign LUT_4[48790] = 32'b00000000000000000010110011111000;
assign LUT_4[48791] = 32'b11111111111111111011111111110000;
assign LUT_4[48792] = 32'b11111111111111111111100101001101;
assign LUT_4[48793] = 32'b11111111111111111000110001000101;
assign LUT_4[48794] = 32'b11111111111111111110111111110001;
assign LUT_4[48795] = 32'b11111111111111111000001011101001;
assign LUT_4[48796] = 32'b11111111111111111100100101101001;
assign LUT_4[48797] = 32'b11111111111111110101110001100001;
assign LUT_4[48798] = 32'b11111111111111111100000000001101;
assign LUT_4[48799] = 32'b11111111111111110101001100000101;
assign LUT_4[48800] = 32'b00000000000000000111000010010001;
assign LUT_4[48801] = 32'b00000000000000000000001110001001;
assign LUT_4[48802] = 32'b00000000000000000110011100110101;
assign LUT_4[48803] = 32'b11111111111111111111101000101101;
assign LUT_4[48804] = 32'b00000000000000000100000010101101;
assign LUT_4[48805] = 32'b11111111111111111101001110100101;
assign LUT_4[48806] = 32'b00000000000000000011011101010001;
assign LUT_4[48807] = 32'b11111111111111111100101001001001;
assign LUT_4[48808] = 32'b00000000000000000000001110100110;
assign LUT_4[48809] = 32'b11111111111111111001011010011110;
assign LUT_4[48810] = 32'b11111111111111111111101001001010;
assign LUT_4[48811] = 32'b11111111111111111000110101000010;
assign LUT_4[48812] = 32'b11111111111111111101001111000010;
assign LUT_4[48813] = 32'b11111111111111110110011010111010;
assign LUT_4[48814] = 32'b11111111111111111100101001100110;
assign LUT_4[48815] = 32'b11111111111111110101110101011110;
assign LUT_4[48816] = 32'b00000000000000000100110011111111;
assign LUT_4[48817] = 32'b11111111111111111101111111110111;
assign LUT_4[48818] = 32'b00000000000000000100001110100011;
assign LUT_4[48819] = 32'b11111111111111111101011010011011;
assign LUT_4[48820] = 32'b00000000000000000001110100011011;
assign LUT_4[48821] = 32'b11111111111111111011000000010011;
assign LUT_4[48822] = 32'b00000000000000000001001110111111;
assign LUT_4[48823] = 32'b11111111111111111010011010110111;
assign LUT_4[48824] = 32'b11111111111111111110000000010100;
assign LUT_4[48825] = 32'b11111111111111110111001100001100;
assign LUT_4[48826] = 32'b11111111111111111101011010111000;
assign LUT_4[48827] = 32'b11111111111111110110100110110000;
assign LUT_4[48828] = 32'b11111111111111111011000000110000;
assign LUT_4[48829] = 32'b11111111111111110100001100101000;
assign LUT_4[48830] = 32'b11111111111111111010011011010100;
assign LUT_4[48831] = 32'b11111111111111110011100111001100;
assign LUT_4[48832] = 32'b00000000000000001001111110011110;
assign LUT_4[48833] = 32'b00000000000000000011001010010110;
assign LUT_4[48834] = 32'b00000000000000001001011001000010;
assign LUT_4[48835] = 32'b00000000000000000010100100111010;
assign LUT_4[48836] = 32'b00000000000000000110111110111010;
assign LUT_4[48837] = 32'b00000000000000000000001010110010;
assign LUT_4[48838] = 32'b00000000000000000110011001011110;
assign LUT_4[48839] = 32'b11111111111111111111100101010110;
assign LUT_4[48840] = 32'b00000000000000000011001010110011;
assign LUT_4[48841] = 32'b11111111111111111100010110101011;
assign LUT_4[48842] = 32'b00000000000000000010100101010111;
assign LUT_4[48843] = 32'b11111111111111111011110001001111;
assign LUT_4[48844] = 32'b00000000000000000000001011001111;
assign LUT_4[48845] = 32'b11111111111111111001010111000111;
assign LUT_4[48846] = 32'b11111111111111111111100101110011;
assign LUT_4[48847] = 32'b11111111111111111000110001101011;
assign LUT_4[48848] = 32'b00000000000000000111110000001100;
assign LUT_4[48849] = 32'b00000000000000000000111100000100;
assign LUT_4[48850] = 32'b00000000000000000111001010110000;
assign LUT_4[48851] = 32'b00000000000000000000010110101000;
assign LUT_4[48852] = 32'b00000000000000000100110000101000;
assign LUT_4[48853] = 32'b11111111111111111101111100100000;
assign LUT_4[48854] = 32'b00000000000000000100001011001100;
assign LUT_4[48855] = 32'b11111111111111111101010111000100;
assign LUT_4[48856] = 32'b00000000000000000000111100100001;
assign LUT_4[48857] = 32'b11111111111111111010001000011001;
assign LUT_4[48858] = 32'b00000000000000000000010111000101;
assign LUT_4[48859] = 32'b11111111111111111001100010111101;
assign LUT_4[48860] = 32'b11111111111111111101111100111101;
assign LUT_4[48861] = 32'b11111111111111110111001000110101;
assign LUT_4[48862] = 32'b11111111111111111101010111100001;
assign LUT_4[48863] = 32'b11111111111111110110100011011001;
assign LUT_4[48864] = 32'b00000000000000001000011001100101;
assign LUT_4[48865] = 32'b00000000000000000001100101011101;
assign LUT_4[48866] = 32'b00000000000000000111110100001001;
assign LUT_4[48867] = 32'b00000000000000000001000000000001;
assign LUT_4[48868] = 32'b00000000000000000101011010000001;
assign LUT_4[48869] = 32'b11111111111111111110100101111001;
assign LUT_4[48870] = 32'b00000000000000000100110100100101;
assign LUT_4[48871] = 32'b11111111111111111110000000011101;
assign LUT_4[48872] = 32'b00000000000000000001100101111010;
assign LUT_4[48873] = 32'b11111111111111111010110001110010;
assign LUT_4[48874] = 32'b00000000000000000001000000011110;
assign LUT_4[48875] = 32'b11111111111111111010001100010110;
assign LUT_4[48876] = 32'b11111111111111111110100110010110;
assign LUT_4[48877] = 32'b11111111111111110111110010001110;
assign LUT_4[48878] = 32'b11111111111111111110000000111010;
assign LUT_4[48879] = 32'b11111111111111110111001100110010;
assign LUT_4[48880] = 32'b00000000000000000110001011010011;
assign LUT_4[48881] = 32'b11111111111111111111010111001011;
assign LUT_4[48882] = 32'b00000000000000000101100101110111;
assign LUT_4[48883] = 32'b11111111111111111110110001101111;
assign LUT_4[48884] = 32'b00000000000000000011001011101111;
assign LUT_4[48885] = 32'b11111111111111111100010111100111;
assign LUT_4[48886] = 32'b00000000000000000010100110010011;
assign LUT_4[48887] = 32'b11111111111111111011110010001011;
assign LUT_4[48888] = 32'b11111111111111111111010111101000;
assign LUT_4[48889] = 32'b11111111111111111000100011100000;
assign LUT_4[48890] = 32'b11111111111111111110110010001100;
assign LUT_4[48891] = 32'b11111111111111110111111110000100;
assign LUT_4[48892] = 32'b11111111111111111100011000000100;
assign LUT_4[48893] = 32'b11111111111111110101100011111100;
assign LUT_4[48894] = 32'b11111111111111111011110010101000;
assign LUT_4[48895] = 32'b11111111111111110100111110100000;
assign LUT_4[48896] = 32'b00000000000000001010111100100101;
assign LUT_4[48897] = 32'b00000000000000000100001000011101;
assign LUT_4[48898] = 32'b00000000000000001010010111001001;
assign LUT_4[48899] = 32'b00000000000000000011100011000001;
assign LUT_4[48900] = 32'b00000000000000000111111101000001;
assign LUT_4[48901] = 32'b00000000000000000001001000111001;
assign LUT_4[48902] = 32'b00000000000000000111010111100101;
assign LUT_4[48903] = 32'b00000000000000000000100011011101;
assign LUT_4[48904] = 32'b00000000000000000100001000111010;
assign LUT_4[48905] = 32'b11111111111111111101010100110010;
assign LUT_4[48906] = 32'b00000000000000000011100011011110;
assign LUT_4[48907] = 32'b11111111111111111100101111010110;
assign LUT_4[48908] = 32'b00000000000000000001001001010110;
assign LUT_4[48909] = 32'b11111111111111111010010101001110;
assign LUT_4[48910] = 32'b00000000000000000000100011111010;
assign LUT_4[48911] = 32'b11111111111111111001101111110010;
assign LUT_4[48912] = 32'b00000000000000001000101110010011;
assign LUT_4[48913] = 32'b00000000000000000001111010001011;
assign LUT_4[48914] = 32'b00000000000000001000001000110111;
assign LUT_4[48915] = 32'b00000000000000000001010100101111;
assign LUT_4[48916] = 32'b00000000000000000101101110101111;
assign LUT_4[48917] = 32'b11111111111111111110111010100111;
assign LUT_4[48918] = 32'b00000000000000000101001001010011;
assign LUT_4[48919] = 32'b11111111111111111110010101001011;
assign LUT_4[48920] = 32'b00000000000000000001111010101000;
assign LUT_4[48921] = 32'b11111111111111111011000110100000;
assign LUT_4[48922] = 32'b00000000000000000001010101001100;
assign LUT_4[48923] = 32'b11111111111111111010100001000100;
assign LUT_4[48924] = 32'b11111111111111111110111011000100;
assign LUT_4[48925] = 32'b11111111111111111000000110111100;
assign LUT_4[48926] = 32'b11111111111111111110010101101000;
assign LUT_4[48927] = 32'b11111111111111110111100001100000;
assign LUT_4[48928] = 32'b00000000000000001001010111101100;
assign LUT_4[48929] = 32'b00000000000000000010100011100100;
assign LUT_4[48930] = 32'b00000000000000001000110010010000;
assign LUT_4[48931] = 32'b00000000000000000001111110001000;
assign LUT_4[48932] = 32'b00000000000000000110011000001000;
assign LUT_4[48933] = 32'b11111111111111111111100100000000;
assign LUT_4[48934] = 32'b00000000000000000101110010101100;
assign LUT_4[48935] = 32'b11111111111111111110111110100100;
assign LUT_4[48936] = 32'b00000000000000000010100100000001;
assign LUT_4[48937] = 32'b11111111111111111011101111111001;
assign LUT_4[48938] = 32'b00000000000000000001111110100101;
assign LUT_4[48939] = 32'b11111111111111111011001010011101;
assign LUT_4[48940] = 32'b11111111111111111111100100011101;
assign LUT_4[48941] = 32'b11111111111111111000110000010101;
assign LUT_4[48942] = 32'b11111111111111111110111111000001;
assign LUT_4[48943] = 32'b11111111111111111000001010111001;
assign LUT_4[48944] = 32'b00000000000000000111001001011010;
assign LUT_4[48945] = 32'b00000000000000000000010101010010;
assign LUT_4[48946] = 32'b00000000000000000110100011111110;
assign LUT_4[48947] = 32'b11111111111111111111101111110110;
assign LUT_4[48948] = 32'b00000000000000000100001001110110;
assign LUT_4[48949] = 32'b11111111111111111101010101101110;
assign LUT_4[48950] = 32'b00000000000000000011100100011010;
assign LUT_4[48951] = 32'b11111111111111111100110000010010;
assign LUT_4[48952] = 32'b00000000000000000000010101101111;
assign LUT_4[48953] = 32'b11111111111111111001100001100111;
assign LUT_4[48954] = 32'b11111111111111111111110000010011;
assign LUT_4[48955] = 32'b11111111111111111000111100001011;
assign LUT_4[48956] = 32'b11111111111111111101010110001011;
assign LUT_4[48957] = 32'b11111111111111110110100010000011;
assign LUT_4[48958] = 32'b11111111111111111100110000101111;
assign LUT_4[48959] = 32'b11111111111111110101111100100111;
assign LUT_4[48960] = 32'b00000000000000001100010011111001;
assign LUT_4[48961] = 32'b00000000000000000101011111110001;
assign LUT_4[48962] = 32'b00000000000000001011101110011101;
assign LUT_4[48963] = 32'b00000000000000000100111010010101;
assign LUT_4[48964] = 32'b00000000000000001001010100010101;
assign LUT_4[48965] = 32'b00000000000000000010100000001101;
assign LUT_4[48966] = 32'b00000000000000001000101110111001;
assign LUT_4[48967] = 32'b00000000000000000001111010110001;
assign LUT_4[48968] = 32'b00000000000000000101100000001110;
assign LUT_4[48969] = 32'b11111111111111111110101100000110;
assign LUT_4[48970] = 32'b00000000000000000100111010110010;
assign LUT_4[48971] = 32'b11111111111111111110000110101010;
assign LUT_4[48972] = 32'b00000000000000000010100000101010;
assign LUT_4[48973] = 32'b11111111111111111011101100100010;
assign LUT_4[48974] = 32'b00000000000000000001111011001110;
assign LUT_4[48975] = 32'b11111111111111111011000111000110;
assign LUT_4[48976] = 32'b00000000000000001010000101100111;
assign LUT_4[48977] = 32'b00000000000000000011010001011111;
assign LUT_4[48978] = 32'b00000000000000001001100000001011;
assign LUT_4[48979] = 32'b00000000000000000010101100000011;
assign LUT_4[48980] = 32'b00000000000000000111000110000011;
assign LUT_4[48981] = 32'b00000000000000000000010001111011;
assign LUT_4[48982] = 32'b00000000000000000110100000100111;
assign LUT_4[48983] = 32'b11111111111111111111101100011111;
assign LUT_4[48984] = 32'b00000000000000000011010001111100;
assign LUT_4[48985] = 32'b11111111111111111100011101110100;
assign LUT_4[48986] = 32'b00000000000000000010101100100000;
assign LUT_4[48987] = 32'b11111111111111111011111000011000;
assign LUT_4[48988] = 32'b00000000000000000000010010011000;
assign LUT_4[48989] = 32'b11111111111111111001011110010000;
assign LUT_4[48990] = 32'b11111111111111111111101100111100;
assign LUT_4[48991] = 32'b11111111111111111000111000110100;
assign LUT_4[48992] = 32'b00000000000000001010101111000000;
assign LUT_4[48993] = 32'b00000000000000000011111010111000;
assign LUT_4[48994] = 32'b00000000000000001010001001100100;
assign LUT_4[48995] = 32'b00000000000000000011010101011100;
assign LUT_4[48996] = 32'b00000000000000000111101111011100;
assign LUT_4[48997] = 32'b00000000000000000000111011010100;
assign LUT_4[48998] = 32'b00000000000000000111001010000000;
assign LUT_4[48999] = 32'b00000000000000000000010101111000;
assign LUT_4[49000] = 32'b00000000000000000011111011010101;
assign LUT_4[49001] = 32'b11111111111111111101000111001101;
assign LUT_4[49002] = 32'b00000000000000000011010101111001;
assign LUT_4[49003] = 32'b11111111111111111100100001110001;
assign LUT_4[49004] = 32'b00000000000000000000111011110001;
assign LUT_4[49005] = 32'b11111111111111111010000111101001;
assign LUT_4[49006] = 32'b00000000000000000000010110010101;
assign LUT_4[49007] = 32'b11111111111111111001100010001101;
assign LUT_4[49008] = 32'b00000000000000001000100000101110;
assign LUT_4[49009] = 32'b00000000000000000001101100100110;
assign LUT_4[49010] = 32'b00000000000000000111111011010010;
assign LUT_4[49011] = 32'b00000000000000000001000111001010;
assign LUT_4[49012] = 32'b00000000000000000101100001001010;
assign LUT_4[49013] = 32'b11111111111111111110101101000010;
assign LUT_4[49014] = 32'b00000000000000000100111011101110;
assign LUT_4[49015] = 32'b11111111111111111110000111100110;
assign LUT_4[49016] = 32'b00000000000000000001101101000011;
assign LUT_4[49017] = 32'b11111111111111111010111000111011;
assign LUT_4[49018] = 32'b00000000000000000001000111100111;
assign LUT_4[49019] = 32'b11111111111111111010010011011111;
assign LUT_4[49020] = 32'b11111111111111111110101101011111;
assign LUT_4[49021] = 32'b11111111111111110111111001010111;
assign LUT_4[49022] = 32'b11111111111111111110001000000011;
assign LUT_4[49023] = 32'b11111111111111110111010011111011;
assign LUT_4[49024] = 32'b00000000000000001101100010101101;
assign LUT_4[49025] = 32'b00000000000000000110101110100101;
assign LUT_4[49026] = 32'b00000000000000001100111101010001;
assign LUT_4[49027] = 32'b00000000000000000110001001001001;
assign LUT_4[49028] = 32'b00000000000000001010100011001001;
assign LUT_4[49029] = 32'b00000000000000000011101111000001;
assign LUT_4[49030] = 32'b00000000000000001001111101101101;
assign LUT_4[49031] = 32'b00000000000000000011001001100101;
assign LUT_4[49032] = 32'b00000000000000000110101111000010;
assign LUT_4[49033] = 32'b11111111111111111111111010111010;
assign LUT_4[49034] = 32'b00000000000000000110001001100110;
assign LUT_4[49035] = 32'b11111111111111111111010101011110;
assign LUT_4[49036] = 32'b00000000000000000011101111011110;
assign LUT_4[49037] = 32'b11111111111111111100111011010110;
assign LUT_4[49038] = 32'b00000000000000000011001010000010;
assign LUT_4[49039] = 32'b11111111111111111100010101111010;
assign LUT_4[49040] = 32'b00000000000000001011010100011011;
assign LUT_4[49041] = 32'b00000000000000000100100000010011;
assign LUT_4[49042] = 32'b00000000000000001010101110111111;
assign LUT_4[49043] = 32'b00000000000000000011111010110111;
assign LUT_4[49044] = 32'b00000000000000001000010100110111;
assign LUT_4[49045] = 32'b00000000000000000001100000101111;
assign LUT_4[49046] = 32'b00000000000000000111101111011011;
assign LUT_4[49047] = 32'b00000000000000000000111011010011;
assign LUT_4[49048] = 32'b00000000000000000100100000110000;
assign LUT_4[49049] = 32'b11111111111111111101101100101000;
assign LUT_4[49050] = 32'b00000000000000000011111011010100;
assign LUT_4[49051] = 32'b11111111111111111101000111001100;
assign LUT_4[49052] = 32'b00000000000000000001100001001100;
assign LUT_4[49053] = 32'b11111111111111111010101101000100;
assign LUT_4[49054] = 32'b00000000000000000000111011110000;
assign LUT_4[49055] = 32'b11111111111111111010000111101000;
assign LUT_4[49056] = 32'b00000000000000001011111101110100;
assign LUT_4[49057] = 32'b00000000000000000101001001101100;
assign LUT_4[49058] = 32'b00000000000000001011011000011000;
assign LUT_4[49059] = 32'b00000000000000000100100100010000;
assign LUT_4[49060] = 32'b00000000000000001000111110010000;
assign LUT_4[49061] = 32'b00000000000000000010001010001000;
assign LUT_4[49062] = 32'b00000000000000001000011000110100;
assign LUT_4[49063] = 32'b00000000000000000001100100101100;
assign LUT_4[49064] = 32'b00000000000000000101001010001001;
assign LUT_4[49065] = 32'b11111111111111111110010110000001;
assign LUT_4[49066] = 32'b00000000000000000100100100101101;
assign LUT_4[49067] = 32'b11111111111111111101110000100101;
assign LUT_4[49068] = 32'b00000000000000000010001010100101;
assign LUT_4[49069] = 32'b11111111111111111011010110011101;
assign LUT_4[49070] = 32'b00000000000000000001100101001001;
assign LUT_4[49071] = 32'b11111111111111111010110001000001;
assign LUT_4[49072] = 32'b00000000000000001001101111100010;
assign LUT_4[49073] = 32'b00000000000000000010111011011010;
assign LUT_4[49074] = 32'b00000000000000001001001010000110;
assign LUT_4[49075] = 32'b00000000000000000010010101111110;
assign LUT_4[49076] = 32'b00000000000000000110101111111110;
assign LUT_4[49077] = 32'b11111111111111111111111011110110;
assign LUT_4[49078] = 32'b00000000000000000110001010100010;
assign LUT_4[49079] = 32'b11111111111111111111010110011010;
assign LUT_4[49080] = 32'b00000000000000000010111011110111;
assign LUT_4[49081] = 32'b11111111111111111100000111101111;
assign LUT_4[49082] = 32'b00000000000000000010010110011011;
assign LUT_4[49083] = 32'b11111111111111111011100010010011;
assign LUT_4[49084] = 32'b11111111111111111111111100010011;
assign LUT_4[49085] = 32'b11111111111111111001001000001011;
assign LUT_4[49086] = 32'b11111111111111111111010110110111;
assign LUT_4[49087] = 32'b11111111111111111000100010101111;
assign LUT_4[49088] = 32'b00000000000000001110111010000001;
assign LUT_4[49089] = 32'b00000000000000001000000101111001;
assign LUT_4[49090] = 32'b00000000000000001110010100100101;
assign LUT_4[49091] = 32'b00000000000000000111100000011101;
assign LUT_4[49092] = 32'b00000000000000001011111010011101;
assign LUT_4[49093] = 32'b00000000000000000101000110010101;
assign LUT_4[49094] = 32'b00000000000000001011010101000001;
assign LUT_4[49095] = 32'b00000000000000000100100000111001;
assign LUT_4[49096] = 32'b00000000000000001000000110010110;
assign LUT_4[49097] = 32'b00000000000000000001010010001110;
assign LUT_4[49098] = 32'b00000000000000000111100000111010;
assign LUT_4[49099] = 32'b00000000000000000000101100110010;
assign LUT_4[49100] = 32'b00000000000000000101000110110010;
assign LUT_4[49101] = 32'b11111111111111111110010010101010;
assign LUT_4[49102] = 32'b00000000000000000100100001010110;
assign LUT_4[49103] = 32'b11111111111111111101101101001110;
assign LUT_4[49104] = 32'b00000000000000001100101011101111;
assign LUT_4[49105] = 32'b00000000000000000101110111100111;
assign LUT_4[49106] = 32'b00000000000000001100000110010011;
assign LUT_4[49107] = 32'b00000000000000000101010010001011;
assign LUT_4[49108] = 32'b00000000000000001001101100001011;
assign LUT_4[49109] = 32'b00000000000000000010111000000011;
assign LUT_4[49110] = 32'b00000000000000001001000110101111;
assign LUT_4[49111] = 32'b00000000000000000010010010100111;
assign LUT_4[49112] = 32'b00000000000000000101111000000100;
assign LUT_4[49113] = 32'b11111111111111111111000011111100;
assign LUT_4[49114] = 32'b00000000000000000101010010101000;
assign LUT_4[49115] = 32'b11111111111111111110011110100000;
assign LUT_4[49116] = 32'b00000000000000000010111000100000;
assign LUT_4[49117] = 32'b11111111111111111100000100011000;
assign LUT_4[49118] = 32'b00000000000000000010010011000100;
assign LUT_4[49119] = 32'b11111111111111111011011110111100;
assign LUT_4[49120] = 32'b00000000000000001101010101001000;
assign LUT_4[49121] = 32'b00000000000000000110100001000000;
assign LUT_4[49122] = 32'b00000000000000001100101111101100;
assign LUT_4[49123] = 32'b00000000000000000101111011100100;
assign LUT_4[49124] = 32'b00000000000000001010010101100100;
assign LUT_4[49125] = 32'b00000000000000000011100001011100;
assign LUT_4[49126] = 32'b00000000000000001001110000001000;
assign LUT_4[49127] = 32'b00000000000000000010111100000000;
assign LUT_4[49128] = 32'b00000000000000000110100001011101;
assign LUT_4[49129] = 32'b11111111111111111111101101010101;
assign LUT_4[49130] = 32'b00000000000000000101111100000001;
assign LUT_4[49131] = 32'b11111111111111111111000111111001;
assign LUT_4[49132] = 32'b00000000000000000011100001111001;
assign LUT_4[49133] = 32'b11111111111111111100101101110001;
assign LUT_4[49134] = 32'b00000000000000000010111100011101;
assign LUT_4[49135] = 32'b11111111111111111100001000010101;
assign LUT_4[49136] = 32'b00000000000000001011000110110110;
assign LUT_4[49137] = 32'b00000000000000000100010010101110;
assign LUT_4[49138] = 32'b00000000000000001010100001011010;
assign LUT_4[49139] = 32'b00000000000000000011101101010010;
assign LUT_4[49140] = 32'b00000000000000001000000111010010;
assign LUT_4[49141] = 32'b00000000000000000001010011001010;
assign LUT_4[49142] = 32'b00000000000000000111100001110110;
assign LUT_4[49143] = 32'b00000000000000000000101101101110;
assign LUT_4[49144] = 32'b00000000000000000100010011001011;
assign LUT_4[49145] = 32'b11111111111111111101011111000011;
assign LUT_4[49146] = 32'b00000000000000000011101101101111;
assign LUT_4[49147] = 32'b11111111111111111100111001100111;
assign LUT_4[49148] = 32'b00000000000000000001010011100111;
assign LUT_4[49149] = 32'b11111111111111111010011111011111;
assign LUT_4[49150] = 32'b00000000000000000000101110001011;
assign LUT_4[49151] = 32'b11111111111111111001111010000011;
assign LUT_4[49152] = 32'b00000000000000001100110001100000;
assign LUT_4[49153] = 32'b00000000000000000101111101011000;
assign LUT_4[49154] = 32'b00000000000000001100001100000100;
assign LUT_4[49155] = 32'b00000000000000000101010111111100;
assign LUT_4[49156] = 32'b00000000000000001001110001111100;
assign LUT_4[49157] = 32'b00000000000000000010111101110100;
assign LUT_4[49158] = 32'b00000000000000001001001100100000;
assign LUT_4[49159] = 32'b00000000000000000010011000011000;
assign LUT_4[49160] = 32'b00000000000000000101111101110101;
assign LUT_4[49161] = 32'b11111111111111111111001001101101;
assign LUT_4[49162] = 32'b00000000000000000101011000011001;
assign LUT_4[49163] = 32'b11111111111111111110100100010001;
assign LUT_4[49164] = 32'b00000000000000000010111110010001;
assign LUT_4[49165] = 32'b11111111111111111100001010001001;
assign LUT_4[49166] = 32'b00000000000000000010011000110101;
assign LUT_4[49167] = 32'b11111111111111111011100100101101;
assign LUT_4[49168] = 32'b00000000000000001010100011001110;
assign LUT_4[49169] = 32'b00000000000000000011101111000110;
assign LUT_4[49170] = 32'b00000000000000001001111101110010;
assign LUT_4[49171] = 32'b00000000000000000011001001101010;
assign LUT_4[49172] = 32'b00000000000000000111100011101010;
assign LUT_4[49173] = 32'b00000000000000000000101111100010;
assign LUT_4[49174] = 32'b00000000000000000110111110001110;
assign LUT_4[49175] = 32'b00000000000000000000001010000110;
assign LUT_4[49176] = 32'b00000000000000000011101111100011;
assign LUT_4[49177] = 32'b11111111111111111100111011011011;
assign LUT_4[49178] = 32'b00000000000000000011001010000111;
assign LUT_4[49179] = 32'b11111111111111111100010101111111;
assign LUT_4[49180] = 32'b00000000000000000000101111111111;
assign LUT_4[49181] = 32'b11111111111111111001111011110111;
assign LUT_4[49182] = 32'b00000000000000000000001010100011;
assign LUT_4[49183] = 32'b11111111111111111001010110011011;
assign LUT_4[49184] = 32'b00000000000000001011001100100111;
assign LUT_4[49185] = 32'b00000000000000000100011000011111;
assign LUT_4[49186] = 32'b00000000000000001010100111001011;
assign LUT_4[49187] = 32'b00000000000000000011110011000011;
assign LUT_4[49188] = 32'b00000000000000001000001101000011;
assign LUT_4[49189] = 32'b00000000000000000001011000111011;
assign LUT_4[49190] = 32'b00000000000000000111100111100111;
assign LUT_4[49191] = 32'b00000000000000000000110011011111;
assign LUT_4[49192] = 32'b00000000000000000100011000111100;
assign LUT_4[49193] = 32'b11111111111111111101100100110100;
assign LUT_4[49194] = 32'b00000000000000000011110011100000;
assign LUT_4[49195] = 32'b11111111111111111100111111011000;
assign LUT_4[49196] = 32'b00000000000000000001011001011000;
assign LUT_4[49197] = 32'b11111111111111111010100101010000;
assign LUT_4[49198] = 32'b00000000000000000000110011111100;
assign LUT_4[49199] = 32'b11111111111111111001111111110100;
assign LUT_4[49200] = 32'b00000000000000001000111110010101;
assign LUT_4[49201] = 32'b00000000000000000010001010001101;
assign LUT_4[49202] = 32'b00000000000000001000011000111001;
assign LUT_4[49203] = 32'b00000000000000000001100100110001;
assign LUT_4[49204] = 32'b00000000000000000101111110110001;
assign LUT_4[49205] = 32'b11111111111111111111001010101001;
assign LUT_4[49206] = 32'b00000000000000000101011001010101;
assign LUT_4[49207] = 32'b11111111111111111110100101001101;
assign LUT_4[49208] = 32'b00000000000000000010001010101010;
assign LUT_4[49209] = 32'b11111111111111111011010110100010;
assign LUT_4[49210] = 32'b00000000000000000001100101001110;
assign LUT_4[49211] = 32'b11111111111111111010110001000110;
assign LUT_4[49212] = 32'b11111111111111111111001011000110;
assign LUT_4[49213] = 32'b11111111111111111000010110111110;
assign LUT_4[49214] = 32'b11111111111111111110100101101010;
assign LUT_4[49215] = 32'b11111111111111110111110001100010;
assign LUT_4[49216] = 32'b00000000000000001110001000110100;
assign LUT_4[49217] = 32'b00000000000000000111010100101100;
assign LUT_4[49218] = 32'b00000000000000001101100011011000;
assign LUT_4[49219] = 32'b00000000000000000110101111010000;
assign LUT_4[49220] = 32'b00000000000000001011001001010000;
assign LUT_4[49221] = 32'b00000000000000000100010101001000;
assign LUT_4[49222] = 32'b00000000000000001010100011110100;
assign LUT_4[49223] = 32'b00000000000000000011101111101100;
assign LUT_4[49224] = 32'b00000000000000000111010101001001;
assign LUT_4[49225] = 32'b00000000000000000000100001000001;
assign LUT_4[49226] = 32'b00000000000000000110101111101101;
assign LUT_4[49227] = 32'b11111111111111111111111011100101;
assign LUT_4[49228] = 32'b00000000000000000100010101100101;
assign LUT_4[49229] = 32'b11111111111111111101100001011101;
assign LUT_4[49230] = 32'b00000000000000000011110000001001;
assign LUT_4[49231] = 32'b11111111111111111100111100000001;
assign LUT_4[49232] = 32'b00000000000000001011111010100010;
assign LUT_4[49233] = 32'b00000000000000000101000110011010;
assign LUT_4[49234] = 32'b00000000000000001011010101000110;
assign LUT_4[49235] = 32'b00000000000000000100100000111110;
assign LUT_4[49236] = 32'b00000000000000001000111010111110;
assign LUT_4[49237] = 32'b00000000000000000010000110110110;
assign LUT_4[49238] = 32'b00000000000000001000010101100010;
assign LUT_4[49239] = 32'b00000000000000000001100001011010;
assign LUT_4[49240] = 32'b00000000000000000101000110110111;
assign LUT_4[49241] = 32'b11111111111111111110010010101111;
assign LUT_4[49242] = 32'b00000000000000000100100001011011;
assign LUT_4[49243] = 32'b11111111111111111101101101010011;
assign LUT_4[49244] = 32'b00000000000000000010000111010011;
assign LUT_4[49245] = 32'b11111111111111111011010011001011;
assign LUT_4[49246] = 32'b00000000000000000001100001110111;
assign LUT_4[49247] = 32'b11111111111111111010101101101111;
assign LUT_4[49248] = 32'b00000000000000001100100011111011;
assign LUT_4[49249] = 32'b00000000000000000101101111110011;
assign LUT_4[49250] = 32'b00000000000000001011111110011111;
assign LUT_4[49251] = 32'b00000000000000000101001010010111;
assign LUT_4[49252] = 32'b00000000000000001001100100010111;
assign LUT_4[49253] = 32'b00000000000000000010110000001111;
assign LUT_4[49254] = 32'b00000000000000001000111110111011;
assign LUT_4[49255] = 32'b00000000000000000010001010110011;
assign LUT_4[49256] = 32'b00000000000000000101110000010000;
assign LUT_4[49257] = 32'b11111111111111111110111100001000;
assign LUT_4[49258] = 32'b00000000000000000101001010110100;
assign LUT_4[49259] = 32'b11111111111111111110010110101100;
assign LUT_4[49260] = 32'b00000000000000000010110000101100;
assign LUT_4[49261] = 32'b11111111111111111011111100100100;
assign LUT_4[49262] = 32'b00000000000000000010001011010000;
assign LUT_4[49263] = 32'b11111111111111111011010111001000;
assign LUT_4[49264] = 32'b00000000000000001010010101101001;
assign LUT_4[49265] = 32'b00000000000000000011100001100001;
assign LUT_4[49266] = 32'b00000000000000001001110000001101;
assign LUT_4[49267] = 32'b00000000000000000010111100000101;
assign LUT_4[49268] = 32'b00000000000000000111010110000101;
assign LUT_4[49269] = 32'b00000000000000000000100001111101;
assign LUT_4[49270] = 32'b00000000000000000110110000101001;
assign LUT_4[49271] = 32'b11111111111111111111111100100001;
assign LUT_4[49272] = 32'b00000000000000000011100001111110;
assign LUT_4[49273] = 32'b11111111111111111100101101110110;
assign LUT_4[49274] = 32'b00000000000000000010111100100010;
assign LUT_4[49275] = 32'b11111111111111111100001000011010;
assign LUT_4[49276] = 32'b00000000000000000000100010011010;
assign LUT_4[49277] = 32'b11111111111111111001101110010010;
assign LUT_4[49278] = 32'b11111111111111111111111100111110;
assign LUT_4[49279] = 32'b11111111111111111001001000110110;
assign LUT_4[49280] = 32'b00000000000000001111010111101000;
assign LUT_4[49281] = 32'b00000000000000001000100011100000;
assign LUT_4[49282] = 32'b00000000000000001110110010001100;
assign LUT_4[49283] = 32'b00000000000000000111111110000100;
assign LUT_4[49284] = 32'b00000000000000001100011000000100;
assign LUT_4[49285] = 32'b00000000000000000101100011111100;
assign LUT_4[49286] = 32'b00000000000000001011110010101000;
assign LUT_4[49287] = 32'b00000000000000000100111110100000;
assign LUT_4[49288] = 32'b00000000000000001000100011111101;
assign LUT_4[49289] = 32'b00000000000000000001101111110101;
assign LUT_4[49290] = 32'b00000000000000000111111110100001;
assign LUT_4[49291] = 32'b00000000000000000001001010011001;
assign LUT_4[49292] = 32'b00000000000000000101100100011001;
assign LUT_4[49293] = 32'b11111111111111111110110000010001;
assign LUT_4[49294] = 32'b00000000000000000100111110111101;
assign LUT_4[49295] = 32'b11111111111111111110001010110101;
assign LUT_4[49296] = 32'b00000000000000001101001001010110;
assign LUT_4[49297] = 32'b00000000000000000110010101001110;
assign LUT_4[49298] = 32'b00000000000000001100100011111010;
assign LUT_4[49299] = 32'b00000000000000000101101111110010;
assign LUT_4[49300] = 32'b00000000000000001010001001110010;
assign LUT_4[49301] = 32'b00000000000000000011010101101010;
assign LUT_4[49302] = 32'b00000000000000001001100100010110;
assign LUT_4[49303] = 32'b00000000000000000010110000001110;
assign LUT_4[49304] = 32'b00000000000000000110010101101011;
assign LUT_4[49305] = 32'b11111111111111111111100001100011;
assign LUT_4[49306] = 32'b00000000000000000101110000001111;
assign LUT_4[49307] = 32'b11111111111111111110111100000111;
assign LUT_4[49308] = 32'b00000000000000000011010110000111;
assign LUT_4[49309] = 32'b11111111111111111100100001111111;
assign LUT_4[49310] = 32'b00000000000000000010110000101011;
assign LUT_4[49311] = 32'b11111111111111111011111100100011;
assign LUT_4[49312] = 32'b00000000000000001101110010101111;
assign LUT_4[49313] = 32'b00000000000000000110111110100111;
assign LUT_4[49314] = 32'b00000000000000001101001101010011;
assign LUT_4[49315] = 32'b00000000000000000110011001001011;
assign LUT_4[49316] = 32'b00000000000000001010110011001011;
assign LUT_4[49317] = 32'b00000000000000000011111111000011;
assign LUT_4[49318] = 32'b00000000000000001010001101101111;
assign LUT_4[49319] = 32'b00000000000000000011011001100111;
assign LUT_4[49320] = 32'b00000000000000000110111111000100;
assign LUT_4[49321] = 32'b00000000000000000000001010111100;
assign LUT_4[49322] = 32'b00000000000000000110011001101000;
assign LUT_4[49323] = 32'b11111111111111111111100101100000;
assign LUT_4[49324] = 32'b00000000000000000011111111100000;
assign LUT_4[49325] = 32'b11111111111111111101001011011000;
assign LUT_4[49326] = 32'b00000000000000000011011010000100;
assign LUT_4[49327] = 32'b11111111111111111100100101111100;
assign LUT_4[49328] = 32'b00000000000000001011100100011101;
assign LUT_4[49329] = 32'b00000000000000000100110000010101;
assign LUT_4[49330] = 32'b00000000000000001010111111000001;
assign LUT_4[49331] = 32'b00000000000000000100001010111001;
assign LUT_4[49332] = 32'b00000000000000001000100100111001;
assign LUT_4[49333] = 32'b00000000000000000001110000110001;
assign LUT_4[49334] = 32'b00000000000000000111111111011101;
assign LUT_4[49335] = 32'b00000000000000000001001011010101;
assign LUT_4[49336] = 32'b00000000000000000100110000110010;
assign LUT_4[49337] = 32'b11111111111111111101111100101010;
assign LUT_4[49338] = 32'b00000000000000000100001011010110;
assign LUT_4[49339] = 32'b11111111111111111101010111001110;
assign LUT_4[49340] = 32'b00000000000000000001110001001110;
assign LUT_4[49341] = 32'b11111111111111111010111101000110;
assign LUT_4[49342] = 32'b00000000000000000001001011110010;
assign LUT_4[49343] = 32'b11111111111111111010010111101010;
assign LUT_4[49344] = 32'b00000000000000010000101110111100;
assign LUT_4[49345] = 32'b00000000000000001001111010110100;
assign LUT_4[49346] = 32'b00000000000000010000001001100000;
assign LUT_4[49347] = 32'b00000000000000001001010101011000;
assign LUT_4[49348] = 32'b00000000000000001101101111011000;
assign LUT_4[49349] = 32'b00000000000000000110111011010000;
assign LUT_4[49350] = 32'b00000000000000001101001001111100;
assign LUT_4[49351] = 32'b00000000000000000110010101110100;
assign LUT_4[49352] = 32'b00000000000000001001111011010001;
assign LUT_4[49353] = 32'b00000000000000000011000111001001;
assign LUT_4[49354] = 32'b00000000000000001001010101110101;
assign LUT_4[49355] = 32'b00000000000000000010100001101101;
assign LUT_4[49356] = 32'b00000000000000000110111011101101;
assign LUT_4[49357] = 32'b00000000000000000000000111100101;
assign LUT_4[49358] = 32'b00000000000000000110010110010001;
assign LUT_4[49359] = 32'b11111111111111111111100010001001;
assign LUT_4[49360] = 32'b00000000000000001110100000101010;
assign LUT_4[49361] = 32'b00000000000000000111101100100010;
assign LUT_4[49362] = 32'b00000000000000001101111011001110;
assign LUT_4[49363] = 32'b00000000000000000111000111000110;
assign LUT_4[49364] = 32'b00000000000000001011100001000110;
assign LUT_4[49365] = 32'b00000000000000000100101100111110;
assign LUT_4[49366] = 32'b00000000000000001010111011101010;
assign LUT_4[49367] = 32'b00000000000000000100000111100010;
assign LUT_4[49368] = 32'b00000000000000000111101100111111;
assign LUT_4[49369] = 32'b00000000000000000000111000110111;
assign LUT_4[49370] = 32'b00000000000000000111000111100011;
assign LUT_4[49371] = 32'b00000000000000000000010011011011;
assign LUT_4[49372] = 32'b00000000000000000100101101011011;
assign LUT_4[49373] = 32'b11111111111111111101111001010011;
assign LUT_4[49374] = 32'b00000000000000000100000111111111;
assign LUT_4[49375] = 32'b11111111111111111101010011110111;
assign LUT_4[49376] = 32'b00000000000000001111001010000011;
assign LUT_4[49377] = 32'b00000000000000001000010101111011;
assign LUT_4[49378] = 32'b00000000000000001110100100100111;
assign LUT_4[49379] = 32'b00000000000000000111110000011111;
assign LUT_4[49380] = 32'b00000000000000001100001010011111;
assign LUT_4[49381] = 32'b00000000000000000101010110010111;
assign LUT_4[49382] = 32'b00000000000000001011100101000011;
assign LUT_4[49383] = 32'b00000000000000000100110000111011;
assign LUT_4[49384] = 32'b00000000000000001000010110011000;
assign LUT_4[49385] = 32'b00000000000000000001100010010000;
assign LUT_4[49386] = 32'b00000000000000000111110000111100;
assign LUT_4[49387] = 32'b00000000000000000000111100110100;
assign LUT_4[49388] = 32'b00000000000000000101010110110100;
assign LUT_4[49389] = 32'b11111111111111111110100010101100;
assign LUT_4[49390] = 32'b00000000000000000100110001011000;
assign LUT_4[49391] = 32'b11111111111111111101111101010000;
assign LUT_4[49392] = 32'b00000000000000001100111011110001;
assign LUT_4[49393] = 32'b00000000000000000110000111101001;
assign LUT_4[49394] = 32'b00000000000000001100010110010101;
assign LUT_4[49395] = 32'b00000000000000000101100010001101;
assign LUT_4[49396] = 32'b00000000000000001001111100001101;
assign LUT_4[49397] = 32'b00000000000000000011001000000101;
assign LUT_4[49398] = 32'b00000000000000001001010110110001;
assign LUT_4[49399] = 32'b00000000000000000010100010101001;
assign LUT_4[49400] = 32'b00000000000000000110001000000110;
assign LUT_4[49401] = 32'b11111111111111111111010011111110;
assign LUT_4[49402] = 32'b00000000000000000101100010101010;
assign LUT_4[49403] = 32'b11111111111111111110101110100010;
assign LUT_4[49404] = 32'b00000000000000000011001000100010;
assign LUT_4[49405] = 32'b11111111111111111100010100011010;
assign LUT_4[49406] = 32'b00000000000000000010100011000110;
assign LUT_4[49407] = 32'b11111111111111111011101110111110;
assign LUT_4[49408] = 32'b00000000000000010001101101000011;
assign LUT_4[49409] = 32'b00000000000000001010111000111011;
assign LUT_4[49410] = 32'b00000000000000010001000111100111;
assign LUT_4[49411] = 32'b00000000000000001010010011011111;
assign LUT_4[49412] = 32'b00000000000000001110101101011111;
assign LUT_4[49413] = 32'b00000000000000000111111001010111;
assign LUT_4[49414] = 32'b00000000000000001110001000000011;
assign LUT_4[49415] = 32'b00000000000000000111010011111011;
assign LUT_4[49416] = 32'b00000000000000001010111001011000;
assign LUT_4[49417] = 32'b00000000000000000100000101010000;
assign LUT_4[49418] = 32'b00000000000000001010010011111100;
assign LUT_4[49419] = 32'b00000000000000000011011111110100;
assign LUT_4[49420] = 32'b00000000000000000111111001110100;
assign LUT_4[49421] = 32'b00000000000000000001000101101100;
assign LUT_4[49422] = 32'b00000000000000000111010100011000;
assign LUT_4[49423] = 32'b00000000000000000000100000010000;
assign LUT_4[49424] = 32'b00000000000000001111011110110001;
assign LUT_4[49425] = 32'b00000000000000001000101010101001;
assign LUT_4[49426] = 32'b00000000000000001110111001010101;
assign LUT_4[49427] = 32'b00000000000000001000000101001101;
assign LUT_4[49428] = 32'b00000000000000001100011111001101;
assign LUT_4[49429] = 32'b00000000000000000101101011000101;
assign LUT_4[49430] = 32'b00000000000000001011111001110001;
assign LUT_4[49431] = 32'b00000000000000000101000101101001;
assign LUT_4[49432] = 32'b00000000000000001000101011000110;
assign LUT_4[49433] = 32'b00000000000000000001110110111110;
assign LUT_4[49434] = 32'b00000000000000001000000101101010;
assign LUT_4[49435] = 32'b00000000000000000001010001100010;
assign LUT_4[49436] = 32'b00000000000000000101101011100010;
assign LUT_4[49437] = 32'b11111111111111111110110111011010;
assign LUT_4[49438] = 32'b00000000000000000101000110000110;
assign LUT_4[49439] = 32'b11111111111111111110010001111110;
assign LUT_4[49440] = 32'b00000000000000010000001000001010;
assign LUT_4[49441] = 32'b00000000000000001001010100000010;
assign LUT_4[49442] = 32'b00000000000000001111100010101110;
assign LUT_4[49443] = 32'b00000000000000001000101110100110;
assign LUT_4[49444] = 32'b00000000000000001101001000100110;
assign LUT_4[49445] = 32'b00000000000000000110010100011110;
assign LUT_4[49446] = 32'b00000000000000001100100011001010;
assign LUT_4[49447] = 32'b00000000000000000101101111000010;
assign LUT_4[49448] = 32'b00000000000000001001010100011111;
assign LUT_4[49449] = 32'b00000000000000000010100000010111;
assign LUT_4[49450] = 32'b00000000000000001000101111000011;
assign LUT_4[49451] = 32'b00000000000000000001111010111011;
assign LUT_4[49452] = 32'b00000000000000000110010100111011;
assign LUT_4[49453] = 32'b11111111111111111111100000110011;
assign LUT_4[49454] = 32'b00000000000000000101101111011111;
assign LUT_4[49455] = 32'b11111111111111111110111011010111;
assign LUT_4[49456] = 32'b00000000000000001101111001111000;
assign LUT_4[49457] = 32'b00000000000000000111000101110000;
assign LUT_4[49458] = 32'b00000000000000001101010100011100;
assign LUT_4[49459] = 32'b00000000000000000110100000010100;
assign LUT_4[49460] = 32'b00000000000000001010111010010100;
assign LUT_4[49461] = 32'b00000000000000000100000110001100;
assign LUT_4[49462] = 32'b00000000000000001010010100111000;
assign LUT_4[49463] = 32'b00000000000000000011100000110000;
assign LUT_4[49464] = 32'b00000000000000000111000110001101;
assign LUT_4[49465] = 32'b00000000000000000000010010000101;
assign LUT_4[49466] = 32'b00000000000000000110100000110001;
assign LUT_4[49467] = 32'b11111111111111111111101100101001;
assign LUT_4[49468] = 32'b00000000000000000100000110101001;
assign LUT_4[49469] = 32'b11111111111111111101010010100001;
assign LUT_4[49470] = 32'b00000000000000000011100001001101;
assign LUT_4[49471] = 32'b11111111111111111100101101000101;
assign LUT_4[49472] = 32'b00000000000000010011000100010111;
assign LUT_4[49473] = 32'b00000000000000001100010000001111;
assign LUT_4[49474] = 32'b00000000000000010010011110111011;
assign LUT_4[49475] = 32'b00000000000000001011101010110011;
assign LUT_4[49476] = 32'b00000000000000010000000100110011;
assign LUT_4[49477] = 32'b00000000000000001001010000101011;
assign LUT_4[49478] = 32'b00000000000000001111011111010111;
assign LUT_4[49479] = 32'b00000000000000001000101011001111;
assign LUT_4[49480] = 32'b00000000000000001100010000101100;
assign LUT_4[49481] = 32'b00000000000000000101011100100100;
assign LUT_4[49482] = 32'b00000000000000001011101011010000;
assign LUT_4[49483] = 32'b00000000000000000100110111001000;
assign LUT_4[49484] = 32'b00000000000000001001010001001000;
assign LUT_4[49485] = 32'b00000000000000000010011101000000;
assign LUT_4[49486] = 32'b00000000000000001000101011101100;
assign LUT_4[49487] = 32'b00000000000000000001110111100100;
assign LUT_4[49488] = 32'b00000000000000010000110110000101;
assign LUT_4[49489] = 32'b00000000000000001010000001111101;
assign LUT_4[49490] = 32'b00000000000000010000010000101001;
assign LUT_4[49491] = 32'b00000000000000001001011100100001;
assign LUT_4[49492] = 32'b00000000000000001101110110100001;
assign LUT_4[49493] = 32'b00000000000000000111000010011001;
assign LUT_4[49494] = 32'b00000000000000001101010001000101;
assign LUT_4[49495] = 32'b00000000000000000110011100111101;
assign LUT_4[49496] = 32'b00000000000000001010000010011010;
assign LUT_4[49497] = 32'b00000000000000000011001110010010;
assign LUT_4[49498] = 32'b00000000000000001001011100111110;
assign LUT_4[49499] = 32'b00000000000000000010101000110110;
assign LUT_4[49500] = 32'b00000000000000000111000010110110;
assign LUT_4[49501] = 32'b00000000000000000000001110101110;
assign LUT_4[49502] = 32'b00000000000000000110011101011010;
assign LUT_4[49503] = 32'b11111111111111111111101001010010;
assign LUT_4[49504] = 32'b00000000000000010001011111011110;
assign LUT_4[49505] = 32'b00000000000000001010101011010110;
assign LUT_4[49506] = 32'b00000000000000010000111010000010;
assign LUT_4[49507] = 32'b00000000000000001010000101111010;
assign LUT_4[49508] = 32'b00000000000000001110011111111010;
assign LUT_4[49509] = 32'b00000000000000000111101011110010;
assign LUT_4[49510] = 32'b00000000000000001101111010011110;
assign LUT_4[49511] = 32'b00000000000000000111000110010110;
assign LUT_4[49512] = 32'b00000000000000001010101011110011;
assign LUT_4[49513] = 32'b00000000000000000011110111101011;
assign LUT_4[49514] = 32'b00000000000000001010000110010111;
assign LUT_4[49515] = 32'b00000000000000000011010010001111;
assign LUT_4[49516] = 32'b00000000000000000111101100001111;
assign LUT_4[49517] = 32'b00000000000000000000111000000111;
assign LUT_4[49518] = 32'b00000000000000000111000110110011;
assign LUT_4[49519] = 32'b00000000000000000000010010101011;
assign LUT_4[49520] = 32'b00000000000000001111010001001100;
assign LUT_4[49521] = 32'b00000000000000001000011101000100;
assign LUT_4[49522] = 32'b00000000000000001110101011110000;
assign LUT_4[49523] = 32'b00000000000000000111110111101000;
assign LUT_4[49524] = 32'b00000000000000001100010001101000;
assign LUT_4[49525] = 32'b00000000000000000101011101100000;
assign LUT_4[49526] = 32'b00000000000000001011101100001100;
assign LUT_4[49527] = 32'b00000000000000000100111000000100;
assign LUT_4[49528] = 32'b00000000000000001000011101100001;
assign LUT_4[49529] = 32'b00000000000000000001101001011001;
assign LUT_4[49530] = 32'b00000000000000000111111000000101;
assign LUT_4[49531] = 32'b00000000000000000001000011111101;
assign LUT_4[49532] = 32'b00000000000000000101011101111101;
assign LUT_4[49533] = 32'b11111111111111111110101001110101;
assign LUT_4[49534] = 32'b00000000000000000100111000100001;
assign LUT_4[49535] = 32'b11111111111111111110000100011001;
assign LUT_4[49536] = 32'b00000000000000010100010011001011;
assign LUT_4[49537] = 32'b00000000000000001101011111000011;
assign LUT_4[49538] = 32'b00000000000000010011101101101111;
assign LUT_4[49539] = 32'b00000000000000001100111001100111;
assign LUT_4[49540] = 32'b00000000000000010001010011100111;
assign LUT_4[49541] = 32'b00000000000000001010011111011111;
assign LUT_4[49542] = 32'b00000000000000010000101110001011;
assign LUT_4[49543] = 32'b00000000000000001001111010000011;
assign LUT_4[49544] = 32'b00000000000000001101011111100000;
assign LUT_4[49545] = 32'b00000000000000000110101011011000;
assign LUT_4[49546] = 32'b00000000000000001100111010000100;
assign LUT_4[49547] = 32'b00000000000000000110000101111100;
assign LUT_4[49548] = 32'b00000000000000001010011111111100;
assign LUT_4[49549] = 32'b00000000000000000011101011110100;
assign LUT_4[49550] = 32'b00000000000000001001111010100000;
assign LUT_4[49551] = 32'b00000000000000000011000110011000;
assign LUT_4[49552] = 32'b00000000000000010010000100111001;
assign LUT_4[49553] = 32'b00000000000000001011010000110001;
assign LUT_4[49554] = 32'b00000000000000010001011111011101;
assign LUT_4[49555] = 32'b00000000000000001010101011010101;
assign LUT_4[49556] = 32'b00000000000000001111000101010101;
assign LUT_4[49557] = 32'b00000000000000001000010001001101;
assign LUT_4[49558] = 32'b00000000000000001110011111111001;
assign LUT_4[49559] = 32'b00000000000000000111101011110001;
assign LUT_4[49560] = 32'b00000000000000001011010001001110;
assign LUT_4[49561] = 32'b00000000000000000100011101000110;
assign LUT_4[49562] = 32'b00000000000000001010101011110010;
assign LUT_4[49563] = 32'b00000000000000000011110111101010;
assign LUT_4[49564] = 32'b00000000000000001000010001101010;
assign LUT_4[49565] = 32'b00000000000000000001011101100010;
assign LUT_4[49566] = 32'b00000000000000000111101100001110;
assign LUT_4[49567] = 32'b00000000000000000000111000000110;
assign LUT_4[49568] = 32'b00000000000000010010101110010010;
assign LUT_4[49569] = 32'b00000000000000001011111010001010;
assign LUT_4[49570] = 32'b00000000000000010010001000110110;
assign LUT_4[49571] = 32'b00000000000000001011010100101110;
assign LUT_4[49572] = 32'b00000000000000001111101110101110;
assign LUT_4[49573] = 32'b00000000000000001000111010100110;
assign LUT_4[49574] = 32'b00000000000000001111001001010010;
assign LUT_4[49575] = 32'b00000000000000001000010101001010;
assign LUT_4[49576] = 32'b00000000000000001011111010100111;
assign LUT_4[49577] = 32'b00000000000000000101000110011111;
assign LUT_4[49578] = 32'b00000000000000001011010101001011;
assign LUT_4[49579] = 32'b00000000000000000100100001000011;
assign LUT_4[49580] = 32'b00000000000000001000111011000011;
assign LUT_4[49581] = 32'b00000000000000000010000110111011;
assign LUT_4[49582] = 32'b00000000000000001000010101100111;
assign LUT_4[49583] = 32'b00000000000000000001100001011111;
assign LUT_4[49584] = 32'b00000000000000010000100000000000;
assign LUT_4[49585] = 32'b00000000000000001001101011111000;
assign LUT_4[49586] = 32'b00000000000000001111111010100100;
assign LUT_4[49587] = 32'b00000000000000001001000110011100;
assign LUT_4[49588] = 32'b00000000000000001101100000011100;
assign LUT_4[49589] = 32'b00000000000000000110101100010100;
assign LUT_4[49590] = 32'b00000000000000001100111011000000;
assign LUT_4[49591] = 32'b00000000000000000110000110111000;
assign LUT_4[49592] = 32'b00000000000000001001101100010101;
assign LUT_4[49593] = 32'b00000000000000000010111000001101;
assign LUT_4[49594] = 32'b00000000000000001001000110111001;
assign LUT_4[49595] = 32'b00000000000000000010010010110001;
assign LUT_4[49596] = 32'b00000000000000000110101100110001;
assign LUT_4[49597] = 32'b11111111111111111111111000101001;
assign LUT_4[49598] = 32'b00000000000000000110000111010101;
assign LUT_4[49599] = 32'b11111111111111111111010011001101;
assign LUT_4[49600] = 32'b00000000000000010101101010011111;
assign LUT_4[49601] = 32'b00000000000000001110110110010111;
assign LUT_4[49602] = 32'b00000000000000010101000101000011;
assign LUT_4[49603] = 32'b00000000000000001110010000111011;
assign LUT_4[49604] = 32'b00000000000000010010101010111011;
assign LUT_4[49605] = 32'b00000000000000001011110110110011;
assign LUT_4[49606] = 32'b00000000000000010010000101011111;
assign LUT_4[49607] = 32'b00000000000000001011010001010111;
assign LUT_4[49608] = 32'b00000000000000001110110110110100;
assign LUT_4[49609] = 32'b00000000000000001000000010101100;
assign LUT_4[49610] = 32'b00000000000000001110010001011000;
assign LUT_4[49611] = 32'b00000000000000000111011101010000;
assign LUT_4[49612] = 32'b00000000000000001011110111010000;
assign LUT_4[49613] = 32'b00000000000000000101000011001000;
assign LUT_4[49614] = 32'b00000000000000001011010001110100;
assign LUT_4[49615] = 32'b00000000000000000100011101101100;
assign LUT_4[49616] = 32'b00000000000000010011011100001101;
assign LUT_4[49617] = 32'b00000000000000001100101000000101;
assign LUT_4[49618] = 32'b00000000000000010010110110110001;
assign LUT_4[49619] = 32'b00000000000000001100000010101001;
assign LUT_4[49620] = 32'b00000000000000010000011100101001;
assign LUT_4[49621] = 32'b00000000000000001001101000100001;
assign LUT_4[49622] = 32'b00000000000000001111110111001101;
assign LUT_4[49623] = 32'b00000000000000001001000011000101;
assign LUT_4[49624] = 32'b00000000000000001100101000100010;
assign LUT_4[49625] = 32'b00000000000000000101110100011010;
assign LUT_4[49626] = 32'b00000000000000001100000011000110;
assign LUT_4[49627] = 32'b00000000000000000101001110111110;
assign LUT_4[49628] = 32'b00000000000000001001101000111110;
assign LUT_4[49629] = 32'b00000000000000000010110100110110;
assign LUT_4[49630] = 32'b00000000000000001001000011100010;
assign LUT_4[49631] = 32'b00000000000000000010001111011010;
assign LUT_4[49632] = 32'b00000000000000010100000101100110;
assign LUT_4[49633] = 32'b00000000000000001101010001011110;
assign LUT_4[49634] = 32'b00000000000000010011100000001010;
assign LUT_4[49635] = 32'b00000000000000001100101100000010;
assign LUT_4[49636] = 32'b00000000000000010001000110000010;
assign LUT_4[49637] = 32'b00000000000000001010010001111010;
assign LUT_4[49638] = 32'b00000000000000010000100000100110;
assign LUT_4[49639] = 32'b00000000000000001001101100011110;
assign LUT_4[49640] = 32'b00000000000000001101010001111011;
assign LUT_4[49641] = 32'b00000000000000000110011101110011;
assign LUT_4[49642] = 32'b00000000000000001100101100011111;
assign LUT_4[49643] = 32'b00000000000000000101111000010111;
assign LUT_4[49644] = 32'b00000000000000001010010010010111;
assign LUT_4[49645] = 32'b00000000000000000011011110001111;
assign LUT_4[49646] = 32'b00000000000000001001101100111011;
assign LUT_4[49647] = 32'b00000000000000000010111000110011;
assign LUT_4[49648] = 32'b00000000000000010001110111010100;
assign LUT_4[49649] = 32'b00000000000000001011000011001100;
assign LUT_4[49650] = 32'b00000000000000010001010001111000;
assign LUT_4[49651] = 32'b00000000000000001010011101110000;
assign LUT_4[49652] = 32'b00000000000000001110110111110000;
assign LUT_4[49653] = 32'b00000000000000001000000011101000;
assign LUT_4[49654] = 32'b00000000000000001110010010010100;
assign LUT_4[49655] = 32'b00000000000000000111011110001100;
assign LUT_4[49656] = 32'b00000000000000001011000011101001;
assign LUT_4[49657] = 32'b00000000000000000100001111100001;
assign LUT_4[49658] = 32'b00000000000000001010011110001101;
assign LUT_4[49659] = 32'b00000000000000000011101010000101;
assign LUT_4[49660] = 32'b00000000000000001000000100000101;
assign LUT_4[49661] = 32'b00000000000000000001001111111101;
assign LUT_4[49662] = 32'b00000000000000000111011110101001;
assign LUT_4[49663] = 32'b00000000000000000000101010100001;
assign LUT_4[49664] = 32'b00000000000000001011110101101000;
assign LUT_4[49665] = 32'b00000000000000000101000001100000;
assign LUT_4[49666] = 32'b00000000000000001011010000001100;
assign LUT_4[49667] = 32'b00000000000000000100011100000100;
assign LUT_4[49668] = 32'b00000000000000001000110110000100;
assign LUT_4[49669] = 32'b00000000000000000010000001111100;
assign LUT_4[49670] = 32'b00000000000000001000010000101000;
assign LUT_4[49671] = 32'b00000000000000000001011100100000;
assign LUT_4[49672] = 32'b00000000000000000101000001111101;
assign LUT_4[49673] = 32'b11111111111111111110001101110101;
assign LUT_4[49674] = 32'b00000000000000000100011100100001;
assign LUT_4[49675] = 32'b11111111111111111101101000011001;
assign LUT_4[49676] = 32'b00000000000000000010000010011001;
assign LUT_4[49677] = 32'b11111111111111111011001110010001;
assign LUT_4[49678] = 32'b00000000000000000001011100111101;
assign LUT_4[49679] = 32'b11111111111111111010101000110101;
assign LUT_4[49680] = 32'b00000000000000001001100111010110;
assign LUT_4[49681] = 32'b00000000000000000010110011001110;
assign LUT_4[49682] = 32'b00000000000000001001000001111010;
assign LUT_4[49683] = 32'b00000000000000000010001101110010;
assign LUT_4[49684] = 32'b00000000000000000110100111110010;
assign LUT_4[49685] = 32'b11111111111111111111110011101010;
assign LUT_4[49686] = 32'b00000000000000000110000010010110;
assign LUT_4[49687] = 32'b11111111111111111111001110001110;
assign LUT_4[49688] = 32'b00000000000000000010110011101011;
assign LUT_4[49689] = 32'b11111111111111111011111111100011;
assign LUT_4[49690] = 32'b00000000000000000010001110001111;
assign LUT_4[49691] = 32'b11111111111111111011011010000111;
assign LUT_4[49692] = 32'b11111111111111111111110100000111;
assign LUT_4[49693] = 32'b11111111111111111000111111111111;
assign LUT_4[49694] = 32'b11111111111111111111001110101011;
assign LUT_4[49695] = 32'b11111111111111111000011010100011;
assign LUT_4[49696] = 32'b00000000000000001010010000101111;
assign LUT_4[49697] = 32'b00000000000000000011011100100111;
assign LUT_4[49698] = 32'b00000000000000001001101011010011;
assign LUT_4[49699] = 32'b00000000000000000010110111001011;
assign LUT_4[49700] = 32'b00000000000000000111010001001011;
assign LUT_4[49701] = 32'b00000000000000000000011101000011;
assign LUT_4[49702] = 32'b00000000000000000110101011101111;
assign LUT_4[49703] = 32'b11111111111111111111110111100111;
assign LUT_4[49704] = 32'b00000000000000000011011101000100;
assign LUT_4[49705] = 32'b11111111111111111100101000111100;
assign LUT_4[49706] = 32'b00000000000000000010110111101000;
assign LUT_4[49707] = 32'b11111111111111111100000011100000;
assign LUT_4[49708] = 32'b00000000000000000000011101100000;
assign LUT_4[49709] = 32'b11111111111111111001101001011000;
assign LUT_4[49710] = 32'b11111111111111111111111000000100;
assign LUT_4[49711] = 32'b11111111111111111001000011111100;
assign LUT_4[49712] = 32'b00000000000000001000000010011101;
assign LUT_4[49713] = 32'b00000000000000000001001110010101;
assign LUT_4[49714] = 32'b00000000000000000111011101000001;
assign LUT_4[49715] = 32'b00000000000000000000101000111001;
assign LUT_4[49716] = 32'b00000000000000000101000010111001;
assign LUT_4[49717] = 32'b11111111111111111110001110110001;
assign LUT_4[49718] = 32'b00000000000000000100011101011101;
assign LUT_4[49719] = 32'b11111111111111111101101001010101;
assign LUT_4[49720] = 32'b00000000000000000001001110110010;
assign LUT_4[49721] = 32'b11111111111111111010011010101010;
assign LUT_4[49722] = 32'b00000000000000000000101001010110;
assign LUT_4[49723] = 32'b11111111111111111001110101001110;
assign LUT_4[49724] = 32'b11111111111111111110001111001110;
assign LUT_4[49725] = 32'b11111111111111110111011011000110;
assign LUT_4[49726] = 32'b11111111111111111101101001110010;
assign LUT_4[49727] = 32'b11111111111111110110110101101010;
assign LUT_4[49728] = 32'b00000000000000001101001100111100;
assign LUT_4[49729] = 32'b00000000000000000110011000110100;
assign LUT_4[49730] = 32'b00000000000000001100100111100000;
assign LUT_4[49731] = 32'b00000000000000000101110011011000;
assign LUT_4[49732] = 32'b00000000000000001010001101011000;
assign LUT_4[49733] = 32'b00000000000000000011011001010000;
assign LUT_4[49734] = 32'b00000000000000001001100111111100;
assign LUT_4[49735] = 32'b00000000000000000010110011110100;
assign LUT_4[49736] = 32'b00000000000000000110011001010001;
assign LUT_4[49737] = 32'b11111111111111111111100101001001;
assign LUT_4[49738] = 32'b00000000000000000101110011110101;
assign LUT_4[49739] = 32'b11111111111111111110111111101101;
assign LUT_4[49740] = 32'b00000000000000000011011001101101;
assign LUT_4[49741] = 32'b11111111111111111100100101100101;
assign LUT_4[49742] = 32'b00000000000000000010110100010001;
assign LUT_4[49743] = 32'b11111111111111111100000000001001;
assign LUT_4[49744] = 32'b00000000000000001010111110101010;
assign LUT_4[49745] = 32'b00000000000000000100001010100010;
assign LUT_4[49746] = 32'b00000000000000001010011001001110;
assign LUT_4[49747] = 32'b00000000000000000011100101000110;
assign LUT_4[49748] = 32'b00000000000000000111111111000110;
assign LUT_4[49749] = 32'b00000000000000000001001010111110;
assign LUT_4[49750] = 32'b00000000000000000111011001101010;
assign LUT_4[49751] = 32'b00000000000000000000100101100010;
assign LUT_4[49752] = 32'b00000000000000000100001010111111;
assign LUT_4[49753] = 32'b11111111111111111101010110110111;
assign LUT_4[49754] = 32'b00000000000000000011100101100011;
assign LUT_4[49755] = 32'b11111111111111111100110001011011;
assign LUT_4[49756] = 32'b00000000000000000001001011011011;
assign LUT_4[49757] = 32'b11111111111111111010010111010011;
assign LUT_4[49758] = 32'b00000000000000000000100101111111;
assign LUT_4[49759] = 32'b11111111111111111001110001110111;
assign LUT_4[49760] = 32'b00000000000000001011101000000011;
assign LUT_4[49761] = 32'b00000000000000000100110011111011;
assign LUT_4[49762] = 32'b00000000000000001011000010100111;
assign LUT_4[49763] = 32'b00000000000000000100001110011111;
assign LUT_4[49764] = 32'b00000000000000001000101000011111;
assign LUT_4[49765] = 32'b00000000000000000001110100010111;
assign LUT_4[49766] = 32'b00000000000000001000000011000011;
assign LUT_4[49767] = 32'b00000000000000000001001110111011;
assign LUT_4[49768] = 32'b00000000000000000100110100011000;
assign LUT_4[49769] = 32'b11111111111111111110000000010000;
assign LUT_4[49770] = 32'b00000000000000000100001110111100;
assign LUT_4[49771] = 32'b11111111111111111101011010110100;
assign LUT_4[49772] = 32'b00000000000000000001110100110100;
assign LUT_4[49773] = 32'b11111111111111111011000000101100;
assign LUT_4[49774] = 32'b00000000000000000001001111011000;
assign LUT_4[49775] = 32'b11111111111111111010011011010000;
assign LUT_4[49776] = 32'b00000000000000001001011001110001;
assign LUT_4[49777] = 32'b00000000000000000010100101101001;
assign LUT_4[49778] = 32'b00000000000000001000110100010101;
assign LUT_4[49779] = 32'b00000000000000000010000000001101;
assign LUT_4[49780] = 32'b00000000000000000110011010001101;
assign LUT_4[49781] = 32'b11111111111111111111100110000101;
assign LUT_4[49782] = 32'b00000000000000000101110100110001;
assign LUT_4[49783] = 32'b11111111111111111111000000101001;
assign LUT_4[49784] = 32'b00000000000000000010100110000110;
assign LUT_4[49785] = 32'b11111111111111111011110001111110;
assign LUT_4[49786] = 32'b00000000000000000010000000101010;
assign LUT_4[49787] = 32'b11111111111111111011001100100010;
assign LUT_4[49788] = 32'b11111111111111111111100110100010;
assign LUT_4[49789] = 32'b11111111111111111000110010011010;
assign LUT_4[49790] = 32'b11111111111111111111000001000110;
assign LUT_4[49791] = 32'b11111111111111111000001100111110;
assign LUT_4[49792] = 32'b00000000000000001110011011110000;
assign LUT_4[49793] = 32'b00000000000000000111100111101000;
assign LUT_4[49794] = 32'b00000000000000001101110110010100;
assign LUT_4[49795] = 32'b00000000000000000111000010001100;
assign LUT_4[49796] = 32'b00000000000000001011011100001100;
assign LUT_4[49797] = 32'b00000000000000000100101000000100;
assign LUT_4[49798] = 32'b00000000000000001010110110110000;
assign LUT_4[49799] = 32'b00000000000000000100000010101000;
assign LUT_4[49800] = 32'b00000000000000000111101000000101;
assign LUT_4[49801] = 32'b00000000000000000000110011111101;
assign LUT_4[49802] = 32'b00000000000000000111000010101001;
assign LUT_4[49803] = 32'b00000000000000000000001110100001;
assign LUT_4[49804] = 32'b00000000000000000100101000100001;
assign LUT_4[49805] = 32'b11111111111111111101110100011001;
assign LUT_4[49806] = 32'b00000000000000000100000011000101;
assign LUT_4[49807] = 32'b11111111111111111101001110111101;
assign LUT_4[49808] = 32'b00000000000000001100001101011110;
assign LUT_4[49809] = 32'b00000000000000000101011001010110;
assign LUT_4[49810] = 32'b00000000000000001011101000000010;
assign LUT_4[49811] = 32'b00000000000000000100110011111010;
assign LUT_4[49812] = 32'b00000000000000001001001101111010;
assign LUT_4[49813] = 32'b00000000000000000010011001110010;
assign LUT_4[49814] = 32'b00000000000000001000101000011110;
assign LUT_4[49815] = 32'b00000000000000000001110100010110;
assign LUT_4[49816] = 32'b00000000000000000101011001110011;
assign LUT_4[49817] = 32'b11111111111111111110100101101011;
assign LUT_4[49818] = 32'b00000000000000000100110100010111;
assign LUT_4[49819] = 32'b11111111111111111110000000001111;
assign LUT_4[49820] = 32'b00000000000000000010011010001111;
assign LUT_4[49821] = 32'b11111111111111111011100110000111;
assign LUT_4[49822] = 32'b00000000000000000001110100110011;
assign LUT_4[49823] = 32'b11111111111111111011000000101011;
assign LUT_4[49824] = 32'b00000000000000001100110110110111;
assign LUT_4[49825] = 32'b00000000000000000110000010101111;
assign LUT_4[49826] = 32'b00000000000000001100010001011011;
assign LUT_4[49827] = 32'b00000000000000000101011101010011;
assign LUT_4[49828] = 32'b00000000000000001001110111010011;
assign LUT_4[49829] = 32'b00000000000000000011000011001011;
assign LUT_4[49830] = 32'b00000000000000001001010001110111;
assign LUT_4[49831] = 32'b00000000000000000010011101101111;
assign LUT_4[49832] = 32'b00000000000000000110000011001100;
assign LUT_4[49833] = 32'b11111111111111111111001111000100;
assign LUT_4[49834] = 32'b00000000000000000101011101110000;
assign LUT_4[49835] = 32'b11111111111111111110101001101000;
assign LUT_4[49836] = 32'b00000000000000000011000011101000;
assign LUT_4[49837] = 32'b11111111111111111100001111100000;
assign LUT_4[49838] = 32'b00000000000000000010011110001100;
assign LUT_4[49839] = 32'b11111111111111111011101010000100;
assign LUT_4[49840] = 32'b00000000000000001010101000100101;
assign LUT_4[49841] = 32'b00000000000000000011110100011101;
assign LUT_4[49842] = 32'b00000000000000001010000011001001;
assign LUT_4[49843] = 32'b00000000000000000011001111000001;
assign LUT_4[49844] = 32'b00000000000000000111101001000001;
assign LUT_4[49845] = 32'b00000000000000000000110100111001;
assign LUT_4[49846] = 32'b00000000000000000111000011100101;
assign LUT_4[49847] = 32'b00000000000000000000001111011101;
assign LUT_4[49848] = 32'b00000000000000000011110100111010;
assign LUT_4[49849] = 32'b11111111111111111101000000110010;
assign LUT_4[49850] = 32'b00000000000000000011001111011110;
assign LUT_4[49851] = 32'b11111111111111111100011011010110;
assign LUT_4[49852] = 32'b00000000000000000000110101010110;
assign LUT_4[49853] = 32'b11111111111111111010000001001110;
assign LUT_4[49854] = 32'b00000000000000000000001111111010;
assign LUT_4[49855] = 32'b11111111111111111001011011110010;
assign LUT_4[49856] = 32'b00000000000000001111110011000100;
assign LUT_4[49857] = 32'b00000000000000001000111110111100;
assign LUT_4[49858] = 32'b00000000000000001111001101101000;
assign LUT_4[49859] = 32'b00000000000000001000011001100000;
assign LUT_4[49860] = 32'b00000000000000001100110011100000;
assign LUT_4[49861] = 32'b00000000000000000101111111011000;
assign LUT_4[49862] = 32'b00000000000000001100001110000100;
assign LUT_4[49863] = 32'b00000000000000000101011001111100;
assign LUT_4[49864] = 32'b00000000000000001000111111011001;
assign LUT_4[49865] = 32'b00000000000000000010001011010001;
assign LUT_4[49866] = 32'b00000000000000001000011001111101;
assign LUT_4[49867] = 32'b00000000000000000001100101110101;
assign LUT_4[49868] = 32'b00000000000000000101111111110101;
assign LUT_4[49869] = 32'b11111111111111111111001011101101;
assign LUT_4[49870] = 32'b00000000000000000101011010011001;
assign LUT_4[49871] = 32'b11111111111111111110100110010001;
assign LUT_4[49872] = 32'b00000000000000001101100100110010;
assign LUT_4[49873] = 32'b00000000000000000110110000101010;
assign LUT_4[49874] = 32'b00000000000000001100111111010110;
assign LUT_4[49875] = 32'b00000000000000000110001011001110;
assign LUT_4[49876] = 32'b00000000000000001010100101001110;
assign LUT_4[49877] = 32'b00000000000000000011110001000110;
assign LUT_4[49878] = 32'b00000000000000001001111111110010;
assign LUT_4[49879] = 32'b00000000000000000011001011101010;
assign LUT_4[49880] = 32'b00000000000000000110110001000111;
assign LUT_4[49881] = 32'b11111111111111111111111100111111;
assign LUT_4[49882] = 32'b00000000000000000110001011101011;
assign LUT_4[49883] = 32'b11111111111111111111010111100011;
assign LUT_4[49884] = 32'b00000000000000000011110001100011;
assign LUT_4[49885] = 32'b11111111111111111100111101011011;
assign LUT_4[49886] = 32'b00000000000000000011001100000111;
assign LUT_4[49887] = 32'b11111111111111111100010111111111;
assign LUT_4[49888] = 32'b00000000000000001110001110001011;
assign LUT_4[49889] = 32'b00000000000000000111011010000011;
assign LUT_4[49890] = 32'b00000000000000001101101000101111;
assign LUT_4[49891] = 32'b00000000000000000110110100100111;
assign LUT_4[49892] = 32'b00000000000000001011001110100111;
assign LUT_4[49893] = 32'b00000000000000000100011010011111;
assign LUT_4[49894] = 32'b00000000000000001010101001001011;
assign LUT_4[49895] = 32'b00000000000000000011110101000011;
assign LUT_4[49896] = 32'b00000000000000000111011010100000;
assign LUT_4[49897] = 32'b00000000000000000000100110011000;
assign LUT_4[49898] = 32'b00000000000000000110110101000100;
assign LUT_4[49899] = 32'b00000000000000000000000000111100;
assign LUT_4[49900] = 32'b00000000000000000100011010111100;
assign LUT_4[49901] = 32'b11111111111111111101100110110100;
assign LUT_4[49902] = 32'b00000000000000000011110101100000;
assign LUT_4[49903] = 32'b11111111111111111101000001011000;
assign LUT_4[49904] = 32'b00000000000000001011111111111001;
assign LUT_4[49905] = 32'b00000000000000000101001011110001;
assign LUT_4[49906] = 32'b00000000000000001011011010011101;
assign LUT_4[49907] = 32'b00000000000000000100100110010101;
assign LUT_4[49908] = 32'b00000000000000001001000000010101;
assign LUT_4[49909] = 32'b00000000000000000010001100001101;
assign LUT_4[49910] = 32'b00000000000000001000011010111001;
assign LUT_4[49911] = 32'b00000000000000000001100110110001;
assign LUT_4[49912] = 32'b00000000000000000101001100001110;
assign LUT_4[49913] = 32'b11111111111111111110011000000110;
assign LUT_4[49914] = 32'b00000000000000000100100110110010;
assign LUT_4[49915] = 32'b11111111111111111101110010101010;
assign LUT_4[49916] = 32'b00000000000000000010001100101010;
assign LUT_4[49917] = 32'b11111111111111111011011000100010;
assign LUT_4[49918] = 32'b00000000000000000001100111001110;
assign LUT_4[49919] = 32'b11111111111111111010110011000110;
assign LUT_4[49920] = 32'b00000000000000010000110001001011;
assign LUT_4[49921] = 32'b00000000000000001001111101000011;
assign LUT_4[49922] = 32'b00000000000000010000001011101111;
assign LUT_4[49923] = 32'b00000000000000001001010111100111;
assign LUT_4[49924] = 32'b00000000000000001101110001100111;
assign LUT_4[49925] = 32'b00000000000000000110111101011111;
assign LUT_4[49926] = 32'b00000000000000001101001100001011;
assign LUT_4[49927] = 32'b00000000000000000110011000000011;
assign LUT_4[49928] = 32'b00000000000000001001111101100000;
assign LUT_4[49929] = 32'b00000000000000000011001001011000;
assign LUT_4[49930] = 32'b00000000000000001001011000000100;
assign LUT_4[49931] = 32'b00000000000000000010100011111100;
assign LUT_4[49932] = 32'b00000000000000000110111101111100;
assign LUT_4[49933] = 32'b00000000000000000000001001110100;
assign LUT_4[49934] = 32'b00000000000000000110011000100000;
assign LUT_4[49935] = 32'b11111111111111111111100100011000;
assign LUT_4[49936] = 32'b00000000000000001110100010111001;
assign LUT_4[49937] = 32'b00000000000000000111101110110001;
assign LUT_4[49938] = 32'b00000000000000001101111101011101;
assign LUT_4[49939] = 32'b00000000000000000111001001010101;
assign LUT_4[49940] = 32'b00000000000000001011100011010101;
assign LUT_4[49941] = 32'b00000000000000000100101111001101;
assign LUT_4[49942] = 32'b00000000000000001010111101111001;
assign LUT_4[49943] = 32'b00000000000000000100001001110001;
assign LUT_4[49944] = 32'b00000000000000000111101111001110;
assign LUT_4[49945] = 32'b00000000000000000000111011000110;
assign LUT_4[49946] = 32'b00000000000000000111001001110010;
assign LUT_4[49947] = 32'b00000000000000000000010101101010;
assign LUT_4[49948] = 32'b00000000000000000100101111101010;
assign LUT_4[49949] = 32'b11111111111111111101111011100010;
assign LUT_4[49950] = 32'b00000000000000000100001010001110;
assign LUT_4[49951] = 32'b11111111111111111101010110000110;
assign LUT_4[49952] = 32'b00000000000000001111001100010010;
assign LUT_4[49953] = 32'b00000000000000001000011000001010;
assign LUT_4[49954] = 32'b00000000000000001110100110110110;
assign LUT_4[49955] = 32'b00000000000000000111110010101110;
assign LUT_4[49956] = 32'b00000000000000001100001100101110;
assign LUT_4[49957] = 32'b00000000000000000101011000100110;
assign LUT_4[49958] = 32'b00000000000000001011100111010010;
assign LUT_4[49959] = 32'b00000000000000000100110011001010;
assign LUT_4[49960] = 32'b00000000000000001000011000100111;
assign LUT_4[49961] = 32'b00000000000000000001100100011111;
assign LUT_4[49962] = 32'b00000000000000000111110011001011;
assign LUT_4[49963] = 32'b00000000000000000000111111000011;
assign LUT_4[49964] = 32'b00000000000000000101011001000011;
assign LUT_4[49965] = 32'b11111111111111111110100100111011;
assign LUT_4[49966] = 32'b00000000000000000100110011100111;
assign LUT_4[49967] = 32'b11111111111111111101111111011111;
assign LUT_4[49968] = 32'b00000000000000001100111110000000;
assign LUT_4[49969] = 32'b00000000000000000110001001111000;
assign LUT_4[49970] = 32'b00000000000000001100011000100100;
assign LUT_4[49971] = 32'b00000000000000000101100100011100;
assign LUT_4[49972] = 32'b00000000000000001001111110011100;
assign LUT_4[49973] = 32'b00000000000000000011001010010100;
assign LUT_4[49974] = 32'b00000000000000001001011001000000;
assign LUT_4[49975] = 32'b00000000000000000010100100111000;
assign LUT_4[49976] = 32'b00000000000000000110001010010101;
assign LUT_4[49977] = 32'b11111111111111111111010110001101;
assign LUT_4[49978] = 32'b00000000000000000101100100111001;
assign LUT_4[49979] = 32'b11111111111111111110110000110001;
assign LUT_4[49980] = 32'b00000000000000000011001010110001;
assign LUT_4[49981] = 32'b11111111111111111100010110101001;
assign LUT_4[49982] = 32'b00000000000000000010100101010101;
assign LUT_4[49983] = 32'b11111111111111111011110001001101;
assign LUT_4[49984] = 32'b00000000000000010010001000011111;
assign LUT_4[49985] = 32'b00000000000000001011010100010111;
assign LUT_4[49986] = 32'b00000000000000010001100011000011;
assign LUT_4[49987] = 32'b00000000000000001010101110111011;
assign LUT_4[49988] = 32'b00000000000000001111001000111011;
assign LUT_4[49989] = 32'b00000000000000001000010100110011;
assign LUT_4[49990] = 32'b00000000000000001110100011011111;
assign LUT_4[49991] = 32'b00000000000000000111101111010111;
assign LUT_4[49992] = 32'b00000000000000001011010100110100;
assign LUT_4[49993] = 32'b00000000000000000100100000101100;
assign LUT_4[49994] = 32'b00000000000000001010101111011000;
assign LUT_4[49995] = 32'b00000000000000000011111011010000;
assign LUT_4[49996] = 32'b00000000000000001000010101010000;
assign LUT_4[49997] = 32'b00000000000000000001100001001000;
assign LUT_4[49998] = 32'b00000000000000000111101111110100;
assign LUT_4[49999] = 32'b00000000000000000000111011101100;
assign LUT_4[50000] = 32'b00000000000000001111111010001101;
assign LUT_4[50001] = 32'b00000000000000001001000110000101;
assign LUT_4[50002] = 32'b00000000000000001111010100110001;
assign LUT_4[50003] = 32'b00000000000000001000100000101001;
assign LUT_4[50004] = 32'b00000000000000001100111010101001;
assign LUT_4[50005] = 32'b00000000000000000110000110100001;
assign LUT_4[50006] = 32'b00000000000000001100010101001101;
assign LUT_4[50007] = 32'b00000000000000000101100001000101;
assign LUT_4[50008] = 32'b00000000000000001001000110100010;
assign LUT_4[50009] = 32'b00000000000000000010010010011010;
assign LUT_4[50010] = 32'b00000000000000001000100001000110;
assign LUT_4[50011] = 32'b00000000000000000001101100111110;
assign LUT_4[50012] = 32'b00000000000000000110000110111110;
assign LUT_4[50013] = 32'b11111111111111111111010010110110;
assign LUT_4[50014] = 32'b00000000000000000101100001100010;
assign LUT_4[50015] = 32'b11111111111111111110101101011010;
assign LUT_4[50016] = 32'b00000000000000010000100011100110;
assign LUT_4[50017] = 32'b00000000000000001001101111011110;
assign LUT_4[50018] = 32'b00000000000000001111111110001010;
assign LUT_4[50019] = 32'b00000000000000001001001010000010;
assign LUT_4[50020] = 32'b00000000000000001101100100000010;
assign LUT_4[50021] = 32'b00000000000000000110101111111010;
assign LUT_4[50022] = 32'b00000000000000001100111110100110;
assign LUT_4[50023] = 32'b00000000000000000110001010011110;
assign LUT_4[50024] = 32'b00000000000000001001101111111011;
assign LUT_4[50025] = 32'b00000000000000000010111011110011;
assign LUT_4[50026] = 32'b00000000000000001001001010011111;
assign LUT_4[50027] = 32'b00000000000000000010010110010111;
assign LUT_4[50028] = 32'b00000000000000000110110000010111;
assign LUT_4[50029] = 32'b11111111111111111111111100001111;
assign LUT_4[50030] = 32'b00000000000000000110001010111011;
assign LUT_4[50031] = 32'b11111111111111111111010110110011;
assign LUT_4[50032] = 32'b00000000000000001110010101010100;
assign LUT_4[50033] = 32'b00000000000000000111100001001100;
assign LUT_4[50034] = 32'b00000000000000001101101111111000;
assign LUT_4[50035] = 32'b00000000000000000110111011110000;
assign LUT_4[50036] = 32'b00000000000000001011010101110000;
assign LUT_4[50037] = 32'b00000000000000000100100001101000;
assign LUT_4[50038] = 32'b00000000000000001010110000010100;
assign LUT_4[50039] = 32'b00000000000000000011111100001100;
assign LUT_4[50040] = 32'b00000000000000000111100001101001;
assign LUT_4[50041] = 32'b00000000000000000000101101100001;
assign LUT_4[50042] = 32'b00000000000000000110111100001101;
assign LUT_4[50043] = 32'b00000000000000000000001000000101;
assign LUT_4[50044] = 32'b00000000000000000100100010000101;
assign LUT_4[50045] = 32'b11111111111111111101101101111101;
assign LUT_4[50046] = 32'b00000000000000000011111100101001;
assign LUT_4[50047] = 32'b11111111111111111101001000100001;
assign LUT_4[50048] = 32'b00000000000000010011010111010011;
assign LUT_4[50049] = 32'b00000000000000001100100011001011;
assign LUT_4[50050] = 32'b00000000000000010010110001110111;
assign LUT_4[50051] = 32'b00000000000000001011111101101111;
assign LUT_4[50052] = 32'b00000000000000010000010111101111;
assign LUT_4[50053] = 32'b00000000000000001001100011100111;
assign LUT_4[50054] = 32'b00000000000000001111110010010011;
assign LUT_4[50055] = 32'b00000000000000001000111110001011;
assign LUT_4[50056] = 32'b00000000000000001100100011101000;
assign LUT_4[50057] = 32'b00000000000000000101101111100000;
assign LUT_4[50058] = 32'b00000000000000001011111110001100;
assign LUT_4[50059] = 32'b00000000000000000101001010000100;
assign LUT_4[50060] = 32'b00000000000000001001100100000100;
assign LUT_4[50061] = 32'b00000000000000000010101111111100;
assign LUT_4[50062] = 32'b00000000000000001000111110101000;
assign LUT_4[50063] = 32'b00000000000000000010001010100000;
assign LUT_4[50064] = 32'b00000000000000010001001001000001;
assign LUT_4[50065] = 32'b00000000000000001010010100111001;
assign LUT_4[50066] = 32'b00000000000000010000100011100101;
assign LUT_4[50067] = 32'b00000000000000001001101111011101;
assign LUT_4[50068] = 32'b00000000000000001110001001011101;
assign LUT_4[50069] = 32'b00000000000000000111010101010101;
assign LUT_4[50070] = 32'b00000000000000001101100100000001;
assign LUT_4[50071] = 32'b00000000000000000110101111111001;
assign LUT_4[50072] = 32'b00000000000000001010010101010110;
assign LUT_4[50073] = 32'b00000000000000000011100001001110;
assign LUT_4[50074] = 32'b00000000000000001001101111111010;
assign LUT_4[50075] = 32'b00000000000000000010111011110010;
assign LUT_4[50076] = 32'b00000000000000000111010101110010;
assign LUT_4[50077] = 32'b00000000000000000000100001101010;
assign LUT_4[50078] = 32'b00000000000000000110110000010110;
assign LUT_4[50079] = 32'b11111111111111111111111100001110;
assign LUT_4[50080] = 32'b00000000000000010001110010011010;
assign LUT_4[50081] = 32'b00000000000000001010111110010010;
assign LUT_4[50082] = 32'b00000000000000010001001100111110;
assign LUT_4[50083] = 32'b00000000000000001010011000110110;
assign LUT_4[50084] = 32'b00000000000000001110110010110110;
assign LUT_4[50085] = 32'b00000000000000000111111110101110;
assign LUT_4[50086] = 32'b00000000000000001110001101011010;
assign LUT_4[50087] = 32'b00000000000000000111011001010010;
assign LUT_4[50088] = 32'b00000000000000001010111110101111;
assign LUT_4[50089] = 32'b00000000000000000100001010100111;
assign LUT_4[50090] = 32'b00000000000000001010011001010011;
assign LUT_4[50091] = 32'b00000000000000000011100101001011;
assign LUT_4[50092] = 32'b00000000000000000111111111001011;
assign LUT_4[50093] = 32'b00000000000000000001001011000011;
assign LUT_4[50094] = 32'b00000000000000000111011001101111;
assign LUT_4[50095] = 32'b00000000000000000000100101100111;
assign LUT_4[50096] = 32'b00000000000000001111100100001000;
assign LUT_4[50097] = 32'b00000000000000001000110000000000;
assign LUT_4[50098] = 32'b00000000000000001110111110101100;
assign LUT_4[50099] = 32'b00000000000000001000001010100100;
assign LUT_4[50100] = 32'b00000000000000001100100100100100;
assign LUT_4[50101] = 32'b00000000000000000101110000011100;
assign LUT_4[50102] = 32'b00000000000000001011111111001000;
assign LUT_4[50103] = 32'b00000000000000000101001011000000;
assign LUT_4[50104] = 32'b00000000000000001000110000011101;
assign LUT_4[50105] = 32'b00000000000000000001111100010101;
assign LUT_4[50106] = 32'b00000000000000001000001011000001;
assign LUT_4[50107] = 32'b00000000000000000001010110111001;
assign LUT_4[50108] = 32'b00000000000000000101110000111001;
assign LUT_4[50109] = 32'b11111111111111111110111100110001;
assign LUT_4[50110] = 32'b00000000000000000101001011011101;
assign LUT_4[50111] = 32'b11111111111111111110010111010101;
assign LUT_4[50112] = 32'b00000000000000010100101110100111;
assign LUT_4[50113] = 32'b00000000000000001101111010011111;
assign LUT_4[50114] = 32'b00000000000000010100001001001011;
assign LUT_4[50115] = 32'b00000000000000001101010101000011;
assign LUT_4[50116] = 32'b00000000000000010001101111000011;
assign LUT_4[50117] = 32'b00000000000000001010111010111011;
assign LUT_4[50118] = 32'b00000000000000010001001001100111;
assign LUT_4[50119] = 32'b00000000000000001010010101011111;
assign LUT_4[50120] = 32'b00000000000000001101111010111100;
assign LUT_4[50121] = 32'b00000000000000000111000110110100;
assign LUT_4[50122] = 32'b00000000000000001101010101100000;
assign LUT_4[50123] = 32'b00000000000000000110100001011000;
assign LUT_4[50124] = 32'b00000000000000001010111011011000;
assign LUT_4[50125] = 32'b00000000000000000100000111010000;
assign LUT_4[50126] = 32'b00000000000000001010010101111100;
assign LUT_4[50127] = 32'b00000000000000000011100001110100;
assign LUT_4[50128] = 32'b00000000000000010010100000010101;
assign LUT_4[50129] = 32'b00000000000000001011101100001101;
assign LUT_4[50130] = 32'b00000000000000010001111010111001;
assign LUT_4[50131] = 32'b00000000000000001011000110110001;
assign LUT_4[50132] = 32'b00000000000000001111100000110001;
assign LUT_4[50133] = 32'b00000000000000001000101100101001;
assign LUT_4[50134] = 32'b00000000000000001110111011010101;
assign LUT_4[50135] = 32'b00000000000000001000000111001101;
assign LUT_4[50136] = 32'b00000000000000001011101100101010;
assign LUT_4[50137] = 32'b00000000000000000100111000100010;
assign LUT_4[50138] = 32'b00000000000000001011000111001110;
assign LUT_4[50139] = 32'b00000000000000000100010011000110;
assign LUT_4[50140] = 32'b00000000000000001000101101000110;
assign LUT_4[50141] = 32'b00000000000000000001111000111110;
assign LUT_4[50142] = 32'b00000000000000001000000111101010;
assign LUT_4[50143] = 32'b00000000000000000001010011100010;
assign LUT_4[50144] = 32'b00000000000000010011001001101110;
assign LUT_4[50145] = 32'b00000000000000001100010101100110;
assign LUT_4[50146] = 32'b00000000000000010010100100010010;
assign LUT_4[50147] = 32'b00000000000000001011110000001010;
assign LUT_4[50148] = 32'b00000000000000010000001010001010;
assign LUT_4[50149] = 32'b00000000000000001001010110000010;
assign LUT_4[50150] = 32'b00000000000000001111100100101110;
assign LUT_4[50151] = 32'b00000000000000001000110000100110;
assign LUT_4[50152] = 32'b00000000000000001100010110000011;
assign LUT_4[50153] = 32'b00000000000000000101100001111011;
assign LUT_4[50154] = 32'b00000000000000001011110000100111;
assign LUT_4[50155] = 32'b00000000000000000100111100011111;
assign LUT_4[50156] = 32'b00000000000000001001010110011111;
assign LUT_4[50157] = 32'b00000000000000000010100010010111;
assign LUT_4[50158] = 32'b00000000000000001000110001000011;
assign LUT_4[50159] = 32'b00000000000000000001111100111011;
assign LUT_4[50160] = 32'b00000000000000010000111011011100;
assign LUT_4[50161] = 32'b00000000000000001010000111010100;
assign LUT_4[50162] = 32'b00000000000000010000010110000000;
assign LUT_4[50163] = 32'b00000000000000001001100001111000;
assign LUT_4[50164] = 32'b00000000000000001101111011111000;
assign LUT_4[50165] = 32'b00000000000000000111000111110000;
assign LUT_4[50166] = 32'b00000000000000001101010110011100;
assign LUT_4[50167] = 32'b00000000000000000110100010010100;
assign LUT_4[50168] = 32'b00000000000000001010000111110001;
assign LUT_4[50169] = 32'b00000000000000000011010011101001;
assign LUT_4[50170] = 32'b00000000000000001001100010010101;
assign LUT_4[50171] = 32'b00000000000000000010101110001101;
assign LUT_4[50172] = 32'b00000000000000000111001000001101;
assign LUT_4[50173] = 32'b00000000000000000000010100000101;
assign LUT_4[50174] = 32'b00000000000000000110100010110001;
assign LUT_4[50175] = 32'b11111111111111111111101110101001;
assign LUT_4[50176] = 32'b00000000000000001110011011111111;
assign LUT_4[50177] = 32'b00000000000000000111100111110111;
assign LUT_4[50178] = 32'b00000000000000001101110110100011;
assign LUT_4[50179] = 32'b00000000000000000111000010011011;
assign LUT_4[50180] = 32'b00000000000000001011011100011011;
assign LUT_4[50181] = 32'b00000000000000000100101000010011;
assign LUT_4[50182] = 32'b00000000000000001010110110111111;
assign LUT_4[50183] = 32'b00000000000000000100000010110111;
assign LUT_4[50184] = 32'b00000000000000000111101000010100;
assign LUT_4[50185] = 32'b00000000000000000000110100001100;
assign LUT_4[50186] = 32'b00000000000000000111000010111000;
assign LUT_4[50187] = 32'b00000000000000000000001110110000;
assign LUT_4[50188] = 32'b00000000000000000100101000110000;
assign LUT_4[50189] = 32'b11111111111111111101110100101000;
assign LUT_4[50190] = 32'b00000000000000000100000011010100;
assign LUT_4[50191] = 32'b11111111111111111101001111001100;
assign LUT_4[50192] = 32'b00000000000000001100001101101101;
assign LUT_4[50193] = 32'b00000000000000000101011001100101;
assign LUT_4[50194] = 32'b00000000000000001011101000010001;
assign LUT_4[50195] = 32'b00000000000000000100110100001001;
assign LUT_4[50196] = 32'b00000000000000001001001110001001;
assign LUT_4[50197] = 32'b00000000000000000010011010000001;
assign LUT_4[50198] = 32'b00000000000000001000101000101101;
assign LUT_4[50199] = 32'b00000000000000000001110100100101;
assign LUT_4[50200] = 32'b00000000000000000101011010000010;
assign LUT_4[50201] = 32'b11111111111111111110100101111010;
assign LUT_4[50202] = 32'b00000000000000000100110100100110;
assign LUT_4[50203] = 32'b11111111111111111110000000011110;
assign LUT_4[50204] = 32'b00000000000000000010011010011110;
assign LUT_4[50205] = 32'b11111111111111111011100110010110;
assign LUT_4[50206] = 32'b00000000000000000001110101000010;
assign LUT_4[50207] = 32'b11111111111111111011000000111010;
assign LUT_4[50208] = 32'b00000000000000001100110111000110;
assign LUT_4[50209] = 32'b00000000000000000110000010111110;
assign LUT_4[50210] = 32'b00000000000000001100010001101010;
assign LUT_4[50211] = 32'b00000000000000000101011101100010;
assign LUT_4[50212] = 32'b00000000000000001001110111100010;
assign LUT_4[50213] = 32'b00000000000000000011000011011010;
assign LUT_4[50214] = 32'b00000000000000001001010010000110;
assign LUT_4[50215] = 32'b00000000000000000010011101111110;
assign LUT_4[50216] = 32'b00000000000000000110000011011011;
assign LUT_4[50217] = 32'b11111111111111111111001111010011;
assign LUT_4[50218] = 32'b00000000000000000101011101111111;
assign LUT_4[50219] = 32'b11111111111111111110101001110111;
assign LUT_4[50220] = 32'b00000000000000000011000011110111;
assign LUT_4[50221] = 32'b11111111111111111100001111101111;
assign LUT_4[50222] = 32'b00000000000000000010011110011011;
assign LUT_4[50223] = 32'b11111111111111111011101010010011;
assign LUT_4[50224] = 32'b00000000000000001010101000110100;
assign LUT_4[50225] = 32'b00000000000000000011110100101100;
assign LUT_4[50226] = 32'b00000000000000001010000011011000;
assign LUT_4[50227] = 32'b00000000000000000011001111010000;
assign LUT_4[50228] = 32'b00000000000000000111101001010000;
assign LUT_4[50229] = 32'b00000000000000000000110101001000;
assign LUT_4[50230] = 32'b00000000000000000111000011110100;
assign LUT_4[50231] = 32'b00000000000000000000001111101100;
assign LUT_4[50232] = 32'b00000000000000000011110101001001;
assign LUT_4[50233] = 32'b11111111111111111101000001000001;
assign LUT_4[50234] = 32'b00000000000000000011001111101101;
assign LUT_4[50235] = 32'b11111111111111111100011011100101;
assign LUT_4[50236] = 32'b00000000000000000000110101100101;
assign LUT_4[50237] = 32'b11111111111111111010000001011101;
assign LUT_4[50238] = 32'b00000000000000000000010000001001;
assign LUT_4[50239] = 32'b11111111111111111001011100000001;
assign LUT_4[50240] = 32'b00000000000000001111110011010011;
assign LUT_4[50241] = 32'b00000000000000001000111111001011;
assign LUT_4[50242] = 32'b00000000000000001111001101110111;
assign LUT_4[50243] = 32'b00000000000000001000011001101111;
assign LUT_4[50244] = 32'b00000000000000001100110011101111;
assign LUT_4[50245] = 32'b00000000000000000101111111100111;
assign LUT_4[50246] = 32'b00000000000000001100001110010011;
assign LUT_4[50247] = 32'b00000000000000000101011010001011;
assign LUT_4[50248] = 32'b00000000000000001000111111101000;
assign LUT_4[50249] = 32'b00000000000000000010001011100000;
assign LUT_4[50250] = 32'b00000000000000001000011010001100;
assign LUT_4[50251] = 32'b00000000000000000001100110000100;
assign LUT_4[50252] = 32'b00000000000000000110000000000100;
assign LUT_4[50253] = 32'b11111111111111111111001011111100;
assign LUT_4[50254] = 32'b00000000000000000101011010101000;
assign LUT_4[50255] = 32'b11111111111111111110100110100000;
assign LUT_4[50256] = 32'b00000000000000001101100101000001;
assign LUT_4[50257] = 32'b00000000000000000110110000111001;
assign LUT_4[50258] = 32'b00000000000000001100111111100101;
assign LUT_4[50259] = 32'b00000000000000000110001011011101;
assign LUT_4[50260] = 32'b00000000000000001010100101011101;
assign LUT_4[50261] = 32'b00000000000000000011110001010101;
assign LUT_4[50262] = 32'b00000000000000001010000000000001;
assign LUT_4[50263] = 32'b00000000000000000011001011111001;
assign LUT_4[50264] = 32'b00000000000000000110110001010110;
assign LUT_4[50265] = 32'b11111111111111111111111101001110;
assign LUT_4[50266] = 32'b00000000000000000110001011111010;
assign LUT_4[50267] = 32'b11111111111111111111010111110010;
assign LUT_4[50268] = 32'b00000000000000000011110001110010;
assign LUT_4[50269] = 32'b11111111111111111100111101101010;
assign LUT_4[50270] = 32'b00000000000000000011001100010110;
assign LUT_4[50271] = 32'b11111111111111111100011000001110;
assign LUT_4[50272] = 32'b00000000000000001110001110011010;
assign LUT_4[50273] = 32'b00000000000000000111011010010010;
assign LUT_4[50274] = 32'b00000000000000001101101000111110;
assign LUT_4[50275] = 32'b00000000000000000110110100110110;
assign LUT_4[50276] = 32'b00000000000000001011001110110110;
assign LUT_4[50277] = 32'b00000000000000000100011010101110;
assign LUT_4[50278] = 32'b00000000000000001010101001011010;
assign LUT_4[50279] = 32'b00000000000000000011110101010010;
assign LUT_4[50280] = 32'b00000000000000000111011010101111;
assign LUT_4[50281] = 32'b00000000000000000000100110100111;
assign LUT_4[50282] = 32'b00000000000000000110110101010011;
assign LUT_4[50283] = 32'b00000000000000000000000001001011;
assign LUT_4[50284] = 32'b00000000000000000100011011001011;
assign LUT_4[50285] = 32'b11111111111111111101100111000011;
assign LUT_4[50286] = 32'b00000000000000000011110101101111;
assign LUT_4[50287] = 32'b11111111111111111101000001100111;
assign LUT_4[50288] = 32'b00000000000000001100000000001000;
assign LUT_4[50289] = 32'b00000000000000000101001100000000;
assign LUT_4[50290] = 32'b00000000000000001011011010101100;
assign LUT_4[50291] = 32'b00000000000000000100100110100100;
assign LUT_4[50292] = 32'b00000000000000001001000000100100;
assign LUT_4[50293] = 32'b00000000000000000010001100011100;
assign LUT_4[50294] = 32'b00000000000000001000011011001000;
assign LUT_4[50295] = 32'b00000000000000000001100111000000;
assign LUT_4[50296] = 32'b00000000000000000101001100011101;
assign LUT_4[50297] = 32'b11111111111111111110011000010101;
assign LUT_4[50298] = 32'b00000000000000000100100111000001;
assign LUT_4[50299] = 32'b11111111111111111101110010111001;
assign LUT_4[50300] = 32'b00000000000000000010001100111001;
assign LUT_4[50301] = 32'b11111111111111111011011000110001;
assign LUT_4[50302] = 32'b00000000000000000001100111011101;
assign LUT_4[50303] = 32'b11111111111111111010110011010101;
assign LUT_4[50304] = 32'b00000000000000010001000010000111;
assign LUT_4[50305] = 32'b00000000000000001010001101111111;
assign LUT_4[50306] = 32'b00000000000000010000011100101011;
assign LUT_4[50307] = 32'b00000000000000001001101000100011;
assign LUT_4[50308] = 32'b00000000000000001110000010100011;
assign LUT_4[50309] = 32'b00000000000000000111001110011011;
assign LUT_4[50310] = 32'b00000000000000001101011101000111;
assign LUT_4[50311] = 32'b00000000000000000110101000111111;
assign LUT_4[50312] = 32'b00000000000000001010001110011100;
assign LUT_4[50313] = 32'b00000000000000000011011010010100;
assign LUT_4[50314] = 32'b00000000000000001001101001000000;
assign LUT_4[50315] = 32'b00000000000000000010110100111000;
assign LUT_4[50316] = 32'b00000000000000000111001110111000;
assign LUT_4[50317] = 32'b00000000000000000000011010110000;
assign LUT_4[50318] = 32'b00000000000000000110101001011100;
assign LUT_4[50319] = 32'b11111111111111111111110101010100;
assign LUT_4[50320] = 32'b00000000000000001110110011110101;
assign LUT_4[50321] = 32'b00000000000000000111111111101101;
assign LUT_4[50322] = 32'b00000000000000001110001110011001;
assign LUT_4[50323] = 32'b00000000000000000111011010010001;
assign LUT_4[50324] = 32'b00000000000000001011110100010001;
assign LUT_4[50325] = 32'b00000000000000000101000000001001;
assign LUT_4[50326] = 32'b00000000000000001011001110110101;
assign LUT_4[50327] = 32'b00000000000000000100011010101101;
assign LUT_4[50328] = 32'b00000000000000001000000000001010;
assign LUT_4[50329] = 32'b00000000000000000001001100000010;
assign LUT_4[50330] = 32'b00000000000000000111011010101110;
assign LUT_4[50331] = 32'b00000000000000000000100110100110;
assign LUT_4[50332] = 32'b00000000000000000101000000100110;
assign LUT_4[50333] = 32'b11111111111111111110001100011110;
assign LUT_4[50334] = 32'b00000000000000000100011011001010;
assign LUT_4[50335] = 32'b11111111111111111101100111000010;
assign LUT_4[50336] = 32'b00000000000000001111011101001110;
assign LUT_4[50337] = 32'b00000000000000001000101001000110;
assign LUT_4[50338] = 32'b00000000000000001110110111110010;
assign LUT_4[50339] = 32'b00000000000000001000000011101010;
assign LUT_4[50340] = 32'b00000000000000001100011101101010;
assign LUT_4[50341] = 32'b00000000000000000101101001100010;
assign LUT_4[50342] = 32'b00000000000000001011111000001110;
assign LUT_4[50343] = 32'b00000000000000000101000100000110;
assign LUT_4[50344] = 32'b00000000000000001000101001100011;
assign LUT_4[50345] = 32'b00000000000000000001110101011011;
assign LUT_4[50346] = 32'b00000000000000001000000100000111;
assign LUT_4[50347] = 32'b00000000000000000001001111111111;
assign LUT_4[50348] = 32'b00000000000000000101101001111111;
assign LUT_4[50349] = 32'b11111111111111111110110101110111;
assign LUT_4[50350] = 32'b00000000000000000101000100100011;
assign LUT_4[50351] = 32'b11111111111111111110010000011011;
assign LUT_4[50352] = 32'b00000000000000001101001110111100;
assign LUT_4[50353] = 32'b00000000000000000110011010110100;
assign LUT_4[50354] = 32'b00000000000000001100101001100000;
assign LUT_4[50355] = 32'b00000000000000000101110101011000;
assign LUT_4[50356] = 32'b00000000000000001010001111011000;
assign LUT_4[50357] = 32'b00000000000000000011011011010000;
assign LUT_4[50358] = 32'b00000000000000001001101001111100;
assign LUT_4[50359] = 32'b00000000000000000010110101110100;
assign LUT_4[50360] = 32'b00000000000000000110011011010001;
assign LUT_4[50361] = 32'b11111111111111111111100111001001;
assign LUT_4[50362] = 32'b00000000000000000101110101110101;
assign LUT_4[50363] = 32'b11111111111111111111000001101101;
assign LUT_4[50364] = 32'b00000000000000000011011011101101;
assign LUT_4[50365] = 32'b11111111111111111100100111100101;
assign LUT_4[50366] = 32'b00000000000000000010110110010001;
assign LUT_4[50367] = 32'b11111111111111111100000010001001;
assign LUT_4[50368] = 32'b00000000000000010010011001011011;
assign LUT_4[50369] = 32'b00000000000000001011100101010011;
assign LUT_4[50370] = 32'b00000000000000010001110011111111;
assign LUT_4[50371] = 32'b00000000000000001010111111110111;
assign LUT_4[50372] = 32'b00000000000000001111011001110111;
assign LUT_4[50373] = 32'b00000000000000001000100101101111;
assign LUT_4[50374] = 32'b00000000000000001110110100011011;
assign LUT_4[50375] = 32'b00000000000000001000000000010011;
assign LUT_4[50376] = 32'b00000000000000001011100101110000;
assign LUT_4[50377] = 32'b00000000000000000100110001101000;
assign LUT_4[50378] = 32'b00000000000000001011000000010100;
assign LUT_4[50379] = 32'b00000000000000000100001100001100;
assign LUT_4[50380] = 32'b00000000000000001000100110001100;
assign LUT_4[50381] = 32'b00000000000000000001110010000100;
assign LUT_4[50382] = 32'b00000000000000001000000000110000;
assign LUT_4[50383] = 32'b00000000000000000001001100101000;
assign LUT_4[50384] = 32'b00000000000000010000001011001001;
assign LUT_4[50385] = 32'b00000000000000001001010111000001;
assign LUT_4[50386] = 32'b00000000000000001111100101101101;
assign LUT_4[50387] = 32'b00000000000000001000110001100101;
assign LUT_4[50388] = 32'b00000000000000001101001011100101;
assign LUT_4[50389] = 32'b00000000000000000110010111011101;
assign LUT_4[50390] = 32'b00000000000000001100100110001001;
assign LUT_4[50391] = 32'b00000000000000000101110010000001;
assign LUT_4[50392] = 32'b00000000000000001001010111011110;
assign LUT_4[50393] = 32'b00000000000000000010100011010110;
assign LUT_4[50394] = 32'b00000000000000001000110010000010;
assign LUT_4[50395] = 32'b00000000000000000001111101111010;
assign LUT_4[50396] = 32'b00000000000000000110010111111010;
assign LUT_4[50397] = 32'b11111111111111111111100011110010;
assign LUT_4[50398] = 32'b00000000000000000101110010011110;
assign LUT_4[50399] = 32'b11111111111111111110111110010110;
assign LUT_4[50400] = 32'b00000000000000010000110100100010;
assign LUT_4[50401] = 32'b00000000000000001010000000011010;
assign LUT_4[50402] = 32'b00000000000000010000001111000110;
assign LUT_4[50403] = 32'b00000000000000001001011010111110;
assign LUT_4[50404] = 32'b00000000000000001101110100111110;
assign LUT_4[50405] = 32'b00000000000000000111000000110110;
assign LUT_4[50406] = 32'b00000000000000001101001111100010;
assign LUT_4[50407] = 32'b00000000000000000110011011011010;
assign LUT_4[50408] = 32'b00000000000000001010000000110111;
assign LUT_4[50409] = 32'b00000000000000000011001100101111;
assign LUT_4[50410] = 32'b00000000000000001001011011011011;
assign LUT_4[50411] = 32'b00000000000000000010100111010011;
assign LUT_4[50412] = 32'b00000000000000000111000001010011;
assign LUT_4[50413] = 32'b00000000000000000000001101001011;
assign LUT_4[50414] = 32'b00000000000000000110011011110111;
assign LUT_4[50415] = 32'b11111111111111111111100111101111;
assign LUT_4[50416] = 32'b00000000000000001110100110010000;
assign LUT_4[50417] = 32'b00000000000000000111110010001000;
assign LUT_4[50418] = 32'b00000000000000001110000000110100;
assign LUT_4[50419] = 32'b00000000000000000111001100101100;
assign LUT_4[50420] = 32'b00000000000000001011100110101100;
assign LUT_4[50421] = 32'b00000000000000000100110010100100;
assign LUT_4[50422] = 32'b00000000000000001011000001010000;
assign LUT_4[50423] = 32'b00000000000000000100001101001000;
assign LUT_4[50424] = 32'b00000000000000000111110010100101;
assign LUT_4[50425] = 32'b00000000000000000000111110011101;
assign LUT_4[50426] = 32'b00000000000000000111001101001001;
assign LUT_4[50427] = 32'b00000000000000000000011001000001;
assign LUT_4[50428] = 32'b00000000000000000100110011000001;
assign LUT_4[50429] = 32'b11111111111111111101111110111001;
assign LUT_4[50430] = 32'b00000000000000000100001101100101;
assign LUT_4[50431] = 32'b11111111111111111101011001011101;
assign LUT_4[50432] = 32'b00000000000000010011010111100010;
assign LUT_4[50433] = 32'b00000000000000001100100011011010;
assign LUT_4[50434] = 32'b00000000000000010010110010000110;
assign LUT_4[50435] = 32'b00000000000000001011111101111110;
assign LUT_4[50436] = 32'b00000000000000010000010111111110;
assign LUT_4[50437] = 32'b00000000000000001001100011110110;
assign LUT_4[50438] = 32'b00000000000000001111110010100010;
assign LUT_4[50439] = 32'b00000000000000001000111110011010;
assign LUT_4[50440] = 32'b00000000000000001100100011110111;
assign LUT_4[50441] = 32'b00000000000000000101101111101111;
assign LUT_4[50442] = 32'b00000000000000001011111110011011;
assign LUT_4[50443] = 32'b00000000000000000101001010010011;
assign LUT_4[50444] = 32'b00000000000000001001100100010011;
assign LUT_4[50445] = 32'b00000000000000000010110000001011;
assign LUT_4[50446] = 32'b00000000000000001000111110110111;
assign LUT_4[50447] = 32'b00000000000000000010001010101111;
assign LUT_4[50448] = 32'b00000000000000010001001001010000;
assign LUT_4[50449] = 32'b00000000000000001010010101001000;
assign LUT_4[50450] = 32'b00000000000000010000100011110100;
assign LUT_4[50451] = 32'b00000000000000001001101111101100;
assign LUT_4[50452] = 32'b00000000000000001110001001101100;
assign LUT_4[50453] = 32'b00000000000000000111010101100100;
assign LUT_4[50454] = 32'b00000000000000001101100100010000;
assign LUT_4[50455] = 32'b00000000000000000110110000001000;
assign LUT_4[50456] = 32'b00000000000000001010010101100101;
assign LUT_4[50457] = 32'b00000000000000000011100001011101;
assign LUT_4[50458] = 32'b00000000000000001001110000001001;
assign LUT_4[50459] = 32'b00000000000000000010111100000001;
assign LUT_4[50460] = 32'b00000000000000000111010110000001;
assign LUT_4[50461] = 32'b00000000000000000000100001111001;
assign LUT_4[50462] = 32'b00000000000000000110110000100101;
assign LUT_4[50463] = 32'b11111111111111111111111100011101;
assign LUT_4[50464] = 32'b00000000000000010001110010101001;
assign LUT_4[50465] = 32'b00000000000000001010111110100001;
assign LUT_4[50466] = 32'b00000000000000010001001101001101;
assign LUT_4[50467] = 32'b00000000000000001010011001000101;
assign LUT_4[50468] = 32'b00000000000000001110110011000101;
assign LUT_4[50469] = 32'b00000000000000000111111110111101;
assign LUT_4[50470] = 32'b00000000000000001110001101101001;
assign LUT_4[50471] = 32'b00000000000000000111011001100001;
assign LUT_4[50472] = 32'b00000000000000001010111110111110;
assign LUT_4[50473] = 32'b00000000000000000100001010110110;
assign LUT_4[50474] = 32'b00000000000000001010011001100010;
assign LUT_4[50475] = 32'b00000000000000000011100101011010;
assign LUT_4[50476] = 32'b00000000000000000111111111011010;
assign LUT_4[50477] = 32'b00000000000000000001001011010010;
assign LUT_4[50478] = 32'b00000000000000000111011001111110;
assign LUT_4[50479] = 32'b00000000000000000000100101110110;
assign LUT_4[50480] = 32'b00000000000000001111100100010111;
assign LUT_4[50481] = 32'b00000000000000001000110000001111;
assign LUT_4[50482] = 32'b00000000000000001110111110111011;
assign LUT_4[50483] = 32'b00000000000000001000001010110011;
assign LUT_4[50484] = 32'b00000000000000001100100100110011;
assign LUT_4[50485] = 32'b00000000000000000101110000101011;
assign LUT_4[50486] = 32'b00000000000000001011111111010111;
assign LUT_4[50487] = 32'b00000000000000000101001011001111;
assign LUT_4[50488] = 32'b00000000000000001000110000101100;
assign LUT_4[50489] = 32'b00000000000000000001111100100100;
assign LUT_4[50490] = 32'b00000000000000001000001011010000;
assign LUT_4[50491] = 32'b00000000000000000001010111001000;
assign LUT_4[50492] = 32'b00000000000000000101110001001000;
assign LUT_4[50493] = 32'b11111111111111111110111101000000;
assign LUT_4[50494] = 32'b00000000000000000101001011101100;
assign LUT_4[50495] = 32'b11111111111111111110010111100100;
assign LUT_4[50496] = 32'b00000000000000010100101110110110;
assign LUT_4[50497] = 32'b00000000000000001101111010101110;
assign LUT_4[50498] = 32'b00000000000000010100001001011010;
assign LUT_4[50499] = 32'b00000000000000001101010101010010;
assign LUT_4[50500] = 32'b00000000000000010001101111010010;
assign LUT_4[50501] = 32'b00000000000000001010111011001010;
assign LUT_4[50502] = 32'b00000000000000010001001001110110;
assign LUT_4[50503] = 32'b00000000000000001010010101101110;
assign LUT_4[50504] = 32'b00000000000000001101111011001011;
assign LUT_4[50505] = 32'b00000000000000000111000111000011;
assign LUT_4[50506] = 32'b00000000000000001101010101101111;
assign LUT_4[50507] = 32'b00000000000000000110100001100111;
assign LUT_4[50508] = 32'b00000000000000001010111011100111;
assign LUT_4[50509] = 32'b00000000000000000100000111011111;
assign LUT_4[50510] = 32'b00000000000000001010010110001011;
assign LUT_4[50511] = 32'b00000000000000000011100010000011;
assign LUT_4[50512] = 32'b00000000000000010010100000100100;
assign LUT_4[50513] = 32'b00000000000000001011101100011100;
assign LUT_4[50514] = 32'b00000000000000010001111011001000;
assign LUT_4[50515] = 32'b00000000000000001011000111000000;
assign LUT_4[50516] = 32'b00000000000000001111100001000000;
assign LUT_4[50517] = 32'b00000000000000001000101100111000;
assign LUT_4[50518] = 32'b00000000000000001110111011100100;
assign LUT_4[50519] = 32'b00000000000000001000000111011100;
assign LUT_4[50520] = 32'b00000000000000001011101100111001;
assign LUT_4[50521] = 32'b00000000000000000100111000110001;
assign LUT_4[50522] = 32'b00000000000000001011000111011101;
assign LUT_4[50523] = 32'b00000000000000000100010011010101;
assign LUT_4[50524] = 32'b00000000000000001000101101010101;
assign LUT_4[50525] = 32'b00000000000000000001111001001101;
assign LUT_4[50526] = 32'b00000000000000001000000111111001;
assign LUT_4[50527] = 32'b00000000000000000001010011110001;
assign LUT_4[50528] = 32'b00000000000000010011001001111101;
assign LUT_4[50529] = 32'b00000000000000001100010101110101;
assign LUT_4[50530] = 32'b00000000000000010010100100100001;
assign LUT_4[50531] = 32'b00000000000000001011110000011001;
assign LUT_4[50532] = 32'b00000000000000010000001010011001;
assign LUT_4[50533] = 32'b00000000000000001001010110010001;
assign LUT_4[50534] = 32'b00000000000000001111100100111101;
assign LUT_4[50535] = 32'b00000000000000001000110000110101;
assign LUT_4[50536] = 32'b00000000000000001100010110010010;
assign LUT_4[50537] = 32'b00000000000000000101100010001010;
assign LUT_4[50538] = 32'b00000000000000001011110000110110;
assign LUT_4[50539] = 32'b00000000000000000100111100101110;
assign LUT_4[50540] = 32'b00000000000000001001010110101110;
assign LUT_4[50541] = 32'b00000000000000000010100010100110;
assign LUT_4[50542] = 32'b00000000000000001000110001010010;
assign LUT_4[50543] = 32'b00000000000000000001111101001010;
assign LUT_4[50544] = 32'b00000000000000010000111011101011;
assign LUT_4[50545] = 32'b00000000000000001010000111100011;
assign LUT_4[50546] = 32'b00000000000000010000010110001111;
assign LUT_4[50547] = 32'b00000000000000001001100010000111;
assign LUT_4[50548] = 32'b00000000000000001101111100000111;
assign LUT_4[50549] = 32'b00000000000000000111000111111111;
assign LUT_4[50550] = 32'b00000000000000001101010110101011;
assign LUT_4[50551] = 32'b00000000000000000110100010100011;
assign LUT_4[50552] = 32'b00000000000000001010001000000000;
assign LUT_4[50553] = 32'b00000000000000000011010011111000;
assign LUT_4[50554] = 32'b00000000000000001001100010100100;
assign LUT_4[50555] = 32'b00000000000000000010101110011100;
assign LUT_4[50556] = 32'b00000000000000000111001000011100;
assign LUT_4[50557] = 32'b00000000000000000000010100010100;
assign LUT_4[50558] = 32'b00000000000000000110100011000000;
assign LUT_4[50559] = 32'b11111111111111111111101110111000;
assign LUT_4[50560] = 32'b00000000000000010101111101101010;
assign LUT_4[50561] = 32'b00000000000000001111001001100010;
assign LUT_4[50562] = 32'b00000000000000010101011000001110;
assign LUT_4[50563] = 32'b00000000000000001110100100000110;
assign LUT_4[50564] = 32'b00000000000000010010111110000110;
assign LUT_4[50565] = 32'b00000000000000001100001001111110;
assign LUT_4[50566] = 32'b00000000000000010010011000101010;
assign LUT_4[50567] = 32'b00000000000000001011100100100010;
assign LUT_4[50568] = 32'b00000000000000001111001001111111;
assign LUT_4[50569] = 32'b00000000000000001000010101110111;
assign LUT_4[50570] = 32'b00000000000000001110100100100011;
assign LUT_4[50571] = 32'b00000000000000000111110000011011;
assign LUT_4[50572] = 32'b00000000000000001100001010011011;
assign LUT_4[50573] = 32'b00000000000000000101010110010011;
assign LUT_4[50574] = 32'b00000000000000001011100100111111;
assign LUT_4[50575] = 32'b00000000000000000100110000110111;
assign LUT_4[50576] = 32'b00000000000000010011101111011000;
assign LUT_4[50577] = 32'b00000000000000001100111011010000;
assign LUT_4[50578] = 32'b00000000000000010011001001111100;
assign LUT_4[50579] = 32'b00000000000000001100010101110100;
assign LUT_4[50580] = 32'b00000000000000010000101111110100;
assign LUT_4[50581] = 32'b00000000000000001001111011101100;
assign LUT_4[50582] = 32'b00000000000000010000001010011000;
assign LUT_4[50583] = 32'b00000000000000001001010110010000;
assign LUT_4[50584] = 32'b00000000000000001100111011101101;
assign LUT_4[50585] = 32'b00000000000000000110000111100101;
assign LUT_4[50586] = 32'b00000000000000001100010110010001;
assign LUT_4[50587] = 32'b00000000000000000101100010001001;
assign LUT_4[50588] = 32'b00000000000000001001111100001001;
assign LUT_4[50589] = 32'b00000000000000000011001000000001;
assign LUT_4[50590] = 32'b00000000000000001001010110101101;
assign LUT_4[50591] = 32'b00000000000000000010100010100101;
assign LUT_4[50592] = 32'b00000000000000010100011000110001;
assign LUT_4[50593] = 32'b00000000000000001101100100101001;
assign LUT_4[50594] = 32'b00000000000000010011110011010101;
assign LUT_4[50595] = 32'b00000000000000001100111111001101;
assign LUT_4[50596] = 32'b00000000000000010001011001001101;
assign LUT_4[50597] = 32'b00000000000000001010100101000101;
assign LUT_4[50598] = 32'b00000000000000010000110011110001;
assign LUT_4[50599] = 32'b00000000000000001001111111101001;
assign LUT_4[50600] = 32'b00000000000000001101100101000110;
assign LUT_4[50601] = 32'b00000000000000000110110000111110;
assign LUT_4[50602] = 32'b00000000000000001100111111101010;
assign LUT_4[50603] = 32'b00000000000000000110001011100010;
assign LUT_4[50604] = 32'b00000000000000001010100101100010;
assign LUT_4[50605] = 32'b00000000000000000011110001011010;
assign LUT_4[50606] = 32'b00000000000000001010000000000110;
assign LUT_4[50607] = 32'b00000000000000000011001011111110;
assign LUT_4[50608] = 32'b00000000000000010010001010011111;
assign LUT_4[50609] = 32'b00000000000000001011010110010111;
assign LUT_4[50610] = 32'b00000000000000010001100101000011;
assign LUT_4[50611] = 32'b00000000000000001010110000111011;
assign LUT_4[50612] = 32'b00000000000000001111001010111011;
assign LUT_4[50613] = 32'b00000000000000001000010110110011;
assign LUT_4[50614] = 32'b00000000000000001110100101011111;
assign LUT_4[50615] = 32'b00000000000000000111110001010111;
assign LUT_4[50616] = 32'b00000000000000001011010110110100;
assign LUT_4[50617] = 32'b00000000000000000100100010101100;
assign LUT_4[50618] = 32'b00000000000000001010110001011000;
assign LUT_4[50619] = 32'b00000000000000000011111101010000;
assign LUT_4[50620] = 32'b00000000000000001000010111010000;
assign LUT_4[50621] = 32'b00000000000000000001100011001000;
assign LUT_4[50622] = 32'b00000000000000000111110001110100;
assign LUT_4[50623] = 32'b00000000000000000000111101101100;
assign LUT_4[50624] = 32'b00000000000000010111010100111110;
assign LUT_4[50625] = 32'b00000000000000010000100000110110;
assign LUT_4[50626] = 32'b00000000000000010110101111100010;
assign LUT_4[50627] = 32'b00000000000000001111111011011010;
assign LUT_4[50628] = 32'b00000000000000010100010101011010;
assign LUT_4[50629] = 32'b00000000000000001101100001010010;
assign LUT_4[50630] = 32'b00000000000000010011101111111110;
assign LUT_4[50631] = 32'b00000000000000001100111011110110;
assign LUT_4[50632] = 32'b00000000000000010000100001010011;
assign LUT_4[50633] = 32'b00000000000000001001101101001011;
assign LUT_4[50634] = 32'b00000000000000001111111011110111;
assign LUT_4[50635] = 32'b00000000000000001001000111101111;
assign LUT_4[50636] = 32'b00000000000000001101100001101111;
assign LUT_4[50637] = 32'b00000000000000000110101101100111;
assign LUT_4[50638] = 32'b00000000000000001100111100010011;
assign LUT_4[50639] = 32'b00000000000000000110001000001011;
assign LUT_4[50640] = 32'b00000000000000010101000110101100;
assign LUT_4[50641] = 32'b00000000000000001110010010100100;
assign LUT_4[50642] = 32'b00000000000000010100100001010000;
assign LUT_4[50643] = 32'b00000000000000001101101101001000;
assign LUT_4[50644] = 32'b00000000000000010010000111001000;
assign LUT_4[50645] = 32'b00000000000000001011010011000000;
assign LUT_4[50646] = 32'b00000000000000010001100001101100;
assign LUT_4[50647] = 32'b00000000000000001010101101100100;
assign LUT_4[50648] = 32'b00000000000000001110010011000001;
assign LUT_4[50649] = 32'b00000000000000000111011110111001;
assign LUT_4[50650] = 32'b00000000000000001101101101100101;
assign LUT_4[50651] = 32'b00000000000000000110111001011101;
assign LUT_4[50652] = 32'b00000000000000001011010011011101;
assign LUT_4[50653] = 32'b00000000000000000100011111010101;
assign LUT_4[50654] = 32'b00000000000000001010101110000001;
assign LUT_4[50655] = 32'b00000000000000000011111001111001;
assign LUT_4[50656] = 32'b00000000000000010101110000000101;
assign LUT_4[50657] = 32'b00000000000000001110111011111101;
assign LUT_4[50658] = 32'b00000000000000010101001010101001;
assign LUT_4[50659] = 32'b00000000000000001110010110100001;
assign LUT_4[50660] = 32'b00000000000000010010110000100001;
assign LUT_4[50661] = 32'b00000000000000001011111100011001;
assign LUT_4[50662] = 32'b00000000000000010010001011000101;
assign LUT_4[50663] = 32'b00000000000000001011010110111101;
assign LUT_4[50664] = 32'b00000000000000001110111100011010;
assign LUT_4[50665] = 32'b00000000000000001000001000010010;
assign LUT_4[50666] = 32'b00000000000000001110010110111110;
assign LUT_4[50667] = 32'b00000000000000000111100010110110;
assign LUT_4[50668] = 32'b00000000000000001011111100110110;
assign LUT_4[50669] = 32'b00000000000000000101001000101110;
assign LUT_4[50670] = 32'b00000000000000001011010111011010;
assign LUT_4[50671] = 32'b00000000000000000100100011010010;
assign LUT_4[50672] = 32'b00000000000000010011100001110011;
assign LUT_4[50673] = 32'b00000000000000001100101101101011;
assign LUT_4[50674] = 32'b00000000000000010010111100010111;
assign LUT_4[50675] = 32'b00000000000000001100001000001111;
assign LUT_4[50676] = 32'b00000000000000010000100010001111;
assign LUT_4[50677] = 32'b00000000000000001001101110000111;
assign LUT_4[50678] = 32'b00000000000000001111111100110011;
assign LUT_4[50679] = 32'b00000000000000001001001000101011;
assign LUT_4[50680] = 32'b00000000000000001100101110001000;
assign LUT_4[50681] = 32'b00000000000000000101111010000000;
assign LUT_4[50682] = 32'b00000000000000001100001000101100;
assign LUT_4[50683] = 32'b00000000000000000101010100100100;
assign LUT_4[50684] = 32'b00000000000000001001101110100100;
assign LUT_4[50685] = 32'b00000000000000000010111010011100;
assign LUT_4[50686] = 32'b00000000000000001001001001001000;
assign LUT_4[50687] = 32'b00000000000000000010010101000000;
assign LUT_4[50688] = 32'b00000000000000001101100000000111;
assign LUT_4[50689] = 32'b00000000000000000110101011111111;
assign LUT_4[50690] = 32'b00000000000000001100111010101011;
assign LUT_4[50691] = 32'b00000000000000000110000110100011;
assign LUT_4[50692] = 32'b00000000000000001010100000100011;
assign LUT_4[50693] = 32'b00000000000000000011101100011011;
assign LUT_4[50694] = 32'b00000000000000001001111011000111;
assign LUT_4[50695] = 32'b00000000000000000011000110111111;
assign LUT_4[50696] = 32'b00000000000000000110101100011100;
assign LUT_4[50697] = 32'b11111111111111111111111000010100;
assign LUT_4[50698] = 32'b00000000000000000110000111000000;
assign LUT_4[50699] = 32'b11111111111111111111010010111000;
assign LUT_4[50700] = 32'b00000000000000000011101100111000;
assign LUT_4[50701] = 32'b11111111111111111100111000110000;
assign LUT_4[50702] = 32'b00000000000000000011000111011100;
assign LUT_4[50703] = 32'b11111111111111111100010011010100;
assign LUT_4[50704] = 32'b00000000000000001011010001110101;
assign LUT_4[50705] = 32'b00000000000000000100011101101101;
assign LUT_4[50706] = 32'b00000000000000001010101100011001;
assign LUT_4[50707] = 32'b00000000000000000011111000010001;
assign LUT_4[50708] = 32'b00000000000000001000010010010001;
assign LUT_4[50709] = 32'b00000000000000000001011110001001;
assign LUT_4[50710] = 32'b00000000000000000111101100110101;
assign LUT_4[50711] = 32'b00000000000000000000111000101101;
assign LUT_4[50712] = 32'b00000000000000000100011110001010;
assign LUT_4[50713] = 32'b11111111111111111101101010000010;
assign LUT_4[50714] = 32'b00000000000000000011111000101110;
assign LUT_4[50715] = 32'b11111111111111111101000100100110;
assign LUT_4[50716] = 32'b00000000000000000001011110100110;
assign LUT_4[50717] = 32'b11111111111111111010101010011110;
assign LUT_4[50718] = 32'b00000000000000000000111001001010;
assign LUT_4[50719] = 32'b11111111111111111010000101000010;
assign LUT_4[50720] = 32'b00000000000000001011111011001110;
assign LUT_4[50721] = 32'b00000000000000000101000111000110;
assign LUT_4[50722] = 32'b00000000000000001011010101110010;
assign LUT_4[50723] = 32'b00000000000000000100100001101010;
assign LUT_4[50724] = 32'b00000000000000001000111011101010;
assign LUT_4[50725] = 32'b00000000000000000010000111100010;
assign LUT_4[50726] = 32'b00000000000000001000010110001110;
assign LUT_4[50727] = 32'b00000000000000000001100010000110;
assign LUT_4[50728] = 32'b00000000000000000101000111100011;
assign LUT_4[50729] = 32'b11111111111111111110010011011011;
assign LUT_4[50730] = 32'b00000000000000000100100010000111;
assign LUT_4[50731] = 32'b11111111111111111101101101111111;
assign LUT_4[50732] = 32'b00000000000000000010000111111111;
assign LUT_4[50733] = 32'b11111111111111111011010011110111;
assign LUT_4[50734] = 32'b00000000000000000001100010100011;
assign LUT_4[50735] = 32'b11111111111111111010101110011011;
assign LUT_4[50736] = 32'b00000000000000001001101100111100;
assign LUT_4[50737] = 32'b00000000000000000010111000110100;
assign LUT_4[50738] = 32'b00000000000000001001000111100000;
assign LUT_4[50739] = 32'b00000000000000000010010011011000;
assign LUT_4[50740] = 32'b00000000000000000110101101011000;
assign LUT_4[50741] = 32'b11111111111111111111111001010000;
assign LUT_4[50742] = 32'b00000000000000000110000111111100;
assign LUT_4[50743] = 32'b11111111111111111111010011110100;
assign LUT_4[50744] = 32'b00000000000000000010111001010001;
assign LUT_4[50745] = 32'b11111111111111111100000101001001;
assign LUT_4[50746] = 32'b00000000000000000010010011110101;
assign LUT_4[50747] = 32'b11111111111111111011011111101101;
assign LUT_4[50748] = 32'b11111111111111111111111001101101;
assign LUT_4[50749] = 32'b11111111111111111001000101100101;
assign LUT_4[50750] = 32'b11111111111111111111010100010001;
assign LUT_4[50751] = 32'b11111111111111111000100000001001;
assign LUT_4[50752] = 32'b00000000000000001110110111011011;
assign LUT_4[50753] = 32'b00000000000000001000000011010011;
assign LUT_4[50754] = 32'b00000000000000001110010001111111;
assign LUT_4[50755] = 32'b00000000000000000111011101110111;
assign LUT_4[50756] = 32'b00000000000000001011110111110111;
assign LUT_4[50757] = 32'b00000000000000000101000011101111;
assign LUT_4[50758] = 32'b00000000000000001011010010011011;
assign LUT_4[50759] = 32'b00000000000000000100011110010011;
assign LUT_4[50760] = 32'b00000000000000001000000011110000;
assign LUT_4[50761] = 32'b00000000000000000001001111101000;
assign LUT_4[50762] = 32'b00000000000000000111011110010100;
assign LUT_4[50763] = 32'b00000000000000000000101010001100;
assign LUT_4[50764] = 32'b00000000000000000101000100001100;
assign LUT_4[50765] = 32'b11111111111111111110010000000100;
assign LUT_4[50766] = 32'b00000000000000000100011110110000;
assign LUT_4[50767] = 32'b11111111111111111101101010101000;
assign LUT_4[50768] = 32'b00000000000000001100101001001001;
assign LUT_4[50769] = 32'b00000000000000000101110101000001;
assign LUT_4[50770] = 32'b00000000000000001100000011101101;
assign LUT_4[50771] = 32'b00000000000000000101001111100101;
assign LUT_4[50772] = 32'b00000000000000001001101001100101;
assign LUT_4[50773] = 32'b00000000000000000010110101011101;
assign LUT_4[50774] = 32'b00000000000000001001000100001001;
assign LUT_4[50775] = 32'b00000000000000000010010000000001;
assign LUT_4[50776] = 32'b00000000000000000101110101011110;
assign LUT_4[50777] = 32'b11111111111111111111000001010110;
assign LUT_4[50778] = 32'b00000000000000000101010000000010;
assign LUT_4[50779] = 32'b11111111111111111110011011111010;
assign LUT_4[50780] = 32'b00000000000000000010110101111010;
assign LUT_4[50781] = 32'b11111111111111111100000001110010;
assign LUT_4[50782] = 32'b00000000000000000010010000011110;
assign LUT_4[50783] = 32'b11111111111111111011011100010110;
assign LUT_4[50784] = 32'b00000000000000001101010010100010;
assign LUT_4[50785] = 32'b00000000000000000110011110011010;
assign LUT_4[50786] = 32'b00000000000000001100101101000110;
assign LUT_4[50787] = 32'b00000000000000000101111000111110;
assign LUT_4[50788] = 32'b00000000000000001010010010111110;
assign LUT_4[50789] = 32'b00000000000000000011011110110110;
assign LUT_4[50790] = 32'b00000000000000001001101101100010;
assign LUT_4[50791] = 32'b00000000000000000010111001011010;
assign LUT_4[50792] = 32'b00000000000000000110011110110111;
assign LUT_4[50793] = 32'b11111111111111111111101010101111;
assign LUT_4[50794] = 32'b00000000000000000101111001011011;
assign LUT_4[50795] = 32'b11111111111111111111000101010011;
assign LUT_4[50796] = 32'b00000000000000000011011111010011;
assign LUT_4[50797] = 32'b11111111111111111100101011001011;
assign LUT_4[50798] = 32'b00000000000000000010111001110111;
assign LUT_4[50799] = 32'b11111111111111111100000101101111;
assign LUT_4[50800] = 32'b00000000000000001011000100010000;
assign LUT_4[50801] = 32'b00000000000000000100010000001000;
assign LUT_4[50802] = 32'b00000000000000001010011110110100;
assign LUT_4[50803] = 32'b00000000000000000011101010101100;
assign LUT_4[50804] = 32'b00000000000000001000000100101100;
assign LUT_4[50805] = 32'b00000000000000000001010000100100;
assign LUT_4[50806] = 32'b00000000000000000111011111010000;
assign LUT_4[50807] = 32'b00000000000000000000101011001000;
assign LUT_4[50808] = 32'b00000000000000000100010000100101;
assign LUT_4[50809] = 32'b11111111111111111101011100011101;
assign LUT_4[50810] = 32'b00000000000000000011101011001001;
assign LUT_4[50811] = 32'b11111111111111111100110111000001;
assign LUT_4[50812] = 32'b00000000000000000001010001000001;
assign LUT_4[50813] = 32'b11111111111111111010011100111001;
assign LUT_4[50814] = 32'b00000000000000000000101011100101;
assign LUT_4[50815] = 32'b11111111111111111001110111011101;
assign LUT_4[50816] = 32'b00000000000000010000000110001111;
assign LUT_4[50817] = 32'b00000000000000001001010010000111;
assign LUT_4[50818] = 32'b00000000000000001111100000110011;
assign LUT_4[50819] = 32'b00000000000000001000101100101011;
assign LUT_4[50820] = 32'b00000000000000001101000110101011;
assign LUT_4[50821] = 32'b00000000000000000110010010100011;
assign LUT_4[50822] = 32'b00000000000000001100100001001111;
assign LUT_4[50823] = 32'b00000000000000000101101101000111;
assign LUT_4[50824] = 32'b00000000000000001001010010100100;
assign LUT_4[50825] = 32'b00000000000000000010011110011100;
assign LUT_4[50826] = 32'b00000000000000001000101101001000;
assign LUT_4[50827] = 32'b00000000000000000001111001000000;
assign LUT_4[50828] = 32'b00000000000000000110010011000000;
assign LUT_4[50829] = 32'b11111111111111111111011110111000;
assign LUT_4[50830] = 32'b00000000000000000101101101100100;
assign LUT_4[50831] = 32'b11111111111111111110111001011100;
assign LUT_4[50832] = 32'b00000000000000001101110111111101;
assign LUT_4[50833] = 32'b00000000000000000111000011110101;
assign LUT_4[50834] = 32'b00000000000000001101010010100001;
assign LUT_4[50835] = 32'b00000000000000000110011110011001;
assign LUT_4[50836] = 32'b00000000000000001010111000011001;
assign LUT_4[50837] = 32'b00000000000000000100000100010001;
assign LUT_4[50838] = 32'b00000000000000001010010010111101;
assign LUT_4[50839] = 32'b00000000000000000011011110110101;
assign LUT_4[50840] = 32'b00000000000000000111000100010010;
assign LUT_4[50841] = 32'b00000000000000000000010000001010;
assign LUT_4[50842] = 32'b00000000000000000110011110110110;
assign LUT_4[50843] = 32'b11111111111111111111101010101110;
assign LUT_4[50844] = 32'b00000000000000000100000100101110;
assign LUT_4[50845] = 32'b11111111111111111101010000100110;
assign LUT_4[50846] = 32'b00000000000000000011011111010010;
assign LUT_4[50847] = 32'b11111111111111111100101011001010;
assign LUT_4[50848] = 32'b00000000000000001110100001010110;
assign LUT_4[50849] = 32'b00000000000000000111101101001110;
assign LUT_4[50850] = 32'b00000000000000001101111011111010;
assign LUT_4[50851] = 32'b00000000000000000111000111110010;
assign LUT_4[50852] = 32'b00000000000000001011100001110010;
assign LUT_4[50853] = 32'b00000000000000000100101101101010;
assign LUT_4[50854] = 32'b00000000000000001010111100010110;
assign LUT_4[50855] = 32'b00000000000000000100001000001110;
assign LUT_4[50856] = 32'b00000000000000000111101101101011;
assign LUT_4[50857] = 32'b00000000000000000000111001100011;
assign LUT_4[50858] = 32'b00000000000000000111001000001111;
assign LUT_4[50859] = 32'b00000000000000000000010100000111;
assign LUT_4[50860] = 32'b00000000000000000100101110000111;
assign LUT_4[50861] = 32'b11111111111111111101111001111111;
assign LUT_4[50862] = 32'b00000000000000000100001000101011;
assign LUT_4[50863] = 32'b11111111111111111101010100100011;
assign LUT_4[50864] = 32'b00000000000000001100010011000100;
assign LUT_4[50865] = 32'b00000000000000000101011110111100;
assign LUT_4[50866] = 32'b00000000000000001011101101101000;
assign LUT_4[50867] = 32'b00000000000000000100111001100000;
assign LUT_4[50868] = 32'b00000000000000001001010011100000;
assign LUT_4[50869] = 32'b00000000000000000010011111011000;
assign LUT_4[50870] = 32'b00000000000000001000101110000100;
assign LUT_4[50871] = 32'b00000000000000000001111001111100;
assign LUT_4[50872] = 32'b00000000000000000101011111011001;
assign LUT_4[50873] = 32'b11111111111111111110101011010001;
assign LUT_4[50874] = 32'b00000000000000000100111001111101;
assign LUT_4[50875] = 32'b11111111111111111110000101110101;
assign LUT_4[50876] = 32'b00000000000000000010011111110101;
assign LUT_4[50877] = 32'b11111111111111111011101011101101;
assign LUT_4[50878] = 32'b00000000000000000001111010011001;
assign LUT_4[50879] = 32'b11111111111111111011000110010001;
assign LUT_4[50880] = 32'b00000000000000010001011101100011;
assign LUT_4[50881] = 32'b00000000000000001010101001011011;
assign LUT_4[50882] = 32'b00000000000000010000111000000111;
assign LUT_4[50883] = 32'b00000000000000001010000011111111;
assign LUT_4[50884] = 32'b00000000000000001110011101111111;
assign LUT_4[50885] = 32'b00000000000000000111101001110111;
assign LUT_4[50886] = 32'b00000000000000001101111000100011;
assign LUT_4[50887] = 32'b00000000000000000111000100011011;
assign LUT_4[50888] = 32'b00000000000000001010101001111000;
assign LUT_4[50889] = 32'b00000000000000000011110101110000;
assign LUT_4[50890] = 32'b00000000000000001010000100011100;
assign LUT_4[50891] = 32'b00000000000000000011010000010100;
assign LUT_4[50892] = 32'b00000000000000000111101010010100;
assign LUT_4[50893] = 32'b00000000000000000000110110001100;
assign LUT_4[50894] = 32'b00000000000000000111000100111000;
assign LUT_4[50895] = 32'b00000000000000000000010000110000;
assign LUT_4[50896] = 32'b00000000000000001111001111010001;
assign LUT_4[50897] = 32'b00000000000000001000011011001001;
assign LUT_4[50898] = 32'b00000000000000001110101001110101;
assign LUT_4[50899] = 32'b00000000000000000111110101101101;
assign LUT_4[50900] = 32'b00000000000000001100001111101101;
assign LUT_4[50901] = 32'b00000000000000000101011011100101;
assign LUT_4[50902] = 32'b00000000000000001011101010010001;
assign LUT_4[50903] = 32'b00000000000000000100110110001001;
assign LUT_4[50904] = 32'b00000000000000001000011011100110;
assign LUT_4[50905] = 32'b00000000000000000001100111011110;
assign LUT_4[50906] = 32'b00000000000000000111110110001010;
assign LUT_4[50907] = 32'b00000000000000000001000010000010;
assign LUT_4[50908] = 32'b00000000000000000101011100000010;
assign LUT_4[50909] = 32'b11111111111111111110100111111010;
assign LUT_4[50910] = 32'b00000000000000000100110110100110;
assign LUT_4[50911] = 32'b11111111111111111110000010011110;
assign LUT_4[50912] = 32'b00000000000000001111111000101010;
assign LUT_4[50913] = 32'b00000000000000001001000100100010;
assign LUT_4[50914] = 32'b00000000000000001111010011001110;
assign LUT_4[50915] = 32'b00000000000000001000011111000110;
assign LUT_4[50916] = 32'b00000000000000001100111001000110;
assign LUT_4[50917] = 32'b00000000000000000110000100111110;
assign LUT_4[50918] = 32'b00000000000000001100010011101010;
assign LUT_4[50919] = 32'b00000000000000000101011111100010;
assign LUT_4[50920] = 32'b00000000000000001001000100111111;
assign LUT_4[50921] = 32'b00000000000000000010010000110111;
assign LUT_4[50922] = 32'b00000000000000001000011111100011;
assign LUT_4[50923] = 32'b00000000000000000001101011011011;
assign LUT_4[50924] = 32'b00000000000000000110000101011011;
assign LUT_4[50925] = 32'b11111111111111111111010001010011;
assign LUT_4[50926] = 32'b00000000000000000101011111111111;
assign LUT_4[50927] = 32'b11111111111111111110101011110111;
assign LUT_4[50928] = 32'b00000000000000001101101010011000;
assign LUT_4[50929] = 32'b00000000000000000110110110010000;
assign LUT_4[50930] = 32'b00000000000000001101000100111100;
assign LUT_4[50931] = 32'b00000000000000000110010000110100;
assign LUT_4[50932] = 32'b00000000000000001010101010110100;
assign LUT_4[50933] = 32'b00000000000000000011110110101100;
assign LUT_4[50934] = 32'b00000000000000001010000101011000;
assign LUT_4[50935] = 32'b00000000000000000011010001010000;
assign LUT_4[50936] = 32'b00000000000000000110110110101101;
assign LUT_4[50937] = 32'b00000000000000000000000010100101;
assign LUT_4[50938] = 32'b00000000000000000110010001010001;
assign LUT_4[50939] = 32'b11111111111111111111011101001001;
assign LUT_4[50940] = 32'b00000000000000000011110111001001;
assign LUT_4[50941] = 32'b11111111111111111101000011000001;
assign LUT_4[50942] = 32'b00000000000000000011010001101101;
assign LUT_4[50943] = 32'b11111111111111111100011101100101;
assign LUT_4[50944] = 32'b00000000000000010010011011101010;
assign LUT_4[50945] = 32'b00000000000000001011100111100010;
assign LUT_4[50946] = 32'b00000000000000010001110110001110;
assign LUT_4[50947] = 32'b00000000000000001011000010000110;
assign LUT_4[50948] = 32'b00000000000000001111011100000110;
assign LUT_4[50949] = 32'b00000000000000001000100111111110;
assign LUT_4[50950] = 32'b00000000000000001110110110101010;
assign LUT_4[50951] = 32'b00000000000000001000000010100010;
assign LUT_4[50952] = 32'b00000000000000001011100111111111;
assign LUT_4[50953] = 32'b00000000000000000100110011110111;
assign LUT_4[50954] = 32'b00000000000000001011000010100011;
assign LUT_4[50955] = 32'b00000000000000000100001110011011;
assign LUT_4[50956] = 32'b00000000000000001000101000011011;
assign LUT_4[50957] = 32'b00000000000000000001110100010011;
assign LUT_4[50958] = 32'b00000000000000001000000010111111;
assign LUT_4[50959] = 32'b00000000000000000001001110110111;
assign LUT_4[50960] = 32'b00000000000000010000001101011000;
assign LUT_4[50961] = 32'b00000000000000001001011001010000;
assign LUT_4[50962] = 32'b00000000000000001111100111111100;
assign LUT_4[50963] = 32'b00000000000000001000110011110100;
assign LUT_4[50964] = 32'b00000000000000001101001101110100;
assign LUT_4[50965] = 32'b00000000000000000110011001101100;
assign LUT_4[50966] = 32'b00000000000000001100101000011000;
assign LUT_4[50967] = 32'b00000000000000000101110100010000;
assign LUT_4[50968] = 32'b00000000000000001001011001101101;
assign LUT_4[50969] = 32'b00000000000000000010100101100101;
assign LUT_4[50970] = 32'b00000000000000001000110100010001;
assign LUT_4[50971] = 32'b00000000000000000010000000001001;
assign LUT_4[50972] = 32'b00000000000000000110011010001001;
assign LUT_4[50973] = 32'b11111111111111111111100110000001;
assign LUT_4[50974] = 32'b00000000000000000101110100101101;
assign LUT_4[50975] = 32'b11111111111111111111000000100101;
assign LUT_4[50976] = 32'b00000000000000010000110110110001;
assign LUT_4[50977] = 32'b00000000000000001010000010101001;
assign LUT_4[50978] = 32'b00000000000000010000010001010101;
assign LUT_4[50979] = 32'b00000000000000001001011101001101;
assign LUT_4[50980] = 32'b00000000000000001101110111001101;
assign LUT_4[50981] = 32'b00000000000000000111000011000101;
assign LUT_4[50982] = 32'b00000000000000001101010001110001;
assign LUT_4[50983] = 32'b00000000000000000110011101101001;
assign LUT_4[50984] = 32'b00000000000000001010000011000110;
assign LUT_4[50985] = 32'b00000000000000000011001110111110;
assign LUT_4[50986] = 32'b00000000000000001001011101101010;
assign LUT_4[50987] = 32'b00000000000000000010101001100010;
assign LUT_4[50988] = 32'b00000000000000000111000011100010;
assign LUT_4[50989] = 32'b00000000000000000000001111011010;
assign LUT_4[50990] = 32'b00000000000000000110011110000110;
assign LUT_4[50991] = 32'b11111111111111111111101001111110;
assign LUT_4[50992] = 32'b00000000000000001110101000011111;
assign LUT_4[50993] = 32'b00000000000000000111110100010111;
assign LUT_4[50994] = 32'b00000000000000001110000011000011;
assign LUT_4[50995] = 32'b00000000000000000111001110111011;
assign LUT_4[50996] = 32'b00000000000000001011101000111011;
assign LUT_4[50997] = 32'b00000000000000000100110100110011;
assign LUT_4[50998] = 32'b00000000000000001011000011011111;
assign LUT_4[50999] = 32'b00000000000000000100001111010111;
assign LUT_4[51000] = 32'b00000000000000000111110100110100;
assign LUT_4[51001] = 32'b00000000000000000001000000101100;
assign LUT_4[51002] = 32'b00000000000000000111001111011000;
assign LUT_4[51003] = 32'b00000000000000000000011011010000;
assign LUT_4[51004] = 32'b00000000000000000100110101010000;
assign LUT_4[51005] = 32'b11111111111111111110000001001000;
assign LUT_4[51006] = 32'b00000000000000000100001111110100;
assign LUT_4[51007] = 32'b11111111111111111101011011101100;
assign LUT_4[51008] = 32'b00000000000000010011110010111110;
assign LUT_4[51009] = 32'b00000000000000001100111110110110;
assign LUT_4[51010] = 32'b00000000000000010011001101100010;
assign LUT_4[51011] = 32'b00000000000000001100011001011010;
assign LUT_4[51012] = 32'b00000000000000010000110011011010;
assign LUT_4[51013] = 32'b00000000000000001001111111010010;
assign LUT_4[51014] = 32'b00000000000000010000001101111110;
assign LUT_4[51015] = 32'b00000000000000001001011001110110;
assign LUT_4[51016] = 32'b00000000000000001100111111010011;
assign LUT_4[51017] = 32'b00000000000000000110001011001011;
assign LUT_4[51018] = 32'b00000000000000001100011001110111;
assign LUT_4[51019] = 32'b00000000000000000101100101101111;
assign LUT_4[51020] = 32'b00000000000000001001111111101111;
assign LUT_4[51021] = 32'b00000000000000000011001011100111;
assign LUT_4[51022] = 32'b00000000000000001001011010010011;
assign LUT_4[51023] = 32'b00000000000000000010100110001011;
assign LUT_4[51024] = 32'b00000000000000010001100100101100;
assign LUT_4[51025] = 32'b00000000000000001010110000100100;
assign LUT_4[51026] = 32'b00000000000000010000111111010000;
assign LUT_4[51027] = 32'b00000000000000001010001011001000;
assign LUT_4[51028] = 32'b00000000000000001110100101001000;
assign LUT_4[51029] = 32'b00000000000000000111110001000000;
assign LUT_4[51030] = 32'b00000000000000001101111111101100;
assign LUT_4[51031] = 32'b00000000000000000111001011100100;
assign LUT_4[51032] = 32'b00000000000000001010110001000001;
assign LUT_4[51033] = 32'b00000000000000000011111100111001;
assign LUT_4[51034] = 32'b00000000000000001010001011100101;
assign LUT_4[51035] = 32'b00000000000000000011010111011101;
assign LUT_4[51036] = 32'b00000000000000000111110001011101;
assign LUT_4[51037] = 32'b00000000000000000000111101010101;
assign LUT_4[51038] = 32'b00000000000000000111001100000001;
assign LUT_4[51039] = 32'b00000000000000000000010111111001;
assign LUT_4[51040] = 32'b00000000000000010010001110000101;
assign LUT_4[51041] = 32'b00000000000000001011011001111101;
assign LUT_4[51042] = 32'b00000000000000010001101000101001;
assign LUT_4[51043] = 32'b00000000000000001010110100100001;
assign LUT_4[51044] = 32'b00000000000000001111001110100001;
assign LUT_4[51045] = 32'b00000000000000001000011010011001;
assign LUT_4[51046] = 32'b00000000000000001110101001000101;
assign LUT_4[51047] = 32'b00000000000000000111110100111101;
assign LUT_4[51048] = 32'b00000000000000001011011010011010;
assign LUT_4[51049] = 32'b00000000000000000100100110010010;
assign LUT_4[51050] = 32'b00000000000000001010110100111110;
assign LUT_4[51051] = 32'b00000000000000000100000000110110;
assign LUT_4[51052] = 32'b00000000000000001000011010110110;
assign LUT_4[51053] = 32'b00000000000000000001100110101110;
assign LUT_4[51054] = 32'b00000000000000000111110101011010;
assign LUT_4[51055] = 32'b00000000000000000001000001010010;
assign LUT_4[51056] = 32'b00000000000000001111111111110011;
assign LUT_4[51057] = 32'b00000000000000001001001011101011;
assign LUT_4[51058] = 32'b00000000000000001111011010010111;
assign LUT_4[51059] = 32'b00000000000000001000100110001111;
assign LUT_4[51060] = 32'b00000000000000001101000000001111;
assign LUT_4[51061] = 32'b00000000000000000110001100000111;
assign LUT_4[51062] = 32'b00000000000000001100011010110011;
assign LUT_4[51063] = 32'b00000000000000000101100110101011;
assign LUT_4[51064] = 32'b00000000000000001001001100001000;
assign LUT_4[51065] = 32'b00000000000000000010011000000000;
assign LUT_4[51066] = 32'b00000000000000001000100110101100;
assign LUT_4[51067] = 32'b00000000000000000001110010100100;
assign LUT_4[51068] = 32'b00000000000000000110001100100100;
assign LUT_4[51069] = 32'b11111111111111111111011000011100;
assign LUT_4[51070] = 32'b00000000000000000101100111001000;
assign LUT_4[51071] = 32'b11111111111111111110110011000000;
assign LUT_4[51072] = 32'b00000000000000010101000001110010;
assign LUT_4[51073] = 32'b00000000000000001110001101101010;
assign LUT_4[51074] = 32'b00000000000000010100011100010110;
assign LUT_4[51075] = 32'b00000000000000001101101000001110;
assign LUT_4[51076] = 32'b00000000000000010010000010001110;
assign LUT_4[51077] = 32'b00000000000000001011001110000110;
assign LUT_4[51078] = 32'b00000000000000010001011100110010;
assign LUT_4[51079] = 32'b00000000000000001010101000101010;
assign LUT_4[51080] = 32'b00000000000000001110001110000111;
assign LUT_4[51081] = 32'b00000000000000000111011001111111;
assign LUT_4[51082] = 32'b00000000000000001101101000101011;
assign LUT_4[51083] = 32'b00000000000000000110110100100011;
assign LUT_4[51084] = 32'b00000000000000001011001110100011;
assign LUT_4[51085] = 32'b00000000000000000100011010011011;
assign LUT_4[51086] = 32'b00000000000000001010101001000111;
assign LUT_4[51087] = 32'b00000000000000000011110100111111;
assign LUT_4[51088] = 32'b00000000000000010010110011100000;
assign LUT_4[51089] = 32'b00000000000000001011111111011000;
assign LUT_4[51090] = 32'b00000000000000010010001110000100;
assign LUT_4[51091] = 32'b00000000000000001011011001111100;
assign LUT_4[51092] = 32'b00000000000000001111110011111100;
assign LUT_4[51093] = 32'b00000000000000001000111111110100;
assign LUT_4[51094] = 32'b00000000000000001111001110100000;
assign LUT_4[51095] = 32'b00000000000000001000011010011000;
assign LUT_4[51096] = 32'b00000000000000001011111111110101;
assign LUT_4[51097] = 32'b00000000000000000101001011101101;
assign LUT_4[51098] = 32'b00000000000000001011011010011001;
assign LUT_4[51099] = 32'b00000000000000000100100110010001;
assign LUT_4[51100] = 32'b00000000000000001001000000010001;
assign LUT_4[51101] = 32'b00000000000000000010001100001001;
assign LUT_4[51102] = 32'b00000000000000001000011010110101;
assign LUT_4[51103] = 32'b00000000000000000001100110101101;
assign LUT_4[51104] = 32'b00000000000000010011011100111001;
assign LUT_4[51105] = 32'b00000000000000001100101000110001;
assign LUT_4[51106] = 32'b00000000000000010010110111011101;
assign LUT_4[51107] = 32'b00000000000000001100000011010101;
assign LUT_4[51108] = 32'b00000000000000010000011101010101;
assign LUT_4[51109] = 32'b00000000000000001001101001001101;
assign LUT_4[51110] = 32'b00000000000000001111110111111001;
assign LUT_4[51111] = 32'b00000000000000001001000011110001;
assign LUT_4[51112] = 32'b00000000000000001100101001001110;
assign LUT_4[51113] = 32'b00000000000000000101110101000110;
assign LUT_4[51114] = 32'b00000000000000001100000011110010;
assign LUT_4[51115] = 32'b00000000000000000101001111101010;
assign LUT_4[51116] = 32'b00000000000000001001101001101010;
assign LUT_4[51117] = 32'b00000000000000000010110101100010;
assign LUT_4[51118] = 32'b00000000000000001001000100001110;
assign LUT_4[51119] = 32'b00000000000000000010010000000110;
assign LUT_4[51120] = 32'b00000000000000010001001110100111;
assign LUT_4[51121] = 32'b00000000000000001010011010011111;
assign LUT_4[51122] = 32'b00000000000000010000101001001011;
assign LUT_4[51123] = 32'b00000000000000001001110101000011;
assign LUT_4[51124] = 32'b00000000000000001110001111000011;
assign LUT_4[51125] = 32'b00000000000000000111011010111011;
assign LUT_4[51126] = 32'b00000000000000001101101001100111;
assign LUT_4[51127] = 32'b00000000000000000110110101011111;
assign LUT_4[51128] = 32'b00000000000000001010011010111100;
assign LUT_4[51129] = 32'b00000000000000000011100110110100;
assign LUT_4[51130] = 32'b00000000000000001001110101100000;
assign LUT_4[51131] = 32'b00000000000000000011000001011000;
assign LUT_4[51132] = 32'b00000000000000000111011011011000;
assign LUT_4[51133] = 32'b00000000000000000000100111010000;
assign LUT_4[51134] = 32'b00000000000000000110110101111100;
assign LUT_4[51135] = 32'b00000000000000000000000001110100;
assign LUT_4[51136] = 32'b00000000000000010110011001000110;
assign LUT_4[51137] = 32'b00000000000000001111100100111110;
assign LUT_4[51138] = 32'b00000000000000010101110011101010;
assign LUT_4[51139] = 32'b00000000000000001110111111100010;
assign LUT_4[51140] = 32'b00000000000000010011011001100010;
assign LUT_4[51141] = 32'b00000000000000001100100101011010;
assign LUT_4[51142] = 32'b00000000000000010010110100000110;
assign LUT_4[51143] = 32'b00000000000000001011111111111110;
assign LUT_4[51144] = 32'b00000000000000001111100101011011;
assign LUT_4[51145] = 32'b00000000000000001000110001010011;
assign LUT_4[51146] = 32'b00000000000000001110111111111111;
assign LUT_4[51147] = 32'b00000000000000001000001011110111;
assign LUT_4[51148] = 32'b00000000000000001100100101110111;
assign LUT_4[51149] = 32'b00000000000000000101110001101111;
assign LUT_4[51150] = 32'b00000000000000001100000000011011;
assign LUT_4[51151] = 32'b00000000000000000101001100010011;
assign LUT_4[51152] = 32'b00000000000000010100001010110100;
assign LUT_4[51153] = 32'b00000000000000001101010110101100;
assign LUT_4[51154] = 32'b00000000000000010011100101011000;
assign LUT_4[51155] = 32'b00000000000000001100110001010000;
assign LUT_4[51156] = 32'b00000000000000010001001011010000;
assign LUT_4[51157] = 32'b00000000000000001010010111001000;
assign LUT_4[51158] = 32'b00000000000000010000100101110100;
assign LUT_4[51159] = 32'b00000000000000001001110001101100;
assign LUT_4[51160] = 32'b00000000000000001101010111001001;
assign LUT_4[51161] = 32'b00000000000000000110100011000001;
assign LUT_4[51162] = 32'b00000000000000001100110001101101;
assign LUT_4[51163] = 32'b00000000000000000101111101100101;
assign LUT_4[51164] = 32'b00000000000000001010010111100101;
assign LUT_4[51165] = 32'b00000000000000000011100011011101;
assign LUT_4[51166] = 32'b00000000000000001001110010001001;
assign LUT_4[51167] = 32'b00000000000000000010111110000001;
assign LUT_4[51168] = 32'b00000000000000010100110100001101;
assign LUT_4[51169] = 32'b00000000000000001110000000000101;
assign LUT_4[51170] = 32'b00000000000000010100001110110001;
assign LUT_4[51171] = 32'b00000000000000001101011010101001;
assign LUT_4[51172] = 32'b00000000000000010001110100101001;
assign LUT_4[51173] = 32'b00000000000000001011000000100001;
assign LUT_4[51174] = 32'b00000000000000010001001111001101;
assign LUT_4[51175] = 32'b00000000000000001010011011000101;
assign LUT_4[51176] = 32'b00000000000000001110000000100010;
assign LUT_4[51177] = 32'b00000000000000000111001100011010;
assign LUT_4[51178] = 32'b00000000000000001101011011000110;
assign LUT_4[51179] = 32'b00000000000000000110100110111110;
assign LUT_4[51180] = 32'b00000000000000001011000000111110;
assign LUT_4[51181] = 32'b00000000000000000100001100110110;
assign LUT_4[51182] = 32'b00000000000000001010011011100010;
assign LUT_4[51183] = 32'b00000000000000000011100111011010;
assign LUT_4[51184] = 32'b00000000000000010010100101111011;
assign LUT_4[51185] = 32'b00000000000000001011110001110011;
assign LUT_4[51186] = 32'b00000000000000010010000000011111;
assign LUT_4[51187] = 32'b00000000000000001011001100010111;
assign LUT_4[51188] = 32'b00000000000000001111100110010111;
assign LUT_4[51189] = 32'b00000000000000001000110010001111;
assign LUT_4[51190] = 32'b00000000000000001111000000111011;
assign LUT_4[51191] = 32'b00000000000000001000001100110011;
assign LUT_4[51192] = 32'b00000000000000001011110010010000;
assign LUT_4[51193] = 32'b00000000000000000100111110001000;
assign LUT_4[51194] = 32'b00000000000000001011001100110100;
assign LUT_4[51195] = 32'b00000000000000000100011000101100;
assign LUT_4[51196] = 32'b00000000000000001000110010101100;
assign LUT_4[51197] = 32'b00000000000000000001111110100100;
assign LUT_4[51198] = 32'b00000000000000001000001101010000;
assign LUT_4[51199] = 32'b00000000000000000001011001001000;
assign LUT_4[51200] = 32'b00000000000000001000010000101010;
assign LUT_4[51201] = 32'b00000000000000000001011100100010;
assign LUT_4[51202] = 32'b00000000000000000111101011001110;
assign LUT_4[51203] = 32'b00000000000000000000110111000110;
assign LUT_4[51204] = 32'b00000000000000000101010001000110;
assign LUT_4[51205] = 32'b11111111111111111110011100111110;
assign LUT_4[51206] = 32'b00000000000000000100101011101010;
assign LUT_4[51207] = 32'b11111111111111111101110111100010;
assign LUT_4[51208] = 32'b00000000000000000001011100111111;
assign LUT_4[51209] = 32'b11111111111111111010101000110111;
assign LUT_4[51210] = 32'b00000000000000000000110111100011;
assign LUT_4[51211] = 32'b11111111111111111010000011011011;
assign LUT_4[51212] = 32'b11111111111111111110011101011011;
assign LUT_4[51213] = 32'b11111111111111110111101001010011;
assign LUT_4[51214] = 32'b11111111111111111101110111111111;
assign LUT_4[51215] = 32'b11111111111111110111000011110111;
assign LUT_4[51216] = 32'b00000000000000000110000010011000;
assign LUT_4[51217] = 32'b11111111111111111111001110010000;
assign LUT_4[51218] = 32'b00000000000000000101011100111100;
assign LUT_4[51219] = 32'b11111111111111111110101000110100;
assign LUT_4[51220] = 32'b00000000000000000011000010110100;
assign LUT_4[51221] = 32'b11111111111111111100001110101100;
assign LUT_4[51222] = 32'b00000000000000000010011101011000;
assign LUT_4[51223] = 32'b11111111111111111011101001010000;
assign LUT_4[51224] = 32'b11111111111111111111001110101101;
assign LUT_4[51225] = 32'b11111111111111111000011010100101;
assign LUT_4[51226] = 32'b11111111111111111110101001010001;
assign LUT_4[51227] = 32'b11111111111111110111110101001001;
assign LUT_4[51228] = 32'b11111111111111111100001111001001;
assign LUT_4[51229] = 32'b11111111111111110101011011000001;
assign LUT_4[51230] = 32'b11111111111111111011101001101101;
assign LUT_4[51231] = 32'b11111111111111110100110101100101;
assign LUT_4[51232] = 32'b00000000000000000110101011110001;
assign LUT_4[51233] = 32'b11111111111111111111110111101001;
assign LUT_4[51234] = 32'b00000000000000000110000110010101;
assign LUT_4[51235] = 32'b11111111111111111111010010001101;
assign LUT_4[51236] = 32'b00000000000000000011101100001101;
assign LUT_4[51237] = 32'b11111111111111111100111000000101;
assign LUT_4[51238] = 32'b00000000000000000011000110110001;
assign LUT_4[51239] = 32'b11111111111111111100010010101001;
assign LUT_4[51240] = 32'b11111111111111111111111000000110;
assign LUT_4[51241] = 32'b11111111111111111001000011111110;
assign LUT_4[51242] = 32'b11111111111111111111010010101010;
assign LUT_4[51243] = 32'b11111111111111111000011110100010;
assign LUT_4[51244] = 32'b11111111111111111100111000100010;
assign LUT_4[51245] = 32'b11111111111111110110000100011010;
assign LUT_4[51246] = 32'b11111111111111111100010011000110;
assign LUT_4[51247] = 32'b11111111111111110101011110111110;
assign LUT_4[51248] = 32'b00000000000000000100011101011111;
assign LUT_4[51249] = 32'b11111111111111111101101001010111;
assign LUT_4[51250] = 32'b00000000000000000011111000000011;
assign LUT_4[51251] = 32'b11111111111111111101000011111011;
assign LUT_4[51252] = 32'b00000000000000000001011101111011;
assign LUT_4[51253] = 32'b11111111111111111010101001110011;
assign LUT_4[51254] = 32'b00000000000000000000111000011111;
assign LUT_4[51255] = 32'b11111111111111111010000100010111;
assign LUT_4[51256] = 32'b11111111111111111101101001110100;
assign LUT_4[51257] = 32'b11111111111111110110110101101100;
assign LUT_4[51258] = 32'b11111111111111111101000100011000;
assign LUT_4[51259] = 32'b11111111111111110110010000010000;
assign LUT_4[51260] = 32'b11111111111111111010101010010000;
assign LUT_4[51261] = 32'b11111111111111110011110110001000;
assign LUT_4[51262] = 32'b11111111111111111010000100110100;
assign LUT_4[51263] = 32'b11111111111111110011010000101100;
assign LUT_4[51264] = 32'b00000000000000001001100111111110;
assign LUT_4[51265] = 32'b00000000000000000010110011110110;
assign LUT_4[51266] = 32'b00000000000000001001000010100010;
assign LUT_4[51267] = 32'b00000000000000000010001110011010;
assign LUT_4[51268] = 32'b00000000000000000110101000011010;
assign LUT_4[51269] = 32'b11111111111111111111110100010010;
assign LUT_4[51270] = 32'b00000000000000000110000010111110;
assign LUT_4[51271] = 32'b11111111111111111111001110110110;
assign LUT_4[51272] = 32'b00000000000000000010110100010011;
assign LUT_4[51273] = 32'b11111111111111111100000000001011;
assign LUT_4[51274] = 32'b00000000000000000010001110110111;
assign LUT_4[51275] = 32'b11111111111111111011011010101111;
assign LUT_4[51276] = 32'b11111111111111111111110100101111;
assign LUT_4[51277] = 32'b11111111111111111001000000100111;
assign LUT_4[51278] = 32'b11111111111111111111001111010011;
assign LUT_4[51279] = 32'b11111111111111111000011011001011;
assign LUT_4[51280] = 32'b00000000000000000111011001101100;
assign LUT_4[51281] = 32'b00000000000000000000100101100100;
assign LUT_4[51282] = 32'b00000000000000000110110100010000;
assign LUT_4[51283] = 32'b00000000000000000000000000001000;
assign LUT_4[51284] = 32'b00000000000000000100011010001000;
assign LUT_4[51285] = 32'b11111111111111111101100110000000;
assign LUT_4[51286] = 32'b00000000000000000011110100101100;
assign LUT_4[51287] = 32'b11111111111111111101000000100100;
assign LUT_4[51288] = 32'b00000000000000000000100110000001;
assign LUT_4[51289] = 32'b11111111111111111001110001111001;
assign LUT_4[51290] = 32'b00000000000000000000000000100101;
assign LUT_4[51291] = 32'b11111111111111111001001100011101;
assign LUT_4[51292] = 32'b11111111111111111101100110011101;
assign LUT_4[51293] = 32'b11111111111111110110110010010101;
assign LUT_4[51294] = 32'b11111111111111111101000001000001;
assign LUT_4[51295] = 32'b11111111111111110110001100111001;
assign LUT_4[51296] = 32'b00000000000000001000000011000101;
assign LUT_4[51297] = 32'b00000000000000000001001110111101;
assign LUT_4[51298] = 32'b00000000000000000111011101101001;
assign LUT_4[51299] = 32'b00000000000000000000101001100001;
assign LUT_4[51300] = 32'b00000000000000000101000011100001;
assign LUT_4[51301] = 32'b11111111111111111110001111011001;
assign LUT_4[51302] = 32'b00000000000000000100011110000101;
assign LUT_4[51303] = 32'b11111111111111111101101001111101;
assign LUT_4[51304] = 32'b00000000000000000001001111011010;
assign LUT_4[51305] = 32'b11111111111111111010011011010010;
assign LUT_4[51306] = 32'b00000000000000000000101001111110;
assign LUT_4[51307] = 32'b11111111111111111001110101110110;
assign LUT_4[51308] = 32'b11111111111111111110001111110110;
assign LUT_4[51309] = 32'b11111111111111110111011011101110;
assign LUT_4[51310] = 32'b11111111111111111101101010011010;
assign LUT_4[51311] = 32'b11111111111111110110110110010010;
assign LUT_4[51312] = 32'b00000000000000000101110100110011;
assign LUT_4[51313] = 32'b11111111111111111111000000101011;
assign LUT_4[51314] = 32'b00000000000000000101001111010111;
assign LUT_4[51315] = 32'b11111111111111111110011011001111;
assign LUT_4[51316] = 32'b00000000000000000010110101001111;
assign LUT_4[51317] = 32'b11111111111111111100000001000111;
assign LUT_4[51318] = 32'b00000000000000000010001111110011;
assign LUT_4[51319] = 32'b11111111111111111011011011101011;
assign LUT_4[51320] = 32'b11111111111111111111000001001000;
assign LUT_4[51321] = 32'b11111111111111111000001101000000;
assign LUT_4[51322] = 32'b11111111111111111110011011101100;
assign LUT_4[51323] = 32'b11111111111111110111100111100100;
assign LUT_4[51324] = 32'b11111111111111111100000001100100;
assign LUT_4[51325] = 32'b11111111111111110101001101011100;
assign LUT_4[51326] = 32'b11111111111111111011011100001000;
assign LUT_4[51327] = 32'b11111111111111110100101000000000;
assign LUT_4[51328] = 32'b00000000000000001010110110110010;
assign LUT_4[51329] = 32'b00000000000000000100000010101010;
assign LUT_4[51330] = 32'b00000000000000001010010001010110;
assign LUT_4[51331] = 32'b00000000000000000011011101001110;
assign LUT_4[51332] = 32'b00000000000000000111110111001110;
assign LUT_4[51333] = 32'b00000000000000000001000011000110;
assign LUT_4[51334] = 32'b00000000000000000111010001110010;
assign LUT_4[51335] = 32'b00000000000000000000011101101010;
assign LUT_4[51336] = 32'b00000000000000000100000011000111;
assign LUT_4[51337] = 32'b11111111111111111101001110111111;
assign LUT_4[51338] = 32'b00000000000000000011011101101011;
assign LUT_4[51339] = 32'b11111111111111111100101001100011;
assign LUT_4[51340] = 32'b00000000000000000001000011100011;
assign LUT_4[51341] = 32'b11111111111111111010001111011011;
assign LUT_4[51342] = 32'b00000000000000000000011110000111;
assign LUT_4[51343] = 32'b11111111111111111001101001111111;
assign LUT_4[51344] = 32'b00000000000000001000101000100000;
assign LUT_4[51345] = 32'b00000000000000000001110100011000;
assign LUT_4[51346] = 32'b00000000000000001000000011000100;
assign LUT_4[51347] = 32'b00000000000000000001001110111100;
assign LUT_4[51348] = 32'b00000000000000000101101000111100;
assign LUT_4[51349] = 32'b11111111111111111110110100110100;
assign LUT_4[51350] = 32'b00000000000000000101000011100000;
assign LUT_4[51351] = 32'b11111111111111111110001111011000;
assign LUT_4[51352] = 32'b00000000000000000001110100110101;
assign LUT_4[51353] = 32'b11111111111111111011000000101101;
assign LUT_4[51354] = 32'b00000000000000000001001111011001;
assign LUT_4[51355] = 32'b11111111111111111010011011010001;
assign LUT_4[51356] = 32'b11111111111111111110110101010001;
assign LUT_4[51357] = 32'b11111111111111111000000001001001;
assign LUT_4[51358] = 32'b11111111111111111110001111110101;
assign LUT_4[51359] = 32'b11111111111111110111011011101101;
assign LUT_4[51360] = 32'b00000000000000001001010001111001;
assign LUT_4[51361] = 32'b00000000000000000010011101110001;
assign LUT_4[51362] = 32'b00000000000000001000101100011101;
assign LUT_4[51363] = 32'b00000000000000000001111000010101;
assign LUT_4[51364] = 32'b00000000000000000110010010010101;
assign LUT_4[51365] = 32'b11111111111111111111011110001101;
assign LUT_4[51366] = 32'b00000000000000000101101100111001;
assign LUT_4[51367] = 32'b11111111111111111110111000110001;
assign LUT_4[51368] = 32'b00000000000000000010011110001110;
assign LUT_4[51369] = 32'b11111111111111111011101010000110;
assign LUT_4[51370] = 32'b00000000000000000001111000110010;
assign LUT_4[51371] = 32'b11111111111111111011000100101010;
assign LUT_4[51372] = 32'b11111111111111111111011110101010;
assign LUT_4[51373] = 32'b11111111111111111000101010100010;
assign LUT_4[51374] = 32'b11111111111111111110111001001110;
assign LUT_4[51375] = 32'b11111111111111111000000101000110;
assign LUT_4[51376] = 32'b00000000000000000111000011100111;
assign LUT_4[51377] = 32'b00000000000000000000001111011111;
assign LUT_4[51378] = 32'b00000000000000000110011110001011;
assign LUT_4[51379] = 32'b11111111111111111111101010000011;
assign LUT_4[51380] = 32'b00000000000000000100000100000011;
assign LUT_4[51381] = 32'b11111111111111111101001111111011;
assign LUT_4[51382] = 32'b00000000000000000011011110100111;
assign LUT_4[51383] = 32'b11111111111111111100101010011111;
assign LUT_4[51384] = 32'b00000000000000000000001111111100;
assign LUT_4[51385] = 32'b11111111111111111001011011110100;
assign LUT_4[51386] = 32'b11111111111111111111101010100000;
assign LUT_4[51387] = 32'b11111111111111111000110110011000;
assign LUT_4[51388] = 32'b11111111111111111101010000011000;
assign LUT_4[51389] = 32'b11111111111111110110011100010000;
assign LUT_4[51390] = 32'b11111111111111111100101010111100;
assign LUT_4[51391] = 32'b11111111111111110101110110110100;
assign LUT_4[51392] = 32'b00000000000000001100001110000110;
assign LUT_4[51393] = 32'b00000000000000000101011001111110;
assign LUT_4[51394] = 32'b00000000000000001011101000101010;
assign LUT_4[51395] = 32'b00000000000000000100110100100010;
assign LUT_4[51396] = 32'b00000000000000001001001110100010;
assign LUT_4[51397] = 32'b00000000000000000010011010011010;
assign LUT_4[51398] = 32'b00000000000000001000101001000110;
assign LUT_4[51399] = 32'b00000000000000000001110100111110;
assign LUT_4[51400] = 32'b00000000000000000101011010011011;
assign LUT_4[51401] = 32'b11111111111111111110100110010011;
assign LUT_4[51402] = 32'b00000000000000000100110100111111;
assign LUT_4[51403] = 32'b11111111111111111110000000110111;
assign LUT_4[51404] = 32'b00000000000000000010011010110111;
assign LUT_4[51405] = 32'b11111111111111111011100110101111;
assign LUT_4[51406] = 32'b00000000000000000001110101011011;
assign LUT_4[51407] = 32'b11111111111111111011000001010011;
assign LUT_4[51408] = 32'b00000000000000001001111111110100;
assign LUT_4[51409] = 32'b00000000000000000011001011101100;
assign LUT_4[51410] = 32'b00000000000000001001011010011000;
assign LUT_4[51411] = 32'b00000000000000000010100110010000;
assign LUT_4[51412] = 32'b00000000000000000111000000010000;
assign LUT_4[51413] = 32'b00000000000000000000001100001000;
assign LUT_4[51414] = 32'b00000000000000000110011010110100;
assign LUT_4[51415] = 32'b11111111111111111111100110101100;
assign LUT_4[51416] = 32'b00000000000000000011001100001001;
assign LUT_4[51417] = 32'b11111111111111111100011000000001;
assign LUT_4[51418] = 32'b00000000000000000010100110101101;
assign LUT_4[51419] = 32'b11111111111111111011110010100101;
assign LUT_4[51420] = 32'b00000000000000000000001100100101;
assign LUT_4[51421] = 32'b11111111111111111001011000011101;
assign LUT_4[51422] = 32'b11111111111111111111100111001001;
assign LUT_4[51423] = 32'b11111111111111111000110011000001;
assign LUT_4[51424] = 32'b00000000000000001010101001001101;
assign LUT_4[51425] = 32'b00000000000000000011110101000101;
assign LUT_4[51426] = 32'b00000000000000001010000011110001;
assign LUT_4[51427] = 32'b00000000000000000011001111101001;
assign LUT_4[51428] = 32'b00000000000000000111101001101001;
assign LUT_4[51429] = 32'b00000000000000000000110101100001;
assign LUT_4[51430] = 32'b00000000000000000111000100001101;
assign LUT_4[51431] = 32'b00000000000000000000010000000101;
assign LUT_4[51432] = 32'b00000000000000000011110101100010;
assign LUT_4[51433] = 32'b11111111111111111101000001011010;
assign LUT_4[51434] = 32'b00000000000000000011010000000110;
assign LUT_4[51435] = 32'b11111111111111111100011011111110;
assign LUT_4[51436] = 32'b00000000000000000000110101111110;
assign LUT_4[51437] = 32'b11111111111111111010000001110110;
assign LUT_4[51438] = 32'b00000000000000000000010000100010;
assign LUT_4[51439] = 32'b11111111111111111001011100011010;
assign LUT_4[51440] = 32'b00000000000000001000011010111011;
assign LUT_4[51441] = 32'b00000000000000000001100110110011;
assign LUT_4[51442] = 32'b00000000000000000111110101011111;
assign LUT_4[51443] = 32'b00000000000000000001000001010111;
assign LUT_4[51444] = 32'b00000000000000000101011011010111;
assign LUT_4[51445] = 32'b11111111111111111110100111001111;
assign LUT_4[51446] = 32'b00000000000000000100110101111011;
assign LUT_4[51447] = 32'b11111111111111111110000001110011;
assign LUT_4[51448] = 32'b00000000000000000001100111010000;
assign LUT_4[51449] = 32'b11111111111111111010110011001000;
assign LUT_4[51450] = 32'b00000000000000000001000001110100;
assign LUT_4[51451] = 32'b11111111111111111010001101101100;
assign LUT_4[51452] = 32'b11111111111111111110100111101100;
assign LUT_4[51453] = 32'b11111111111111110111110011100100;
assign LUT_4[51454] = 32'b11111111111111111110000010010000;
assign LUT_4[51455] = 32'b11111111111111110111001110001000;
assign LUT_4[51456] = 32'b00000000000000001101001100001101;
assign LUT_4[51457] = 32'b00000000000000000110011000000101;
assign LUT_4[51458] = 32'b00000000000000001100100110110001;
assign LUT_4[51459] = 32'b00000000000000000101110010101001;
assign LUT_4[51460] = 32'b00000000000000001010001100101001;
assign LUT_4[51461] = 32'b00000000000000000011011000100001;
assign LUT_4[51462] = 32'b00000000000000001001100111001101;
assign LUT_4[51463] = 32'b00000000000000000010110011000101;
assign LUT_4[51464] = 32'b00000000000000000110011000100010;
assign LUT_4[51465] = 32'b11111111111111111111100100011010;
assign LUT_4[51466] = 32'b00000000000000000101110011000110;
assign LUT_4[51467] = 32'b11111111111111111110111110111110;
assign LUT_4[51468] = 32'b00000000000000000011011000111110;
assign LUT_4[51469] = 32'b11111111111111111100100100110110;
assign LUT_4[51470] = 32'b00000000000000000010110011100010;
assign LUT_4[51471] = 32'b11111111111111111011111111011010;
assign LUT_4[51472] = 32'b00000000000000001010111101111011;
assign LUT_4[51473] = 32'b00000000000000000100001001110011;
assign LUT_4[51474] = 32'b00000000000000001010011000011111;
assign LUT_4[51475] = 32'b00000000000000000011100100010111;
assign LUT_4[51476] = 32'b00000000000000000111111110010111;
assign LUT_4[51477] = 32'b00000000000000000001001010001111;
assign LUT_4[51478] = 32'b00000000000000000111011000111011;
assign LUT_4[51479] = 32'b00000000000000000000100100110011;
assign LUT_4[51480] = 32'b00000000000000000100001010010000;
assign LUT_4[51481] = 32'b11111111111111111101010110001000;
assign LUT_4[51482] = 32'b00000000000000000011100100110100;
assign LUT_4[51483] = 32'b11111111111111111100110000101100;
assign LUT_4[51484] = 32'b00000000000000000001001010101100;
assign LUT_4[51485] = 32'b11111111111111111010010110100100;
assign LUT_4[51486] = 32'b00000000000000000000100101010000;
assign LUT_4[51487] = 32'b11111111111111111001110001001000;
assign LUT_4[51488] = 32'b00000000000000001011100111010100;
assign LUT_4[51489] = 32'b00000000000000000100110011001100;
assign LUT_4[51490] = 32'b00000000000000001011000001111000;
assign LUT_4[51491] = 32'b00000000000000000100001101110000;
assign LUT_4[51492] = 32'b00000000000000001000100111110000;
assign LUT_4[51493] = 32'b00000000000000000001110011101000;
assign LUT_4[51494] = 32'b00000000000000001000000010010100;
assign LUT_4[51495] = 32'b00000000000000000001001110001100;
assign LUT_4[51496] = 32'b00000000000000000100110011101001;
assign LUT_4[51497] = 32'b11111111111111111101111111100001;
assign LUT_4[51498] = 32'b00000000000000000100001110001101;
assign LUT_4[51499] = 32'b11111111111111111101011010000101;
assign LUT_4[51500] = 32'b00000000000000000001110100000101;
assign LUT_4[51501] = 32'b11111111111111111010111111111101;
assign LUT_4[51502] = 32'b00000000000000000001001110101001;
assign LUT_4[51503] = 32'b11111111111111111010011010100001;
assign LUT_4[51504] = 32'b00000000000000001001011001000010;
assign LUT_4[51505] = 32'b00000000000000000010100100111010;
assign LUT_4[51506] = 32'b00000000000000001000110011100110;
assign LUT_4[51507] = 32'b00000000000000000001111111011110;
assign LUT_4[51508] = 32'b00000000000000000110011001011110;
assign LUT_4[51509] = 32'b11111111111111111111100101010110;
assign LUT_4[51510] = 32'b00000000000000000101110100000010;
assign LUT_4[51511] = 32'b11111111111111111110111111111010;
assign LUT_4[51512] = 32'b00000000000000000010100101010111;
assign LUT_4[51513] = 32'b11111111111111111011110001001111;
assign LUT_4[51514] = 32'b00000000000000000001111111111011;
assign LUT_4[51515] = 32'b11111111111111111011001011110011;
assign LUT_4[51516] = 32'b11111111111111111111100101110011;
assign LUT_4[51517] = 32'b11111111111111111000110001101011;
assign LUT_4[51518] = 32'b11111111111111111111000000010111;
assign LUT_4[51519] = 32'b11111111111111111000001100001111;
assign LUT_4[51520] = 32'b00000000000000001110100011100001;
assign LUT_4[51521] = 32'b00000000000000000111101111011001;
assign LUT_4[51522] = 32'b00000000000000001101111110000101;
assign LUT_4[51523] = 32'b00000000000000000111001001111101;
assign LUT_4[51524] = 32'b00000000000000001011100011111101;
assign LUT_4[51525] = 32'b00000000000000000100101111110101;
assign LUT_4[51526] = 32'b00000000000000001010111110100001;
assign LUT_4[51527] = 32'b00000000000000000100001010011001;
assign LUT_4[51528] = 32'b00000000000000000111101111110110;
assign LUT_4[51529] = 32'b00000000000000000000111011101110;
assign LUT_4[51530] = 32'b00000000000000000111001010011010;
assign LUT_4[51531] = 32'b00000000000000000000010110010010;
assign LUT_4[51532] = 32'b00000000000000000100110000010010;
assign LUT_4[51533] = 32'b11111111111111111101111100001010;
assign LUT_4[51534] = 32'b00000000000000000100001010110110;
assign LUT_4[51535] = 32'b11111111111111111101010110101110;
assign LUT_4[51536] = 32'b00000000000000001100010101001111;
assign LUT_4[51537] = 32'b00000000000000000101100001000111;
assign LUT_4[51538] = 32'b00000000000000001011101111110011;
assign LUT_4[51539] = 32'b00000000000000000100111011101011;
assign LUT_4[51540] = 32'b00000000000000001001010101101011;
assign LUT_4[51541] = 32'b00000000000000000010100001100011;
assign LUT_4[51542] = 32'b00000000000000001000110000001111;
assign LUT_4[51543] = 32'b00000000000000000001111100000111;
assign LUT_4[51544] = 32'b00000000000000000101100001100100;
assign LUT_4[51545] = 32'b11111111111111111110101101011100;
assign LUT_4[51546] = 32'b00000000000000000100111100001000;
assign LUT_4[51547] = 32'b11111111111111111110001000000000;
assign LUT_4[51548] = 32'b00000000000000000010100010000000;
assign LUT_4[51549] = 32'b11111111111111111011101101111000;
assign LUT_4[51550] = 32'b00000000000000000001111100100100;
assign LUT_4[51551] = 32'b11111111111111111011001000011100;
assign LUT_4[51552] = 32'b00000000000000001100111110101000;
assign LUT_4[51553] = 32'b00000000000000000110001010100000;
assign LUT_4[51554] = 32'b00000000000000001100011001001100;
assign LUT_4[51555] = 32'b00000000000000000101100101000100;
assign LUT_4[51556] = 32'b00000000000000001001111111000100;
assign LUT_4[51557] = 32'b00000000000000000011001010111100;
assign LUT_4[51558] = 32'b00000000000000001001011001101000;
assign LUT_4[51559] = 32'b00000000000000000010100101100000;
assign LUT_4[51560] = 32'b00000000000000000110001010111101;
assign LUT_4[51561] = 32'b11111111111111111111010110110101;
assign LUT_4[51562] = 32'b00000000000000000101100101100001;
assign LUT_4[51563] = 32'b11111111111111111110110001011001;
assign LUT_4[51564] = 32'b00000000000000000011001011011001;
assign LUT_4[51565] = 32'b11111111111111111100010111010001;
assign LUT_4[51566] = 32'b00000000000000000010100101111101;
assign LUT_4[51567] = 32'b11111111111111111011110001110101;
assign LUT_4[51568] = 32'b00000000000000001010110000010110;
assign LUT_4[51569] = 32'b00000000000000000011111100001110;
assign LUT_4[51570] = 32'b00000000000000001010001010111010;
assign LUT_4[51571] = 32'b00000000000000000011010110110010;
assign LUT_4[51572] = 32'b00000000000000000111110000110010;
assign LUT_4[51573] = 32'b00000000000000000000111100101010;
assign LUT_4[51574] = 32'b00000000000000000111001011010110;
assign LUT_4[51575] = 32'b00000000000000000000010111001110;
assign LUT_4[51576] = 32'b00000000000000000011111100101011;
assign LUT_4[51577] = 32'b11111111111111111101001000100011;
assign LUT_4[51578] = 32'b00000000000000000011010111001111;
assign LUT_4[51579] = 32'b11111111111111111100100011000111;
assign LUT_4[51580] = 32'b00000000000000000000111101000111;
assign LUT_4[51581] = 32'b11111111111111111010001000111111;
assign LUT_4[51582] = 32'b00000000000000000000010111101011;
assign LUT_4[51583] = 32'b11111111111111111001100011100011;
assign LUT_4[51584] = 32'b00000000000000001111110010010101;
assign LUT_4[51585] = 32'b00000000000000001000111110001101;
assign LUT_4[51586] = 32'b00000000000000001111001100111001;
assign LUT_4[51587] = 32'b00000000000000001000011000110001;
assign LUT_4[51588] = 32'b00000000000000001100110010110001;
assign LUT_4[51589] = 32'b00000000000000000101111110101001;
assign LUT_4[51590] = 32'b00000000000000001100001101010101;
assign LUT_4[51591] = 32'b00000000000000000101011001001101;
assign LUT_4[51592] = 32'b00000000000000001000111110101010;
assign LUT_4[51593] = 32'b00000000000000000010001010100010;
assign LUT_4[51594] = 32'b00000000000000001000011001001110;
assign LUT_4[51595] = 32'b00000000000000000001100101000110;
assign LUT_4[51596] = 32'b00000000000000000101111111000110;
assign LUT_4[51597] = 32'b11111111111111111111001010111110;
assign LUT_4[51598] = 32'b00000000000000000101011001101010;
assign LUT_4[51599] = 32'b11111111111111111110100101100010;
assign LUT_4[51600] = 32'b00000000000000001101100100000011;
assign LUT_4[51601] = 32'b00000000000000000110101111111011;
assign LUT_4[51602] = 32'b00000000000000001100111110100111;
assign LUT_4[51603] = 32'b00000000000000000110001010011111;
assign LUT_4[51604] = 32'b00000000000000001010100100011111;
assign LUT_4[51605] = 32'b00000000000000000011110000010111;
assign LUT_4[51606] = 32'b00000000000000001001111111000011;
assign LUT_4[51607] = 32'b00000000000000000011001010111011;
assign LUT_4[51608] = 32'b00000000000000000110110000011000;
assign LUT_4[51609] = 32'b11111111111111111111111100010000;
assign LUT_4[51610] = 32'b00000000000000000110001010111100;
assign LUT_4[51611] = 32'b11111111111111111111010110110100;
assign LUT_4[51612] = 32'b00000000000000000011110000110100;
assign LUT_4[51613] = 32'b11111111111111111100111100101100;
assign LUT_4[51614] = 32'b00000000000000000011001011011000;
assign LUT_4[51615] = 32'b11111111111111111100010111010000;
assign LUT_4[51616] = 32'b00000000000000001110001101011100;
assign LUT_4[51617] = 32'b00000000000000000111011001010100;
assign LUT_4[51618] = 32'b00000000000000001101101000000000;
assign LUT_4[51619] = 32'b00000000000000000110110011111000;
assign LUT_4[51620] = 32'b00000000000000001011001101111000;
assign LUT_4[51621] = 32'b00000000000000000100011001110000;
assign LUT_4[51622] = 32'b00000000000000001010101000011100;
assign LUT_4[51623] = 32'b00000000000000000011110100010100;
assign LUT_4[51624] = 32'b00000000000000000111011001110001;
assign LUT_4[51625] = 32'b00000000000000000000100101101001;
assign LUT_4[51626] = 32'b00000000000000000110110100010101;
assign LUT_4[51627] = 32'b00000000000000000000000000001101;
assign LUT_4[51628] = 32'b00000000000000000100011010001101;
assign LUT_4[51629] = 32'b11111111111111111101100110000101;
assign LUT_4[51630] = 32'b00000000000000000011110100110001;
assign LUT_4[51631] = 32'b11111111111111111101000000101001;
assign LUT_4[51632] = 32'b00000000000000001011111111001010;
assign LUT_4[51633] = 32'b00000000000000000101001011000010;
assign LUT_4[51634] = 32'b00000000000000001011011001101110;
assign LUT_4[51635] = 32'b00000000000000000100100101100110;
assign LUT_4[51636] = 32'b00000000000000001000111111100110;
assign LUT_4[51637] = 32'b00000000000000000010001011011110;
assign LUT_4[51638] = 32'b00000000000000001000011010001010;
assign LUT_4[51639] = 32'b00000000000000000001100110000010;
assign LUT_4[51640] = 32'b00000000000000000101001011011111;
assign LUT_4[51641] = 32'b11111111111111111110010111010111;
assign LUT_4[51642] = 32'b00000000000000000100100110000011;
assign LUT_4[51643] = 32'b11111111111111111101110001111011;
assign LUT_4[51644] = 32'b00000000000000000010001011111011;
assign LUT_4[51645] = 32'b11111111111111111011010111110011;
assign LUT_4[51646] = 32'b00000000000000000001100110011111;
assign LUT_4[51647] = 32'b11111111111111111010110010010111;
assign LUT_4[51648] = 32'b00000000000000010001001001101001;
assign LUT_4[51649] = 32'b00000000000000001010010101100001;
assign LUT_4[51650] = 32'b00000000000000010000100100001101;
assign LUT_4[51651] = 32'b00000000000000001001110000000101;
assign LUT_4[51652] = 32'b00000000000000001110001010000101;
assign LUT_4[51653] = 32'b00000000000000000111010101111101;
assign LUT_4[51654] = 32'b00000000000000001101100100101001;
assign LUT_4[51655] = 32'b00000000000000000110110000100001;
assign LUT_4[51656] = 32'b00000000000000001010010101111110;
assign LUT_4[51657] = 32'b00000000000000000011100001110110;
assign LUT_4[51658] = 32'b00000000000000001001110000100010;
assign LUT_4[51659] = 32'b00000000000000000010111100011010;
assign LUT_4[51660] = 32'b00000000000000000111010110011010;
assign LUT_4[51661] = 32'b00000000000000000000100010010010;
assign LUT_4[51662] = 32'b00000000000000000110110000111110;
assign LUT_4[51663] = 32'b11111111111111111111111100110110;
assign LUT_4[51664] = 32'b00000000000000001110111011010111;
assign LUT_4[51665] = 32'b00000000000000001000000111001111;
assign LUT_4[51666] = 32'b00000000000000001110010101111011;
assign LUT_4[51667] = 32'b00000000000000000111100001110011;
assign LUT_4[51668] = 32'b00000000000000001011111011110011;
assign LUT_4[51669] = 32'b00000000000000000101000111101011;
assign LUT_4[51670] = 32'b00000000000000001011010110010111;
assign LUT_4[51671] = 32'b00000000000000000100100010001111;
assign LUT_4[51672] = 32'b00000000000000001000000111101100;
assign LUT_4[51673] = 32'b00000000000000000001010011100100;
assign LUT_4[51674] = 32'b00000000000000000111100010010000;
assign LUT_4[51675] = 32'b00000000000000000000101110001000;
assign LUT_4[51676] = 32'b00000000000000000101001000001000;
assign LUT_4[51677] = 32'b11111111111111111110010100000000;
assign LUT_4[51678] = 32'b00000000000000000100100010101100;
assign LUT_4[51679] = 32'b11111111111111111101101110100100;
assign LUT_4[51680] = 32'b00000000000000001111100100110000;
assign LUT_4[51681] = 32'b00000000000000001000110000101000;
assign LUT_4[51682] = 32'b00000000000000001110111111010100;
assign LUT_4[51683] = 32'b00000000000000001000001011001100;
assign LUT_4[51684] = 32'b00000000000000001100100101001100;
assign LUT_4[51685] = 32'b00000000000000000101110001000100;
assign LUT_4[51686] = 32'b00000000000000001011111111110000;
assign LUT_4[51687] = 32'b00000000000000000101001011101000;
assign LUT_4[51688] = 32'b00000000000000001000110001000101;
assign LUT_4[51689] = 32'b00000000000000000001111100111101;
assign LUT_4[51690] = 32'b00000000000000001000001011101001;
assign LUT_4[51691] = 32'b00000000000000000001010111100001;
assign LUT_4[51692] = 32'b00000000000000000101110001100001;
assign LUT_4[51693] = 32'b11111111111111111110111101011001;
assign LUT_4[51694] = 32'b00000000000000000101001100000101;
assign LUT_4[51695] = 32'b11111111111111111110010111111101;
assign LUT_4[51696] = 32'b00000000000000001101010110011110;
assign LUT_4[51697] = 32'b00000000000000000110100010010110;
assign LUT_4[51698] = 32'b00000000000000001100110001000010;
assign LUT_4[51699] = 32'b00000000000000000101111100111010;
assign LUT_4[51700] = 32'b00000000000000001010010110111010;
assign LUT_4[51701] = 32'b00000000000000000011100010110010;
assign LUT_4[51702] = 32'b00000000000000001001110001011110;
assign LUT_4[51703] = 32'b00000000000000000010111101010110;
assign LUT_4[51704] = 32'b00000000000000000110100010110011;
assign LUT_4[51705] = 32'b11111111111111111111101110101011;
assign LUT_4[51706] = 32'b00000000000000000101111101010111;
assign LUT_4[51707] = 32'b11111111111111111111001001001111;
assign LUT_4[51708] = 32'b00000000000000000011100011001111;
assign LUT_4[51709] = 32'b11111111111111111100101111000111;
assign LUT_4[51710] = 32'b00000000000000000010111101110011;
assign LUT_4[51711] = 32'b11111111111111111100001001101011;
assign LUT_4[51712] = 32'b00000000000000000111010100110010;
assign LUT_4[51713] = 32'b00000000000000000000100000101010;
assign LUT_4[51714] = 32'b00000000000000000110101111010110;
assign LUT_4[51715] = 32'b11111111111111111111111011001110;
assign LUT_4[51716] = 32'b00000000000000000100010101001110;
assign LUT_4[51717] = 32'b11111111111111111101100001000110;
assign LUT_4[51718] = 32'b00000000000000000011101111110010;
assign LUT_4[51719] = 32'b11111111111111111100111011101010;
assign LUT_4[51720] = 32'b00000000000000000000100001000111;
assign LUT_4[51721] = 32'b11111111111111111001101100111111;
assign LUT_4[51722] = 32'b11111111111111111111111011101011;
assign LUT_4[51723] = 32'b11111111111111111001000111100011;
assign LUT_4[51724] = 32'b11111111111111111101100001100011;
assign LUT_4[51725] = 32'b11111111111111110110101101011011;
assign LUT_4[51726] = 32'b11111111111111111100111100000111;
assign LUT_4[51727] = 32'b11111111111111110110000111111111;
assign LUT_4[51728] = 32'b00000000000000000101000110100000;
assign LUT_4[51729] = 32'b11111111111111111110010010011000;
assign LUT_4[51730] = 32'b00000000000000000100100001000100;
assign LUT_4[51731] = 32'b11111111111111111101101100111100;
assign LUT_4[51732] = 32'b00000000000000000010000110111100;
assign LUT_4[51733] = 32'b11111111111111111011010010110100;
assign LUT_4[51734] = 32'b00000000000000000001100001100000;
assign LUT_4[51735] = 32'b11111111111111111010101101011000;
assign LUT_4[51736] = 32'b11111111111111111110010010110101;
assign LUT_4[51737] = 32'b11111111111111110111011110101101;
assign LUT_4[51738] = 32'b11111111111111111101101101011001;
assign LUT_4[51739] = 32'b11111111111111110110111001010001;
assign LUT_4[51740] = 32'b11111111111111111011010011010001;
assign LUT_4[51741] = 32'b11111111111111110100011111001001;
assign LUT_4[51742] = 32'b11111111111111111010101101110101;
assign LUT_4[51743] = 32'b11111111111111110011111001101101;
assign LUT_4[51744] = 32'b00000000000000000101101111111001;
assign LUT_4[51745] = 32'b11111111111111111110111011110001;
assign LUT_4[51746] = 32'b00000000000000000101001010011101;
assign LUT_4[51747] = 32'b11111111111111111110010110010101;
assign LUT_4[51748] = 32'b00000000000000000010110000010101;
assign LUT_4[51749] = 32'b11111111111111111011111100001101;
assign LUT_4[51750] = 32'b00000000000000000010001010111001;
assign LUT_4[51751] = 32'b11111111111111111011010110110001;
assign LUT_4[51752] = 32'b11111111111111111110111100001110;
assign LUT_4[51753] = 32'b11111111111111111000001000000110;
assign LUT_4[51754] = 32'b11111111111111111110010110110010;
assign LUT_4[51755] = 32'b11111111111111110111100010101010;
assign LUT_4[51756] = 32'b11111111111111111011111100101010;
assign LUT_4[51757] = 32'b11111111111111110101001000100010;
assign LUT_4[51758] = 32'b11111111111111111011010111001110;
assign LUT_4[51759] = 32'b11111111111111110100100011000110;
assign LUT_4[51760] = 32'b00000000000000000011100001100111;
assign LUT_4[51761] = 32'b11111111111111111100101101011111;
assign LUT_4[51762] = 32'b00000000000000000010111100001011;
assign LUT_4[51763] = 32'b11111111111111111100001000000011;
assign LUT_4[51764] = 32'b00000000000000000000100010000011;
assign LUT_4[51765] = 32'b11111111111111111001101101111011;
assign LUT_4[51766] = 32'b11111111111111111111111100100111;
assign LUT_4[51767] = 32'b11111111111111111001001000011111;
assign LUT_4[51768] = 32'b11111111111111111100101101111100;
assign LUT_4[51769] = 32'b11111111111111110101111001110100;
assign LUT_4[51770] = 32'b11111111111111111100001000100000;
assign LUT_4[51771] = 32'b11111111111111110101010100011000;
assign LUT_4[51772] = 32'b11111111111111111001101110011000;
assign LUT_4[51773] = 32'b11111111111111110010111010010000;
assign LUT_4[51774] = 32'b11111111111111111001001000111100;
assign LUT_4[51775] = 32'b11111111111111110010010100110100;
assign LUT_4[51776] = 32'b00000000000000001000101100000110;
assign LUT_4[51777] = 32'b00000000000000000001110111111110;
assign LUT_4[51778] = 32'b00000000000000001000000110101010;
assign LUT_4[51779] = 32'b00000000000000000001010010100010;
assign LUT_4[51780] = 32'b00000000000000000101101100100010;
assign LUT_4[51781] = 32'b11111111111111111110111000011010;
assign LUT_4[51782] = 32'b00000000000000000101000111000110;
assign LUT_4[51783] = 32'b11111111111111111110010010111110;
assign LUT_4[51784] = 32'b00000000000000000001111000011011;
assign LUT_4[51785] = 32'b11111111111111111011000100010011;
assign LUT_4[51786] = 32'b00000000000000000001010010111111;
assign LUT_4[51787] = 32'b11111111111111111010011110110111;
assign LUT_4[51788] = 32'b11111111111111111110111000110111;
assign LUT_4[51789] = 32'b11111111111111111000000100101111;
assign LUT_4[51790] = 32'b11111111111111111110010011011011;
assign LUT_4[51791] = 32'b11111111111111110111011111010011;
assign LUT_4[51792] = 32'b00000000000000000110011101110100;
assign LUT_4[51793] = 32'b11111111111111111111101001101100;
assign LUT_4[51794] = 32'b00000000000000000101111000011000;
assign LUT_4[51795] = 32'b11111111111111111111000100010000;
assign LUT_4[51796] = 32'b00000000000000000011011110010000;
assign LUT_4[51797] = 32'b11111111111111111100101010001000;
assign LUT_4[51798] = 32'b00000000000000000010111000110100;
assign LUT_4[51799] = 32'b11111111111111111100000100101100;
assign LUT_4[51800] = 32'b11111111111111111111101010001001;
assign LUT_4[51801] = 32'b11111111111111111000110110000001;
assign LUT_4[51802] = 32'b11111111111111111111000100101101;
assign LUT_4[51803] = 32'b11111111111111111000010000100101;
assign LUT_4[51804] = 32'b11111111111111111100101010100101;
assign LUT_4[51805] = 32'b11111111111111110101110110011101;
assign LUT_4[51806] = 32'b11111111111111111100000101001001;
assign LUT_4[51807] = 32'b11111111111111110101010001000001;
assign LUT_4[51808] = 32'b00000000000000000111000111001101;
assign LUT_4[51809] = 32'b00000000000000000000010011000101;
assign LUT_4[51810] = 32'b00000000000000000110100001110001;
assign LUT_4[51811] = 32'b11111111111111111111101101101001;
assign LUT_4[51812] = 32'b00000000000000000100000111101001;
assign LUT_4[51813] = 32'b11111111111111111101010011100001;
assign LUT_4[51814] = 32'b00000000000000000011100010001101;
assign LUT_4[51815] = 32'b11111111111111111100101110000101;
assign LUT_4[51816] = 32'b00000000000000000000010011100010;
assign LUT_4[51817] = 32'b11111111111111111001011111011010;
assign LUT_4[51818] = 32'b11111111111111111111101110000110;
assign LUT_4[51819] = 32'b11111111111111111000111001111110;
assign LUT_4[51820] = 32'b11111111111111111101010011111110;
assign LUT_4[51821] = 32'b11111111111111110110011111110110;
assign LUT_4[51822] = 32'b11111111111111111100101110100010;
assign LUT_4[51823] = 32'b11111111111111110101111010011010;
assign LUT_4[51824] = 32'b00000000000000000100111000111011;
assign LUT_4[51825] = 32'b11111111111111111110000100110011;
assign LUT_4[51826] = 32'b00000000000000000100010011011111;
assign LUT_4[51827] = 32'b11111111111111111101011111010111;
assign LUT_4[51828] = 32'b00000000000000000001111001010111;
assign LUT_4[51829] = 32'b11111111111111111011000101001111;
assign LUT_4[51830] = 32'b00000000000000000001010011111011;
assign LUT_4[51831] = 32'b11111111111111111010011111110011;
assign LUT_4[51832] = 32'b11111111111111111110000101010000;
assign LUT_4[51833] = 32'b11111111111111110111010001001000;
assign LUT_4[51834] = 32'b11111111111111111101011111110100;
assign LUT_4[51835] = 32'b11111111111111110110101011101100;
assign LUT_4[51836] = 32'b11111111111111111011000101101100;
assign LUT_4[51837] = 32'b11111111111111110100010001100100;
assign LUT_4[51838] = 32'b11111111111111111010100000010000;
assign LUT_4[51839] = 32'b11111111111111110011101100001000;
assign LUT_4[51840] = 32'b00000000000000001001111010111010;
assign LUT_4[51841] = 32'b00000000000000000011000110110010;
assign LUT_4[51842] = 32'b00000000000000001001010101011110;
assign LUT_4[51843] = 32'b00000000000000000010100001010110;
assign LUT_4[51844] = 32'b00000000000000000110111011010110;
assign LUT_4[51845] = 32'b00000000000000000000000111001110;
assign LUT_4[51846] = 32'b00000000000000000110010101111010;
assign LUT_4[51847] = 32'b11111111111111111111100001110010;
assign LUT_4[51848] = 32'b00000000000000000011000111001111;
assign LUT_4[51849] = 32'b11111111111111111100010011000111;
assign LUT_4[51850] = 32'b00000000000000000010100001110011;
assign LUT_4[51851] = 32'b11111111111111111011101101101011;
assign LUT_4[51852] = 32'b00000000000000000000000111101011;
assign LUT_4[51853] = 32'b11111111111111111001010011100011;
assign LUT_4[51854] = 32'b11111111111111111111100010001111;
assign LUT_4[51855] = 32'b11111111111111111000101110000111;
assign LUT_4[51856] = 32'b00000000000000000111101100101000;
assign LUT_4[51857] = 32'b00000000000000000000111000100000;
assign LUT_4[51858] = 32'b00000000000000000111000111001100;
assign LUT_4[51859] = 32'b00000000000000000000010011000100;
assign LUT_4[51860] = 32'b00000000000000000100101101000100;
assign LUT_4[51861] = 32'b11111111111111111101111000111100;
assign LUT_4[51862] = 32'b00000000000000000100000111101000;
assign LUT_4[51863] = 32'b11111111111111111101010011100000;
assign LUT_4[51864] = 32'b00000000000000000000111000111101;
assign LUT_4[51865] = 32'b11111111111111111010000100110101;
assign LUT_4[51866] = 32'b00000000000000000000010011100001;
assign LUT_4[51867] = 32'b11111111111111111001011111011001;
assign LUT_4[51868] = 32'b11111111111111111101111001011001;
assign LUT_4[51869] = 32'b11111111111111110111000101010001;
assign LUT_4[51870] = 32'b11111111111111111101010011111101;
assign LUT_4[51871] = 32'b11111111111111110110011111110101;
assign LUT_4[51872] = 32'b00000000000000001000010110000001;
assign LUT_4[51873] = 32'b00000000000000000001100001111001;
assign LUT_4[51874] = 32'b00000000000000000111110000100101;
assign LUT_4[51875] = 32'b00000000000000000000111100011101;
assign LUT_4[51876] = 32'b00000000000000000101010110011101;
assign LUT_4[51877] = 32'b11111111111111111110100010010101;
assign LUT_4[51878] = 32'b00000000000000000100110001000001;
assign LUT_4[51879] = 32'b11111111111111111101111100111001;
assign LUT_4[51880] = 32'b00000000000000000001100010010110;
assign LUT_4[51881] = 32'b11111111111111111010101110001110;
assign LUT_4[51882] = 32'b00000000000000000000111100111010;
assign LUT_4[51883] = 32'b11111111111111111010001000110010;
assign LUT_4[51884] = 32'b11111111111111111110100010110010;
assign LUT_4[51885] = 32'b11111111111111110111101110101010;
assign LUT_4[51886] = 32'b11111111111111111101111101010110;
assign LUT_4[51887] = 32'b11111111111111110111001001001110;
assign LUT_4[51888] = 32'b00000000000000000110000111101111;
assign LUT_4[51889] = 32'b11111111111111111111010011100111;
assign LUT_4[51890] = 32'b00000000000000000101100010010011;
assign LUT_4[51891] = 32'b11111111111111111110101110001011;
assign LUT_4[51892] = 32'b00000000000000000011001000001011;
assign LUT_4[51893] = 32'b11111111111111111100010100000011;
assign LUT_4[51894] = 32'b00000000000000000010100010101111;
assign LUT_4[51895] = 32'b11111111111111111011101110100111;
assign LUT_4[51896] = 32'b11111111111111111111010100000100;
assign LUT_4[51897] = 32'b11111111111111111000011111111100;
assign LUT_4[51898] = 32'b11111111111111111110101110101000;
assign LUT_4[51899] = 32'b11111111111111110111111010100000;
assign LUT_4[51900] = 32'b11111111111111111100010100100000;
assign LUT_4[51901] = 32'b11111111111111110101100000011000;
assign LUT_4[51902] = 32'b11111111111111111011101111000100;
assign LUT_4[51903] = 32'b11111111111111110100111010111100;
assign LUT_4[51904] = 32'b00000000000000001011010010001110;
assign LUT_4[51905] = 32'b00000000000000000100011110000110;
assign LUT_4[51906] = 32'b00000000000000001010101100110010;
assign LUT_4[51907] = 32'b00000000000000000011111000101010;
assign LUT_4[51908] = 32'b00000000000000001000010010101010;
assign LUT_4[51909] = 32'b00000000000000000001011110100010;
assign LUT_4[51910] = 32'b00000000000000000111101101001110;
assign LUT_4[51911] = 32'b00000000000000000000111001000110;
assign LUT_4[51912] = 32'b00000000000000000100011110100011;
assign LUT_4[51913] = 32'b11111111111111111101101010011011;
assign LUT_4[51914] = 32'b00000000000000000011111001000111;
assign LUT_4[51915] = 32'b11111111111111111101000100111111;
assign LUT_4[51916] = 32'b00000000000000000001011110111111;
assign LUT_4[51917] = 32'b11111111111111111010101010110111;
assign LUT_4[51918] = 32'b00000000000000000000111001100011;
assign LUT_4[51919] = 32'b11111111111111111010000101011011;
assign LUT_4[51920] = 32'b00000000000000001001000011111100;
assign LUT_4[51921] = 32'b00000000000000000010001111110100;
assign LUT_4[51922] = 32'b00000000000000001000011110100000;
assign LUT_4[51923] = 32'b00000000000000000001101010011000;
assign LUT_4[51924] = 32'b00000000000000000110000100011000;
assign LUT_4[51925] = 32'b11111111111111111111010000010000;
assign LUT_4[51926] = 32'b00000000000000000101011110111100;
assign LUT_4[51927] = 32'b11111111111111111110101010110100;
assign LUT_4[51928] = 32'b00000000000000000010010000010001;
assign LUT_4[51929] = 32'b11111111111111111011011100001001;
assign LUT_4[51930] = 32'b00000000000000000001101010110101;
assign LUT_4[51931] = 32'b11111111111111111010110110101101;
assign LUT_4[51932] = 32'b11111111111111111111010000101101;
assign LUT_4[51933] = 32'b11111111111111111000011100100101;
assign LUT_4[51934] = 32'b11111111111111111110101011010001;
assign LUT_4[51935] = 32'b11111111111111110111110111001001;
assign LUT_4[51936] = 32'b00000000000000001001101101010101;
assign LUT_4[51937] = 32'b00000000000000000010111001001101;
assign LUT_4[51938] = 32'b00000000000000001001000111111001;
assign LUT_4[51939] = 32'b00000000000000000010010011110001;
assign LUT_4[51940] = 32'b00000000000000000110101101110001;
assign LUT_4[51941] = 32'b11111111111111111111111001101001;
assign LUT_4[51942] = 32'b00000000000000000110001000010101;
assign LUT_4[51943] = 32'b11111111111111111111010100001101;
assign LUT_4[51944] = 32'b00000000000000000010111001101010;
assign LUT_4[51945] = 32'b11111111111111111100000101100010;
assign LUT_4[51946] = 32'b00000000000000000010010100001110;
assign LUT_4[51947] = 32'b11111111111111111011100000000110;
assign LUT_4[51948] = 32'b11111111111111111111111010000110;
assign LUT_4[51949] = 32'b11111111111111111001000101111110;
assign LUT_4[51950] = 32'b11111111111111111111010100101010;
assign LUT_4[51951] = 32'b11111111111111111000100000100010;
assign LUT_4[51952] = 32'b00000000000000000111011111000011;
assign LUT_4[51953] = 32'b00000000000000000000101010111011;
assign LUT_4[51954] = 32'b00000000000000000110111001100111;
assign LUT_4[51955] = 32'b00000000000000000000000101011111;
assign LUT_4[51956] = 32'b00000000000000000100011111011111;
assign LUT_4[51957] = 32'b11111111111111111101101011010111;
assign LUT_4[51958] = 32'b00000000000000000011111010000011;
assign LUT_4[51959] = 32'b11111111111111111101000101111011;
assign LUT_4[51960] = 32'b00000000000000000000101011011000;
assign LUT_4[51961] = 32'b11111111111111111001110111010000;
assign LUT_4[51962] = 32'b00000000000000000000000101111100;
assign LUT_4[51963] = 32'b11111111111111111001010001110100;
assign LUT_4[51964] = 32'b11111111111111111101101011110100;
assign LUT_4[51965] = 32'b11111111111111110110110111101100;
assign LUT_4[51966] = 32'b11111111111111111101000110011000;
assign LUT_4[51967] = 32'b11111111111111110110010010010000;
assign LUT_4[51968] = 32'b00000000000000001100010000010101;
assign LUT_4[51969] = 32'b00000000000000000101011100001101;
assign LUT_4[51970] = 32'b00000000000000001011101010111001;
assign LUT_4[51971] = 32'b00000000000000000100110110110001;
assign LUT_4[51972] = 32'b00000000000000001001010000110001;
assign LUT_4[51973] = 32'b00000000000000000010011100101001;
assign LUT_4[51974] = 32'b00000000000000001000101011010101;
assign LUT_4[51975] = 32'b00000000000000000001110111001101;
assign LUT_4[51976] = 32'b00000000000000000101011100101010;
assign LUT_4[51977] = 32'b11111111111111111110101000100010;
assign LUT_4[51978] = 32'b00000000000000000100110111001110;
assign LUT_4[51979] = 32'b11111111111111111110000011000110;
assign LUT_4[51980] = 32'b00000000000000000010011101000110;
assign LUT_4[51981] = 32'b11111111111111111011101000111110;
assign LUT_4[51982] = 32'b00000000000000000001110111101010;
assign LUT_4[51983] = 32'b11111111111111111011000011100010;
assign LUT_4[51984] = 32'b00000000000000001010000010000011;
assign LUT_4[51985] = 32'b00000000000000000011001101111011;
assign LUT_4[51986] = 32'b00000000000000001001011100100111;
assign LUT_4[51987] = 32'b00000000000000000010101000011111;
assign LUT_4[51988] = 32'b00000000000000000111000010011111;
assign LUT_4[51989] = 32'b00000000000000000000001110010111;
assign LUT_4[51990] = 32'b00000000000000000110011101000011;
assign LUT_4[51991] = 32'b11111111111111111111101000111011;
assign LUT_4[51992] = 32'b00000000000000000011001110011000;
assign LUT_4[51993] = 32'b11111111111111111100011010010000;
assign LUT_4[51994] = 32'b00000000000000000010101000111100;
assign LUT_4[51995] = 32'b11111111111111111011110100110100;
assign LUT_4[51996] = 32'b00000000000000000000001110110100;
assign LUT_4[51997] = 32'b11111111111111111001011010101100;
assign LUT_4[51998] = 32'b11111111111111111111101001011000;
assign LUT_4[51999] = 32'b11111111111111111000110101010000;
assign LUT_4[52000] = 32'b00000000000000001010101011011100;
assign LUT_4[52001] = 32'b00000000000000000011110111010100;
assign LUT_4[52002] = 32'b00000000000000001010000110000000;
assign LUT_4[52003] = 32'b00000000000000000011010001111000;
assign LUT_4[52004] = 32'b00000000000000000111101011111000;
assign LUT_4[52005] = 32'b00000000000000000000110111110000;
assign LUT_4[52006] = 32'b00000000000000000111000110011100;
assign LUT_4[52007] = 32'b00000000000000000000010010010100;
assign LUT_4[52008] = 32'b00000000000000000011110111110001;
assign LUT_4[52009] = 32'b11111111111111111101000011101001;
assign LUT_4[52010] = 32'b00000000000000000011010010010101;
assign LUT_4[52011] = 32'b11111111111111111100011110001101;
assign LUT_4[52012] = 32'b00000000000000000000111000001101;
assign LUT_4[52013] = 32'b11111111111111111010000100000101;
assign LUT_4[52014] = 32'b00000000000000000000010010110001;
assign LUT_4[52015] = 32'b11111111111111111001011110101001;
assign LUT_4[52016] = 32'b00000000000000001000011101001010;
assign LUT_4[52017] = 32'b00000000000000000001101001000010;
assign LUT_4[52018] = 32'b00000000000000000111110111101110;
assign LUT_4[52019] = 32'b00000000000000000001000011100110;
assign LUT_4[52020] = 32'b00000000000000000101011101100110;
assign LUT_4[52021] = 32'b11111111111111111110101001011110;
assign LUT_4[52022] = 32'b00000000000000000100111000001010;
assign LUT_4[52023] = 32'b11111111111111111110000100000010;
assign LUT_4[52024] = 32'b00000000000000000001101001011111;
assign LUT_4[52025] = 32'b11111111111111111010110101010111;
assign LUT_4[52026] = 32'b00000000000000000001000100000011;
assign LUT_4[52027] = 32'b11111111111111111010001111111011;
assign LUT_4[52028] = 32'b11111111111111111110101001111011;
assign LUT_4[52029] = 32'b11111111111111110111110101110011;
assign LUT_4[52030] = 32'b11111111111111111110000100011111;
assign LUT_4[52031] = 32'b11111111111111110111010000010111;
assign LUT_4[52032] = 32'b00000000000000001101100111101001;
assign LUT_4[52033] = 32'b00000000000000000110110011100001;
assign LUT_4[52034] = 32'b00000000000000001101000010001101;
assign LUT_4[52035] = 32'b00000000000000000110001110000101;
assign LUT_4[52036] = 32'b00000000000000001010101000000101;
assign LUT_4[52037] = 32'b00000000000000000011110011111101;
assign LUT_4[52038] = 32'b00000000000000001010000010101001;
assign LUT_4[52039] = 32'b00000000000000000011001110100001;
assign LUT_4[52040] = 32'b00000000000000000110110011111110;
assign LUT_4[52041] = 32'b11111111111111111111111111110110;
assign LUT_4[52042] = 32'b00000000000000000110001110100010;
assign LUT_4[52043] = 32'b11111111111111111111011010011010;
assign LUT_4[52044] = 32'b00000000000000000011110100011010;
assign LUT_4[52045] = 32'b11111111111111111101000000010010;
assign LUT_4[52046] = 32'b00000000000000000011001110111110;
assign LUT_4[52047] = 32'b11111111111111111100011010110110;
assign LUT_4[52048] = 32'b00000000000000001011011001010111;
assign LUT_4[52049] = 32'b00000000000000000100100101001111;
assign LUT_4[52050] = 32'b00000000000000001010110011111011;
assign LUT_4[52051] = 32'b00000000000000000011111111110011;
assign LUT_4[52052] = 32'b00000000000000001000011001110011;
assign LUT_4[52053] = 32'b00000000000000000001100101101011;
assign LUT_4[52054] = 32'b00000000000000000111110100010111;
assign LUT_4[52055] = 32'b00000000000000000001000000001111;
assign LUT_4[52056] = 32'b00000000000000000100100101101100;
assign LUT_4[52057] = 32'b11111111111111111101110001100100;
assign LUT_4[52058] = 32'b00000000000000000100000000010000;
assign LUT_4[52059] = 32'b11111111111111111101001100001000;
assign LUT_4[52060] = 32'b00000000000000000001100110001000;
assign LUT_4[52061] = 32'b11111111111111111010110010000000;
assign LUT_4[52062] = 32'b00000000000000000001000000101100;
assign LUT_4[52063] = 32'b11111111111111111010001100100100;
assign LUT_4[52064] = 32'b00000000000000001100000010110000;
assign LUT_4[52065] = 32'b00000000000000000101001110101000;
assign LUT_4[52066] = 32'b00000000000000001011011101010100;
assign LUT_4[52067] = 32'b00000000000000000100101001001100;
assign LUT_4[52068] = 32'b00000000000000001001000011001100;
assign LUT_4[52069] = 32'b00000000000000000010001111000100;
assign LUT_4[52070] = 32'b00000000000000001000011101110000;
assign LUT_4[52071] = 32'b00000000000000000001101001101000;
assign LUT_4[52072] = 32'b00000000000000000101001111000101;
assign LUT_4[52073] = 32'b11111111111111111110011010111101;
assign LUT_4[52074] = 32'b00000000000000000100101001101001;
assign LUT_4[52075] = 32'b11111111111111111101110101100001;
assign LUT_4[52076] = 32'b00000000000000000010001111100001;
assign LUT_4[52077] = 32'b11111111111111111011011011011001;
assign LUT_4[52078] = 32'b00000000000000000001101010000101;
assign LUT_4[52079] = 32'b11111111111111111010110101111101;
assign LUT_4[52080] = 32'b00000000000000001001110100011110;
assign LUT_4[52081] = 32'b00000000000000000011000000010110;
assign LUT_4[52082] = 32'b00000000000000001001001111000010;
assign LUT_4[52083] = 32'b00000000000000000010011010111010;
assign LUT_4[52084] = 32'b00000000000000000110110100111010;
assign LUT_4[52085] = 32'b00000000000000000000000000110010;
assign LUT_4[52086] = 32'b00000000000000000110001111011110;
assign LUT_4[52087] = 32'b11111111111111111111011011010110;
assign LUT_4[52088] = 32'b00000000000000000011000000110011;
assign LUT_4[52089] = 32'b11111111111111111100001100101011;
assign LUT_4[52090] = 32'b00000000000000000010011011010111;
assign LUT_4[52091] = 32'b11111111111111111011100111001111;
assign LUT_4[52092] = 32'b00000000000000000000000001001111;
assign LUT_4[52093] = 32'b11111111111111111001001101000111;
assign LUT_4[52094] = 32'b11111111111111111111011011110011;
assign LUT_4[52095] = 32'b11111111111111111000100111101011;
assign LUT_4[52096] = 32'b00000000000000001110110110011101;
assign LUT_4[52097] = 32'b00000000000000001000000010010101;
assign LUT_4[52098] = 32'b00000000000000001110010001000001;
assign LUT_4[52099] = 32'b00000000000000000111011100111001;
assign LUT_4[52100] = 32'b00000000000000001011110110111001;
assign LUT_4[52101] = 32'b00000000000000000101000010110001;
assign LUT_4[52102] = 32'b00000000000000001011010001011101;
assign LUT_4[52103] = 32'b00000000000000000100011101010101;
assign LUT_4[52104] = 32'b00000000000000001000000010110010;
assign LUT_4[52105] = 32'b00000000000000000001001110101010;
assign LUT_4[52106] = 32'b00000000000000000111011101010110;
assign LUT_4[52107] = 32'b00000000000000000000101001001110;
assign LUT_4[52108] = 32'b00000000000000000101000011001110;
assign LUT_4[52109] = 32'b11111111111111111110001111000110;
assign LUT_4[52110] = 32'b00000000000000000100011101110010;
assign LUT_4[52111] = 32'b11111111111111111101101001101010;
assign LUT_4[52112] = 32'b00000000000000001100101000001011;
assign LUT_4[52113] = 32'b00000000000000000101110100000011;
assign LUT_4[52114] = 32'b00000000000000001100000010101111;
assign LUT_4[52115] = 32'b00000000000000000101001110100111;
assign LUT_4[52116] = 32'b00000000000000001001101000100111;
assign LUT_4[52117] = 32'b00000000000000000010110100011111;
assign LUT_4[52118] = 32'b00000000000000001001000011001011;
assign LUT_4[52119] = 32'b00000000000000000010001111000011;
assign LUT_4[52120] = 32'b00000000000000000101110100100000;
assign LUT_4[52121] = 32'b11111111111111111111000000011000;
assign LUT_4[52122] = 32'b00000000000000000101001111000100;
assign LUT_4[52123] = 32'b11111111111111111110011010111100;
assign LUT_4[52124] = 32'b00000000000000000010110100111100;
assign LUT_4[52125] = 32'b11111111111111111100000000110100;
assign LUT_4[52126] = 32'b00000000000000000010001111100000;
assign LUT_4[52127] = 32'b11111111111111111011011011011000;
assign LUT_4[52128] = 32'b00000000000000001101010001100100;
assign LUT_4[52129] = 32'b00000000000000000110011101011100;
assign LUT_4[52130] = 32'b00000000000000001100101100001000;
assign LUT_4[52131] = 32'b00000000000000000101111000000000;
assign LUT_4[52132] = 32'b00000000000000001010010010000000;
assign LUT_4[52133] = 32'b00000000000000000011011101111000;
assign LUT_4[52134] = 32'b00000000000000001001101100100100;
assign LUT_4[52135] = 32'b00000000000000000010111000011100;
assign LUT_4[52136] = 32'b00000000000000000110011101111001;
assign LUT_4[52137] = 32'b11111111111111111111101001110001;
assign LUT_4[52138] = 32'b00000000000000000101111000011101;
assign LUT_4[52139] = 32'b11111111111111111111000100010101;
assign LUT_4[52140] = 32'b00000000000000000011011110010101;
assign LUT_4[52141] = 32'b11111111111111111100101010001101;
assign LUT_4[52142] = 32'b00000000000000000010111000111001;
assign LUT_4[52143] = 32'b11111111111111111100000100110001;
assign LUT_4[52144] = 32'b00000000000000001011000011010010;
assign LUT_4[52145] = 32'b00000000000000000100001111001010;
assign LUT_4[52146] = 32'b00000000000000001010011101110110;
assign LUT_4[52147] = 32'b00000000000000000011101001101110;
assign LUT_4[52148] = 32'b00000000000000001000000011101110;
assign LUT_4[52149] = 32'b00000000000000000001001111100110;
assign LUT_4[52150] = 32'b00000000000000000111011110010010;
assign LUT_4[52151] = 32'b00000000000000000000101010001010;
assign LUT_4[52152] = 32'b00000000000000000100001111100111;
assign LUT_4[52153] = 32'b11111111111111111101011011011111;
assign LUT_4[52154] = 32'b00000000000000000011101010001011;
assign LUT_4[52155] = 32'b11111111111111111100110110000011;
assign LUT_4[52156] = 32'b00000000000000000001010000000011;
assign LUT_4[52157] = 32'b11111111111111111010011011111011;
assign LUT_4[52158] = 32'b00000000000000000000101010100111;
assign LUT_4[52159] = 32'b11111111111111111001110110011111;
assign LUT_4[52160] = 32'b00000000000000010000001101110001;
assign LUT_4[52161] = 32'b00000000000000001001011001101001;
assign LUT_4[52162] = 32'b00000000000000001111101000010101;
assign LUT_4[52163] = 32'b00000000000000001000110100001101;
assign LUT_4[52164] = 32'b00000000000000001101001110001101;
assign LUT_4[52165] = 32'b00000000000000000110011010000101;
assign LUT_4[52166] = 32'b00000000000000001100101000110001;
assign LUT_4[52167] = 32'b00000000000000000101110100101001;
assign LUT_4[52168] = 32'b00000000000000001001011010000110;
assign LUT_4[52169] = 32'b00000000000000000010100101111110;
assign LUT_4[52170] = 32'b00000000000000001000110100101010;
assign LUT_4[52171] = 32'b00000000000000000010000000100010;
assign LUT_4[52172] = 32'b00000000000000000110011010100010;
assign LUT_4[52173] = 32'b11111111111111111111100110011010;
assign LUT_4[52174] = 32'b00000000000000000101110101000110;
assign LUT_4[52175] = 32'b11111111111111111111000000111110;
assign LUT_4[52176] = 32'b00000000000000001101111111011111;
assign LUT_4[52177] = 32'b00000000000000000111001011010111;
assign LUT_4[52178] = 32'b00000000000000001101011010000011;
assign LUT_4[52179] = 32'b00000000000000000110100101111011;
assign LUT_4[52180] = 32'b00000000000000001010111111111011;
assign LUT_4[52181] = 32'b00000000000000000100001011110011;
assign LUT_4[52182] = 32'b00000000000000001010011010011111;
assign LUT_4[52183] = 32'b00000000000000000011100110010111;
assign LUT_4[52184] = 32'b00000000000000000111001011110100;
assign LUT_4[52185] = 32'b00000000000000000000010111101100;
assign LUT_4[52186] = 32'b00000000000000000110100110011000;
assign LUT_4[52187] = 32'b11111111111111111111110010010000;
assign LUT_4[52188] = 32'b00000000000000000100001100010000;
assign LUT_4[52189] = 32'b11111111111111111101011000001000;
assign LUT_4[52190] = 32'b00000000000000000011100110110100;
assign LUT_4[52191] = 32'b11111111111111111100110010101100;
assign LUT_4[52192] = 32'b00000000000000001110101000111000;
assign LUT_4[52193] = 32'b00000000000000000111110100110000;
assign LUT_4[52194] = 32'b00000000000000001110000011011100;
assign LUT_4[52195] = 32'b00000000000000000111001111010100;
assign LUT_4[52196] = 32'b00000000000000001011101001010100;
assign LUT_4[52197] = 32'b00000000000000000100110101001100;
assign LUT_4[52198] = 32'b00000000000000001011000011111000;
assign LUT_4[52199] = 32'b00000000000000000100001111110000;
assign LUT_4[52200] = 32'b00000000000000000111110101001101;
assign LUT_4[52201] = 32'b00000000000000000001000001000101;
assign LUT_4[52202] = 32'b00000000000000000111001111110001;
assign LUT_4[52203] = 32'b00000000000000000000011011101001;
assign LUT_4[52204] = 32'b00000000000000000100110101101001;
assign LUT_4[52205] = 32'b11111111111111111110000001100001;
assign LUT_4[52206] = 32'b00000000000000000100010000001101;
assign LUT_4[52207] = 32'b11111111111111111101011100000101;
assign LUT_4[52208] = 32'b00000000000000001100011010100110;
assign LUT_4[52209] = 32'b00000000000000000101100110011110;
assign LUT_4[52210] = 32'b00000000000000001011110101001010;
assign LUT_4[52211] = 32'b00000000000000000101000001000010;
assign LUT_4[52212] = 32'b00000000000000001001011011000010;
assign LUT_4[52213] = 32'b00000000000000000010100110111010;
assign LUT_4[52214] = 32'b00000000000000001000110101100110;
assign LUT_4[52215] = 32'b00000000000000000010000001011110;
assign LUT_4[52216] = 32'b00000000000000000101100110111011;
assign LUT_4[52217] = 32'b11111111111111111110110010110011;
assign LUT_4[52218] = 32'b00000000000000000101000001011111;
assign LUT_4[52219] = 32'b11111111111111111110001101010111;
assign LUT_4[52220] = 32'b00000000000000000010100111010111;
assign LUT_4[52221] = 32'b11111111111111111011110011001111;
assign LUT_4[52222] = 32'b00000000000000000010000001111011;
assign LUT_4[52223] = 32'b11111111111111111011001101110011;
assign LUT_4[52224] = 32'b00000000000000001001111011001001;
assign LUT_4[52225] = 32'b00000000000000000011000111000001;
assign LUT_4[52226] = 32'b00000000000000001001010101101101;
assign LUT_4[52227] = 32'b00000000000000000010100001100101;
assign LUT_4[52228] = 32'b00000000000000000110111011100101;
assign LUT_4[52229] = 32'b00000000000000000000000111011101;
assign LUT_4[52230] = 32'b00000000000000000110010110001001;
assign LUT_4[52231] = 32'b11111111111111111111100010000001;
assign LUT_4[52232] = 32'b00000000000000000011000111011110;
assign LUT_4[52233] = 32'b11111111111111111100010011010110;
assign LUT_4[52234] = 32'b00000000000000000010100010000010;
assign LUT_4[52235] = 32'b11111111111111111011101101111010;
assign LUT_4[52236] = 32'b00000000000000000000000111111010;
assign LUT_4[52237] = 32'b11111111111111111001010011110010;
assign LUT_4[52238] = 32'b11111111111111111111100010011110;
assign LUT_4[52239] = 32'b11111111111111111000101110010110;
assign LUT_4[52240] = 32'b00000000000000000111101100110111;
assign LUT_4[52241] = 32'b00000000000000000000111000101111;
assign LUT_4[52242] = 32'b00000000000000000111000111011011;
assign LUT_4[52243] = 32'b00000000000000000000010011010011;
assign LUT_4[52244] = 32'b00000000000000000100101101010011;
assign LUT_4[52245] = 32'b11111111111111111101111001001011;
assign LUT_4[52246] = 32'b00000000000000000100000111110111;
assign LUT_4[52247] = 32'b11111111111111111101010011101111;
assign LUT_4[52248] = 32'b00000000000000000000111001001100;
assign LUT_4[52249] = 32'b11111111111111111010000101000100;
assign LUT_4[52250] = 32'b00000000000000000000010011110000;
assign LUT_4[52251] = 32'b11111111111111111001011111101000;
assign LUT_4[52252] = 32'b11111111111111111101111001101000;
assign LUT_4[52253] = 32'b11111111111111110111000101100000;
assign LUT_4[52254] = 32'b11111111111111111101010100001100;
assign LUT_4[52255] = 32'b11111111111111110110100000000100;
assign LUT_4[52256] = 32'b00000000000000001000010110010000;
assign LUT_4[52257] = 32'b00000000000000000001100010001000;
assign LUT_4[52258] = 32'b00000000000000000111110000110100;
assign LUT_4[52259] = 32'b00000000000000000000111100101100;
assign LUT_4[52260] = 32'b00000000000000000101010110101100;
assign LUT_4[52261] = 32'b11111111111111111110100010100100;
assign LUT_4[52262] = 32'b00000000000000000100110001010000;
assign LUT_4[52263] = 32'b11111111111111111101111101001000;
assign LUT_4[52264] = 32'b00000000000000000001100010100101;
assign LUT_4[52265] = 32'b11111111111111111010101110011101;
assign LUT_4[52266] = 32'b00000000000000000000111101001001;
assign LUT_4[52267] = 32'b11111111111111111010001001000001;
assign LUT_4[52268] = 32'b11111111111111111110100011000001;
assign LUT_4[52269] = 32'b11111111111111110111101110111001;
assign LUT_4[52270] = 32'b11111111111111111101111101100101;
assign LUT_4[52271] = 32'b11111111111111110111001001011101;
assign LUT_4[52272] = 32'b00000000000000000110000111111110;
assign LUT_4[52273] = 32'b11111111111111111111010011110110;
assign LUT_4[52274] = 32'b00000000000000000101100010100010;
assign LUT_4[52275] = 32'b11111111111111111110101110011010;
assign LUT_4[52276] = 32'b00000000000000000011001000011010;
assign LUT_4[52277] = 32'b11111111111111111100010100010010;
assign LUT_4[52278] = 32'b00000000000000000010100010111110;
assign LUT_4[52279] = 32'b11111111111111111011101110110110;
assign LUT_4[52280] = 32'b11111111111111111111010100010011;
assign LUT_4[52281] = 32'b11111111111111111000100000001011;
assign LUT_4[52282] = 32'b11111111111111111110101110110111;
assign LUT_4[52283] = 32'b11111111111111110111111010101111;
assign LUT_4[52284] = 32'b11111111111111111100010100101111;
assign LUT_4[52285] = 32'b11111111111111110101100000100111;
assign LUT_4[52286] = 32'b11111111111111111011101111010011;
assign LUT_4[52287] = 32'b11111111111111110100111011001011;
assign LUT_4[52288] = 32'b00000000000000001011010010011101;
assign LUT_4[52289] = 32'b00000000000000000100011110010101;
assign LUT_4[52290] = 32'b00000000000000001010101101000001;
assign LUT_4[52291] = 32'b00000000000000000011111000111001;
assign LUT_4[52292] = 32'b00000000000000001000010010111001;
assign LUT_4[52293] = 32'b00000000000000000001011110110001;
assign LUT_4[52294] = 32'b00000000000000000111101101011101;
assign LUT_4[52295] = 32'b00000000000000000000111001010101;
assign LUT_4[52296] = 32'b00000000000000000100011110110010;
assign LUT_4[52297] = 32'b11111111111111111101101010101010;
assign LUT_4[52298] = 32'b00000000000000000011111001010110;
assign LUT_4[52299] = 32'b11111111111111111101000101001110;
assign LUT_4[52300] = 32'b00000000000000000001011111001110;
assign LUT_4[52301] = 32'b11111111111111111010101011000110;
assign LUT_4[52302] = 32'b00000000000000000000111001110010;
assign LUT_4[52303] = 32'b11111111111111111010000101101010;
assign LUT_4[52304] = 32'b00000000000000001001000100001011;
assign LUT_4[52305] = 32'b00000000000000000010010000000011;
assign LUT_4[52306] = 32'b00000000000000001000011110101111;
assign LUT_4[52307] = 32'b00000000000000000001101010100111;
assign LUT_4[52308] = 32'b00000000000000000110000100100111;
assign LUT_4[52309] = 32'b11111111111111111111010000011111;
assign LUT_4[52310] = 32'b00000000000000000101011111001011;
assign LUT_4[52311] = 32'b11111111111111111110101011000011;
assign LUT_4[52312] = 32'b00000000000000000010010000100000;
assign LUT_4[52313] = 32'b11111111111111111011011100011000;
assign LUT_4[52314] = 32'b00000000000000000001101011000100;
assign LUT_4[52315] = 32'b11111111111111111010110110111100;
assign LUT_4[52316] = 32'b11111111111111111111010000111100;
assign LUT_4[52317] = 32'b11111111111111111000011100110100;
assign LUT_4[52318] = 32'b11111111111111111110101011100000;
assign LUT_4[52319] = 32'b11111111111111110111110111011000;
assign LUT_4[52320] = 32'b00000000000000001001101101100100;
assign LUT_4[52321] = 32'b00000000000000000010111001011100;
assign LUT_4[52322] = 32'b00000000000000001001001000001000;
assign LUT_4[52323] = 32'b00000000000000000010010100000000;
assign LUT_4[52324] = 32'b00000000000000000110101110000000;
assign LUT_4[52325] = 32'b11111111111111111111111001111000;
assign LUT_4[52326] = 32'b00000000000000000110001000100100;
assign LUT_4[52327] = 32'b11111111111111111111010100011100;
assign LUT_4[52328] = 32'b00000000000000000010111001111001;
assign LUT_4[52329] = 32'b11111111111111111100000101110001;
assign LUT_4[52330] = 32'b00000000000000000010010100011101;
assign LUT_4[52331] = 32'b11111111111111111011100000010101;
assign LUT_4[52332] = 32'b11111111111111111111111010010101;
assign LUT_4[52333] = 32'b11111111111111111001000110001101;
assign LUT_4[52334] = 32'b11111111111111111111010100111001;
assign LUT_4[52335] = 32'b11111111111111111000100000110001;
assign LUT_4[52336] = 32'b00000000000000000111011111010010;
assign LUT_4[52337] = 32'b00000000000000000000101011001010;
assign LUT_4[52338] = 32'b00000000000000000110111001110110;
assign LUT_4[52339] = 32'b00000000000000000000000101101110;
assign LUT_4[52340] = 32'b00000000000000000100011111101110;
assign LUT_4[52341] = 32'b11111111111111111101101011100110;
assign LUT_4[52342] = 32'b00000000000000000011111010010010;
assign LUT_4[52343] = 32'b11111111111111111101000110001010;
assign LUT_4[52344] = 32'b00000000000000000000101011100111;
assign LUT_4[52345] = 32'b11111111111111111001110111011111;
assign LUT_4[52346] = 32'b00000000000000000000000110001011;
assign LUT_4[52347] = 32'b11111111111111111001010010000011;
assign LUT_4[52348] = 32'b11111111111111111101101100000011;
assign LUT_4[52349] = 32'b11111111111111110110110111111011;
assign LUT_4[52350] = 32'b11111111111111111101000110100111;
assign LUT_4[52351] = 32'b11111111111111110110010010011111;
assign LUT_4[52352] = 32'b00000000000000001100100001010001;
assign LUT_4[52353] = 32'b00000000000000000101101101001001;
assign LUT_4[52354] = 32'b00000000000000001011111011110101;
assign LUT_4[52355] = 32'b00000000000000000101000111101101;
assign LUT_4[52356] = 32'b00000000000000001001100001101101;
assign LUT_4[52357] = 32'b00000000000000000010101101100101;
assign LUT_4[52358] = 32'b00000000000000001000111100010001;
assign LUT_4[52359] = 32'b00000000000000000010001000001001;
assign LUT_4[52360] = 32'b00000000000000000101101101100110;
assign LUT_4[52361] = 32'b11111111111111111110111001011110;
assign LUT_4[52362] = 32'b00000000000000000101001000001010;
assign LUT_4[52363] = 32'b11111111111111111110010100000010;
assign LUT_4[52364] = 32'b00000000000000000010101110000010;
assign LUT_4[52365] = 32'b11111111111111111011111001111010;
assign LUT_4[52366] = 32'b00000000000000000010001000100110;
assign LUT_4[52367] = 32'b11111111111111111011010100011110;
assign LUT_4[52368] = 32'b00000000000000001010010010111111;
assign LUT_4[52369] = 32'b00000000000000000011011110110111;
assign LUT_4[52370] = 32'b00000000000000001001101101100011;
assign LUT_4[52371] = 32'b00000000000000000010111001011011;
assign LUT_4[52372] = 32'b00000000000000000111010011011011;
assign LUT_4[52373] = 32'b00000000000000000000011111010011;
assign LUT_4[52374] = 32'b00000000000000000110101101111111;
assign LUT_4[52375] = 32'b11111111111111111111111001110111;
assign LUT_4[52376] = 32'b00000000000000000011011111010100;
assign LUT_4[52377] = 32'b11111111111111111100101011001100;
assign LUT_4[52378] = 32'b00000000000000000010111001111000;
assign LUT_4[52379] = 32'b11111111111111111100000101110000;
assign LUT_4[52380] = 32'b00000000000000000000011111110000;
assign LUT_4[52381] = 32'b11111111111111111001101011101000;
assign LUT_4[52382] = 32'b11111111111111111111111010010100;
assign LUT_4[52383] = 32'b11111111111111111001000110001100;
assign LUT_4[52384] = 32'b00000000000000001010111100011000;
assign LUT_4[52385] = 32'b00000000000000000100001000010000;
assign LUT_4[52386] = 32'b00000000000000001010010110111100;
assign LUT_4[52387] = 32'b00000000000000000011100010110100;
assign LUT_4[52388] = 32'b00000000000000000111111100110100;
assign LUT_4[52389] = 32'b00000000000000000001001000101100;
assign LUT_4[52390] = 32'b00000000000000000111010111011000;
assign LUT_4[52391] = 32'b00000000000000000000100011010000;
assign LUT_4[52392] = 32'b00000000000000000100001000101101;
assign LUT_4[52393] = 32'b11111111111111111101010100100101;
assign LUT_4[52394] = 32'b00000000000000000011100011010001;
assign LUT_4[52395] = 32'b11111111111111111100101111001001;
assign LUT_4[52396] = 32'b00000000000000000001001001001001;
assign LUT_4[52397] = 32'b11111111111111111010010101000001;
assign LUT_4[52398] = 32'b00000000000000000000100011101101;
assign LUT_4[52399] = 32'b11111111111111111001101111100101;
assign LUT_4[52400] = 32'b00000000000000001000101110000110;
assign LUT_4[52401] = 32'b00000000000000000001111001111110;
assign LUT_4[52402] = 32'b00000000000000001000001000101010;
assign LUT_4[52403] = 32'b00000000000000000001010100100010;
assign LUT_4[52404] = 32'b00000000000000000101101110100010;
assign LUT_4[52405] = 32'b11111111111111111110111010011010;
assign LUT_4[52406] = 32'b00000000000000000101001001000110;
assign LUT_4[52407] = 32'b11111111111111111110010100111110;
assign LUT_4[52408] = 32'b00000000000000000001111010011011;
assign LUT_4[52409] = 32'b11111111111111111011000110010011;
assign LUT_4[52410] = 32'b00000000000000000001010100111111;
assign LUT_4[52411] = 32'b11111111111111111010100000110111;
assign LUT_4[52412] = 32'b11111111111111111110111010110111;
assign LUT_4[52413] = 32'b11111111111111111000000110101111;
assign LUT_4[52414] = 32'b11111111111111111110010101011011;
assign LUT_4[52415] = 32'b11111111111111110111100001010011;
assign LUT_4[52416] = 32'b00000000000000001101111000100101;
assign LUT_4[52417] = 32'b00000000000000000111000100011101;
assign LUT_4[52418] = 32'b00000000000000001101010011001001;
assign LUT_4[52419] = 32'b00000000000000000110011111000001;
assign LUT_4[52420] = 32'b00000000000000001010111001000001;
assign LUT_4[52421] = 32'b00000000000000000100000100111001;
assign LUT_4[52422] = 32'b00000000000000001010010011100101;
assign LUT_4[52423] = 32'b00000000000000000011011111011101;
assign LUT_4[52424] = 32'b00000000000000000111000100111010;
assign LUT_4[52425] = 32'b00000000000000000000010000110010;
assign LUT_4[52426] = 32'b00000000000000000110011111011110;
assign LUT_4[52427] = 32'b11111111111111111111101011010110;
assign LUT_4[52428] = 32'b00000000000000000100000101010110;
assign LUT_4[52429] = 32'b11111111111111111101010001001110;
assign LUT_4[52430] = 32'b00000000000000000011011111111010;
assign LUT_4[52431] = 32'b11111111111111111100101011110010;
assign LUT_4[52432] = 32'b00000000000000001011101010010011;
assign LUT_4[52433] = 32'b00000000000000000100110110001011;
assign LUT_4[52434] = 32'b00000000000000001011000100110111;
assign LUT_4[52435] = 32'b00000000000000000100010000101111;
assign LUT_4[52436] = 32'b00000000000000001000101010101111;
assign LUT_4[52437] = 32'b00000000000000000001110110100111;
assign LUT_4[52438] = 32'b00000000000000001000000101010011;
assign LUT_4[52439] = 32'b00000000000000000001010001001011;
assign LUT_4[52440] = 32'b00000000000000000100110110101000;
assign LUT_4[52441] = 32'b11111111111111111110000010100000;
assign LUT_4[52442] = 32'b00000000000000000100010001001100;
assign LUT_4[52443] = 32'b11111111111111111101011101000100;
assign LUT_4[52444] = 32'b00000000000000000001110111000100;
assign LUT_4[52445] = 32'b11111111111111111011000010111100;
assign LUT_4[52446] = 32'b00000000000000000001010001101000;
assign LUT_4[52447] = 32'b11111111111111111010011101100000;
assign LUT_4[52448] = 32'b00000000000000001100010011101100;
assign LUT_4[52449] = 32'b00000000000000000101011111100100;
assign LUT_4[52450] = 32'b00000000000000001011101110010000;
assign LUT_4[52451] = 32'b00000000000000000100111010001000;
assign LUT_4[52452] = 32'b00000000000000001001010100001000;
assign LUT_4[52453] = 32'b00000000000000000010100000000000;
assign LUT_4[52454] = 32'b00000000000000001000101110101100;
assign LUT_4[52455] = 32'b00000000000000000001111010100100;
assign LUT_4[52456] = 32'b00000000000000000101100000000001;
assign LUT_4[52457] = 32'b11111111111111111110101011111001;
assign LUT_4[52458] = 32'b00000000000000000100111010100101;
assign LUT_4[52459] = 32'b11111111111111111110000110011101;
assign LUT_4[52460] = 32'b00000000000000000010100000011101;
assign LUT_4[52461] = 32'b11111111111111111011101100010101;
assign LUT_4[52462] = 32'b00000000000000000001111011000001;
assign LUT_4[52463] = 32'b11111111111111111011000110111001;
assign LUT_4[52464] = 32'b00000000000000001010000101011010;
assign LUT_4[52465] = 32'b00000000000000000011010001010010;
assign LUT_4[52466] = 32'b00000000000000001001011111111110;
assign LUT_4[52467] = 32'b00000000000000000010101011110110;
assign LUT_4[52468] = 32'b00000000000000000111000101110110;
assign LUT_4[52469] = 32'b00000000000000000000010001101110;
assign LUT_4[52470] = 32'b00000000000000000110100000011010;
assign LUT_4[52471] = 32'b11111111111111111111101100010010;
assign LUT_4[52472] = 32'b00000000000000000011010001101111;
assign LUT_4[52473] = 32'b11111111111111111100011101100111;
assign LUT_4[52474] = 32'b00000000000000000010101100010011;
assign LUT_4[52475] = 32'b11111111111111111011111000001011;
assign LUT_4[52476] = 32'b00000000000000000000010010001011;
assign LUT_4[52477] = 32'b11111111111111111001011110000011;
assign LUT_4[52478] = 32'b11111111111111111111101100101111;
assign LUT_4[52479] = 32'b11111111111111111000111000100111;
assign LUT_4[52480] = 32'b00000000000000001110110110101100;
assign LUT_4[52481] = 32'b00000000000000001000000010100100;
assign LUT_4[52482] = 32'b00000000000000001110010001010000;
assign LUT_4[52483] = 32'b00000000000000000111011101001000;
assign LUT_4[52484] = 32'b00000000000000001011110111001000;
assign LUT_4[52485] = 32'b00000000000000000101000011000000;
assign LUT_4[52486] = 32'b00000000000000001011010001101100;
assign LUT_4[52487] = 32'b00000000000000000100011101100100;
assign LUT_4[52488] = 32'b00000000000000001000000011000001;
assign LUT_4[52489] = 32'b00000000000000000001001110111001;
assign LUT_4[52490] = 32'b00000000000000000111011101100101;
assign LUT_4[52491] = 32'b00000000000000000000101001011101;
assign LUT_4[52492] = 32'b00000000000000000101000011011101;
assign LUT_4[52493] = 32'b11111111111111111110001111010101;
assign LUT_4[52494] = 32'b00000000000000000100011110000001;
assign LUT_4[52495] = 32'b11111111111111111101101001111001;
assign LUT_4[52496] = 32'b00000000000000001100101000011010;
assign LUT_4[52497] = 32'b00000000000000000101110100010010;
assign LUT_4[52498] = 32'b00000000000000001100000010111110;
assign LUT_4[52499] = 32'b00000000000000000101001110110110;
assign LUT_4[52500] = 32'b00000000000000001001101000110110;
assign LUT_4[52501] = 32'b00000000000000000010110100101110;
assign LUT_4[52502] = 32'b00000000000000001001000011011010;
assign LUT_4[52503] = 32'b00000000000000000010001111010010;
assign LUT_4[52504] = 32'b00000000000000000101110100101111;
assign LUT_4[52505] = 32'b11111111111111111111000000100111;
assign LUT_4[52506] = 32'b00000000000000000101001111010011;
assign LUT_4[52507] = 32'b11111111111111111110011011001011;
assign LUT_4[52508] = 32'b00000000000000000010110101001011;
assign LUT_4[52509] = 32'b11111111111111111100000001000011;
assign LUT_4[52510] = 32'b00000000000000000010001111101111;
assign LUT_4[52511] = 32'b11111111111111111011011011100111;
assign LUT_4[52512] = 32'b00000000000000001101010001110011;
assign LUT_4[52513] = 32'b00000000000000000110011101101011;
assign LUT_4[52514] = 32'b00000000000000001100101100010111;
assign LUT_4[52515] = 32'b00000000000000000101111000001111;
assign LUT_4[52516] = 32'b00000000000000001010010010001111;
assign LUT_4[52517] = 32'b00000000000000000011011110000111;
assign LUT_4[52518] = 32'b00000000000000001001101100110011;
assign LUT_4[52519] = 32'b00000000000000000010111000101011;
assign LUT_4[52520] = 32'b00000000000000000110011110001000;
assign LUT_4[52521] = 32'b11111111111111111111101010000000;
assign LUT_4[52522] = 32'b00000000000000000101111000101100;
assign LUT_4[52523] = 32'b11111111111111111111000100100100;
assign LUT_4[52524] = 32'b00000000000000000011011110100100;
assign LUT_4[52525] = 32'b11111111111111111100101010011100;
assign LUT_4[52526] = 32'b00000000000000000010111001001000;
assign LUT_4[52527] = 32'b11111111111111111100000101000000;
assign LUT_4[52528] = 32'b00000000000000001011000011100001;
assign LUT_4[52529] = 32'b00000000000000000100001111011001;
assign LUT_4[52530] = 32'b00000000000000001010011110000101;
assign LUT_4[52531] = 32'b00000000000000000011101001111101;
assign LUT_4[52532] = 32'b00000000000000001000000011111101;
assign LUT_4[52533] = 32'b00000000000000000001001111110101;
assign LUT_4[52534] = 32'b00000000000000000111011110100001;
assign LUT_4[52535] = 32'b00000000000000000000101010011001;
assign LUT_4[52536] = 32'b00000000000000000100001111110110;
assign LUT_4[52537] = 32'b11111111111111111101011011101110;
assign LUT_4[52538] = 32'b00000000000000000011101010011010;
assign LUT_4[52539] = 32'b11111111111111111100110110010010;
assign LUT_4[52540] = 32'b00000000000000000001010000010010;
assign LUT_4[52541] = 32'b11111111111111111010011100001010;
assign LUT_4[52542] = 32'b00000000000000000000101010110110;
assign LUT_4[52543] = 32'b11111111111111111001110110101110;
assign LUT_4[52544] = 32'b00000000000000010000001110000000;
assign LUT_4[52545] = 32'b00000000000000001001011001111000;
assign LUT_4[52546] = 32'b00000000000000001111101000100100;
assign LUT_4[52547] = 32'b00000000000000001000110100011100;
assign LUT_4[52548] = 32'b00000000000000001101001110011100;
assign LUT_4[52549] = 32'b00000000000000000110011010010100;
assign LUT_4[52550] = 32'b00000000000000001100101001000000;
assign LUT_4[52551] = 32'b00000000000000000101110100111000;
assign LUT_4[52552] = 32'b00000000000000001001011010010101;
assign LUT_4[52553] = 32'b00000000000000000010100110001101;
assign LUT_4[52554] = 32'b00000000000000001000110100111001;
assign LUT_4[52555] = 32'b00000000000000000010000000110001;
assign LUT_4[52556] = 32'b00000000000000000110011010110001;
assign LUT_4[52557] = 32'b11111111111111111111100110101001;
assign LUT_4[52558] = 32'b00000000000000000101110101010101;
assign LUT_4[52559] = 32'b11111111111111111111000001001101;
assign LUT_4[52560] = 32'b00000000000000001101111111101110;
assign LUT_4[52561] = 32'b00000000000000000111001011100110;
assign LUT_4[52562] = 32'b00000000000000001101011010010010;
assign LUT_4[52563] = 32'b00000000000000000110100110001010;
assign LUT_4[52564] = 32'b00000000000000001011000000001010;
assign LUT_4[52565] = 32'b00000000000000000100001100000010;
assign LUT_4[52566] = 32'b00000000000000001010011010101110;
assign LUT_4[52567] = 32'b00000000000000000011100110100110;
assign LUT_4[52568] = 32'b00000000000000000111001100000011;
assign LUT_4[52569] = 32'b00000000000000000000010111111011;
assign LUT_4[52570] = 32'b00000000000000000110100110100111;
assign LUT_4[52571] = 32'b11111111111111111111110010011111;
assign LUT_4[52572] = 32'b00000000000000000100001100011111;
assign LUT_4[52573] = 32'b11111111111111111101011000010111;
assign LUT_4[52574] = 32'b00000000000000000011100111000011;
assign LUT_4[52575] = 32'b11111111111111111100110010111011;
assign LUT_4[52576] = 32'b00000000000000001110101001000111;
assign LUT_4[52577] = 32'b00000000000000000111110100111111;
assign LUT_4[52578] = 32'b00000000000000001110000011101011;
assign LUT_4[52579] = 32'b00000000000000000111001111100011;
assign LUT_4[52580] = 32'b00000000000000001011101001100011;
assign LUT_4[52581] = 32'b00000000000000000100110101011011;
assign LUT_4[52582] = 32'b00000000000000001011000100000111;
assign LUT_4[52583] = 32'b00000000000000000100001111111111;
assign LUT_4[52584] = 32'b00000000000000000111110101011100;
assign LUT_4[52585] = 32'b00000000000000000001000001010100;
assign LUT_4[52586] = 32'b00000000000000000111010000000000;
assign LUT_4[52587] = 32'b00000000000000000000011011111000;
assign LUT_4[52588] = 32'b00000000000000000100110101111000;
assign LUT_4[52589] = 32'b11111111111111111110000001110000;
assign LUT_4[52590] = 32'b00000000000000000100010000011100;
assign LUT_4[52591] = 32'b11111111111111111101011100010100;
assign LUT_4[52592] = 32'b00000000000000001100011010110101;
assign LUT_4[52593] = 32'b00000000000000000101100110101101;
assign LUT_4[52594] = 32'b00000000000000001011110101011001;
assign LUT_4[52595] = 32'b00000000000000000101000001010001;
assign LUT_4[52596] = 32'b00000000000000001001011011010001;
assign LUT_4[52597] = 32'b00000000000000000010100111001001;
assign LUT_4[52598] = 32'b00000000000000001000110101110101;
assign LUT_4[52599] = 32'b00000000000000000010000001101101;
assign LUT_4[52600] = 32'b00000000000000000101100111001010;
assign LUT_4[52601] = 32'b11111111111111111110110011000010;
assign LUT_4[52602] = 32'b00000000000000000101000001101110;
assign LUT_4[52603] = 32'b11111111111111111110001101100110;
assign LUT_4[52604] = 32'b00000000000000000010100111100110;
assign LUT_4[52605] = 32'b11111111111111111011110011011110;
assign LUT_4[52606] = 32'b00000000000000000010000010001010;
assign LUT_4[52607] = 32'b11111111111111111011001110000010;
assign LUT_4[52608] = 32'b00000000000000010001011100110100;
assign LUT_4[52609] = 32'b00000000000000001010101000101100;
assign LUT_4[52610] = 32'b00000000000000010000110111011000;
assign LUT_4[52611] = 32'b00000000000000001010000011010000;
assign LUT_4[52612] = 32'b00000000000000001110011101010000;
assign LUT_4[52613] = 32'b00000000000000000111101001001000;
assign LUT_4[52614] = 32'b00000000000000001101110111110100;
assign LUT_4[52615] = 32'b00000000000000000111000011101100;
assign LUT_4[52616] = 32'b00000000000000001010101001001001;
assign LUT_4[52617] = 32'b00000000000000000011110101000001;
assign LUT_4[52618] = 32'b00000000000000001010000011101101;
assign LUT_4[52619] = 32'b00000000000000000011001111100101;
assign LUT_4[52620] = 32'b00000000000000000111101001100101;
assign LUT_4[52621] = 32'b00000000000000000000110101011101;
assign LUT_4[52622] = 32'b00000000000000000111000100001001;
assign LUT_4[52623] = 32'b00000000000000000000010000000001;
assign LUT_4[52624] = 32'b00000000000000001111001110100010;
assign LUT_4[52625] = 32'b00000000000000001000011010011010;
assign LUT_4[52626] = 32'b00000000000000001110101001000110;
assign LUT_4[52627] = 32'b00000000000000000111110100111110;
assign LUT_4[52628] = 32'b00000000000000001100001110111110;
assign LUT_4[52629] = 32'b00000000000000000101011010110110;
assign LUT_4[52630] = 32'b00000000000000001011101001100010;
assign LUT_4[52631] = 32'b00000000000000000100110101011010;
assign LUT_4[52632] = 32'b00000000000000001000011010110111;
assign LUT_4[52633] = 32'b00000000000000000001100110101111;
assign LUT_4[52634] = 32'b00000000000000000111110101011011;
assign LUT_4[52635] = 32'b00000000000000000001000001010011;
assign LUT_4[52636] = 32'b00000000000000000101011011010011;
assign LUT_4[52637] = 32'b11111111111111111110100111001011;
assign LUT_4[52638] = 32'b00000000000000000100110101110111;
assign LUT_4[52639] = 32'b11111111111111111110000001101111;
assign LUT_4[52640] = 32'b00000000000000001111110111111011;
assign LUT_4[52641] = 32'b00000000000000001001000011110011;
assign LUT_4[52642] = 32'b00000000000000001111010010011111;
assign LUT_4[52643] = 32'b00000000000000001000011110010111;
assign LUT_4[52644] = 32'b00000000000000001100111000010111;
assign LUT_4[52645] = 32'b00000000000000000110000100001111;
assign LUT_4[52646] = 32'b00000000000000001100010010111011;
assign LUT_4[52647] = 32'b00000000000000000101011110110011;
assign LUT_4[52648] = 32'b00000000000000001001000100010000;
assign LUT_4[52649] = 32'b00000000000000000010010000001000;
assign LUT_4[52650] = 32'b00000000000000001000011110110100;
assign LUT_4[52651] = 32'b00000000000000000001101010101100;
assign LUT_4[52652] = 32'b00000000000000000110000100101100;
assign LUT_4[52653] = 32'b11111111111111111111010000100100;
assign LUT_4[52654] = 32'b00000000000000000101011111010000;
assign LUT_4[52655] = 32'b11111111111111111110101011001000;
assign LUT_4[52656] = 32'b00000000000000001101101001101001;
assign LUT_4[52657] = 32'b00000000000000000110110101100001;
assign LUT_4[52658] = 32'b00000000000000001101000100001101;
assign LUT_4[52659] = 32'b00000000000000000110010000000101;
assign LUT_4[52660] = 32'b00000000000000001010101010000101;
assign LUT_4[52661] = 32'b00000000000000000011110101111101;
assign LUT_4[52662] = 32'b00000000000000001010000100101001;
assign LUT_4[52663] = 32'b00000000000000000011010000100001;
assign LUT_4[52664] = 32'b00000000000000000110110101111110;
assign LUT_4[52665] = 32'b00000000000000000000000001110110;
assign LUT_4[52666] = 32'b00000000000000000110010000100010;
assign LUT_4[52667] = 32'b11111111111111111111011100011010;
assign LUT_4[52668] = 32'b00000000000000000011110110011010;
assign LUT_4[52669] = 32'b11111111111111111101000010010010;
assign LUT_4[52670] = 32'b00000000000000000011010000111110;
assign LUT_4[52671] = 32'b11111111111111111100011100110110;
assign LUT_4[52672] = 32'b00000000000000010010110100001000;
assign LUT_4[52673] = 32'b00000000000000001100000000000000;
assign LUT_4[52674] = 32'b00000000000000010010001110101100;
assign LUT_4[52675] = 32'b00000000000000001011011010100100;
assign LUT_4[52676] = 32'b00000000000000001111110100100100;
assign LUT_4[52677] = 32'b00000000000000001001000000011100;
assign LUT_4[52678] = 32'b00000000000000001111001111001000;
assign LUT_4[52679] = 32'b00000000000000001000011011000000;
assign LUT_4[52680] = 32'b00000000000000001100000000011101;
assign LUT_4[52681] = 32'b00000000000000000101001100010101;
assign LUT_4[52682] = 32'b00000000000000001011011011000001;
assign LUT_4[52683] = 32'b00000000000000000100100110111001;
assign LUT_4[52684] = 32'b00000000000000001001000000111001;
assign LUT_4[52685] = 32'b00000000000000000010001100110001;
assign LUT_4[52686] = 32'b00000000000000001000011011011101;
assign LUT_4[52687] = 32'b00000000000000000001100111010101;
assign LUT_4[52688] = 32'b00000000000000010000100101110110;
assign LUT_4[52689] = 32'b00000000000000001001110001101110;
assign LUT_4[52690] = 32'b00000000000000010000000000011010;
assign LUT_4[52691] = 32'b00000000000000001001001100010010;
assign LUT_4[52692] = 32'b00000000000000001101100110010010;
assign LUT_4[52693] = 32'b00000000000000000110110010001010;
assign LUT_4[52694] = 32'b00000000000000001101000000110110;
assign LUT_4[52695] = 32'b00000000000000000110001100101110;
assign LUT_4[52696] = 32'b00000000000000001001110010001011;
assign LUT_4[52697] = 32'b00000000000000000010111110000011;
assign LUT_4[52698] = 32'b00000000000000001001001100101111;
assign LUT_4[52699] = 32'b00000000000000000010011000100111;
assign LUT_4[52700] = 32'b00000000000000000110110010100111;
assign LUT_4[52701] = 32'b11111111111111111111111110011111;
assign LUT_4[52702] = 32'b00000000000000000110001101001011;
assign LUT_4[52703] = 32'b11111111111111111111011001000011;
assign LUT_4[52704] = 32'b00000000000000010001001111001111;
assign LUT_4[52705] = 32'b00000000000000001010011011000111;
assign LUT_4[52706] = 32'b00000000000000010000101001110011;
assign LUT_4[52707] = 32'b00000000000000001001110101101011;
assign LUT_4[52708] = 32'b00000000000000001110001111101011;
assign LUT_4[52709] = 32'b00000000000000000111011011100011;
assign LUT_4[52710] = 32'b00000000000000001101101010001111;
assign LUT_4[52711] = 32'b00000000000000000110110110000111;
assign LUT_4[52712] = 32'b00000000000000001010011011100100;
assign LUT_4[52713] = 32'b00000000000000000011100111011100;
assign LUT_4[52714] = 32'b00000000000000001001110110001000;
assign LUT_4[52715] = 32'b00000000000000000011000010000000;
assign LUT_4[52716] = 32'b00000000000000000111011100000000;
assign LUT_4[52717] = 32'b00000000000000000000100111111000;
assign LUT_4[52718] = 32'b00000000000000000110110110100100;
assign LUT_4[52719] = 32'b00000000000000000000000010011100;
assign LUT_4[52720] = 32'b00000000000000001111000000111101;
assign LUT_4[52721] = 32'b00000000000000001000001100110101;
assign LUT_4[52722] = 32'b00000000000000001110011011100001;
assign LUT_4[52723] = 32'b00000000000000000111100111011001;
assign LUT_4[52724] = 32'b00000000000000001100000001011001;
assign LUT_4[52725] = 32'b00000000000000000101001101010001;
assign LUT_4[52726] = 32'b00000000000000001011011011111101;
assign LUT_4[52727] = 32'b00000000000000000100100111110101;
assign LUT_4[52728] = 32'b00000000000000001000001101010010;
assign LUT_4[52729] = 32'b00000000000000000001011001001010;
assign LUT_4[52730] = 32'b00000000000000000111100111110110;
assign LUT_4[52731] = 32'b00000000000000000000110011101110;
assign LUT_4[52732] = 32'b00000000000000000101001101101110;
assign LUT_4[52733] = 32'b11111111111111111110011001100110;
assign LUT_4[52734] = 32'b00000000000000000100101000010010;
assign LUT_4[52735] = 32'b11111111111111111101110100001010;
assign LUT_4[52736] = 32'b00000000000000001000111111010001;
assign LUT_4[52737] = 32'b00000000000000000010001011001001;
assign LUT_4[52738] = 32'b00000000000000001000011001110101;
assign LUT_4[52739] = 32'b00000000000000000001100101101101;
assign LUT_4[52740] = 32'b00000000000000000101111111101101;
assign LUT_4[52741] = 32'b11111111111111111111001011100101;
assign LUT_4[52742] = 32'b00000000000000000101011010010001;
assign LUT_4[52743] = 32'b11111111111111111110100110001001;
assign LUT_4[52744] = 32'b00000000000000000010001011100110;
assign LUT_4[52745] = 32'b11111111111111111011010111011110;
assign LUT_4[52746] = 32'b00000000000000000001100110001010;
assign LUT_4[52747] = 32'b11111111111111111010110010000010;
assign LUT_4[52748] = 32'b11111111111111111111001100000010;
assign LUT_4[52749] = 32'b11111111111111111000010111111010;
assign LUT_4[52750] = 32'b11111111111111111110100110100110;
assign LUT_4[52751] = 32'b11111111111111110111110010011110;
assign LUT_4[52752] = 32'b00000000000000000110110000111111;
assign LUT_4[52753] = 32'b11111111111111111111111100110111;
assign LUT_4[52754] = 32'b00000000000000000110001011100011;
assign LUT_4[52755] = 32'b11111111111111111111010111011011;
assign LUT_4[52756] = 32'b00000000000000000011110001011011;
assign LUT_4[52757] = 32'b11111111111111111100111101010011;
assign LUT_4[52758] = 32'b00000000000000000011001011111111;
assign LUT_4[52759] = 32'b11111111111111111100010111110111;
assign LUT_4[52760] = 32'b11111111111111111111111101010100;
assign LUT_4[52761] = 32'b11111111111111111001001001001100;
assign LUT_4[52762] = 32'b11111111111111111111010111111000;
assign LUT_4[52763] = 32'b11111111111111111000100011110000;
assign LUT_4[52764] = 32'b11111111111111111100111101110000;
assign LUT_4[52765] = 32'b11111111111111110110001001101000;
assign LUT_4[52766] = 32'b11111111111111111100011000010100;
assign LUT_4[52767] = 32'b11111111111111110101100100001100;
assign LUT_4[52768] = 32'b00000000000000000111011010011000;
assign LUT_4[52769] = 32'b00000000000000000000100110010000;
assign LUT_4[52770] = 32'b00000000000000000110110100111100;
assign LUT_4[52771] = 32'b00000000000000000000000000110100;
assign LUT_4[52772] = 32'b00000000000000000100011010110100;
assign LUT_4[52773] = 32'b11111111111111111101100110101100;
assign LUT_4[52774] = 32'b00000000000000000011110101011000;
assign LUT_4[52775] = 32'b11111111111111111101000001010000;
assign LUT_4[52776] = 32'b00000000000000000000100110101101;
assign LUT_4[52777] = 32'b11111111111111111001110010100101;
assign LUT_4[52778] = 32'b00000000000000000000000001010001;
assign LUT_4[52779] = 32'b11111111111111111001001101001001;
assign LUT_4[52780] = 32'b11111111111111111101100111001001;
assign LUT_4[52781] = 32'b11111111111111110110110011000001;
assign LUT_4[52782] = 32'b11111111111111111101000001101101;
assign LUT_4[52783] = 32'b11111111111111110110001101100101;
assign LUT_4[52784] = 32'b00000000000000000101001100000110;
assign LUT_4[52785] = 32'b11111111111111111110010111111110;
assign LUT_4[52786] = 32'b00000000000000000100100110101010;
assign LUT_4[52787] = 32'b11111111111111111101110010100010;
assign LUT_4[52788] = 32'b00000000000000000010001100100010;
assign LUT_4[52789] = 32'b11111111111111111011011000011010;
assign LUT_4[52790] = 32'b00000000000000000001100111000110;
assign LUT_4[52791] = 32'b11111111111111111010110010111110;
assign LUT_4[52792] = 32'b11111111111111111110011000011011;
assign LUT_4[52793] = 32'b11111111111111110111100100010011;
assign LUT_4[52794] = 32'b11111111111111111101110010111111;
assign LUT_4[52795] = 32'b11111111111111110110111110110111;
assign LUT_4[52796] = 32'b11111111111111111011011000110111;
assign LUT_4[52797] = 32'b11111111111111110100100100101111;
assign LUT_4[52798] = 32'b11111111111111111010110011011011;
assign LUT_4[52799] = 32'b11111111111111110011111111010011;
assign LUT_4[52800] = 32'b00000000000000001010010110100101;
assign LUT_4[52801] = 32'b00000000000000000011100010011101;
assign LUT_4[52802] = 32'b00000000000000001001110001001001;
assign LUT_4[52803] = 32'b00000000000000000010111101000001;
assign LUT_4[52804] = 32'b00000000000000000111010111000001;
assign LUT_4[52805] = 32'b00000000000000000000100010111001;
assign LUT_4[52806] = 32'b00000000000000000110110001100101;
assign LUT_4[52807] = 32'b11111111111111111111111101011101;
assign LUT_4[52808] = 32'b00000000000000000011100010111010;
assign LUT_4[52809] = 32'b11111111111111111100101110110010;
assign LUT_4[52810] = 32'b00000000000000000010111101011110;
assign LUT_4[52811] = 32'b11111111111111111100001001010110;
assign LUT_4[52812] = 32'b00000000000000000000100011010110;
assign LUT_4[52813] = 32'b11111111111111111001101111001110;
assign LUT_4[52814] = 32'b11111111111111111111111101111010;
assign LUT_4[52815] = 32'b11111111111111111001001001110010;
assign LUT_4[52816] = 32'b00000000000000001000001000010011;
assign LUT_4[52817] = 32'b00000000000000000001010100001011;
assign LUT_4[52818] = 32'b00000000000000000111100010110111;
assign LUT_4[52819] = 32'b00000000000000000000101110101111;
assign LUT_4[52820] = 32'b00000000000000000101001000101111;
assign LUT_4[52821] = 32'b11111111111111111110010100100111;
assign LUT_4[52822] = 32'b00000000000000000100100011010011;
assign LUT_4[52823] = 32'b11111111111111111101101111001011;
assign LUT_4[52824] = 32'b00000000000000000001010100101000;
assign LUT_4[52825] = 32'b11111111111111111010100000100000;
assign LUT_4[52826] = 32'b00000000000000000000101111001100;
assign LUT_4[52827] = 32'b11111111111111111001111011000100;
assign LUT_4[52828] = 32'b11111111111111111110010101000100;
assign LUT_4[52829] = 32'b11111111111111110111100000111100;
assign LUT_4[52830] = 32'b11111111111111111101101111101000;
assign LUT_4[52831] = 32'b11111111111111110110111011100000;
assign LUT_4[52832] = 32'b00000000000000001000110001101100;
assign LUT_4[52833] = 32'b00000000000000000001111101100100;
assign LUT_4[52834] = 32'b00000000000000001000001100010000;
assign LUT_4[52835] = 32'b00000000000000000001011000001000;
assign LUT_4[52836] = 32'b00000000000000000101110010001000;
assign LUT_4[52837] = 32'b11111111111111111110111110000000;
assign LUT_4[52838] = 32'b00000000000000000101001100101100;
assign LUT_4[52839] = 32'b11111111111111111110011000100100;
assign LUT_4[52840] = 32'b00000000000000000001111110000001;
assign LUT_4[52841] = 32'b11111111111111111011001001111001;
assign LUT_4[52842] = 32'b00000000000000000001011000100101;
assign LUT_4[52843] = 32'b11111111111111111010100100011101;
assign LUT_4[52844] = 32'b11111111111111111110111110011101;
assign LUT_4[52845] = 32'b11111111111111111000001010010101;
assign LUT_4[52846] = 32'b11111111111111111110011001000001;
assign LUT_4[52847] = 32'b11111111111111110111100100111001;
assign LUT_4[52848] = 32'b00000000000000000110100011011010;
assign LUT_4[52849] = 32'b11111111111111111111101111010010;
assign LUT_4[52850] = 32'b00000000000000000101111101111110;
assign LUT_4[52851] = 32'b11111111111111111111001001110110;
assign LUT_4[52852] = 32'b00000000000000000011100011110110;
assign LUT_4[52853] = 32'b11111111111111111100101111101110;
assign LUT_4[52854] = 32'b00000000000000000010111110011010;
assign LUT_4[52855] = 32'b11111111111111111100001010010010;
assign LUT_4[52856] = 32'b11111111111111111111101111101111;
assign LUT_4[52857] = 32'b11111111111111111000111011100111;
assign LUT_4[52858] = 32'b11111111111111111111001010010011;
assign LUT_4[52859] = 32'b11111111111111111000010110001011;
assign LUT_4[52860] = 32'b11111111111111111100110000001011;
assign LUT_4[52861] = 32'b11111111111111110101111100000011;
assign LUT_4[52862] = 32'b11111111111111111100001010101111;
assign LUT_4[52863] = 32'b11111111111111110101010110100111;
assign LUT_4[52864] = 32'b00000000000000001011100101011001;
assign LUT_4[52865] = 32'b00000000000000000100110001010001;
assign LUT_4[52866] = 32'b00000000000000001010111111111101;
assign LUT_4[52867] = 32'b00000000000000000100001011110101;
assign LUT_4[52868] = 32'b00000000000000001000100101110101;
assign LUT_4[52869] = 32'b00000000000000000001110001101101;
assign LUT_4[52870] = 32'b00000000000000001000000000011001;
assign LUT_4[52871] = 32'b00000000000000000001001100010001;
assign LUT_4[52872] = 32'b00000000000000000100110001101110;
assign LUT_4[52873] = 32'b11111111111111111101111101100110;
assign LUT_4[52874] = 32'b00000000000000000100001100010010;
assign LUT_4[52875] = 32'b11111111111111111101011000001010;
assign LUT_4[52876] = 32'b00000000000000000001110010001010;
assign LUT_4[52877] = 32'b11111111111111111010111110000010;
assign LUT_4[52878] = 32'b00000000000000000001001100101110;
assign LUT_4[52879] = 32'b11111111111111111010011000100110;
assign LUT_4[52880] = 32'b00000000000000001001010111000111;
assign LUT_4[52881] = 32'b00000000000000000010100010111111;
assign LUT_4[52882] = 32'b00000000000000001000110001101011;
assign LUT_4[52883] = 32'b00000000000000000001111101100011;
assign LUT_4[52884] = 32'b00000000000000000110010111100011;
assign LUT_4[52885] = 32'b11111111111111111111100011011011;
assign LUT_4[52886] = 32'b00000000000000000101110010000111;
assign LUT_4[52887] = 32'b11111111111111111110111101111111;
assign LUT_4[52888] = 32'b00000000000000000010100011011100;
assign LUT_4[52889] = 32'b11111111111111111011101111010100;
assign LUT_4[52890] = 32'b00000000000000000001111110000000;
assign LUT_4[52891] = 32'b11111111111111111011001001111000;
assign LUT_4[52892] = 32'b11111111111111111111100011111000;
assign LUT_4[52893] = 32'b11111111111111111000101111110000;
assign LUT_4[52894] = 32'b11111111111111111110111110011100;
assign LUT_4[52895] = 32'b11111111111111111000001010010100;
assign LUT_4[52896] = 32'b00000000000000001010000000100000;
assign LUT_4[52897] = 32'b00000000000000000011001100011000;
assign LUT_4[52898] = 32'b00000000000000001001011011000100;
assign LUT_4[52899] = 32'b00000000000000000010100110111100;
assign LUT_4[52900] = 32'b00000000000000000111000000111100;
assign LUT_4[52901] = 32'b00000000000000000000001100110100;
assign LUT_4[52902] = 32'b00000000000000000110011011100000;
assign LUT_4[52903] = 32'b11111111111111111111100111011000;
assign LUT_4[52904] = 32'b00000000000000000011001100110101;
assign LUT_4[52905] = 32'b11111111111111111100011000101101;
assign LUT_4[52906] = 32'b00000000000000000010100111011001;
assign LUT_4[52907] = 32'b11111111111111111011110011010001;
assign LUT_4[52908] = 32'b00000000000000000000001101010001;
assign LUT_4[52909] = 32'b11111111111111111001011001001001;
assign LUT_4[52910] = 32'b11111111111111111111100111110101;
assign LUT_4[52911] = 32'b11111111111111111000110011101101;
assign LUT_4[52912] = 32'b00000000000000000111110010001110;
assign LUT_4[52913] = 32'b00000000000000000000111110000110;
assign LUT_4[52914] = 32'b00000000000000000111001100110010;
assign LUT_4[52915] = 32'b00000000000000000000011000101010;
assign LUT_4[52916] = 32'b00000000000000000100110010101010;
assign LUT_4[52917] = 32'b11111111111111111101111110100010;
assign LUT_4[52918] = 32'b00000000000000000100001101001110;
assign LUT_4[52919] = 32'b11111111111111111101011001000110;
assign LUT_4[52920] = 32'b00000000000000000000111110100011;
assign LUT_4[52921] = 32'b11111111111111111010001010011011;
assign LUT_4[52922] = 32'b00000000000000000000011001000111;
assign LUT_4[52923] = 32'b11111111111111111001100100111111;
assign LUT_4[52924] = 32'b11111111111111111101111110111111;
assign LUT_4[52925] = 32'b11111111111111110111001010110111;
assign LUT_4[52926] = 32'b11111111111111111101011001100011;
assign LUT_4[52927] = 32'b11111111111111110110100101011011;
assign LUT_4[52928] = 32'b00000000000000001100111100101101;
assign LUT_4[52929] = 32'b00000000000000000110001000100101;
assign LUT_4[52930] = 32'b00000000000000001100010111010001;
assign LUT_4[52931] = 32'b00000000000000000101100011001001;
assign LUT_4[52932] = 32'b00000000000000001001111101001001;
assign LUT_4[52933] = 32'b00000000000000000011001001000001;
assign LUT_4[52934] = 32'b00000000000000001001010111101101;
assign LUT_4[52935] = 32'b00000000000000000010100011100101;
assign LUT_4[52936] = 32'b00000000000000000110001001000010;
assign LUT_4[52937] = 32'b11111111111111111111010100111010;
assign LUT_4[52938] = 32'b00000000000000000101100011100110;
assign LUT_4[52939] = 32'b11111111111111111110101111011110;
assign LUT_4[52940] = 32'b00000000000000000011001001011110;
assign LUT_4[52941] = 32'b11111111111111111100010101010110;
assign LUT_4[52942] = 32'b00000000000000000010100100000010;
assign LUT_4[52943] = 32'b11111111111111111011101111111010;
assign LUT_4[52944] = 32'b00000000000000001010101110011011;
assign LUT_4[52945] = 32'b00000000000000000011111010010011;
assign LUT_4[52946] = 32'b00000000000000001010001000111111;
assign LUT_4[52947] = 32'b00000000000000000011010100110111;
assign LUT_4[52948] = 32'b00000000000000000111101110110111;
assign LUT_4[52949] = 32'b00000000000000000000111010101111;
assign LUT_4[52950] = 32'b00000000000000000111001001011011;
assign LUT_4[52951] = 32'b00000000000000000000010101010011;
assign LUT_4[52952] = 32'b00000000000000000011111010110000;
assign LUT_4[52953] = 32'b11111111111111111101000110101000;
assign LUT_4[52954] = 32'b00000000000000000011010101010100;
assign LUT_4[52955] = 32'b11111111111111111100100001001100;
assign LUT_4[52956] = 32'b00000000000000000000111011001100;
assign LUT_4[52957] = 32'b11111111111111111010000111000100;
assign LUT_4[52958] = 32'b00000000000000000000010101110000;
assign LUT_4[52959] = 32'b11111111111111111001100001101000;
assign LUT_4[52960] = 32'b00000000000000001011010111110100;
assign LUT_4[52961] = 32'b00000000000000000100100011101100;
assign LUT_4[52962] = 32'b00000000000000001010110010011000;
assign LUT_4[52963] = 32'b00000000000000000011111110010000;
assign LUT_4[52964] = 32'b00000000000000001000011000010000;
assign LUT_4[52965] = 32'b00000000000000000001100100001000;
assign LUT_4[52966] = 32'b00000000000000000111110010110100;
assign LUT_4[52967] = 32'b00000000000000000000111110101100;
assign LUT_4[52968] = 32'b00000000000000000100100100001001;
assign LUT_4[52969] = 32'b11111111111111111101110000000001;
assign LUT_4[52970] = 32'b00000000000000000011111110101101;
assign LUT_4[52971] = 32'b11111111111111111101001010100101;
assign LUT_4[52972] = 32'b00000000000000000001100100100101;
assign LUT_4[52973] = 32'b11111111111111111010110000011101;
assign LUT_4[52974] = 32'b00000000000000000000111111001001;
assign LUT_4[52975] = 32'b11111111111111111010001011000001;
assign LUT_4[52976] = 32'b00000000000000001001001001100010;
assign LUT_4[52977] = 32'b00000000000000000010010101011010;
assign LUT_4[52978] = 32'b00000000000000001000100100000110;
assign LUT_4[52979] = 32'b00000000000000000001101111111110;
assign LUT_4[52980] = 32'b00000000000000000110001001111110;
assign LUT_4[52981] = 32'b11111111111111111111010101110110;
assign LUT_4[52982] = 32'b00000000000000000101100100100010;
assign LUT_4[52983] = 32'b11111111111111111110110000011010;
assign LUT_4[52984] = 32'b00000000000000000010010101110111;
assign LUT_4[52985] = 32'b11111111111111111011100001101111;
assign LUT_4[52986] = 32'b00000000000000000001110000011011;
assign LUT_4[52987] = 32'b11111111111111111010111100010011;
assign LUT_4[52988] = 32'b11111111111111111111010110010011;
assign LUT_4[52989] = 32'b11111111111111111000100010001011;
assign LUT_4[52990] = 32'b11111111111111111110110000110111;
assign LUT_4[52991] = 32'b11111111111111110111111100101111;
assign LUT_4[52992] = 32'b00000000000000001101111010110100;
assign LUT_4[52993] = 32'b00000000000000000111000110101100;
assign LUT_4[52994] = 32'b00000000000000001101010101011000;
assign LUT_4[52995] = 32'b00000000000000000110100001010000;
assign LUT_4[52996] = 32'b00000000000000001010111011010000;
assign LUT_4[52997] = 32'b00000000000000000100000111001000;
assign LUT_4[52998] = 32'b00000000000000001010010101110100;
assign LUT_4[52999] = 32'b00000000000000000011100001101100;
assign LUT_4[53000] = 32'b00000000000000000111000111001001;
assign LUT_4[53001] = 32'b00000000000000000000010011000001;
assign LUT_4[53002] = 32'b00000000000000000110100001101101;
assign LUT_4[53003] = 32'b11111111111111111111101101100101;
assign LUT_4[53004] = 32'b00000000000000000100000111100101;
assign LUT_4[53005] = 32'b11111111111111111101010011011101;
assign LUT_4[53006] = 32'b00000000000000000011100010001001;
assign LUT_4[53007] = 32'b11111111111111111100101110000001;
assign LUT_4[53008] = 32'b00000000000000001011101100100010;
assign LUT_4[53009] = 32'b00000000000000000100111000011010;
assign LUT_4[53010] = 32'b00000000000000001011000111000110;
assign LUT_4[53011] = 32'b00000000000000000100010010111110;
assign LUT_4[53012] = 32'b00000000000000001000101100111110;
assign LUT_4[53013] = 32'b00000000000000000001111000110110;
assign LUT_4[53014] = 32'b00000000000000001000000111100010;
assign LUT_4[53015] = 32'b00000000000000000001010011011010;
assign LUT_4[53016] = 32'b00000000000000000100111000110111;
assign LUT_4[53017] = 32'b11111111111111111110000100101111;
assign LUT_4[53018] = 32'b00000000000000000100010011011011;
assign LUT_4[53019] = 32'b11111111111111111101011111010011;
assign LUT_4[53020] = 32'b00000000000000000001111001010011;
assign LUT_4[53021] = 32'b11111111111111111011000101001011;
assign LUT_4[53022] = 32'b00000000000000000001010011110111;
assign LUT_4[53023] = 32'b11111111111111111010011111101111;
assign LUT_4[53024] = 32'b00000000000000001100010101111011;
assign LUT_4[53025] = 32'b00000000000000000101100001110011;
assign LUT_4[53026] = 32'b00000000000000001011110000011111;
assign LUT_4[53027] = 32'b00000000000000000100111100010111;
assign LUT_4[53028] = 32'b00000000000000001001010110010111;
assign LUT_4[53029] = 32'b00000000000000000010100010001111;
assign LUT_4[53030] = 32'b00000000000000001000110000111011;
assign LUT_4[53031] = 32'b00000000000000000001111100110011;
assign LUT_4[53032] = 32'b00000000000000000101100010010000;
assign LUT_4[53033] = 32'b11111111111111111110101110001000;
assign LUT_4[53034] = 32'b00000000000000000100111100110100;
assign LUT_4[53035] = 32'b11111111111111111110001000101100;
assign LUT_4[53036] = 32'b00000000000000000010100010101100;
assign LUT_4[53037] = 32'b11111111111111111011101110100100;
assign LUT_4[53038] = 32'b00000000000000000001111101010000;
assign LUT_4[53039] = 32'b11111111111111111011001001001000;
assign LUT_4[53040] = 32'b00000000000000001010000111101001;
assign LUT_4[53041] = 32'b00000000000000000011010011100001;
assign LUT_4[53042] = 32'b00000000000000001001100010001101;
assign LUT_4[53043] = 32'b00000000000000000010101110000101;
assign LUT_4[53044] = 32'b00000000000000000111001000000101;
assign LUT_4[53045] = 32'b00000000000000000000010011111101;
assign LUT_4[53046] = 32'b00000000000000000110100010101001;
assign LUT_4[53047] = 32'b11111111111111111111101110100001;
assign LUT_4[53048] = 32'b00000000000000000011010011111110;
assign LUT_4[53049] = 32'b11111111111111111100011111110110;
assign LUT_4[53050] = 32'b00000000000000000010101110100010;
assign LUT_4[53051] = 32'b11111111111111111011111010011010;
assign LUT_4[53052] = 32'b00000000000000000000010100011010;
assign LUT_4[53053] = 32'b11111111111111111001100000010010;
assign LUT_4[53054] = 32'b11111111111111111111101110111110;
assign LUT_4[53055] = 32'b11111111111111111000111010110110;
assign LUT_4[53056] = 32'b00000000000000001111010010001000;
assign LUT_4[53057] = 32'b00000000000000001000011110000000;
assign LUT_4[53058] = 32'b00000000000000001110101100101100;
assign LUT_4[53059] = 32'b00000000000000000111111000100100;
assign LUT_4[53060] = 32'b00000000000000001100010010100100;
assign LUT_4[53061] = 32'b00000000000000000101011110011100;
assign LUT_4[53062] = 32'b00000000000000001011101101001000;
assign LUT_4[53063] = 32'b00000000000000000100111001000000;
assign LUT_4[53064] = 32'b00000000000000001000011110011101;
assign LUT_4[53065] = 32'b00000000000000000001101010010101;
assign LUT_4[53066] = 32'b00000000000000000111111001000001;
assign LUT_4[53067] = 32'b00000000000000000001000100111001;
assign LUT_4[53068] = 32'b00000000000000000101011110111001;
assign LUT_4[53069] = 32'b11111111111111111110101010110001;
assign LUT_4[53070] = 32'b00000000000000000100111001011101;
assign LUT_4[53071] = 32'b11111111111111111110000101010101;
assign LUT_4[53072] = 32'b00000000000000001101000011110110;
assign LUT_4[53073] = 32'b00000000000000000110001111101110;
assign LUT_4[53074] = 32'b00000000000000001100011110011010;
assign LUT_4[53075] = 32'b00000000000000000101101010010010;
assign LUT_4[53076] = 32'b00000000000000001010000100010010;
assign LUT_4[53077] = 32'b00000000000000000011010000001010;
assign LUT_4[53078] = 32'b00000000000000001001011110110110;
assign LUT_4[53079] = 32'b00000000000000000010101010101110;
assign LUT_4[53080] = 32'b00000000000000000110010000001011;
assign LUT_4[53081] = 32'b11111111111111111111011100000011;
assign LUT_4[53082] = 32'b00000000000000000101101010101111;
assign LUT_4[53083] = 32'b11111111111111111110110110100111;
assign LUT_4[53084] = 32'b00000000000000000011010000100111;
assign LUT_4[53085] = 32'b11111111111111111100011100011111;
assign LUT_4[53086] = 32'b00000000000000000010101011001011;
assign LUT_4[53087] = 32'b11111111111111111011110111000011;
assign LUT_4[53088] = 32'b00000000000000001101101101001111;
assign LUT_4[53089] = 32'b00000000000000000110111001000111;
assign LUT_4[53090] = 32'b00000000000000001101000111110011;
assign LUT_4[53091] = 32'b00000000000000000110010011101011;
assign LUT_4[53092] = 32'b00000000000000001010101101101011;
assign LUT_4[53093] = 32'b00000000000000000011111001100011;
assign LUT_4[53094] = 32'b00000000000000001010001000001111;
assign LUT_4[53095] = 32'b00000000000000000011010100000111;
assign LUT_4[53096] = 32'b00000000000000000110111001100100;
assign LUT_4[53097] = 32'b00000000000000000000000101011100;
assign LUT_4[53098] = 32'b00000000000000000110010100001000;
assign LUT_4[53099] = 32'b11111111111111111111100000000000;
assign LUT_4[53100] = 32'b00000000000000000011111010000000;
assign LUT_4[53101] = 32'b11111111111111111101000101111000;
assign LUT_4[53102] = 32'b00000000000000000011010100100100;
assign LUT_4[53103] = 32'b11111111111111111100100000011100;
assign LUT_4[53104] = 32'b00000000000000001011011110111101;
assign LUT_4[53105] = 32'b00000000000000000100101010110101;
assign LUT_4[53106] = 32'b00000000000000001010111001100001;
assign LUT_4[53107] = 32'b00000000000000000100000101011001;
assign LUT_4[53108] = 32'b00000000000000001000011111011001;
assign LUT_4[53109] = 32'b00000000000000000001101011010001;
assign LUT_4[53110] = 32'b00000000000000000111111001111101;
assign LUT_4[53111] = 32'b00000000000000000001000101110101;
assign LUT_4[53112] = 32'b00000000000000000100101011010010;
assign LUT_4[53113] = 32'b11111111111111111101110111001010;
assign LUT_4[53114] = 32'b00000000000000000100000101110110;
assign LUT_4[53115] = 32'b11111111111111111101010001101110;
assign LUT_4[53116] = 32'b00000000000000000001101011101110;
assign LUT_4[53117] = 32'b11111111111111111010110111100110;
assign LUT_4[53118] = 32'b00000000000000000001000110010010;
assign LUT_4[53119] = 32'b11111111111111111010010010001010;
assign LUT_4[53120] = 32'b00000000000000010000100000111100;
assign LUT_4[53121] = 32'b00000000000000001001101100110100;
assign LUT_4[53122] = 32'b00000000000000001111111011100000;
assign LUT_4[53123] = 32'b00000000000000001001000111011000;
assign LUT_4[53124] = 32'b00000000000000001101100001011000;
assign LUT_4[53125] = 32'b00000000000000000110101101010000;
assign LUT_4[53126] = 32'b00000000000000001100111011111100;
assign LUT_4[53127] = 32'b00000000000000000110000111110100;
assign LUT_4[53128] = 32'b00000000000000001001101101010001;
assign LUT_4[53129] = 32'b00000000000000000010111001001001;
assign LUT_4[53130] = 32'b00000000000000001001000111110101;
assign LUT_4[53131] = 32'b00000000000000000010010011101101;
assign LUT_4[53132] = 32'b00000000000000000110101101101101;
assign LUT_4[53133] = 32'b11111111111111111111111001100101;
assign LUT_4[53134] = 32'b00000000000000000110001000010001;
assign LUT_4[53135] = 32'b11111111111111111111010100001001;
assign LUT_4[53136] = 32'b00000000000000001110010010101010;
assign LUT_4[53137] = 32'b00000000000000000111011110100010;
assign LUT_4[53138] = 32'b00000000000000001101101101001110;
assign LUT_4[53139] = 32'b00000000000000000110111001000110;
assign LUT_4[53140] = 32'b00000000000000001011010011000110;
assign LUT_4[53141] = 32'b00000000000000000100011110111110;
assign LUT_4[53142] = 32'b00000000000000001010101101101010;
assign LUT_4[53143] = 32'b00000000000000000011111001100010;
assign LUT_4[53144] = 32'b00000000000000000111011110111111;
assign LUT_4[53145] = 32'b00000000000000000000101010110111;
assign LUT_4[53146] = 32'b00000000000000000110111001100011;
assign LUT_4[53147] = 32'b00000000000000000000000101011011;
assign LUT_4[53148] = 32'b00000000000000000100011111011011;
assign LUT_4[53149] = 32'b11111111111111111101101011010011;
assign LUT_4[53150] = 32'b00000000000000000011111001111111;
assign LUT_4[53151] = 32'b11111111111111111101000101110111;
assign LUT_4[53152] = 32'b00000000000000001110111100000011;
assign LUT_4[53153] = 32'b00000000000000001000000111111011;
assign LUT_4[53154] = 32'b00000000000000001110010110100111;
assign LUT_4[53155] = 32'b00000000000000000111100010011111;
assign LUT_4[53156] = 32'b00000000000000001011111100011111;
assign LUT_4[53157] = 32'b00000000000000000101001000010111;
assign LUT_4[53158] = 32'b00000000000000001011010111000011;
assign LUT_4[53159] = 32'b00000000000000000100100010111011;
assign LUT_4[53160] = 32'b00000000000000001000001000011000;
assign LUT_4[53161] = 32'b00000000000000000001010100010000;
assign LUT_4[53162] = 32'b00000000000000000111100010111100;
assign LUT_4[53163] = 32'b00000000000000000000101110110100;
assign LUT_4[53164] = 32'b00000000000000000101001000110100;
assign LUT_4[53165] = 32'b11111111111111111110010100101100;
assign LUT_4[53166] = 32'b00000000000000000100100011011000;
assign LUT_4[53167] = 32'b11111111111111111101101111010000;
assign LUT_4[53168] = 32'b00000000000000001100101101110001;
assign LUT_4[53169] = 32'b00000000000000000101111001101001;
assign LUT_4[53170] = 32'b00000000000000001100001000010101;
assign LUT_4[53171] = 32'b00000000000000000101010100001101;
assign LUT_4[53172] = 32'b00000000000000001001101110001101;
assign LUT_4[53173] = 32'b00000000000000000010111010000101;
assign LUT_4[53174] = 32'b00000000000000001001001000110001;
assign LUT_4[53175] = 32'b00000000000000000010010100101001;
assign LUT_4[53176] = 32'b00000000000000000101111010000110;
assign LUT_4[53177] = 32'b11111111111111111111000101111110;
assign LUT_4[53178] = 32'b00000000000000000101010100101010;
assign LUT_4[53179] = 32'b11111111111111111110100000100010;
assign LUT_4[53180] = 32'b00000000000000000010111010100010;
assign LUT_4[53181] = 32'b11111111111111111100000110011010;
assign LUT_4[53182] = 32'b00000000000000000010010101000110;
assign LUT_4[53183] = 32'b11111111111111111011100000111110;
assign LUT_4[53184] = 32'b00000000000000010001111000010000;
assign LUT_4[53185] = 32'b00000000000000001011000100001000;
assign LUT_4[53186] = 32'b00000000000000010001010010110100;
assign LUT_4[53187] = 32'b00000000000000001010011110101100;
assign LUT_4[53188] = 32'b00000000000000001110111000101100;
assign LUT_4[53189] = 32'b00000000000000001000000100100100;
assign LUT_4[53190] = 32'b00000000000000001110010011010000;
assign LUT_4[53191] = 32'b00000000000000000111011111001000;
assign LUT_4[53192] = 32'b00000000000000001011000100100101;
assign LUT_4[53193] = 32'b00000000000000000100010000011101;
assign LUT_4[53194] = 32'b00000000000000001010011111001001;
assign LUT_4[53195] = 32'b00000000000000000011101011000001;
assign LUT_4[53196] = 32'b00000000000000001000000101000001;
assign LUT_4[53197] = 32'b00000000000000000001010000111001;
assign LUT_4[53198] = 32'b00000000000000000111011111100101;
assign LUT_4[53199] = 32'b00000000000000000000101011011101;
assign LUT_4[53200] = 32'b00000000000000001111101001111110;
assign LUT_4[53201] = 32'b00000000000000001000110101110110;
assign LUT_4[53202] = 32'b00000000000000001111000100100010;
assign LUT_4[53203] = 32'b00000000000000001000010000011010;
assign LUT_4[53204] = 32'b00000000000000001100101010011010;
assign LUT_4[53205] = 32'b00000000000000000101110110010010;
assign LUT_4[53206] = 32'b00000000000000001100000100111110;
assign LUT_4[53207] = 32'b00000000000000000101010000110110;
assign LUT_4[53208] = 32'b00000000000000001000110110010011;
assign LUT_4[53209] = 32'b00000000000000000010000010001011;
assign LUT_4[53210] = 32'b00000000000000001000010000110111;
assign LUT_4[53211] = 32'b00000000000000000001011100101111;
assign LUT_4[53212] = 32'b00000000000000000101110110101111;
assign LUT_4[53213] = 32'b11111111111111111111000010100111;
assign LUT_4[53214] = 32'b00000000000000000101010001010011;
assign LUT_4[53215] = 32'b11111111111111111110011101001011;
assign LUT_4[53216] = 32'b00000000000000010000010011010111;
assign LUT_4[53217] = 32'b00000000000000001001011111001111;
assign LUT_4[53218] = 32'b00000000000000001111101101111011;
assign LUT_4[53219] = 32'b00000000000000001000111001110011;
assign LUT_4[53220] = 32'b00000000000000001101010011110011;
assign LUT_4[53221] = 32'b00000000000000000110011111101011;
assign LUT_4[53222] = 32'b00000000000000001100101110010111;
assign LUT_4[53223] = 32'b00000000000000000101111010001111;
assign LUT_4[53224] = 32'b00000000000000001001011111101100;
assign LUT_4[53225] = 32'b00000000000000000010101011100100;
assign LUT_4[53226] = 32'b00000000000000001000111010010000;
assign LUT_4[53227] = 32'b00000000000000000010000110001000;
assign LUT_4[53228] = 32'b00000000000000000110100000001000;
assign LUT_4[53229] = 32'b11111111111111111111101100000000;
assign LUT_4[53230] = 32'b00000000000000000101111010101100;
assign LUT_4[53231] = 32'b11111111111111111111000110100100;
assign LUT_4[53232] = 32'b00000000000000001110000101000101;
assign LUT_4[53233] = 32'b00000000000000000111010000111101;
assign LUT_4[53234] = 32'b00000000000000001101011111101001;
assign LUT_4[53235] = 32'b00000000000000000110101011100001;
assign LUT_4[53236] = 32'b00000000000000001011000101100001;
assign LUT_4[53237] = 32'b00000000000000000100010001011001;
assign LUT_4[53238] = 32'b00000000000000001010100000000101;
assign LUT_4[53239] = 32'b00000000000000000011101011111101;
assign LUT_4[53240] = 32'b00000000000000000111010001011010;
assign LUT_4[53241] = 32'b00000000000000000000011101010010;
assign LUT_4[53242] = 32'b00000000000000000110101011111110;
assign LUT_4[53243] = 32'b11111111111111111111110111110110;
assign LUT_4[53244] = 32'b00000000000000000100010001110110;
assign LUT_4[53245] = 32'b11111111111111111101011101101110;
assign LUT_4[53246] = 32'b00000000000000000011101100011010;
assign LUT_4[53247] = 32'b11111111111111111100111000010010;
assign LUT_4[53248] = 32'b00000000000000001001000001010001;
assign LUT_4[53249] = 32'b00000000000000000010001101001001;
assign LUT_4[53250] = 32'b00000000000000001000011011110101;
assign LUT_4[53251] = 32'b00000000000000000001100111101101;
assign LUT_4[53252] = 32'b00000000000000000110000001101101;
assign LUT_4[53253] = 32'b11111111111111111111001101100101;
assign LUT_4[53254] = 32'b00000000000000000101011100010001;
assign LUT_4[53255] = 32'b11111111111111111110101000001001;
assign LUT_4[53256] = 32'b00000000000000000010001101100110;
assign LUT_4[53257] = 32'b11111111111111111011011001011110;
assign LUT_4[53258] = 32'b00000000000000000001101000001010;
assign LUT_4[53259] = 32'b11111111111111111010110100000010;
assign LUT_4[53260] = 32'b11111111111111111111001110000010;
assign LUT_4[53261] = 32'b11111111111111111000011001111010;
assign LUT_4[53262] = 32'b11111111111111111110101000100110;
assign LUT_4[53263] = 32'b11111111111111110111110100011110;
assign LUT_4[53264] = 32'b00000000000000000110110010111111;
assign LUT_4[53265] = 32'b11111111111111111111111110110111;
assign LUT_4[53266] = 32'b00000000000000000110001101100011;
assign LUT_4[53267] = 32'b11111111111111111111011001011011;
assign LUT_4[53268] = 32'b00000000000000000011110011011011;
assign LUT_4[53269] = 32'b11111111111111111100111111010011;
assign LUT_4[53270] = 32'b00000000000000000011001101111111;
assign LUT_4[53271] = 32'b11111111111111111100011001110111;
assign LUT_4[53272] = 32'b11111111111111111111111111010100;
assign LUT_4[53273] = 32'b11111111111111111001001011001100;
assign LUT_4[53274] = 32'b11111111111111111111011001111000;
assign LUT_4[53275] = 32'b11111111111111111000100101110000;
assign LUT_4[53276] = 32'b11111111111111111100111111110000;
assign LUT_4[53277] = 32'b11111111111111110110001011101000;
assign LUT_4[53278] = 32'b11111111111111111100011010010100;
assign LUT_4[53279] = 32'b11111111111111110101100110001100;
assign LUT_4[53280] = 32'b00000000000000000111011100011000;
assign LUT_4[53281] = 32'b00000000000000000000101000010000;
assign LUT_4[53282] = 32'b00000000000000000110110110111100;
assign LUT_4[53283] = 32'b00000000000000000000000010110100;
assign LUT_4[53284] = 32'b00000000000000000100011100110100;
assign LUT_4[53285] = 32'b11111111111111111101101000101100;
assign LUT_4[53286] = 32'b00000000000000000011110111011000;
assign LUT_4[53287] = 32'b11111111111111111101000011010000;
assign LUT_4[53288] = 32'b00000000000000000000101000101101;
assign LUT_4[53289] = 32'b11111111111111111001110100100101;
assign LUT_4[53290] = 32'b00000000000000000000000011010001;
assign LUT_4[53291] = 32'b11111111111111111001001111001001;
assign LUT_4[53292] = 32'b11111111111111111101101001001001;
assign LUT_4[53293] = 32'b11111111111111110110110101000001;
assign LUT_4[53294] = 32'b11111111111111111101000011101101;
assign LUT_4[53295] = 32'b11111111111111110110001111100101;
assign LUT_4[53296] = 32'b00000000000000000101001110000110;
assign LUT_4[53297] = 32'b11111111111111111110011001111110;
assign LUT_4[53298] = 32'b00000000000000000100101000101010;
assign LUT_4[53299] = 32'b11111111111111111101110100100010;
assign LUT_4[53300] = 32'b00000000000000000010001110100010;
assign LUT_4[53301] = 32'b11111111111111111011011010011010;
assign LUT_4[53302] = 32'b00000000000000000001101001000110;
assign LUT_4[53303] = 32'b11111111111111111010110100111110;
assign LUT_4[53304] = 32'b11111111111111111110011010011011;
assign LUT_4[53305] = 32'b11111111111111110111100110010011;
assign LUT_4[53306] = 32'b11111111111111111101110100111111;
assign LUT_4[53307] = 32'b11111111111111110111000000110111;
assign LUT_4[53308] = 32'b11111111111111111011011010110111;
assign LUT_4[53309] = 32'b11111111111111110100100110101111;
assign LUT_4[53310] = 32'b11111111111111111010110101011011;
assign LUT_4[53311] = 32'b11111111111111110100000001010011;
assign LUT_4[53312] = 32'b00000000000000001010011000100101;
assign LUT_4[53313] = 32'b00000000000000000011100100011101;
assign LUT_4[53314] = 32'b00000000000000001001110011001001;
assign LUT_4[53315] = 32'b00000000000000000010111111000001;
assign LUT_4[53316] = 32'b00000000000000000111011001000001;
assign LUT_4[53317] = 32'b00000000000000000000100100111001;
assign LUT_4[53318] = 32'b00000000000000000110110011100101;
assign LUT_4[53319] = 32'b11111111111111111111111111011101;
assign LUT_4[53320] = 32'b00000000000000000011100100111010;
assign LUT_4[53321] = 32'b11111111111111111100110000110010;
assign LUT_4[53322] = 32'b00000000000000000010111111011110;
assign LUT_4[53323] = 32'b11111111111111111100001011010110;
assign LUT_4[53324] = 32'b00000000000000000000100101010110;
assign LUT_4[53325] = 32'b11111111111111111001110001001110;
assign LUT_4[53326] = 32'b11111111111111111111111111111010;
assign LUT_4[53327] = 32'b11111111111111111001001011110010;
assign LUT_4[53328] = 32'b00000000000000001000001010010011;
assign LUT_4[53329] = 32'b00000000000000000001010110001011;
assign LUT_4[53330] = 32'b00000000000000000111100100110111;
assign LUT_4[53331] = 32'b00000000000000000000110000101111;
assign LUT_4[53332] = 32'b00000000000000000101001010101111;
assign LUT_4[53333] = 32'b11111111111111111110010110100111;
assign LUT_4[53334] = 32'b00000000000000000100100101010011;
assign LUT_4[53335] = 32'b11111111111111111101110001001011;
assign LUT_4[53336] = 32'b00000000000000000001010110101000;
assign LUT_4[53337] = 32'b11111111111111111010100010100000;
assign LUT_4[53338] = 32'b00000000000000000000110001001100;
assign LUT_4[53339] = 32'b11111111111111111001111101000100;
assign LUT_4[53340] = 32'b11111111111111111110010111000100;
assign LUT_4[53341] = 32'b11111111111111110111100010111100;
assign LUT_4[53342] = 32'b11111111111111111101110001101000;
assign LUT_4[53343] = 32'b11111111111111110110111101100000;
assign LUT_4[53344] = 32'b00000000000000001000110011101100;
assign LUT_4[53345] = 32'b00000000000000000001111111100100;
assign LUT_4[53346] = 32'b00000000000000001000001110010000;
assign LUT_4[53347] = 32'b00000000000000000001011010001000;
assign LUT_4[53348] = 32'b00000000000000000101110100001000;
assign LUT_4[53349] = 32'b11111111111111111111000000000000;
assign LUT_4[53350] = 32'b00000000000000000101001110101100;
assign LUT_4[53351] = 32'b11111111111111111110011010100100;
assign LUT_4[53352] = 32'b00000000000000000010000000000001;
assign LUT_4[53353] = 32'b11111111111111111011001011111001;
assign LUT_4[53354] = 32'b00000000000000000001011010100101;
assign LUT_4[53355] = 32'b11111111111111111010100110011101;
assign LUT_4[53356] = 32'b11111111111111111111000000011101;
assign LUT_4[53357] = 32'b11111111111111111000001100010101;
assign LUT_4[53358] = 32'b11111111111111111110011011000001;
assign LUT_4[53359] = 32'b11111111111111110111100110111001;
assign LUT_4[53360] = 32'b00000000000000000110100101011010;
assign LUT_4[53361] = 32'b11111111111111111111110001010010;
assign LUT_4[53362] = 32'b00000000000000000101111111111110;
assign LUT_4[53363] = 32'b11111111111111111111001011110110;
assign LUT_4[53364] = 32'b00000000000000000011100101110110;
assign LUT_4[53365] = 32'b11111111111111111100110001101110;
assign LUT_4[53366] = 32'b00000000000000000011000000011010;
assign LUT_4[53367] = 32'b11111111111111111100001100010010;
assign LUT_4[53368] = 32'b11111111111111111111110001101111;
assign LUT_4[53369] = 32'b11111111111111111000111101100111;
assign LUT_4[53370] = 32'b11111111111111111111001100010011;
assign LUT_4[53371] = 32'b11111111111111111000011000001011;
assign LUT_4[53372] = 32'b11111111111111111100110010001011;
assign LUT_4[53373] = 32'b11111111111111110101111110000011;
assign LUT_4[53374] = 32'b11111111111111111100001100101111;
assign LUT_4[53375] = 32'b11111111111111110101011000100111;
assign LUT_4[53376] = 32'b00000000000000001011100111011001;
assign LUT_4[53377] = 32'b00000000000000000100110011010001;
assign LUT_4[53378] = 32'b00000000000000001011000001111101;
assign LUT_4[53379] = 32'b00000000000000000100001101110101;
assign LUT_4[53380] = 32'b00000000000000001000100111110101;
assign LUT_4[53381] = 32'b00000000000000000001110011101101;
assign LUT_4[53382] = 32'b00000000000000001000000010011001;
assign LUT_4[53383] = 32'b00000000000000000001001110010001;
assign LUT_4[53384] = 32'b00000000000000000100110011101110;
assign LUT_4[53385] = 32'b11111111111111111101111111100110;
assign LUT_4[53386] = 32'b00000000000000000100001110010010;
assign LUT_4[53387] = 32'b11111111111111111101011010001010;
assign LUT_4[53388] = 32'b00000000000000000001110100001010;
assign LUT_4[53389] = 32'b11111111111111111011000000000010;
assign LUT_4[53390] = 32'b00000000000000000001001110101110;
assign LUT_4[53391] = 32'b11111111111111111010011010100110;
assign LUT_4[53392] = 32'b00000000000000001001011001000111;
assign LUT_4[53393] = 32'b00000000000000000010100100111111;
assign LUT_4[53394] = 32'b00000000000000001000110011101011;
assign LUT_4[53395] = 32'b00000000000000000001111111100011;
assign LUT_4[53396] = 32'b00000000000000000110011001100011;
assign LUT_4[53397] = 32'b11111111111111111111100101011011;
assign LUT_4[53398] = 32'b00000000000000000101110100000111;
assign LUT_4[53399] = 32'b11111111111111111110111111111111;
assign LUT_4[53400] = 32'b00000000000000000010100101011100;
assign LUT_4[53401] = 32'b11111111111111111011110001010100;
assign LUT_4[53402] = 32'b00000000000000000010000000000000;
assign LUT_4[53403] = 32'b11111111111111111011001011111000;
assign LUT_4[53404] = 32'b11111111111111111111100101111000;
assign LUT_4[53405] = 32'b11111111111111111000110001110000;
assign LUT_4[53406] = 32'b11111111111111111111000000011100;
assign LUT_4[53407] = 32'b11111111111111111000001100010100;
assign LUT_4[53408] = 32'b00000000000000001010000010100000;
assign LUT_4[53409] = 32'b00000000000000000011001110011000;
assign LUT_4[53410] = 32'b00000000000000001001011101000100;
assign LUT_4[53411] = 32'b00000000000000000010101000111100;
assign LUT_4[53412] = 32'b00000000000000000111000010111100;
assign LUT_4[53413] = 32'b00000000000000000000001110110100;
assign LUT_4[53414] = 32'b00000000000000000110011101100000;
assign LUT_4[53415] = 32'b11111111111111111111101001011000;
assign LUT_4[53416] = 32'b00000000000000000011001110110101;
assign LUT_4[53417] = 32'b11111111111111111100011010101101;
assign LUT_4[53418] = 32'b00000000000000000010101001011001;
assign LUT_4[53419] = 32'b11111111111111111011110101010001;
assign LUT_4[53420] = 32'b00000000000000000000001111010001;
assign LUT_4[53421] = 32'b11111111111111111001011011001001;
assign LUT_4[53422] = 32'b11111111111111111111101001110101;
assign LUT_4[53423] = 32'b11111111111111111000110101101101;
assign LUT_4[53424] = 32'b00000000000000000111110100001110;
assign LUT_4[53425] = 32'b00000000000000000001000000000110;
assign LUT_4[53426] = 32'b00000000000000000111001110110010;
assign LUT_4[53427] = 32'b00000000000000000000011010101010;
assign LUT_4[53428] = 32'b00000000000000000100110100101010;
assign LUT_4[53429] = 32'b11111111111111111110000000100010;
assign LUT_4[53430] = 32'b00000000000000000100001111001110;
assign LUT_4[53431] = 32'b11111111111111111101011011000110;
assign LUT_4[53432] = 32'b00000000000000000001000000100011;
assign LUT_4[53433] = 32'b11111111111111111010001100011011;
assign LUT_4[53434] = 32'b00000000000000000000011011000111;
assign LUT_4[53435] = 32'b11111111111111111001100110111111;
assign LUT_4[53436] = 32'b11111111111111111110000000111111;
assign LUT_4[53437] = 32'b11111111111111110111001100110111;
assign LUT_4[53438] = 32'b11111111111111111101011011100011;
assign LUT_4[53439] = 32'b11111111111111110110100111011011;
assign LUT_4[53440] = 32'b00000000000000001100111110101101;
assign LUT_4[53441] = 32'b00000000000000000110001010100101;
assign LUT_4[53442] = 32'b00000000000000001100011001010001;
assign LUT_4[53443] = 32'b00000000000000000101100101001001;
assign LUT_4[53444] = 32'b00000000000000001001111111001001;
assign LUT_4[53445] = 32'b00000000000000000011001011000001;
assign LUT_4[53446] = 32'b00000000000000001001011001101101;
assign LUT_4[53447] = 32'b00000000000000000010100101100101;
assign LUT_4[53448] = 32'b00000000000000000110001011000010;
assign LUT_4[53449] = 32'b11111111111111111111010110111010;
assign LUT_4[53450] = 32'b00000000000000000101100101100110;
assign LUT_4[53451] = 32'b11111111111111111110110001011110;
assign LUT_4[53452] = 32'b00000000000000000011001011011110;
assign LUT_4[53453] = 32'b11111111111111111100010111010110;
assign LUT_4[53454] = 32'b00000000000000000010100110000010;
assign LUT_4[53455] = 32'b11111111111111111011110001111010;
assign LUT_4[53456] = 32'b00000000000000001010110000011011;
assign LUT_4[53457] = 32'b00000000000000000011111100010011;
assign LUT_4[53458] = 32'b00000000000000001010001010111111;
assign LUT_4[53459] = 32'b00000000000000000011010110110111;
assign LUT_4[53460] = 32'b00000000000000000111110000110111;
assign LUT_4[53461] = 32'b00000000000000000000111100101111;
assign LUT_4[53462] = 32'b00000000000000000111001011011011;
assign LUT_4[53463] = 32'b00000000000000000000010111010011;
assign LUT_4[53464] = 32'b00000000000000000011111100110000;
assign LUT_4[53465] = 32'b11111111111111111101001000101000;
assign LUT_4[53466] = 32'b00000000000000000011010111010100;
assign LUT_4[53467] = 32'b11111111111111111100100011001100;
assign LUT_4[53468] = 32'b00000000000000000000111101001100;
assign LUT_4[53469] = 32'b11111111111111111010001001000100;
assign LUT_4[53470] = 32'b00000000000000000000010111110000;
assign LUT_4[53471] = 32'b11111111111111111001100011101000;
assign LUT_4[53472] = 32'b00000000000000001011011001110100;
assign LUT_4[53473] = 32'b00000000000000000100100101101100;
assign LUT_4[53474] = 32'b00000000000000001010110100011000;
assign LUT_4[53475] = 32'b00000000000000000100000000010000;
assign LUT_4[53476] = 32'b00000000000000001000011010010000;
assign LUT_4[53477] = 32'b00000000000000000001100110001000;
assign LUT_4[53478] = 32'b00000000000000000111110100110100;
assign LUT_4[53479] = 32'b00000000000000000001000000101100;
assign LUT_4[53480] = 32'b00000000000000000100100110001001;
assign LUT_4[53481] = 32'b11111111111111111101110010000001;
assign LUT_4[53482] = 32'b00000000000000000100000000101101;
assign LUT_4[53483] = 32'b11111111111111111101001100100101;
assign LUT_4[53484] = 32'b00000000000000000001100110100101;
assign LUT_4[53485] = 32'b11111111111111111010110010011101;
assign LUT_4[53486] = 32'b00000000000000000001000001001001;
assign LUT_4[53487] = 32'b11111111111111111010001101000001;
assign LUT_4[53488] = 32'b00000000000000001001001011100010;
assign LUT_4[53489] = 32'b00000000000000000010010111011010;
assign LUT_4[53490] = 32'b00000000000000001000100110000110;
assign LUT_4[53491] = 32'b00000000000000000001110001111110;
assign LUT_4[53492] = 32'b00000000000000000110001011111110;
assign LUT_4[53493] = 32'b11111111111111111111010111110110;
assign LUT_4[53494] = 32'b00000000000000000101100110100010;
assign LUT_4[53495] = 32'b11111111111111111110110010011010;
assign LUT_4[53496] = 32'b00000000000000000010010111110111;
assign LUT_4[53497] = 32'b11111111111111111011100011101111;
assign LUT_4[53498] = 32'b00000000000000000001110010011011;
assign LUT_4[53499] = 32'b11111111111111111010111110010011;
assign LUT_4[53500] = 32'b11111111111111111111011000010011;
assign LUT_4[53501] = 32'b11111111111111111000100100001011;
assign LUT_4[53502] = 32'b11111111111111111110110010110111;
assign LUT_4[53503] = 32'b11111111111111110111111110101111;
assign LUT_4[53504] = 32'b00000000000000001101111100110100;
assign LUT_4[53505] = 32'b00000000000000000111001000101100;
assign LUT_4[53506] = 32'b00000000000000001101010111011000;
assign LUT_4[53507] = 32'b00000000000000000110100011010000;
assign LUT_4[53508] = 32'b00000000000000001010111101010000;
assign LUT_4[53509] = 32'b00000000000000000100001001001000;
assign LUT_4[53510] = 32'b00000000000000001010010111110100;
assign LUT_4[53511] = 32'b00000000000000000011100011101100;
assign LUT_4[53512] = 32'b00000000000000000111001001001001;
assign LUT_4[53513] = 32'b00000000000000000000010101000001;
assign LUT_4[53514] = 32'b00000000000000000110100011101101;
assign LUT_4[53515] = 32'b11111111111111111111101111100101;
assign LUT_4[53516] = 32'b00000000000000000100001001100101;
assign LUT_4[53517] = 32'b11111111111111111101010101011101;
assign LUT_4[53518] = 32'b00000000000000000011100100001001;
assign LUT_4[53519] = 32'b11111111111111111100110000000001;
assign LUT_4[53520] = 32'b00000000000000001011101110100010;
assign LUT_4[53521] = 32'b00000000000000000100111010011010;
assign LUT_4[53522] = 32'b00000000000000001011001001000110;
assign LUT_4[53523] = 32'b00000000000000000100010100111110;
assign LUT_4[53524] = 32'b00000000000000001000101110111110;
assign LUT_4[53525] = 32'b00000000000000000001111010110110;
assign LUT_4[53526] = 32'b00000000000000001000001001100010;
assign LUT_4[53527] = 32'b00000000000000000001010101011010;
assign LUT_4[53528] = 32'b00000000000000000100111010110111;
assign LUT_4[53529] = 32'b11111111111111111110000110101111;
assign LUT_4[53530] = 32'b00000000000000000100010101011011;
assign LUT_4[53531] = 32'b11111111111111111101100001010011;
assign LUT_4[53532] = 32'b00000000000000000001111011010011;
assign LUT_4[53533] = 32'b11111111111111111011000111001011;
assign LUT_4[53534] = 32'b00000000000000000001010101110111;
assign LUT_4[53535] = 32'b11111111111111111010100001101111;
assign LUT_4[53536] = 32'b00000000000000001100010111111011;
assign LUT_4[53537] = 32'b00000000000000000101100011110011;
assign LUT_4[53538] = 32'b00000000000000001011110010011111;
assign LUT_4[53539] = 32'b00000000000000000100111110010111;
assign LUT_4[53540] = 32'b00000000000000001001011000010111;
assign LUT_4[53541] = 32'b00000000000000000010100100001111;
assign LUT_4[53542] = 32'b00000000000000001000110010111011;
assign LUT_4[53543] = 32'b00000000000000000001111110110011;
assign LUT_4[53544] = 32'b00000000000000000101100100010000;
assign LUT_4[53545] = 32'b11111111111111111110110000001000;
assign LUT_4[53546] = 32'b00000000000000000100111110110100;
assign LUT_4[53547] = 32'b11111111111111111110001010101100;
assign LUT_4[53548] = 32'b00000000000000000010100100101100;
assign LUT_4[53549] = 32'b11111111111111111011110000100100;
assign LUT_4[53550] = 32'b00000000000000000001111111010000;
assign LUT_4[53551] = 32'b11111111111111111011001011001000;
assign LUT_4[53552] = 32'b00000000000000001010001001101001;
assign LUT_4[53553] = 32'b00000000000000000011010101100001;
assign LUT_4[53554] = 32'b00000000000000001001100100001101;
assign LUT_4[53555] = 32'b00000000000000000010110000000101;
assign LUT_4[53556] = 32'b00000000000000000111001010000101;
assign LUT_4[53557] = 32'b00000000000000000000010101111101;
assign LUT_4[53558] = 32'b00000000000000000110100100101001;
assign LUT_4[53559] = 32'b11111111111111111111110000100001;
assign LUT_4[53560] = 32'b00000000000000000011010101111110;
assign LUT_4[53561] = 32'b11111111111111111100100001110110;
assign LUT_4[53562] = 32'b00000000000000000010110000100010;
assign LUT_4[53563] = 32'b11111111111111111011111100011010;
assign LUT_4[53564] = 32'b00000000000000000000010110011010;
assign LUT_4[53565] = 32'b11111111111111111001100010010010;
assign LUT_4[53566] = 32'b11111111111111111111110000111110;
assign LUT_4[53567] = 32'b11111111111111111000111100110110;
assign LUT_4[53568] = 32'b00000000000000001111010100001000;
assign LUT_4[53569] = 32'b00000000000000001000100000000000;
assign LUT_4[53570] = 32'b00000000000000001110101110101100;
assign LUT_4[53571] = 32'b00000000000000000111111010100100;
assign LUT_4[53572] = 32'b00000000000000001100010100100100;
assign LUT_4[53573] = 32'b00000000000000000101100000011100;
assign LUT_4[53574] = 32'b00000000000000001011101111001000;
assign LUT_4[53575] = 32'b00000000000000000100111011000000;
assign LUT_4[53576] = 32'b00000000000000001000100000011101;
assign LUT_4[53577] = 32'b00000000000000000001101100010101;
assign LUT_4[53578] = 32'b00000000000000000111111011000001;
assign LUT_4[53579] = 32'b00000000000000000001000110111001;
assign LUT_4[53580] = 32'b00000000000000000101100000111001;
assign LUT_4[53581] = 32'b11111111111111111110101100110001;
assign LUT_4[53582] = 32'b00000000000000000100111011011101;
assign LUT_4[53583] = 32'b11111111111111111110000111010101;
assign LUT_4[53584] = 32'b00000000000000001101000101110110;
assign LUT_4[53585] = 32'b00000000000000000110010001101110;
assign LUT_4[53586] = 32'b00000000000000001100100000011010;
assign LUT_4[53587] = 32'b00000000000000000101101100010010;
assign LUT_4[53588] = 32'b00000000000000001010000110010010;
assign LUT_4[53589] = 32'b00000000000000000011010010001010;
assign LUT_4[53590] = 32'b00000000000000001001100000110110;
assign LUT_4[53591] = 32'b00000000000000000010101100101110;
assign LUT_4[53592] = 32'b00000000000000000110010010001011;
assign LUT_4[53593] = 32'b11111111111111111111011110000011;
assign LUT_4[53594] = 32'b00000000000000000101101100101111;
assign LUT_4[53595] = 32'b11111111111111111110111000100111;
assign LUT_4[53596] = 32'b00000000000000000011010010100111;
assign LUT_4[53597] = 32'b11111111111111111100011110011111;
assign LUT_4[53598] = 32'b00000000000000000010101101001011;
assign LUT_4[53599] = 32'b11111111111111111011111001000011;
assign LUT_4[53600] = 32'b00000000000000001101101111001111;
assign LUT_4[53601] = 32'b00000000000000000110111011000111;
assign LUT_4[53602] = 32'b00000000000000001101001001110011;
assign LUT_4[53603] = 32'b00000000000000000110010101101011;
assign LUT_4[53604] = 32'b00000000000000001010101111101011;
assign LUT_4[53605] = 32'b00000000000000000011111011100011;
assign LUT_4[53606] = 32'b00000000000000001010001010001111;
assign LUT_4[53607] = 32'b00000000000000000011010110000111;
assign LUT_4[53608] = 32'b00000000000000000110111011100100;
assign LUT_4[53609] = 32'b00000000000000000000000111011100;
assign LUT_4[53610] = 32'b00000000000000000110010110001000;
assign LUT_4[53611] = 32'b11111111111111111111100010000000;
assign LUT_4[53612] = 32'b00000000000000000011111100000000;
assign LUT_4[53613] = 32'b11111111111111111101000111111000;
assign LUT_4[53614] = 32'b00000000000000000011010110100100;
assign LUT_4[53615] = 32'b11111111111111111100100010011100;
assign LUT_4[53616] = 32'b00000000000000001011100000111101;
assign LUT_4[53617] = 32'b00000000000000000100101100110101;
assign LUT_4[53618] = 32'b00000000000000001010111011100001;
assign LUT_4[53619] = 32'b00000000000000000100000111011001;
assign LUT_4[53620] = 32'b00000000000000001000100001011001;
assign LUT_4[53621] = 32'b00000000000000000001101101010001;
assign LUT_4[53622] = 32'b00000000000000000111111011111101;
assign LUT_4[53623] = 32'b00000000000000000001000111110101;
assign LUT_4[53624] = 32'b00000000000000000100101101010010;
assign LUT_4[53625] = 32'b11111111111111111101111001001010;
assign LUT_4[53626] = 32'b00000000000000000100000111110110;
assign LUT_4[53627] = 32'b11111111111111111101010011101110;
assign LUT_4[53628] = 32'b00000000000000000001101101101110;
assign LUT_4[53629] = 32'b11111111111111111010111001100110;
assign LUT_4[53630] = 32'b00000000000000000001001000010010;
assign LUT_4[53631] = 32'b11111111111111111010010100001010;
assign LUT_4[53632] = 32'b00000000000000010000100010111100;
assign LUT_4[53633] = 32'b00000000000000001001101110110100;
assign LUT_4[53634] = 32'b00000000000000001111111101100000;
assign LUT_4[53635] = 32'b00000000000000001001001001011000;
assign LUT_4[53636] = 32'b00000000000000001101100011011000;
assign LUT_4[53637] = 32'b00000000000000000110101111010000;
assign LUT_4[53638] = 32'b00000000000000001100111101111100;
assign LUT_4[53639] = 32'b00000000000000000110001001110100;
assign LUT_4[53640] = 32'b00000000000000001001101111010001;
assign LUT_4[53641] = 32'b00000000000000000010111011001001;
assign LUT_4[53642] = 32'b00000000000000001001001001110101;
assign LUT_4[53643] = 32'b00000000000000000010010101101101;
assign LUT_4[53644] = 32'b00000000000000000110101111101101;
assign LUT_4[53645] = 32'b11111111111111111111111011100101;
assign LUT_4[53646] = 32'b00000000000000000110001010010001;
assign LUT_4[53647] = 32'b11111111111111111111010110001001;
assign LUT_4[53648] = 32'b00000000000000001110010100101010;
assign LUT_4[53649] = 32'b00000000000000000111100000100010;
assign LUT_4[53650] = 32'b00000000000000001101101111001110;
assign LUT_4[53651] = 32'b00000000000000000110111011000110;
assign LUT_4[53652] = 32'b00000000000000001011010101000110;
assign LUT_4[53653] = 32'b00000000000000000100100000111110;
assign LUT_4[53654] = 32'b00000000000000001010101111101010;
assign LUT_4[53655] = 32'b00000000000000000011111011100010;
assign LUT_4[53656] = 32'b00000000000000000111100000111111;
assign LUT_4[53657] = 32'b00000000000000000000101100110111;
assign LUT_4[53658] = 32'b00000000000000000110111011100011;
assign LUT_4[53659] = 32'b00000000000000000000000111011011;
assign LUT_4[53660] = 32'b00000000000000000100100001011011;
assign LUT_4[53661] = 32'b11111111111111111101101101010011;
assign LUT_4[53662] = 32'b00000000000000000011111011111111;
assign LUT_4[53663] = 32'b11111111111111111101000111110111;
assign LUT_4[53664] = 32'b00000000000000001110111110000011;
assign LUT_4[53665] = 32'b00000000000000001000001001111011;
assign LUT_4[53666] = 32'b00000000000000001110011000100111;
assign LUT_4[53667] = 32'b00000000000000000111100100011111;
assign LUT_4[53668] = 32'b00000000000000001011111110011111;
assign LUT_4[53669] = 32'b00000000000000000101001010010111;
assign LUT_4[53670] = 32'b00000000000000001011011001000011;
assign LUT_4[53671] = 32'b00000000000000000100100100111011;
assign LUT_4[53672] = 32'b00000000000000001000001010011000;
assign LUT_4[53673] = 32'b00000000000000000001010110010000;
assign LUT_4[53674] = 32'b00000000000000000111100100111100;
assign LUT_4[53675] = 32'b00000000000000000000110000110100;
assign LUT_4[53676] = 32'b00000000000000000101001010110100;
assign LUT_4[53677] = 32'b11111111111111111110010110101100;
assign LUT_4[53678] = 32'b00000000000000000100100101011000;
assign LUT_4[53679] = 32'b11111111111111111101110001010000;
assign LUT_4[53680] = 32'b00000000000000001100101111110001;
assign LUT_4[53681] = 32'b00000000000000000101111011101001;
assign LUT_4[53682] = 32'b00000000000000001100001010010101;
assign LUT_4[53683] = 32'b00000000000000000101010110001101;
assign LUT_4[53684] = 32'b00000000000000001001110000001101;
assign LUT_4[53685] = 32'b00000000000000000010111100000101;
assign LUT_4[53686] = 32'b00000000000000001001001010110001;
assign LUT_4[53687] = 32'b00000000000000000010010110101001;
assign LUT_4[53688] = 32'b00000000000000000101111100000110;
assign LUT_4[53689] = 32'b11111111111111111111000111111110;
assign LUT_4[53690] = 32'b00000000000000000101010110101010;
assign LUT_4[53691] = 32'b11111111111111111110100010100010;
assign LUT_4[53692] = 32'b00000000000000000010111100100010;
assign LUT_4[53693] = 32'b11111111111111111100001000011010;
assign LUT_4[53694] = 32'b00000000000000000010010111000110;
assign LUT_4[53695] = 32'b11111111111111111011100010111110;
assign LUT_4[53696] = 32'b00000000000000010001111010010000;
assign LUT_4[53697] = 32'b00000000000000001011000110001000;
assign LUT_4[53698] = 32'b00000000000000010001010100110100;
assign LUT_4[53699] = 32'b00000000000000001010100000101100;
assign LUT_4[53700] = 32'b00000000000000001110111010101100;
assign LUT_4[53701] = 32'b00000000000000001000000110100100;
assign LUT_4[53702] = 32'b00000000000000001110010101010000;
assign LUT_4[53703] = 32'b00000000000000000111100001001000;
assign LUT_4[53704] = 32'b00000000000000001011000110100101;
assign LUT_4[53705] = 32'b00000000000000000100010010011101;
assign LUT_4[53706] = 32'b00000000000000001010100001001001;
assign LUT_4[53707] = 32'b00000000000000000011101101000001;
assign LUT_4[53708] = 32'b00000000000000001000000111000001;
assign LUT_4[53709] = 32'b00000000000000000001010010111001;
assign LUT_4[53710] = 32'b00000000000000000111100001100101;
assign LUT_4[53711] = 32'b00000000000000000000101101011101;
assign LUT_4[53712] = 32'b00000000000000001111101011111110;
assign LUT_4[53713] = 32'b00000000000000001000110111110110;
assign LUT_4[53714] = 32'b00000000000000001111000110100010;
assign LUT_4[53715] = 32'b00000000000000001000010010011010;
assign LUT_4[53716] = 32'b00000000000000001100101100011010;
assign LUT_4[53717] = 32'b00000000000000000101111000010010;
assign LUT_4[53718] = 32'b00000000000000001100000110111110;
assign LUT_4[53719] = 32'b00000000000000000101010010110110;
assign LUT_4[53720] = 32'b00000000000000001000111000010011;
assign LUT_4[53721] = 32'b00000000000000000010000100001011;
assign LUT_4[53722] = 32'b00000000000000001000010010110111;
assign LUT_4[53723] = 32'b00000000000000000001011110101111;
assign LUT_4[53724] = 32'b00000000000000000101111000101111;
assign LUT_4[53725] = 32'b11111111111111111111000100100111;
assign LUT_4[53726] = 32'b00000000000000000101010011010011;
assign LUT_4[53727] = 32'b11111111111111111110011111001011;
assign LUT_4[53728] = 32'b00000000000000010000010101010111;
assign LUT_4[53729] = 32'b00000000000000001001100001001111;
assign LUT_4[53730] = 32'b00000000000000001111101111111011;
assign LUT_4[53731] = 32'b00000000000000001000111011110011;
assign LUT_4[53732] = 32'b00000000000000001101010101110011;
assign LUT_4[53733] = 32'b00000000000000000110100001101011;
assign LUT_4[53734] = 32'b00000000000000001100110000010111;
assign LUT_4[53735] = 32'b00000000000000000101111100001111;
assign LUT_4[53736] = 32'b00000000000000001001100001101100;
assign LUT_4[53737] = 32'b00000000000000000010101101100100;
assign LUT_4[53738] = 32'b00000000000000001000111100010000;
assign LUT_4[53739] = 32'b00000000000000000010001000001000;
assign LUT_4[53740] = 32'b00000000000000000110100010001000;
assign LUT_4[53741] = 32'b11111111111111111111101110000000;
assign LUT_4[53742] = 32'b00000000000000000101111100101100;
assign LUT_4[53743] = 32'b11111111111111111111001000100100;
assign LUT_4[53744] = 32'b00000000000000001110000111000101;
assign LUT_4[53745] = 32'b00000000000000000111010010111101;
assign LUT_4[53746] = 32'b00000000000000001101100001101001;
assign LUT_4[53747] = 32'b00000000000000000110101101100001;
assign LUT_4[53748] = 32'b00000000000000001011000111100001;
assign LUT_4[53749] = 32'b00000000000000000100010011011001;
assign LUT_4[53750] = 32'b00000000000000001010100010000101;
assign LUT_4[53751] = 32'b00000000000000000011101101111101;
assign LUT_4[53752] = 32'b00000000000000000111010011011010;
assign LUT_4[53753] = 32'b00000000000000000000011111010010;
assign LUT_4[53754] = 32'b00000000000000000110101101111110;
assign LUT_4[53755] = 32'b11111111111111111111111001110110;
assign LUT_4[53756] = 32'b00000000000000000100010011110110;
assign LUT_4[53757] = 32'b11111111111111111101011111101110;
assign LUT_4[53758] = 32'b00000000000000000011101110011010;
assign LUT_4[53759] = 32'b11111111111111111100111010010010;
assign LUT_4[53760] = 32'b00000000000000001000000101011001;
assign LUT_4[53761] = 32'b00000000000000000001010001010001;
assign LUT_4[53762] = 32'b00000000000000000111011111111101;
assign LUT_4[53763] = 32'b00000000000000000000101011110101;
assign LUT_4[53764] = 32'b00000000000000000101000101110101;
assign LUT_4[53765] = 32'b11111111111111111110010001101101;
assign LUT_4[53766] = 32'b00000000000000000100100000011001;
assign LUT_4[53767] = 32'b11111111111111111101101100010001;
assign LUT_4[53768] = 32'b00000000000000000001010001101110;
assign LUT_4[53769] = 32'b11111111111111111010011101100110;
assign LUT_4[53770] = 32'b00000000000000000000101100010010;
assign LUT_4[53771] = 32'b11111111111111111001111000001010;
assign LUT_4[53772] = 32'b11111111111111111110010010001010;
assign LUT_4[53773] = 32'b11111111111111110111011110000010;
assign LUT_4[53774] = 32'b11111111111111111101101100101110;
assign LUT_4[53775] = 32'b11111111111111110110111000100110;
assign LUT_4[53776] = 32'b00000000000000000101110111000111;
assign LUT_4[53777] = 32'b11111111111111111111000010111111;
assign LUT_4[53778] = 32'b00000000000000000101010001101011;
assign LUT_4[53779] = 32'b11111111111111111110011101100011;
assign LUT_4[53780] = 32'b00000000000000000010110111100011;
assign LUT_4[53781] = 32'b11111111111111111100000011011011;
assign LUT_4[53782] = 32'b00000000000000000010010010000111;
assign LUT_4[53783] = 32'b11111111111111111011011101111111;
assign LUT_4[53784] = 32'b11111111111111111111000011011100;
assign LUT_4[53785] = 32'b11111111111111111000001111010100;
assign LUT_4[53786] = 32'b11111111111111111110011110000000;
assign LUT_4[53787] = 32'b11111111111111110111101001111000;
assign LUT_4[53788] = 32'b11111111111111111100000011111000;
assign LUT_4[53789] = 32'b11111111111111110101001111110000;
assign LUT_4[53790] = 32'b11111111111111111011011110011100;
assign LUT_4[53791] = 32'b11111111111111110100101010010100;
assign LUT_4[53792] = 32'b00000000000000000110100000100000;
assign LUT_4[53793] = 32'b11111111111111111111101100011000;
assign LUT_4[53794] = 32'b00000000000000000101111011000100;
assign LUT_4[53795] = 32'b11111111111111111111000110111100;
assign LUT_4[53796] = 32'b00000000000000000011100000111100;
assign LUT_4[53797] = 32'b11111111111111111100101100110100;
assign LUT_4[53798] = 32'b00000000000000000010111011100000;
assign LUT_4[53799] = 32'b11111111111111111100000111011000;
assign LUT_4[53800] = 32'b11111111111111111111101100110101;
assign LUT_4[53801] = 32'b11111111111111111000111000101101;
assign LUT_4[53802] = 32'b11111111111111111111000111011001;
assign LUT_4[53803] = 32'b11111111111111111000010011010001;
assign LUT_4[53804] = 32'b11111111111111111100101101010001;
assign LUT_4[53805] = 32'b11111111111111110101111001001001;
assign LUT_4[53806] = 32'b11111111111111111100000111110101;
assign LUT_4[53807] = 32'b11111111111111110101010011101101;
assign LUT_4[53808] = 32'b00000000000000000100010010001110;
assign LUT_4[53809] = 32'b11111111111111111101011110000110;
assign LUT_4[53810] = 32'b00000000000000000011101100110010;
assign LUT_4[53811] = 32'b11111111111111111100111000101010;
assign LUT_4[53812] = 32'b00000000000000000001010010101010;
assign LUT_4[53813] = 32'b11111111111111111010011110100010;
assign LUT_4[53814] = 32'b00000000000000000000101101001110;
assign LUT_4[53815] = 32'b11111111111111111001111001000110;
assign LUT_4[53816] = 32'b11111111111111111101011110100011;
assign LUT_4[53817] = 32'b11111111111111110110101010011011;
assign LUT_4[53818] = 32'b11111111111111111100111001000111;
assign LUT_4[53819] = 32'b11111111111111110110000100111111;
assign LUT_4[53820] = 32'b11111111111111111010011110111111;
assign LUT_4[53821] = 32'b11111111111111110011101010110111;
assign LUT_4[53822] = 32'b11111111111111111001111001100011;
assign LUT_4[53823] = 32'b11111111111111110011000101011011;
assign LUT_4[53824] = 32'b00000000000000001001011100101101;
assign LUT_4[53825] = 32'b00000000000000000010101000100101;
assign LUT_4[53826] = 32'b00000000000000001000110111010001;
assign LUT_4[53827] = 32'b00000000000000000010000011001001;
assign LUT_4[53828] = 32'b00000000000000000110011101001001;
assign LUT_4[53829] = 32'b11111111111111111111101001000001;
assign LUT_4[53830] = 32'b00000000000000000101110111101101;
assign LUT_4[53831] = 32'b11111111111111111111000011100101;
assign LUT_4[53832] = 32'b00000000000000000010101001000010;
assign LUT_4[53833] = 32'b11111111111111111011110100111010;
assign LUT_4[53834] = 32'b00000000000000000010000011100110;
assign LUT_4[53835] = 32'b11111111111111111011001111011110;
assign LUT_4[53836] = 32'b11111111111111111111101001011110;
assign LUT_4[53837] = 32'b11111111111111111000110101010110;
assign LUT_4[53838] = 32'b11111111111111111111000100000010;
assign LUT_4[53839] = 32'b11111111111111111000001111111010;
assign LUT_4[53840] = 32'b00000000000000000111001110011011;
assign LUT_4[53841] = 32'b00000000000000000000011010010011;
assign LUT_4[53842] = 32'b00000000000000000110101000111111;
assign LUT_4[53843] = 32'b11111111111111111111110100110111;
assign LUT_4[53844] = 32'b00000000000000000100001110110111;
assign LUT_4[53845] = 32'b11111111111111111101011010101111;
assign LUT_4[53846] = 32'b00000000000000000011101001011011;
assign LUT_4[53847] = 32'b11111111111111111100110101010011;
assign LUT_4[53848] = 32'b00000000000000000000011010110000;
assign LUT_4[53849] = 32'b11111111111111111001100110101000;
assign LUT_4[53850] = 32'b11111111111111111111110101010100;
assign LUT_4[53851] = 32'b11111111111111111001000001001100;
assign LUT_4[53852] = 32'b11111111111111111101011011001100;
assign LUT_4[53853] = 32'b11111111111111110110100111000100;
assign LUT_4[53854] = 32'b11111111111111111100110101110000;
assign LUT_4[53855] = 32'b11111111111111110110000001101000;
assign LUT_4[53856] = 32'b00000000000000000111110111110100;
assign LUT_4[53857] = 32'b00000000000000000001000011101100;
assign LUT_4[53858] = 32'b00000000000000000111010010011000;
assign LUT_4[53859] = 32'b00000000000000000000011110010000;
assign LUT_4[53860] = 32'b00000000000000000100111000010000;
assign LUT_4[53861] = 32'b11111111111111111110000100001000;
assign LUT_4[53862] = 32'b00000000000000000100010010110100;
assign LUT_4[53863] = 32'b11111111111111111101011110101100;
assign LUT_4[53864] = 32'b00000000000000000001000100001001;
assign LUT_4[53865] = 32'b11111111111111111010010000000001;
assign LUT_4[53866] = 32'b00000000000000000000011110101101;
assign LUT_4[53867] = 32'b11111111111111111001101010100101;
assign LUT_4[53868] = 32'b11111111111111111110000100100101;
assign LUT_4[53869] = 32'b11111111111111110111010000011101;
assign LUT_4[53870] = 32'b11111111111111111101011111001001;
assign LUT_4[53871] = 32'b11111111111111110110101011000001;
assign LUT_4[53872] = 32'b00000000000000000101101001100010;
assign LUT_4[53873] = 32'b11111111111111111110110101011010;
assign LUT_4[53874] = 32'b00000000000000000101000100000110;
assign LUT_4[53875] = 32'b11111111111111111110001111111110;
assign LUT_4[53876] = 32'b00000000000000000010101001111110;
assign LUT_4[53877] = 32'b11111111111111111011110101110110;
assign LUT_4[53878] = 32'b00000000000000000010000100100010;
assign LUT_4[53879] = 32'b11111111111111111011010000011010;
assign LUT_4[53880] = 32'b11111111111111111110110101110111;
assign LUT_4[53881] = 32'b11111111111111111000000001101111;
assign LUT_4[53882] = 32'b11111111111111111110010000011011;
assign LUT_4[53883] = 32'b11111111111111110111011100010011;
assign LUT_4[53884] = 32'b11111111111111111011110110010011;
assign LUT_4[53885] = 32'b11111111111111110101000010001011;
assign LUT_4[53886] = 32'b11111111111111111011010000110111;
assign LUT_4[53887] = 32'b11111111111111110100011100101111;
assign LUT_4[53888] = 32'b00000000000000001010101011100001;
assign LUT_4[53889] = 32'b00000000000000000011110111011001;
assign LUT_4[53890] = 32'b00000000000000001010000110000101;
assign LUT_4[53891] = 32'b00000000000000000011010001111101;
assign LUT_4[53892] = 32'b00000000000000000111101011111101;
assign LUT_4[53893] = 32'b00000000000000000000110111110101;
assign LUT_4[53894] = 32'b00000000000000000111000110100001;
assign LUT_4[53895] = 32'b00000000000000000000010010011001;
assign LUT_4[53896] = 32'b00000000000000000011110111110110;
assign LUT_4[53897] = 32'b11111111111111111101000011101110;
assign LUT_4[53898] = 32'b00000000000000000011010010011010;
assign LUT_4[53899] = 32'b11111111111111111100011110010010;
assign LUT_4[53900] = 32'b00000000000000000000111000010010;
assign LUT_4[53901] = 32'b11111111111111111010000100001010;
assign LUT_4[53902] = 32'b00000000000000000000010010110110;
assign LUT_4[53903] = 32'b11111111111111111001011110101110;
assign LUT_4[53904] = 32'b00000000000000001000011101001111;
assign LUT_4[53905] = 32'b00000000000000000001101001000111;
assign LUT_4[53906] = 32'b00000000000000000111110111110011;
assign LUT_4[53907] = 32'b00000000000000000001000011101011;
assign LUT_4[53908] = 32'b00000000000000000101011101101011;
assign LUT_4[53909] = 32'b11111111111111111110101001100011;
assign LUT_4[53910] = 32'b00000000000000000100111000001111;
assign LUT_4[53911] = 32'b11111111111111111110000100000111;
assign LUT_4[53912] = 32'b00000000000000000001101001100100;
assign LUT_4[53913] = 32'b11111111111111111010110101011100;
assign LUT_4[53914] = 32'b00000000000000000001000100001000;
assign LUT_4[53915] = 32'b11111111111111111010010000000000;
assign LUT_4[53916] = 32'b11111111111111111110101010000000;
assign LUT_4[53917] = 32'b11111111111111110111110101111000;
assign LUT_4[53918] = 32'b11111111111111111110000100100100;
assign LUT_4[53919] = 32'b11111111111111110111010000011100;
assign LUT_4[53920] = 32'b00000000000000001001000110101000;
assign LUT_4[53921] = 32'b00000000000000000010010010100000;
assign LUT_4[53922] = 32'b00000000000000001000100001001100;
assign LUT_4[53923] = 32'b00000000000000000001101101000100;
assign LUT_4[53924] = 32'b00000000000000000110000111000100;
assign LUT_4[53925] = 32'b11111111111111111111010010111100;
assign LUT_4[53926] = 32'b00000000000000000101100001101000;
assign LUT_4[53927] = 32'b11111111111111111110101101100000;
assign LUT_4[53928] = 32'b00000000000000000010010010111101;
assign LUT_4[53929] = 32'b11111111111111111011011110110101;
assign LUT_4[53930] = 32'b00000000000000000001101101100001;
assign LUT_4[53931] = 32'b11111111111111111010111001011001;
assign LUT_4[53932] = 32'b11111111111111111111010011011001;
assign LUT_4[53933] = 32'b11111111111111111000011111010001;
assign LUT_4[53934] = 32'b11111111111111111110101101111101;
assign LUT_4[53935] = 32'b11111111111111110111111001110101;
assign LUT_4[53936] = 32'b00000000000000000110111000010110;
assign LUT_4[53937] = 32'b00000000000000000000000100001110;
assign LUT_4[53938] = 32'b00000000000000000110010010111010;
assign LUT_4[53939] = 32'b11111111111111111111011110110010;
assign LUT_4[53940] = 32'b00000000000000000011111000110010;
assign LUT_4[53941] = 32'b11111111111111111101000100101010;
assign LUT_4[53942] = 32'b00000000000000000011010011010110;
assign LUT_4[53943] = 32'b11111111111111111100011111001110;
assign LUT_4[53944] = 32'b00000000000000000000000100101011;
assign LUT_4[53945] = 32'b11111111111111111001010000100011;
assign LUT_4[53946] = 32'b11111111111111111111011111001111;
assign LUT_4[53947] = 32'b11111111111111111000101011000111;
assign LUT_4[53948] = 32'b11111111111111111101000101000111;
assign LUT_4[53949] = 32'b11111111111111110110010000111111;
assign LUT_4[53950] = 32'b11111111111111111100011111101011;
assign LUT_4[53951] = 32'b11111111111111110101101011100011;
assign LUT_4[53952] = 32'b00000000000000001100000010110101;
assign LUT_4[53953] = 32'b00000000000000000101001110101101;
assign LUT_4[53954] = 32'b00000000000000001011011101011001;
assign LUT_4[53955] = 32'b00000000000000000100101001010001;
assign LUT_4[53956] = 32'b00000000000000001001000011010001;
assign LUT_4[53957] = 32'b00000000000000000010001111001001;
assign LUT_4[53958] = 32'b00000000000000001000011101110101;
assign LUT_4[53959] = 32'b00000000000000000001101001101101;
assign LUT_4[53960] = 32'b00000000000000000101001111001010;
assign LUT_4[53961] = 32'b11111111111111111110011011000010;
assign LUT_4[53962] = 32'b00000000000000000100101001101110;
assign LUT_4[53963] = 32'b11111111111111111101110101100110;
assign LUT_4[53964] = 32'b00000000000000000010001111100110;
assign LUT_4[53965] = 32'b11111111111111111011011011011110;
assign LUT_4[53966] = 32'b00000000000000000001101010001010;
assign LUT_4[53967] = 32'b11111111111111111010110110000010;
assign LUT_4[53968] = 32'b00000000000000001001110100100011;
assign LUT_4[53969] = 32'b00000000000000000011000000011011;
assign LUT_4[53970] = 32'b00000000000000001001001111000111;
assign LUT_4[53971] = 32'b00000000000000000010011010111111;
assign LUT_4[53972] = 32'b00000000000000000110110100111111;
assign LUT_4[53973] = 32'b00000000000000000000000000110111;
assign LUT_4[53974] = 32'b00000000000000000110001111100011;
assign LUT_4[53975] = 32'b11111111111111111111011011011011;
assign LUT_4[53976] = 32'b00000000000000000011000000111000;
assign LUT_4[53977] = 32'b11111111111111111100001100110000;
assign LUT_4[53978] = 32'b00000000000000000010011011011100;
assign LUT_4[53979] = 32'b11111111111111111011100111010100;
assign LUT_4[53980] = 32'b00000000000000000000000001010100;
assign LUT_4[53981] = 32'b11111111111111111001001101001100;
assign LUT_4[53982] = 32'b11111111111111111111011011111000;
assign LUT_4[53983] = 32'b11111111111111111000100111110000;
assign LUT_4[53984] = 32'b00000000000000001010011101111100;
assign LUT_4[53985] = 32'b00000000000000000011101001110100;
assign LUT_4[53986] = 32'b00000000000000001001111000100000;
assign LUT_4[53987] = 32'b00000000000000000011000100011000;
assign LUT_4[53988] = 32'b00000000000000000111011110011000;
assign LUT_4[53989] = 32'b00000000000000000000101010010000;
assign LUT_4[53990] = 32'b00000000000000000110111000111100;
assign LUT_4[53991] = 32'b00000000000000000000000100110100;
assign LUT_4[53992] = 32'b00000000000000000011101010010001;
assign LUT_4[53993] = 32'b11111111111111111100110110001001;
assign LUT_4[53994] = 32'b00000000000000000011000100110101;
assign LUT_4[53995] = 32'b11111111111111111100010000101101;
assign LUT_4[53996] = 32'b00000000000000000000101010101101;
assign LUT_4[53997] = 32'b11111111111111111001110110100101;
assign LUT_4[53998] = 32'b00000000000000000000000101010001;
assign LUT_4[53999] = 32'b11111111111111111001010001001001;
assign LUT_4[54000] = 32'b00000000000000001000001111101010;
assign LUT_4[54001] = 32'b00000000000000000001011011100010;
assign LUT_4[54002] = 32'b00000000000000000111101010001110;
assign LUT_4[54003] = 32'b00000000000000000000110110000110;
assign LUT_4[54004] = 32'b00000000000000000101010000000110;
assign LUT_4[54005] = 32'b11111111111111111110011011111110;
assign LUT_4[54006] = 32'b00000000000000000100101010101010;
assign LUT_4[54007] = 32'b11111111111111111101110110100010;
assign LUT_4[54008] = 32'b00000000000000000001011011111111;
assign LUT_4[54009] = 32'b11111111111111111010100111110111;
assign LUT_4[54010] = 32'b00000000000000000000110110100011;
assign LUT_4[54011] = 32'b11111111111111111010000010011011;
assign LUT_4[54012] = 32'b11111111111111111110011100011011;
assign LUT_4[54013] = 32'b11111111111111110111101000010011;
assign LUT_4[54014] = 32'b11111111111111111101110110111111;
assign LUT_4[54015] = 32'b11111111111111110111000010110111;
assign LUT_4[54016] = 32'b00000000000000001101000000111100;
assign LUT_4[54017] = 32'b00000000000000000110001100110100;
assign LUT_4[54018] = 32'b00000000000000001100011011100000;
assign LUT_4[54019] = 32'b00000000000000000101100111011000;
assign LUT_4[54020] = 32'b00000000000000001010000001011000;
assign LUT_4[54021] = 32'b00000000000000000011001101010000;
assign LUT_4[54022] = 32'b00000000000000001001011011111100;
assign LUT_4[54023] = 32'b00000000000000000010100111110100;
assign LUT_4[54024] = 32'b00000000000000000110001101010001;
assign LUT_4[54025] = 32'b11111111111111111111011001001001;
assign LUT_4[54026] = 32'b00000000000000000101100111110101;
assign LUT_4[54027] = 32'b11111111111111111110110011101101;
assign LUT_4[54028] = 32'b00000000000000000011001101101101;
assign LUT_4[54029] = 32'b11111111111111111100011001100101;
assign LUT_4[54030] = 32'b00000000000000000010101000010001;
assign LUT_4[54031] = 32'b11111111111111111011110100001001;
assign LUT_4[54032] = 32'b00000000000000001010110010101010;
assign LUT_4[54033] = 32'b00000000000000000011111110100010;
assign LUT_4[54034] = 32'b00000000000000001010001101001110;
assign LUT_4[54035] = 32'b00000000000000000011011001000110;
assign LUT_4[54036] = 32'b00000000000000000111110011000110;
assign LUT_4[54037] = 32'b00000000000000000000111110111110;
assign LUT_4[54038] = 32'b00000000000000000111001101101010;
assign LUT_4[54039] = 32'b00000000000000000000011001100010;
assign LUT_4[54040] = 32'b00000000000000000011111110111111;
assign LUT_4[54041] = 32'b11111111111111111101001010110111;
assign LUT_4[54042] = 32'b00000000000000000011011001100011;
assign LUT_4[54043] = 32'b11111111111111111100100101011011;
assign LUT_4[54044] = 32'b00000000000000000000111111011011;
assign LUT_4[54045] = 32'b11111111111111111010001011010011;
assign LUT_4[54046] = 32'b00000000000000000000011001111111;
assign LUT_4[54047] = 32'b11111111111111111001100101110111;
assign LUT_4[54048] = 32'b00000000000000001011011100000011;
assign LUT_4[54049] = 32'b00000000000000000100100111111011;
assign LUT_4[54050] = 32'b00000000000000001010110110100111;
assign LUT_4[54051] = 32'b00000000000000000100000010011111;
assign LUT_4[54052] = 32'b00000000000000001000011100011111;
assign LUT_4[54053] = 32'b00000000000000000001101000010111;
assign LUT_4[54054] = 32'b00000000000000000111110111000011;
assign LUT_4[54055] = 32'b00000000000000000001000010111011;
assign LUT_4[54056] = 32'b00000000000000000100101000011000;
assign LUT_4[54057] = 32'b11111111111111111101110100010000;
assign LUT_4[54058] = 32'b00000000000000000100000010111100;
assign LUT_4[54059] = 32'b11111111111111111101001110110100;
assign LUT_4[54060] = 32'b00000000000000000001101000110100;
assign LUT_4[54061] = 32'b11111111111111111010110100101100;
assign LUT_4[54062] = 32'b00000000000000000001000011011000;
assign LUT_4[54063] = 32'b11111111111111111010001111010000;
assign LUT_4[54064] = 32'b00000000000000001001001101110001;
assign LUT_4[54065] = 32'b00000000000000000010011001101001;
assign LUT_4[54066] = 32'b00000000000000001000101000010101;
assign LUT_4[54067] = 32'b00000000000000000001110100001101;
assign LUT_4[54068] = 32'b00000000000000000110001110001101;
assign LUT_4[54069] = 32'b11111111111111111111011010000101;
assign LUT_4[54070] = 32'b00000000000000000101101000110001;
assign LUT_4[54071] = 32'b11111111111111111110110100101001;
assign LUT_4[54072] = 32'b00000000000000000010011010000110;
assign LUT_4[54073] = 32'b11111111111111111011100101111110;
assign LUT_4[54074] = 32'b00000000000000000001110100101010;
assign LUT_4[54075] = 32'b11111111111111111011000000100010;
assign LUT_4[54076] = 32'b11111111111111111111011010100010;
assign LUT_4[54077] = 32'b11111111111111111000100110011010;
assign LUT_4[54078] = 32'b11111111111111111110110101000110;
assign LUT_4[54079] = 32'b11111111111111111000000000111110;
assign LUT_4[54080] = 32'b00000000000000001110011000010000;
assign LUT_4[54081] = 32'b00000000000000000111100100001000;
assign LUT_4[54082] = 32'b00000000000000001101110010110100;
assign LUT_4[54083] = 32'b00000000000000000110111110101100;
assign LUT_4[54084] = 32'b00000000000000001011011000101100;
assign LUT_4[54085] = 32'b00000000000000000100100100100100;
assign LUT_4[54086] = 32'b00000000000000001010110011010000;
assign LUT_4[54087] = 32'b00000000000000000011111111001000;
assign LUT_4[54088] = 32'b00000000000000000111100100100101;
assign LUT_4[54089] = 32'b00000000000000000000110000011101;
assign LUT_4[54090] = 32'b00000000000000000110111111001001;
assign LUT_4[54091] = 32'b00000000000000000000001011000001;
assign LUT_4[54092] = 32'b00000000000000000100100101000001;
assign LUT_4[54093] = 32'b11111111111111111101110000111001;
assign LUT_4[54094] = 32'b00000000000000000011111111100101;
assign LUT_4[54095] = 32'b11111111111111111101001011011101;
assign LUT_4[54096] = 32'b00000000000000001100001001111110;
assign LUT_4[54097] = 32'b00000000000000000101010101110110;
assign LUT_4[54098] = 32'b00000000000000001011100100100010;
assign LUT_4[54099] = 32'b00000000000000000100110000011010;
assign LUT_4[54100] = 32'b00000000000000001001001010011010;
assign LUT_4[54101] = 32'b00000000000000000010010110010010;
assign LUT_4[54102] = 32'b00000000000000001000100100111110;
assign LUT_4[54103] = 32'b00000000000000000001110000110110;
assign LUT_4[54104] = 32'b00000000000000000101010110010011;
assign LUT_4[54105] = 32'b11111111111111111110100010001011;
assign LUT_4[54106] = 32'b00000000000000000100110000110111;
assign LUT_4[54107] = 32'b11111111111111111101111100101111;
assign LUT_4[54108] = 32'b00000000000000000010010110101111;
assign LUT_4[54109] = 32'b11111111111111111011100010100111;
assign LUT_4[54110] = 32'b00000000000000000001110001010011;
assign LUT_4[54111] = 32'b11111111111111111010111101001011;
assign LUT_4[54112] = 32'b00000000000000001100110011010111;
assign LUT_4[54113] = 32'b00000000000000000101111111001111;
assign LUT_4[54114] = 32'b00000000000000001100001101111011;
assign LUT_4[54115] = 32'b00000000000000000101011001110011;
assign LUT_4[54116] = 32'b00000000000000001001110011110011;
assign LUT_4[54117] = 32'b00000000000000000010111111101011;
assign LUT_4[54118] = 32'b00000000000000001001001110010111;
assign LUT_4[54119] = 32'b00000000000000000010011010001111;
assign LUT_4[54120] = 32'b00000000000000000101111111101100;
assign LUT_4[54121] = 32'b11111111111111111111001011100100;
assign LUT_4[54122] = 32'b00000000000000000101011010010000;
assign LUT_4[54123] = 32'b11111111111111111110100110001000;
assign LUT_4[54124] = 32'b00000000000000000011000000001000;
assign LUT_4[54125] = 32'b11111111111111111100001100000000;
assign LUT_4[54126] = 32'b00000000000000000010011010101100;
assign LUT_4[54127] = 32'b11111111111111111011100110100100;
assign LUT_4[54128] = 32'b00000000000000001010100101000101;
assign LUT_4[54129] = 32'b00000000000000000011110000111101;
assign LUT_4[54130] = 32'b00000000000000001001111111101001;
assign LUT_4[54131] = 32'b00000000000000000011001011100001;
assign LUT_4[54132] = 32'b00000000000000000111100101100001;
assign LUT_4[54133] = 32'b00000000000000000000110001011001;
assign LUT_4[54134] = 32'b00000000000000000111000000000101;
assign LUT_4[54135] = 32'b00000000000000000000001011111101;
assign LUT_4[54136] = 32'b00000000000000000011110001011010;
assign LUT_4[54137] = 32'b11111111111111111100111101010010;
assign LUT_4[54138] = 32'b00000000000000000011001011111110;
assign LUT_4[54139] = 32'b11111111111111111100010111110110;
assign LUT_4[54140] = 32'b00000000000000000000110001110110;
assign LUT_4[54141] = 32'b11111111111111111001111101101110;
assign LUT_4[54142] = 32'b00000000000000000000001100011010;
assign LUT_4[54143] = 32'b11111111111111111001011000010010;
assign LUT_4[54144] = 32'b00000000000000001111100111000100;
assign LUT_4[54145] = 32'b00000000000000001000110010111100;
assign LUT_4[54146] = 32'b00000000000000001111000001101000;
assign LUT_4[54147] = 32'b00000000000000001000001101100000;
assign LUT_4[54148] = 32'b00000000000000001100100111100000;
assign LUT_4[54149] = 32'b00000000000000000101110011011000;
assign LUT_4[54150] = 32'b00000000000000001100000010000100;
assign LUT_4[54151] = 32'b00000000000000000101001101111100;
assign LUT_4[54152] = 32'b00000000000000001000110011011001;
assign LUT_4[54153] = 32'b00000000000000000001111111010001;
assign LUT_4[54154] = 32'b00000000000000001000001101111101;
assign LUT_4[54155] = 32'b00000000000000000001011001110101;
assign LUT_4[54156] = 32'b00000000000000000101110011110101;
assign LUT_4[54157] = 32'b11111111111111111110111111101101;
assign LUT_4[54158] = 32'b00000000000000000101001110011001;
assign LUT_4[54159] = 32'b11111111111111111110011010010001;
assign LUT_4[54160] = 32'b00000000000000001101011000110010;
assign LUT_4[54161] = 32'b00000000000000000110100100101010;
assign LUT_4[54162] = 32'b00000000000000001100110011010110;
assign LUT_4[54163] = 32'b00000000000000000101111111001110;
assign LUT_4[54164] = 32'b00000000000000001010011001001110;
assign LUT_4[54165] = 32'b00000000000000000011100101000110;
assign LUT_4[54166] = 32'b00000000000000001001110011110010;
assign LUT_4[54167] = 32'b00000000000000000010111111101010;
assign LUT_4[54168] = 32'b00000000000000000110100101000111;
assign LUT_4[54169] = 32'b11111111111111111111110000111111;
assign LUT_4[54170] = 32'b00000000000000000101111111101011;
assign LUT_4[54171] = 32'b11111111111111111111001011100011;
assign LUT_4[54172] = 32'b00000000000000000011100101100011;
assign LUT_4[54173] = 32'b11111111111111111100110001011011;
assign LUT_4[54174] = 32'b00000000000000000011000000000111;
assign LUT_4[54175] = 32'b11111111111111111100001011111111;
assign LUT_4[54176] = 32'b00000000000000001110000010001011;
assign LUT_4[54177] = 32'b00000000000000000111001110000011;
assign LUT_4[54178] = 32'b00000000000000001101011100101111;
assign LUT_4[54179] = 32'b00000000000000000110101000100111;
assign LUT_4[54180] = 32'b00000000000000001011000010100111;
assign LUT_4[54181] = 32'b00000000000000000100001110011111;
assign LUT_4[54182] = 32'b00000000000000001010011101001011;
assign LUT_4[54183] = 32'b00000000000000000011101001000011;
assign LUT_4[54184] = 32'b00000000000000000111001110100000;
assign LUT_4[54185] = 32'b00000000000000000000011010011000;
assign LUT_4[54186] = 32'b00000000000000000110101001000100;
assign LUT_4[54187] = 32'b11111111111111111111110100111100;
assign LUT_4[54188] = 32'b00000000000000000100001110111100;
assign LUT_4[54189] = 32'b11111111111111111101011010110100;
assign LUT_4[54190] = 32'b00000000000000000011101001100000;
assign LUT_4[54191] = 32'b11111111111111111100110101011000;
assign LUT_4[54192] = 32'b00000000000000001011110011111001;
assign LUT_4[54193] = 32'b00000000000000000100111111110001;
assign LUT_4[54194] = 32'b00000000000000001011001110011101;
assign LUT_4[54195] = 32'b00000000000000000100011010010101;
assign LUT_4[54196] = 32'b00000000000000001000110100010101;
assign LUT_4[54197] = 32'b00000000000000000010000000001101;
assign LUT_4[54198] = 32'b00000000000000001000001110111001;
assign LUT_4[54199] = 32'b00000000000000000001011010110001;
assign LUT_4[54200] = 32'b00000000000000000101000000001110;
assign LUT_4[54201] = 32'b11111111111111111110001100000110;
assign LUT_4[54202] = 32'b00000000000000000100011010110010;
assign LUT_4[54203] = 32'b11111111111111111101100110101010;
assign LUT_4[54204] = 32'b00000000000000000010000000101010;
assign LUT_4[54205] = 32'b11111111111111111011001100100010;
assign LUT_4[54206] = 32'b00000000000000000001011011001110;
assign LUT_4[54207] = 32'b11111111111111111010100111000110;
assign LUT_4[54208] = 32'b00000000000000010000111110011000;
assign LUT_4[54209] = 32'b00000000000000001010001010010000;
assign LUT_4[54210] = 32'b00000000000000010000011000111100;
assign LUT_4[54211] = 32'b00000000000000001001100100110100;
assign LUT_4[54212] = 32'b00000000000000001101111110110100;
assign LUT_4[54213] = 32'b00000000000000000111001010101100;
assign LUT_4[54214] = 32'b00000000000000001101011001011000;
assign LUT_4[54215] = 32'b00000000000000000110100101010000;
assign LUT_4[54216] = 32'b00000000000000001010001010101101;
assign LUT_4[54217] = 32'b00000000000000000011010110100101;
assign LUT_4[54218] = 32'b00000000000000001001100101010001;
assign LUT_4[54219] = 32'b00000000000000000010110001001001;
assign LUT_4[54220] = 32'b00000000000000000111001011001001;
assign LUT_4[54221] = 32'b00000000000000000000010111000001;
assign LUT_4[54222] = 32'b00000000000000000110100101101101;
assign LUT_4[54223] = 32'b11111111111111111111110001100101;
assign LUT_4[54224] = 32'b00000000000000001110110000000110;
assign LUT_4[54225] = 32'b00000000000000000111111011111110;
assign LUT_4[54226] = 32'b00000000000000001110001010101010;
assign LUT_4[54227] = 32'b00000000000000000111010110100010;
assign LUT_4[54228] = 32'b00000000000000001011110000100010;
assign LUT_4[54229] = 32'b00000000000000000100111100011010;
assign LUT_4[54230] = 32'b00000000000000001011001011000110;
assign LUT_4[54231] = 32'b00000000000000000100010110111110;
assign LUT_4[54232] = 32'b00000000000000000111111100011011;
assign LUT_4[54233] = 32'b00000000000000000001001000010011;
assign LUT_4[54234] = 32'b00000000000000000111010110111111;
assign LUT_4[54235] = 32'b00000000000000000000100010110111;
assign LUT_4[54236] = 32'b00000000000000000100111100110111;
assign LUT_4[54237] = 32'b11111111111111111110001000101111;
assign LUT_4[54238] = 32'b00000000000000000100010111011011;
assign LUT_4[54239] = 32'b11111111111111111101100011010011;
assign LUT_4[54240] = 32'b00000000000000001111011001011111;
assign LUT_4[54241] = 32'b00000000000000001000100101010111;
assign LUT_4[54242] = 32'b00000000000000001110110100000011;
assign LUT_4[54243] = 32'b00000000000000000111111111111011;
assign LUT_4[54244] = 32'b00000000000000001100011001111011;
assign LUT_4[54245] = 32'b00000000000000000101100101110011;
assign LUT_4[54246] = 32'b00000000000000001011110100011111;
assign LUT_4[54247] = 32'b00000000000000000101000000010111;
assign LUT_4[54248] = 32'b00000000000000001000100101110100;
assign LUT_4[54249] = 32'b00000000000000000001110001101100;
assign LUT_4[54250] = 32'b00000000000000001000000000011000;
assign LUT_4[54251] = 32'b00000000000000000001001100010000;
assign LUT_4[54252] = 32'b00000000000000000101100110010000;
assign LUT_4[54253] = 32'b11111111111111111110110010001000;
assign LUT_4[54254] = 32'b00000000000000000101000000110100;
assign LUT_4[54255] = 32'b11111111111111111110001100101100;
assign LUT_4[54256] = 32'b00000000000000001101001011001101;
assign LUT_4[54257] = 32'b00000000000000000110010111000101;
assign LUT_4[54258] = 32'b00000000000000001100100101110001;
assign LUT_4[54259] = 32'b00000000000000000101110001101001;
assign LUT_4[54260] = 32'b00000000000000001010001011101001;
assign LUT_4[54261] = 32'b00000000000000000011010111100001;
assign LUT_4[54262] = 32'b00000000000000001001100110001101;
assign LUT_4[54263] = 32'b00000000000000000010110010000101;
assign LUT_4[54264] = 32'b00000000000000000110010111100010;
assign LUT_4[54265] = 32'b11111111111111111111100011011010;
assign LUT_4[54266] = 32'b00000000000000000101110010000110;
assign LUT_4[54267] = 32'b11111111111111111110111101111110;
assign LUT_4[54268] = 32'b00000000000000000011010111111110;
assign LUT_4[54269] = 32'b11111111111111111100100011110110;
assign LUT_4[54270] = 32'b00000000000000000010110010100010;
assign LUT_4[54271] = 32'b11111111111111111011111110011010;
assign LUT_4[54272] = 32'b00000000000000001010101011110000;
assign LUT_4[54273] = 32'b00000000000000000011110111101000;
assign LUT_4[54274] = 32'b00000000000000001010000110010100;
assign LUT_4[54275] = 32'b00000000000000000011010010001100;
assign LUT_4[54276] = 32'b00000000000000000111101100001100;
assign LUT_4[54277] = 32'b00000000000000000000111000000100;
assign LUT_4[54278] = 32'b00000000000000000111000110110000;
assign LUT_4[54279] = 32'b00000000000000000000010010101000;
assign LUT_4[54280] = 32'b00000000000000000011111000000101;
assign LUT_4[54281] = 32'b11111111111111111101000011111101;
assign LUT_4[54282] = 32'b00000000000000000011010010101001;
assign LUT_4[54283] = 32'b11111111111111111100011110100001;
assign LUT_4[54284] = 32'b00000000000000000000111000100001;
assign LUT_4[54285] = 32'b11111111111111111010000100011001;
assign LUT_4[54286] = 32'b00000000000000000000010011000101;
assign LUT_4[54287] = 32'b11111111111111111001011110111101;
assign LUT_4[54288] = 32'b00000000000000001000011101011110;
assign LUT_4[54289] = 32'b00000000000000000001101001010110;
assign LUT_4[54290] = 32'b00000000000000000111111000000010;
assign LUT_4[54291] = 32'b00000000000000000001000011111010;
assign LUT_4[54292] = 32'b00000000000000000101011101111010;
assign LUT_4[54293] = 32'b11111111111111111110101001110010;
assign LUT_4[54294] = 32'b00000000000000000100111000011110;
assign LUT_4[54295] = 32'b11111111111111111110000100010110;
assign LUT_4[54296] = 32'b00000000000000000001101001110011;
assign LUT_4[54297] = 32'b11111111111111111010110101101011;
assign LUT_4[54298] = 32'b00000000000000000001000100010111;
assign LUT_4[54299] = 32'b11111111111111111010010000001111;
assign LUT_4[54300] = 32'b11111111111111111110101010001111;
assign LUT_4[54301] = 32'b11111111111111110111110110000111;
assign LUT_4[54302] = 32'b11111111111111111110000100110011;
assign LUT_4[54303] = 32'b11111111111111110111010000101011;
assign LUT_4[54304] = 32'b00000000000000001001000110110111;
assign LUT_4[54305] = 32'b00000000000000000010010010101111;
assign LUT_4[54306] = 32'b00000000000000001000100001011011;
assign LUT_4[54307] = 32'b00000000000000000001101101010011;
assign LUT_4[54308] = 32'b00000000000000000110000111010011;
assign LUT_4[54309] = 32'b11111111111111111111010011001011;
assign LUT_4[54310] = 32'b00000000000000000101100001110111;
assign LUT_4[54311] = 32'b11111111111111111110101101101111;
assign LUT_4[54312] = 32'b00000000000000000010010011001100;
assign LUT_4[54313] = 32'b11111111111111111011011111000100;
assign LUT_4[54314] = 32'b00000000000000000001101101110000;
assign LUT_4[54315] = 32'b11111111111111111010111001101000;
assign LUT_4[54316] = 32'b11111111111111111111010011101000;
assign LUT_4[54317] = 32'b11111111111111111000011111100000;
assign LUT_4[54318] = 32'b11111111111111111110101110001100;
assign LUT_4[54319] = 32'b11111111111111110111111010000100;
assign LUT_4[54320] = 32'b00000000000000000110111000100101;
assign LUT_4[54321] = 32'b00000000000000000000000100011101;
assign LUT_4[54322] = 32'b00000000000000000110010011001001;
assign LUT_4[54323] = 32'b11111111111111111111011111000001;
assign LUT_4[54324] = 32'b00000000000000000011111001000001;
assign LUT_4[54325] = 32'b11111111111111111101000100111001;
assign LUT_4[54326] = 32'b00000000000000000011010011100101;
assign LUT_4[54327] = 32'b11111111111111111100011111011101;
assign LUT_4[54328] = 32'b00000000000000000000000100111010;
assign LUT_4[54329] = 32'b11111111111111111001010000110010;
assign LUT_4[54330] = 32'b11111111111111111111011111011110;
assign LUT_4[54331] = 32'b11111111111111111000101011010110;
assign LUT_4[54332] = 32'b11111111111111111101000101010110;
assign LUT_4[54333] = 32'b11111111111111110110010001001110;
assign LUT_4[54334] = 32'b11111111111111111100011111111010;
assign LUT_4[54335] = 32'b11111111111111110101101011110010;
assign LUT_4[54336] = 32'b00000000000000001100000011000100;
assign LUT_4[54337] = 32'b00000000000000000101001110111100;
assign LUT_4[54338] = 32'b00000000000000001011011101101000;
assign LUT_4[54339] = 32'b00000000000000000100101001100000;
assign LUT_4[54340] = 32'b00000000000000001001000011100000;
assign LUT_4[54341] = 32'b00000000000000000010001111011000;
assign LUT_4[54342] = 32'b00000000000000001000011110000100;
assign LUT_4[54343] = 32'b00000000000000000001101001111100;
assign LUT_4[54344] = 32'b00000000000000000101001111011001;
assign LUT_4[54345] = 32'b11111111111111111110011011010001;
assign LUT_4[54346] = 32'b00000000000000000100101001111101;
assign LUT_4[54347] = 32'b11111111111111111101110101110101;
assign LUT_4[54348] = 32'b00000000000000000010001111110101;
assign LUT_4[54349] = 32'b11111111111111111011011011101101;
assign LUT_4[54350] = 32'b00000000000000000001101010011001;
assign LUT_4[54351] = 32'b11111111111111111010110110010001;
assign LUT_4[54352] = 32'b00000000000000001001110100110010;
assign LUT_4[54353] = 32'b00000000000000000011000000101010;
assign LUT_4[54354] = 32'b00000000000000001001001111010110;
assign LUT_4[54355] = 32'b00000000000000000010011011001110;
assign LUT_4[54356] = 32'b00000000000000000110110101001110;
assign LUT_4[54357] = 32'b00000000000000000000000001000110;
assign LUT_4[54358] = 32'b00000000000000000110001111110010;
assign LUT_4[54359] = 32'b11111111111111111111011011101010;
assign LUT_4[54360] = 32'b00000000000000000011000001000111;
assign LUT_4[54361] = 32'b11111111111111111100001100111111;
assign LUT_4[54362] = 32'b00000000000000000010011011101011;
assign LUT_4[54363] = 32'b11111111111111111011100111100011;
assign LUT_4[54364] = 32'b00000000000000000000000001100011;
assign LUT_4[54365] = 32'b11111111111111111001001101011011;
assign LUT_4[54366] = 32'b11111111111111111111011100000111;
assign LUT_4[54367] = 32'b11111111111111111000100111111111;
assign LUT_4[54368] = 32'b00000000000000001010011110001011;
assign LUT_4[54369] = 32'b00000000000000000011101010000011;
assign LUT_4[54370] = 32'b00000000000000001001111000101111;
assign LUT_4[54371] = 32'b00000000000000000011000100100111;
assign LUT_4[54372] = 32'b00000000000000000111011110100111;
assign LUT_4[54373] = 32'b00000000000000000000101010011111;
assign LUT_4[54374] = 32'b00000000000000000110111001001011;
assign LUT_4[54375] = 32'b00000000000000000000000101000011;
assign LUT_4[54376] = 32'b00000000000000000011101010100000;
assign LUT_4[54377] = 32'b11111111111111111100110110011000;
assign LUT_4[54378] = 32'b00000000000000000011000101000100;
assign LUT_4[54379] = 32'b11111111111111111100010000111100;
assign LUT_4[54380] = 32'b00000000000000000000101010111100;
assign LUT_4[54381] = 32'b11111111111111111001110110110100;
assign LUT_4[54382] = 32'b00000000000000000000000101100000;
assign LUT_4[54383] = 32'b11111111111111111001010001011000;
assign LUT_4[54384] = 32'b00000000000000001000001111111001;
assign LUT_4[54385] = 32'b00000000000000000001011011110001;
assign LUT_4[54386] = 32'b00000000000000000111101010011101;
assign LUT_4[54387] = 32'b00000000000000000000110110010101;
assign LUT_4[54388] = 32'b00000000000000000101010000010101;
assign LUT_4[54389] = 32'b11111111111111111110011100001101;
assign LUT_4[54390] = 32'b00000000000000000100101010111001;
assign LUT_4[54391] = 32'b11111111111111111101110110110001;
assign LUT_4[54392] = 32'b00000000000000000001011100001110;
assign LUT_4[54393] = 32'b11111111111111111010101000000110;
assign LUT_4[54394] = 32'b00000000000000000000110110110010;
assign LUT_4[54395] = 32'b11111111111111111010000010101010;
assign LUT_4[54396] = 32'b11111111111111111110011100101010;
assign LUT_4[54397] = 32'b11111111111111110111101000100010;
assign LUT_4[54398] = 32'b11111111111111111101110111001110;
assign LUT_4[54399] = 32'b11111111111111110111000011000110;
assign LUT_4[54400] = 32'b00000000000000001101010001111000;
assign LUT_4[54401] = 32'b00000000000000000110011101110000;
assign LUT_4[54402] = 32'b00000000000000001100101100011100;
assign LUT_4[54403] = 32'b00000000000000000101111000010100;
assign LUT_4[54404] = 32'b00000000000000001010010010010100;
assign LUT_4[54405] = 32'b00000000000000000011011110001100;
assign LUT_4[54406] = 32'b00000000000000001001101100111000;
assign LUT_4[54407] = 32'b00000000000000000010111000110000;
assign LUT_4[54408] = 32'b00000000000000000110011110001101;
assign LUT_4[54409] = 32'b11111111111111111111101010000101;
assign LUT_4[54410] = 32'b00000000000000000101111000110001;
assign LUT_4[54411] = 32'b11111111111111111111000100101001;
assign LUT_4[54412] = 32'b00000000000000000011011110101001;
assign LUT_4[54413] = 32'b11111111111111111100101010100001;
assign LUT_4[54414] = 32'b00000000000000000010111001001101;
assign LUT_4[54415] = 32'b11111111111111111100000101000101;
assign LUT_4[54416] = 32'b00000000000000001011000011100110;
assign LUT_4[54417] = 32'b00000000000000000100001111011110;
assign LUT_4[54418] = 32'b00000000000000001010011110001010;
assign LUT_4[54419] = 32'b00000000000000000011101010000010;
assign LUT_4[54420] = 32'b00000000000000001000000100000010;
assign LUT_4[54421] = 32'b00000000000000000001001111111010;
assign LUT_4[54422] = 32'b00000000000000000111011110100110;
assign LUT_4[54423] = 32'b00000000000000000000101010011110;
assign LUT_4[54424] = 32'b00000000000000000100001111111011;
assign LUT_4[54425] = 32'b11111111111111111101011011110011;
assign LUT_4[54426] = 32'b00000000000000000011101010011111;
assign LUT_4[54427] = 32'b11111111111111111100110110010111;
assign LUT_4[54428] = 32'b00000000000000000001010000010111;
assign LUT_4[54429] = 32'b11111111111111111010011100001111;
assign LUT_4[54430] = 32'b00000000000000000000101010111011;
assign LUT_4[54431] = 32'b11111111111111111001110110110011;
assign LUT_4[54432] = 32'b00000000000000001011101100111111;
assign LUT_4[54433] = 32'b00000000000000000100111000110111;
assign LUT_4[54434] = 32'b00000000000000001011000111100011;
assign LUT_4[54435] = 32'b00000000000000000100010011011011;
assign LUT_4[54436] = 32'b00000000000000001000101101011011;
assign LUT_4[54437] = 32'b00000000000000000001111001010011;
assign LUT_4[54438] = 32'b00000000000000001000000111111111;
assign LUT_4[54439] = 32'b00000000000000000001010011110111;
assign LUT_4[54440] = 32'b00000000000000000100111001010100;
assign LUT_4[54441] = 32'b11111111111111111110000101001100;
assign LUT_4[54442] = 32'b00000000000000000100010011111000;
assign LUT_4[54443] = 32'b11111111111111111101011111110000;
assign LUT_4[54444] = 32'b00000000000000000001111001110000;
assign LUT_4[54445] = 32'b11111111111111111011000101101000;
assign LUT_4[54446] = 32'b00000000000000000001010100010100;
assign LUT_4[54447] = 32'b11111111111111111010100000001100;
assign LUT_4[54448] = 32'b00000000000000001001011110101101;
assign LUT_4[54449] = 32'b00000000000000000010101010100101;
assign LUT_4[54450] = 32'b00000000000000001000111001010001;
assign LUT_4[54451] = 32'b00000000000000000010000101001001;
assign LUT_4[54452] = 32'b00000000000000000110011111001001;
assign LUT_4[54453] = 32'b11111111111111111111101011000001;
assign LUT_4[54454] = 32'b00000000000000000101111001101101;
assign LUT_4[54455] = 32'b11111111111111111111000101100101;
assign LUT_4[54456] = 32'b00000000000000000010101011000010;
assign LUT_4[54457] = 32'b11111111111111111011110110111010;
assign LUT_4[54458] = 32'b00000000000000000010000101100110;
assign LUT_4[54459] = 32'b11111111111111111011010001011110;
assign LUT_4[54460] = 32'b11111111111111111111101011011110;
assign LUT_4[54461] = 32'b11111111111111111000110111010110;
assign LUT_4[54462] = 32'b11111111111111111111000110000010;
assign LUT_4[54463] = 32'b11111111111111111000010001111010;
assign LUT_4[54464] = 32'b00000000000000001110101001001100;
assign LUT_4[54465] = 32'b00000000000000000111110101000100;
assign LUT_4[54466] = 32'b00000000000000001110000011110000;
assign LUT_4[54467] = 32'b00000000000000000111001111101000;
assign LUT_4[54468] = 32'b00000000000000001011101001101000;
assign LUT_4[54469] = 32'b00000000000000000100110101100000;
assign LUT_4[54470] = 32'b00000000000000001011000100001100;
assign LUT_4[54471] = 32'b00000000000000000100010000000100;
assign LUT_4[54472] = 32'b00000000000000000111110101100001;
assign LUT_4[54473] = 32'b00000000000000000001000001011001;
assign LUT_4[54474] = 32'b00000000000000000111010000000101;
assign LUT_4[54475] = 32'b00000000000000000000011011111101;
assign LUT_4[54476] = 32'b00000000000000000100110101111101;
assign LUT_4[54477] = 32'b11111111111111111110000001110101;
assign LUT_4[54478] = 32'b00000000000000000100010000100001;
assign LUT_4[54479] = 32'b11111111111111111101011100011001;
assign LUT_4[54480] = 32'b00000000000000001100011010111010;
assign LUT_4[54481] = 32'b00000000000000000101100110110010;
assign LUT_4[54482] = 32'b00000000000000001011110101011110;
assign LUT_4[54483] = 32'b00000000000000000101000001010110;
assign LUT_4[54484] = 32'b00000000000000001001011011010110;
assign LUT_4[54485] = 32'b00000000000000000010100111001110;
assign LUT_4[54486] = 32'b00000000000000001000110101111010;
assign LUT_4[54487] = 32'b00000000000000000010000001110010;
assign LUT_4[54488] = 32'b00000000000000000101100111001111;
assign LUT_4[54489] = 32'b11111111111111111110110011000111;
assign LUT_4[54490] = 32'b00000000000000000101000001110011;
assign LUT_4[54491] = 32'b11111111111111111110001101101011;
assign LUT_4[54492] = 32'b00000000000000000010100111101011;
assign LUT_4[54493] = 32'b11111111111111111011110011100011;
assign LUT_4[54494] = 32'b00000000000000000010000010001111;
assign LUT_4[54495] = 32'b11111111111111111011001110000111;
assign LUT_4[54496] = 32'b00000000000000001101000100010011;
assign LUT_4[54497] = 32'b00000000000000000110010000001011;
assign LUT_4[54498] = 32'b00000000000000001100011110110111;
assign LUT_4[54499] = 32'b00000000000000000101101010101111;
assign LUT_4[54500] = 32'b00000000000000001010000100101111;
assign LUT_4[54501] = 32'b00000000000000000011010000100111;
assign LUT_4[54502] = 32'b00000000000000001001011111010011;
assign LUT_4[54503] = 32'b00000000000000000010101011001011;
assign LUT_4[54504] = 32'b00000000000000000110010000101000;
assign LUT_4[54505] = 32'b11111111111111111111011100100000;
assign LUT_4[54506] = 32'b00000000000000000101101011001100;
assign LUT_4[54507] = 32'b11111111111111111110110111000100;
assign LUT_4[54508] = 32'b00000000000000000011010001000100;
assign LUT_4[54509] = 32'b11111111111111111100011100111100;
assign LUT_4[54510] = 32'b00000000000000000010101011101000;
assign LUT_4[54511] = 32'b11111111111111111011110111100000;
assign LUT_4[54512] = 32'b00000000000000001010110110000001;
assign LUT_4[54513] = 32'b00000000000000000100000001111001;
assign LUT_4[54514] = 32'b00000000000000001010010000100101;
assign LUT_4[54515] = 32'b00000000000000000011011100011101;
assign LUT_4[54516] = 32'b00000000000000000111110110011101;
assign LUT_4[54517] = 32'b00000000000000000001000010010101;
assign LUT_4[54518] = 32'b00000000000000000111010001000001;
assign LUT_4[54519] = 32'b00000000000000000000011100111001;
assign LUT_4[54520] = 32'b00000000000000000100000010010110;
assign LUT_4[54521] = 32'b11111111111111111101001110001110;
assign LUT_4[54522] = 32'b00000000000000000011011100111010;
assign LUT_4[54523] = 32'b11111111111111111100101000110010;
assign LUT_4[54524] = 32'b00000000000000000001000010110010;
assign LUT_4[54525] = 32'b11111111111111111010001110101010;
assign LUT_4[54526] = 32'b00000000000000000000011101010110;
assign LUT_4[54527] = 32'b11111111111111111001101001001110;
assign LUT_4[54528] = 32'b00000000000000001111100111010011;
assign LUT_4[54529] = 32'b00000000000000001000110011001011;
assign LUT_4[54530] = 32'b00000000000000001111000001110111;
assign LUT_4[54531] = 32'b00000000000000001000001101101111;
assign LUT_4[54532] = 32'b00000000000000001100100111101111;
assign LUT_4[54533] = 32'b00000000000000000101110011100111;
assign LUT_4[54534] = 32'b00000000000000001100000010010011;
assign LUT_4[54535] = 32'b00000000000000000101001110001011;
assign LUT_4[54536] = 32'b00000000000000001000110011101000;
assign LUT_4[54537] = 32'b00000000000000000001111111100000;
assign LUT_4[54538] = 32'b00000000000000001000001110001100;
assign LUT_4[54539] = 32'b00000000000000000001011010000100;
assign LUT_4[54540] = 32'b00000000000000000101110100000100;
assign LUT_4[54541] = 32'b11111111111111111110111111111100;
assign LUT_4[54542] = 32'b00000000000000000101001110101000;
assign LUT_4[54543] = 32'b11111111111111111110011010100000;
assign LUT_4[54544] = 32'b00000000000000001101011001000001;
assign LUT_4[54545] = 32'b00000000000000000110100100111001;
assign LUT_4[54546] = 32'b00000000000000001100110011100101;
assign LUT_4[54547] = 32'b00000000000000000101111111011101;
assign LUT_4[54548] = 32'b00000000000000001010011001011101;
assign LUT_4[54549] = 32'b00000000000000000011100101010101;
assign LUT_4[54550] = 32'b00000000000000001001110100000001;
assign LUT_4[54551] = 32'b00000000000000000010111111111001;
assign LUT_4[54552] = 32'b00000000000000000110100101010110;
assign LUT_4[54553] = 32'b11111111111111111111110001001110;
assign LUT_4[54554] = 32'b00000000000000000101111111111010;
assign LUT_4[54555] = 32'b11111111111111111111001011110010;
assign LUT_4[54556] = 32'b00000000000000000011100101110010;
assign LUT_4[54557] = 32'b11111111111111111100110001101010;
assign LUT_4[54558] = 32'b00000000000000000011000000010110;
assign LUT_4[54559] = 32'b11111111111111111100001100001110;
assign LUT_4[54560] = 32'b00000000000000001110000010011010;
assign LUT_4[54561] = 32'b00000000000000000111001110010010;
assign LUT_4[54562] = 32'b00000000000000001101011100111110;
assign LUT_4[54563] = 32'b00000000000000000110101000110110;
assign LUT_4[54564] = 32'b00000000000000001011000010110110;
assign LUT_4[54565] = 32'b00000000000000000100001110101110;
assign LUT_4[54566] = 32'b00000000000000001010011101011010;
assign LUT_4[54567] = 32'b00000000000000000011101001010010;
assign LUT_4[54568] = 32'b00000000000000000111001110101111;
assign LUT_4[54569] = 32'b00000000000000000000011010100111;
assign LUT_4[54570] = 32'b00000000000000000110101001010011;
assign LUT_4[54571] = 32'b11111111111111111111110101001011;
assign LUT_4[54572] = 32'b00000000000000000100001111001011;
assign LUT_4[54573] = 32'b11111111111111111101011011000011;
assign LUT_4[54574] = 32'b00000000000000000011101001101111;
assign LUT_4[54575] = 32'b11111111111111111100110101100111;
assign LUT_4[54576] = 32'b00000000000000001011110100001000;
assign LUT_4[54577] = 32'b00000000000000000101000000000000;
assign LUT_4[54578] = 32'b00000000000000001011001110101100;
assign LUT_4[54579] = 32'b00000000000000000100011010100100;
assign LUT_4[54580] = 32'b00000000000000001000110100100100;
assign LUT_4[54581] = 32'b00000000000000000010000000011100;
assign LUT_4[54582] = 32'b00000000000000001000001111001000;
assign LUT_4[54583] = 32'b00000000000000000001011011000000;
assign LUT_4[54584] = 32'b00000000000000000101000000011101;
assign LUT_4[54585] = 32'b11111111111111111110001100010101;
assign LUT_4[54586] = 32'b00000000000000000100011011000001;
assign LUT_4[54587] = 32'b11111111111111111101100110111001;
assign LUT_4[54588] = 32'b00000000000000000010000000111001;
assign LUT_4[54589] = 32'b11111111111111111011001100110001;
assign LUT_4[54590] = 32'b00000000000000000001011011011101;
assign LUT_4[54591] = 32'b11111111111111111010100111010101;
assign LUT_4[54592] = 32'b00000000000000010000111110100111;
assign LUT_4[54593] = 32'b00000000000000001010001010011111;
assign LUT_4[54594] = 32'b00000000000000010000011001001011;
assign LUT_4[54595] = 32'b00000000000000001001100101000011;
assign LUT_4[54596] = 32'b00000000000000001101111111000011;
assign LUT_4[54597] = 32'b00000000000000000111001010111011;
assign LUT_4[54598] = 32'b00000000000000001101011001100111;
assign LUT_4[54599] = 32'b00000000000000000110100101011111;
assign LUT_4[54600] = 32'b00000000000000001010001010111100;
assign LUT_4[54601] = 32'b00000000000000000011010110110100;
assign LUT_4[54602] = 32'b00000000000000001001100101100000;
assign LUT_4[54603] = 32'b00000000000000000010110001011000;
assign LUT_4[54604] = 32'b00000000000000000111001011011000;
assign LUT_4[54605] = 32'b00000000000000000000010111010000;
assign LUT_4[54606] = 32'b00000000000000000110100101111100;
assign LUT_4[54607] = 32'b11111111111111111111110001110100;
assign LUT_4[54608] = 32'b00000000000000001110110000010101;
assign LUT_4[54609] = 32'b00000000000000000111111100001101;
assign LUT_4[54610] = 32'b00000000000000001110001010111001;
assign LUT_4[54611] = 32'b00000000000000000111010110110001;
assign LUT_4[54612] = 32'b00000000000000001011110000110001;
assign LUT_4[54613] = 32'b00000000000000000100111100101001;
assign LUT_4[54614] = 32'b00000000000000001011001011010101;
assign LUT_4[54615] = 32'b00000000000000000100010111001101;
assign LUT_4[54616] = 32'b00000000000000000111111100101010;
assign LUT_4[54617] = 32'b00000000000000000001001000100010;
assign LUT_4[54618] = 32'b00000000000000000111010111001110;
assign LUT_4[54619] = 32'b00000000000000000000100011000110;
assign LUT_4[54620] = 32'b00000000000000000100111101000110;
assign LUT_4[54621] = 32'b11111111111111111110001000111110;
assign LUT_4[54622] = 32'b00000000000000000100010111101010;
assign LUT_4[54623] = 32'b11111111111111111101100011100010;
assign LUT_4[54624] = 32'b00000000000000001111011001101110;
assign LUT_4[54625] = 32'b00000000000000001000100101100110;
assign LUT_4[54626] = 32'b00000000000000001110110100010010;
assign LUT_4[54627] = 32'b00000000000000001000000000001010;
assign LUT_4[54628] = 32'b00000000000000001100011010001010;
assign LUT_4[54629] = 32'b00000000000000000101100110000010;
assign LUT_4[54630] = 32'b00000000000000001011110100101110;
assign LUT_4[54631] = 32'b00000000000000000101000000100110;
assign LUT_4[54632] = 32'b00000000000000001000100110000011;
assign LUT_4[54633] = 32'b00000000000000000001110001111011;
assign LUT_4[54634] = 32'b00000000000000001000000000100111;
assign LUT_4[54635] = 32'b00000000000000000001001100011111;
assign LUT_4[54636] = 32'b00000000000000000101100110011111;
assign LUT_4[54637] = 32'b11111111111111111110110010010111;
assign LUT_4[54638] = 32'b00000000000000000101000001000011;
assign LUT_4[54639] = 32'b11111111111111111110001100111011;
assign LUT_4[54640] = 32'b00000000000000001101001011011100;
assign LUT_4[54641] = 32'b00000000000000000110010111010100;
assign LUT_4[54642] = 32'b00000000000000001100100110000000;
assign LUT_4[54643] = 32'b00000000000000000101110001111000;
assign LUT_4[54644] = 32'b00000000000000001010001011111000;
assign LUT_4[54645] = 32'b00000000000000000011010111110000;
assign LUT_4[54646] = 32'b00000000000000001001100110011100;
assign LUT_4[54647] = 32'b00000000000000000010110010010100;
assign LUT_4[54648] = 32'b00000000000000000110010111110001;
assign LUT_4[54649] = 32'b11111111111111111111100011101001;
assign LUT_4[54650] = 32'b00000000000000000101110010010101;
assign LUT_4[54651] = 32'b11111111111111111110111110001101;
assign LUT_4[54652] = 32'b00000000000000000011011000001101;
assign LUT_4[54653] = 32'b11111111111111111100100100000101;
assign LUT_4[54654] = 32'b00000000000000000010110010110001;
assign LUT_4[54655] = 32'b11111111111111111011111110101001;
assign LUT_4[54656] = 32'b00000000000000010010001101011011;
assign LUT_4[54657] = 32'b00000000000000001011011001010011;
assign LUT_4[54658] = 32'b00000000000000010001100111111111;
assign LUT_4[54659] = 32'b00000000000000001010110011110111;
assign LUT_4[54660] = 32'b00000000000000001111001101110111;
assign LUT_4[54661] = 32'b00000000000000001000011001101111;
assign LUT_4[54662] = 32'b00000000000000001110101000011011;
assign LUT_4[54663] = 32'b00000000000000000111110100010011;
assign LUT_4[54664] = 32'b00000000000000001011011001110000;
assign LUT_4[54665] = 32'b00000000000000000100100101101000;
assign LUT_4[54666] = 32'b00000000000000001010110100010100;
assign LUT_4[54667] = 32'b00000000000000000100000000001100;
assign LUT_4[54668] = 32'b00000000000000001000011010001100;
assign LUT_4[54669] = 32'b00000000000000000001100110000100;
assign LUT_4[54670] = 32'b00000000000000000111110100110000;
assign LUT_4[54671] = 32'b00000000000000000001000000101000;
assign LUT_4[54672] = 32'b00000000000000001111111111001001;
assign LUT_4[54673] = 32'b00000000000000001001001011000001;
assign LUT_4[54674] = 32'b00000000000000001111011001101101;
assign LUT_4[54675] = 32'b00000000000000001000100101100101;
assign LUT_4[54676] = 32'b00000000000000001100111111100101;
assign LUT_4[54677] = 32'b00000000000000000110001011011101;
assign LUT_4[54678] = 32'b00000000000000001100011010001001;
assign LUT_4[54679] = 32'b00000000000000000101100110000001;
assign LUT_4[54680] = 32'b00000000000000001001001011011110;
assign LUT_4[54681] = 32'b00000000000000000010010111010110;
assign LUT_4[54682] = 32'b00000000000000001000100110000010;
assign LUT_4[54683] = 32'b00000000000000000001110001111010;
assign LUT_4[54684] = 32'b00000000000000000110001011111010;
assign LUT_4[54685] = 32'b11111111111111111111010111110010;
assign LUT_4[54686] = 32'b00000000000000000101100110011110;
assign LUT_4[54687] = 32'b11111111111111111110110010010110;
assign LUT_4[54688] = 32'b00000000000000010000101000100010;
assign LUT_4[54689] = 32'b00000000000000001001110100011010;
assign LUT_4[54690] = 32'b00000000000000010000000011000110;
assign LUT_4[54691] = 32'b00000000000000001001001110111110;
assign LUT_4[54692] = 32'b00000000000000001101101000111110;
assign LUT_4[54693] = 32'b00000000000000000110110100110110;
assign LUT_4[54694] = 32'b00000000000000001101000011100010;
assign LUT_4[54695] = 32'b00000000000000000110001111011010;
assign LUT_4[54696] = 32'b00000000000000001001110100110111;
assign LUT_4[54697] = 32'b00000000000000000011000000101111;
assign LUT_4[54698] = 32'b00000000000000001001001111011011;
assign LUT_4[54699] = 32'b00000000000000000010011011010011;
assign LUT_4[54700] = 32'b00000000000000000110110101010011;
assign LUT_4[54701] = 32'b00000000000000000000000001001011;
assign LUT_4[54702] = 32'b00000000000000000110001111110111;
assign LUT_4[54703] = 32'b11111111111111111111011011101111;
assign LUT_4[54704] = 32'b00000000000000001110011010010000;
assign LUT_4[54705] = 32'b00000000000000000111100110001000;
assign LUT_4[54706] = 32'b00000000000000001101110100110100;
assign LUT_4[54707] = 32'b00000000000000000111000000101100;
assign LUT_4[54708] = 32'b00000000000000001011011010101100;
assign LUT_4[54709] = 32'b00000000000000000100100110100100;
assign LUT_4[54710] = 32'b00000000000000001010110101010000;
assign LUT_4[54711] = 32'b00000000000000000100000001001000;
assign LUT_4[54712] = 32'b00000000000000000111100110100101;
assign LUT_4[54713] = 32'b00000000000000000000110010011101;
assign LUT_4[54714] = 32'b00000000000000000111000001001001;
assign LUT_4[54715] = 32'b00000000000000000000001101000001;
assign LUT_4[54716] = 32'b00000000000000000100100111000001;
assign LUT_4[54717] = 32'b11111111111111111101110010111001;
assign LUT_4[54718] = 32'b00000000000000000100000001100101;
assign LUT_4[54719] = 32'b11111111111111111101001101011101;
assign LUT_4[54720] = 32'b00000000000000010011100100101111;
assign LUT_4[54721] = 32'b00000000000000001100110000100111;
assign LUT_4[54722] = 32'b00000000000000010010111111010011;
assign LUT_4[54723] = 32'b00000000000000001100001011001011;
assign LUT_4[54724] = 32'b00000000000000010000100101001011;
assign LUT_4[54725] = 32'b00000000000000001001110001000011;
assign LUT_4[54726] = 32'b00000000000000001111111111101111;
assign LUT_4[54727] = 32'b00000000000000001001001011100111;
assign LUT_4[54728] = 32'b00000000000000001100110001000100;
assign LUT_4[54729] = 32'b00000000000000000101111100111100;
assign LUT_4[54730] = 32'b00000000000000001100001011101000;
assign LUT_4[54731] = 32'b00000000000000000101010111100000;
assign LUT_4[54732] = 32'b00000000000000001001110001100000;
assign LUT_4[54733] = 32'b00000000000000000010111101011000;
assign LUT_4[54734] = 32'b00000000000000001001001100000100;
assign LUT_4[54735] = 32'b00000000000000000010010111111100;
assign LUT_4[54736] = 32'b00000000000000010001010110011101;
assign LUT_4[54737] = 32'b00000000000000001010100010010101;
assign LUT_4[54738] = 32'b00000000000000010000110001000001;
assign LUT_4[54739] = 32'b00000000000000001001111100111001;
assign LUT_4[54740] = 32'b00000000000000001110010110111001;
assign LUT_4[54741] = 32'b00000000000000000111100010110001;
assign LUT_4[54742] = 32'b00000000000000001101110001011101;
assign LUT_4[54743] = 32'b00000000000000000110111101010101;
assign LUT_4[54744] = 32'b00000000000000001010100010110010;
assign LUT_4[54745] = 32'b00000000000000000011101110101010;
assign LUT_4[54746] = 32'b00000000000000001001111101010110;
assign LUT_4[54747] = 32'b00000000000000000011001001001110;
assign LUT_4[54748] = 32'b00000000000000000111100011001110;
assign LUT_4[54749] = 32'b00000000000000000000101111000110;
assign LUT_4[54750] = 32'b00000000000000000110111101110010;
assign LUT_4[54751] = 32'b00000000000000000000001001101010;
assign LUT_4[54752] = 32'b00000000000000010001111111110110;
assign LUT_4[54753] = 32'b00000000000000001011001011101110;
assign LUT_4[54754] = 32'b00000000000000010001011010011010;
assign LUT_4[54755] = 32'b00000000000000001010100110010010;
assign LUT_4[54756] = 32'b00000000000000001111000000010010;
assign LUT_4[54757] = 32'b00000000000000001000001100001010;
assign LUT_4[54758] = 32'b00000000000000001110011010110110;
assign LUT_4[54759] = 32'b00000000000000000111100110101110;
assign LUT_4[54760] = 32'b00000000000000001011001100001011;
assign LUT_4[54761] = 32'b00000000000000000100011000000011;
assign LUT_4[54762] = 32'b00000000000000001010100110101111;
assign LUT_4[54763] = 32'b00000000000000000011110010100111;
assign LUT_4[54764] = 32'b00000000000000001000001100100111;
assign LUT_4[54765] = 32'b00000000000000000001011000011111;
assign LUT_4[54766] = 32'b00000000000000000111100111001011;
assign LUT_4[54767] = 32'b00000000000000000000110011000011;
assign LUT_4[54768] = 32'b00000000000000001111110001100100;
assign LUT_4[54769] = 32'b00000000000000001000111101011100;
assign LUT_4[54770] = 32'b00000000000000001111001100001000;
assign LUT_4[54771] = 32'b00000000000000001000011000000000;
assign LUT_4[54772] = 32'b00000000000000001100110010000000;
assign LUT_4[54773] = 32'b00000000000000000101111101111000;
assign LUT_4[54774] = 32'b00000000000000001100001100100100;
assign LUT_4[54775] = 32'b00000000000000000101011000011100;
assign LUT_4[54776] = 32'b00000000000000001000111101111001;
assign LUT_4[54777] = 32'b00000000000000000010001001110001;
assign LUT_4[54778] = 32'b00000000000000001000011000011101;
assign LUT_4[54779] = 32'b00000000000000000001100100010101;
assign LUT_4[54780] = 32'b00000000000000000101111110010101;
assign LUT_4[54781] = 32'b11111111111111111111001010001101;
assign LUT_4[54782] = 32'b00000000000000000101011000111001;
assign LUT_4[54783] = 32'b11111111111111111110100100110001;
assign LUT_4[54784] = 32'b00000000000000001001101111111000;
assign LUT_4[54785] = 32'b00000000000000000010111011110000;
assign LUT_4[54786] = 32'b00000000000000001001001010011100;
assign LUT_4[54787] = 32'b00000000000000000010010110010100;
assign LUT_4[54788] = 32'b00000000000000000110110000010100;
assign LUT_4[54789] = 32'b11111111111111111111111100001100;
assign LUT_4[54790] = 32'b00000000000000000110001010111000;
assign LUT_4[54791] = 32'b11111111111111111111010110110000;
assign LUT_4[54792] = 32'b00000000000000000010111100001101;
assign LUT_4[54793] = 32'b11111111111111111100001000000101;
assign LUT_4[54794] = 32'b00000000000000000010010110110001;
assign LUT_4[54795] = 32'b11111111111111111011100010101001;
assign LUT_4[54796] = 32'b11111111111111111111111100101001;
assign LUT_4[54797] = 32'b11111111111111111001001000100001;
assign LUT_4[54798] = 32'b11111111111111111111010111001101;
assign LUT_4[54799] = 32'b11111111111111111000100011000101;
assign LUT_4[54800] = 32'b00000000000000000111100001100110;
assign LUT_4[54801] = 32'b00000000000000000000101101011110;
assign LUT_4[54802] = 32'b00000000000000000110111100001010;
assign LUT_4[54803] = 32'b00000000000000000000001000000010;
assign LUT_4[54804] = 32'b00000000000000000100100010000010;
assign LUT_4[54805] = 32'b11111111111111111101101101111010;
assign LUT_4[54806] = 32'b00000000000000000011111100100110;
assign LUT_4[54807] = 32'b11111111111111111101001000011110;
assign LUT_4[54808] = 32'b00000000000000000000101101111011;
assign LUT_4[54809] = 32'b11111111111111111001111001110011;
assign LUT_4[54810] = 32'b00000000000000000000001000011111;
assign LUT_4[54811] = 32'b11111111111111111001010100010111;
assign LUT_4[54812] = 32'b11111111111111111101101110010111;
assign LUT_4[54813] = 32'b11111111111111110110111010001111;
assign LUT_4[54814] = 32'b11111111111111111101001000111011;
assign LUT_4[54815] = 32'b11111111111111110110010100110011;
assign LUT_4[54816] = 32'b00000000000000001000001010111111;
assign LUT_4[54817] = 32'b00000000000000000001010110110111;
assign LUT_4[54818] = 32'b00000000000000000111100101100011;
assign LUT_4[54819] = 32'b00000000000000000000110001011011;
assign LUT_4[54820] = 32'b00000000000000000101001011011011;
assign LUT_4[54821] = 32'b11111111111111111110010111010011;
assign LUT_4[54822] = 32'b00000000000000000100100101111111;
assign LUT_4[54823] = 32'b11111111111111111101110001110111;
assign LUT_4[54824] = 32'b00000000000000000001010111010100;
assign LUT_4[54825] = 32'b11111111111111111010100011001100;
assign LUT_4[54826] = 32'b00000000000000000000110001111000;
assign LUT_4[54827] = 32'b11111111111111111001111101110000;
assign LUT_4[54828] = 32'b11111111111111111110010111110000;
assign LUT_4[54829] = 32'b11111111111111110111100011101000;
assign LUT_4[54830] = 32'b11111111111111111101110010010100;
assign LUT_4[54831] = 32'b11111111111111110110111110001100;
assign LUT_4[54832] = 32'b00000000000000000101111100101101;
assign LUT_4[54833] = 32'b11111111111111111111001000100101;
assign LUT_4[54834] = 32'b00000000000000000101010111010001;
assign LUT_4[54835] = 32'b11111111111111111110100011001001;
assign LUT_4[54836] = 32'b00000000000000000010111101001001;
assign LUT_4[54837] = 32'b11111111111111111100001001000001;
assign LUT_4[54838] = 32'b00000000000000000010010111101101;
assign LUT_4[54839] = 32'b11111111111111111011100011100101;
assign LUT_4[54840] = 32'b11111111111111111111001001000010;
assign LUT_4[54841] = 32'b11111111111111111000010100111010;
assign LUT_4[54842] = 32'b11111111111111111110100011100110;
assign LUT_4[54843] = 32'b11111111111111110111101111011110;
assign LUT_4[54844] = 32'b11111111111111111100001001011110;
assign LUT_4[54845] = 32'b11111111111111110101010101010110;
assign LUT_4[54846] = 32'b11111111111111111011100100000010;
assign LUT_4[54847] = 32'b11111111111111110100101111111010;
assign LUT_4[54848] = 32'b00000000000000001011000111001100;
assign LUT_4[54849] = 32'b00000000000000000100010011000100;
assign LUT_4[54850] = 32'b00000000000000001010100001110000;
assign LUT_4[54851] = 32'b00000000000000000011101101101000;
assign LUT_4[54852] = 32'b00000000000000001000000111101000;
assign LUT_4[54853] = 32'b00000000000000000001010011100000;
assign LUT_4[54854] = 32'b00000000000000000111100010001100;
assign LUT_4[54855] = 32'b00000000000000000000101110000100;
assign LUT_4[54856] = 32'b00000000000000000100010011100001;
assign LUT_4[54857] = 32'b11111111111111111101011111011001;
assign LUT_4[54858] = 32'b00000000000000000011101110000101;
assign LUT_4[54859] = 32'b11111111111111111100111001111101;
assign LUT_4[54860] = 32'b00000000000000000001010011111101;
assign LUT_4[54861] = 32'b11111111111111111010011111110101;
assign LUT_4[54862] = 32'b00000000000000000000101110100001;
assign LUT_4[54863] = 32'b11111111111111111001111010011001;
assign LUT_4[54864] = 32'b00000000000000001000111000111010;
assign LUT_4[54865] = 32'b00000000000000000010000100110010;
assign LUT_4[54866] = 32'b00000000000000001000010011011110;
assign LUT_4[54867] = 32'b00000000000000000001011111010110;
assign LUT_4[54868] = 32'b00000000000000000101111001010110;
assign LUT_4[54869] = 32'b11111111111111111111000101001110;
assign LUT_4[54870] = 32'b00000000000000000101010011111010;
assign LUT_4[54871] = 32'b11111111111111111110011111110010;
assign LUT_4[54872] = 32'b00000000000000000010000101001111;
assign LUT_4[54873] = 32'b11111111111111111011010001000111;
assign LUT_4[54874] = 32'b00000000000000000001011111110011;
assign LUT_4[54875] = 32'b11111111111111111010101011101011;
assign LUT_4[54876] = 32'b11111111111111111111000101101011;
assign LUT_4[54877] = 32'b11111111111111111000010001100011;
assign LUT_4[54878] = 32'b11111111111111111110100000001111;
assign LUT_4[54879] = 32'b11111111111111110111101100000111;
assign LUT_4[54880] = 32'b00000000000000001001100010010011;
assign LUT_4[54881] = 32'b00000000000000000010101110001011;
assign LUT_4[54882] = 32'b00000000000000001000111100110111;
assign LUT_4[54883] = 32'b00000000000000000010001000101111;
assign LUT_4[54884] = 32'b00000000000000000110100010101111;
assign LUT_4[54885] = 32'b11111111111111111111101110100111;
assign LUT_4[54886] = 32'b00000000000000000101111101010011;
assign LUT_4[54887] = 32'b11111111111111111111001001001011;
assign LUT_4[54888] = 32'b00000000000000000010101110101000;
assign LUT_4[54889] = 32'b11111111111111111011111010100000;
assign LUT_4[54890] = 32'b00000000000000000010001001001100;
assign LUT_4[54891] = 32'b11111111111111111011010101000100;
assign LUT_4[54892] = 32'b11111111111111111111101111000100;
assign LUT_4[54893] = 32'b11111111111111111000111010111100;
assign LUT_4[54894] = 32'b11111111111111111111001001101000;
assign LUT_4[54895] = 32'b11111111111111111000010101100000;
assign LUT_4[54896] = 32'b00000000000000000111010100000001;
assign LUT_4[54897] = 32'b00000000000000000000011111111001;
assign LUT_4[54898] = 32'b00000000000000000110101110100101;
assign LUT_4[54899] = 32'b11111111111111111111111010011101;
assign LUT_4[54900] = 32'b00000000000000000100010100011101;
assign LUT_4[54901] = 32'b11111111111111111101100000010101;
assign LUT_4[54902] = 32'b00000000000000000011101111000001;
assign LUT_4[54903] = 32'b11111111111111111100111010111001;
assign LUT_4[54904] = 32'b00000000000000000000100000010110;
assign LUT_4[54905] = 32'b11111111111111111001101100001110;
assign LUT_4[54906] = 32'b11111111111111111111111010111010;
assign LUT_4[54907] = 32'b11111111111111111001000110110010;
assign LUT_4[54908] = 32'b11111111111111111101100000110010;
assign LUT_4[54909] = 32'b11111111111111110110101100101010;
assign LUT_4[54910] = 32'b11111111111111111100111011010110;
assign LUT_4[54911] = 32'b11111111111111110110000111001110;
assign LUT_4[54912] = 32'b00000000000000001100010110000000;
assign LUT_4[54913] = 32'b00000000000000000101100001111000;
assign LUT_4[54914] = 32'b00000000000000001011110000100100;
assign LUT_4[54915] = 32'b00000000000000000100111100011100;
assign LUT_4[54916] = 32'b00000000000000001001010110011100;
assign LUT_4[54917] = 32'b00000000000000000010100010010100;
assign LUT_4[54918] = 32'b00000000000000001000110001000000;
assign LUT_4[54919] = 32'b00000000000000000001111100111000;
assign LUT_4[54920] = 32'b00000000000000000101100010010101;
assign LUT_4[54921] = 32'b11111111111111111110101110001101;
assign LUT_4[54922] = 32'b00000000000000000100111100111001;
assign LUT_4[54923] = 32'b11111111111111111110001000110001;
assign LUT_4[54924] = 32'b00000000000000000010100010110001;
assign LUT_4[54925] = 32'b11111111111111111011101110101001;
assign LUT_4[54926] = 32'b00000000000000000001111101010101;
assign LUT_4[54927] = 32'b11111111111111111011001001001101;
assign LUT_4[54928] = 32'b00000000000000001010000111101110;
assign LUT_4[54929] = 32'b00000000000000000011010011100110;
assign LUT_4[54930] = 32'b00000000000000001001100010010010;
assign LUT_4[54931] = 32'b00000000000000000010101110001010;
assign LUT_4[54932] = 32'b00000000000000000111001000001010;
assign LUT_4[54933] = 32'b00000000000000000000010100000010;
assign LUT_4[54934] = 32'b00000000000000000110100010101110;
assign LUT_4[54935] = 32'b11111111111111111111101110100110;
assign LUT_4[54936] = 32'b00000000000000000011010100000011;
assign LUT_4[54937] = 32'b11111111111111111100011111111011;
assign LUT_4[54938] = 32'b00000000000000000010101110100111;
assign LUT_4[54939] = 32'b11111111111111111011111010011111;
assign LUT_4[54940] = 32'b00000000000000000000010100011111;
assign LUT_4[54941] = 32'b11111111111111111001100000010111;
assign LUT_4[54942] = 32'b11111111111111111111101111000011;
assign LUT_4[54943] = 32'b11111111111111111000111010111011;
assign LUT_4[54944] = 32'b00000000000000001010110001000111;
assign LUT_4[54945] = 32'b00000000000000000011111100111111;
assign LUT_4[54946] = 32'b00000000000000001010001011101011;
assign LUT_4[54947] = 32'b00000000000000000011010111100011;
assign LUT_4[54948] = 32'b00000000000000000111110001100011;
assign LUT_4[54949] = 32'b00000000000000000000111101011011;
assign LUT_4[54950] = 32'b00000000000000000111001100000111;
assign LUT_4[54951] = 32'b00000000000000000000010111111111;
assign LUT_4[54952] = 32'b00000000000000000011111101011100;
assign LUT_4[54953] = 32'b11111111111111111101001001010100;
assign LUT_4[54954] = 32'b00000000000000000011011000000000;
assign LUT_4[54955] = 32'b11111111111111111100100011111000;
assign LUT_4[54956] = 32'b00000000000000000000111101111000;
assign LUT_4[54957] = 32'b11111111111111111010001001110000;
assign LUT_4[54958] = 32'b00000000000000000000011000011100;
assign LUT_4[54959] = 32'b11111111111111111001100100010100;
assign LUT_4[54960] = 32'b00000000000000001000100010110101;
assign LUT_4[54961] = 32'b00000000000000000001101110101101;
assign LUT_4[54962] = 32'b00000000000000000111111101011001;
assign LUT_4[54963] = 32'b00000000000000000001001001010001;
assign LUT_4[54964] = 32'b00000000000000000101100011010001;
assign LUT_4[54965] = 32'b11111111111111111110101111001001;
assign LUT_4[54966] = 32'b00000000000000000100111101110101;
assign LUT_4[54967] = 32'b11111111111111111110001001101101;
assign LUT_4[54968] = 32'b00000000000000000001101111001010;
assign LUT_4[54969] = 32'b11111111111111111010111011000010;
assign LUT_4[54970] = 32'b00000000000000000001001001101110;
assign LUT_4[54971] = 32'b11111111111111111010010101100110;
assign LUT_4[54972] = 32'b11111111111111111110101111100110;
assign LUT_4[54973] = 32'b11111111111111110111111011011110;
assign LUT_4[54974] = 32'b11111111111111111110001010001010;
assign LUT_4[54975] = 32'b11111111111111110111010110000010;
assign LUT_4[54976] = 32'b00000000000000001101101101010100;
assign LUT_4[54977] = 32'b00000000000000000110111001001100;
assign LUT_4[54978] = 32'b00000000000000001101000111111000;
assign LUT_4[54979] = 32'b00000000000000000110010011110000;
assign LUT_4[54980] = 32'b00000000000000001010101101110000;
assign LUT_4[54981] = 32'b00000000000000000011111001101000;
assign LUT_4[54982] = 32'b00000000000000001010001000010100;
assign LUT_4[54983] = 32'b00000000000000000011010100001100;
assign LUT_4[54984] = 32'b00000000000000000110111001101001;
assign LUT_4[54985] = 32'b00000000000000000000000101100001;
assign LUT_4[54986] = 32'b00000000000000000110010100001101;
assign LUT_4[54987] = 32'b11111111111111111111100000000101;
assign LUT_4[54988] = 32'b00000000000000000011111010000101;
assign LUT_4[54989] = 32'b11111111111111111101000101111101;
assign LUT_4[54990] = 32'b00000000000000000011010100101001;
assign LUT_4[54991] = 32'b11111111111111111100100000100001;
assign LUT_4[54992] = 32'b00000000000000001011011111000010;
assign LUT_4[54993] = 32'b00000000000000000100101010111010;
assign LUT_4[54994] = 32'b00000000000000001010111001100110;
assign LUT_4[54995] = 32'b00000000000000000100000101011110;
assign LUT_4[54996] = 32'b00000000000000001000011111011110;
assign LUT_4[54997] = 32'b00000000000000000001101011010110;
assign LUT_4[54998] = 32'b00000000000000000111111010000010;
assign LUT_4[54999] = 32'b00000000000000000001000101111010;
assign LUT_4[55000] = 32'b00000000000000000100101011010111;
assign LUT_4[55001] = 32'b11111111111111111101110111001111;
assign LUT_4[55002] = 32'b00000000000000000100000101111011;
assign LUT_4[55003] = 32'b11111111111111111101010001110011;
assign LUT_4[55004] = 32'b00000000000000000001101011110011;
assign LUT_4[55005] = 32'b11111111111111111010110111101011;
assign LUT_4[55006] = 32'b00000000000000000001000110010111;
assign LUT_4[55007] = 32'b11111111111111111010010010001111;
assign LUT_4[55008] = 32'b00000000000000001100001000011011;
assign LUT_4[55009] = 32'b00000000000000000101010100010011;
assign LUT_4[55010] = 32'b00000000000000001011100010111111;
assign LUT_4[55011] = 32'b00000000000000000100101110110111;
assign LUT_4[55012] = 32'b00000000000000001001001000110111;
assign LUT_4[55013] = 32'b00000000000000000010010100101111;
assign LUT_4[55014] = 32'b00000000000000001000100011011011;
assign LUT_4[55015] = 32'b00000000000000000001101111010011;
assign LUT_4[55016] = 32'b00000000000000000101010100110000;
assign LUT_4[55017] = 32'b11111111111111111110100000101000;
assign LUT_4[55018] = 32'b00000000000000000100101111010100;
assign LUT_4[55019] = 32'b11111111111111111101111011001100;
assign LUT_4[55020] = 32'b00000000000000000010010101001100;
assign LUT_4[55021] = 32'b11111111111111111011100001000100;
assign LUT_4[55022] = 32'b00000000000000000001101111110000;
assign LUT_4[55023] = 32'b11111111111111111010111011101000;
assign LUT_4[55024] = 32'b00000000000000001001111010001001;
assign LUT_4[55025] = 32'b00000000000000000011000110000001;
assign LUT_4[55026] = 32'b00000000000000001001010100101101;
assign LUT_4[55027] = 32'b00000000000000000010100000100101;
assign LUT_4[55028] = 32'b00000000000000000110111010100101;
assign LUT_4[55029] = 32'b00000000000000000000000110011101;
assign LUT_4[55030] = 32'b00000000000000000110010101001001;
assign LUT_4[55031] = 32'b11111111111111111111100001000001;
assign LUT_4[55032] = 32'b00000000000000000011000110011110;
assign LUT_4[55033] = 32'b11111111111111111100010010010110;
assign LUT_4[55034] = 32'b00000000000000000010100001000010;
assign LUT_4[55035] = 32'b11111111111111111011101100111010;
assign LUT_4[55036] = 32'b00000000000000000000000110111010;
assign LUT_4[55037] = 32'b11111111111111111001010010110010;
assign LUT_4[55038] = 32'b11111111111111111111100001011110;
assign LUT_4[55039] = 32'b11111111111111111000101101010110;
assign LUT_4[55040] = 32'b00000000000000001110101011011011;
assign LUT_4[55041] = 32'b00000000000000000111110111010011;
assign LUT_4[55042] = 32'b00000000000000001110000101111111;
assign LUT_4[55043] = 32'b00000000000000000111010001110111;
assign LUT_4[55044] = 32'b00000000000000001011101011110111;
assign LUT_4[55045] = 32'b00000000000000000100110111101111;
assign LUT_4[55046] = 32'b00000000000000001011000110011011;
assign LUT_4[55047] = 32'b00000000000000000100010010010011;
assign LUT_4[55048] = 32'b00000000000000000111110111110000;
assign LUT_4[55049] = 32'b00000000000000000001000011101000;
assign LUT_4[55050] = 32'b00000000000000000111010010010100;
assign LUT_4[55051] = 32'b00000000000000000000011110001100;
assign LUT_4[55052] = 32'b00000000000000000100111000001100;
assign LUT_4[55053] = 32'b11111111111111111110000100000100;
assign LUT_4[55054] = 32'b00000000000000000100010010110000;
assign LUT_4[55055] = 32'b11111111111111111101011110101000;
assign LUT_4[55056] = 32'b00000000000000001100011101001001;
assign LUT_4[55057] = 32'b00000000000000000101101001000001;
assign LUT_4[55058] = 32'b00000000000000001011110111101101;
assign LUT_4[55059] = 32'b00000000000000000101000011100101;
assign LUT_4[55060] = 32'b00000000000000001001011101100101;
assign LUT_4[55061] = 32'b00000000000000000010101001011101;
assign LUT_4[55062] = 32'b00000000000000001000111000001001;
assign LUT_4[55063] = 32'b00000000000000000010000100000001;
assign LUT_4[55064] = 32'b00000000000000000101101001011110;
assign LUT_4[55065] = 32'b11111111111111111110110101010110;
assign LUT_4[55066] = 32'b00000000000000000101000100000010;
assign LUT_4[55067] = 32'b11111111111111111110001111111010;
assign LUT_4[55068] = 32'b00000000000000000010101001111010;
assign LUT_4[55069] = 32'b11111111111111111011110101110010;
assign LUT_4[55070] = 32'b00000000000000000010000100011110;
assign LUT_4[55071] = 32'b11111111111111111011010000010110;
assign LUT_4[55072] = 32'b00000000000000001101000110100010;
assign LUT_4[55073] = 32'b00000000000000000110010010011010;
assign LUT_4[55074] = 32'b00000000000000001100100001000110;
assign LUT_4[55075] = 32'b00000000000000000101101100111110;
assign LUT_4[55076] = 32'b00000000000000001010000110111110;
assign LUT_4[55077] = 32'b00000000000000000011010010110110;
assign LUT_4[55078] = 32'b00000000000000001001100001100010;
assign LUT_4[55079] = 32'b00000000000000000010101101011010;
assign LUT_4[55080] = 32'b00000000000000000110010010110111;
assign LUT_4[55081] = 32'b11111111111111111111011110101111;
assign LUT_4[55082] = 32'b00000000000000000101101101011011;
assign LUT_4[55083] = 32'b11111111111111111110111001010011;
assign LUT_4[55084] = 32'b00000000000000000011010011010011;
assign LUT_4[55085] = 32'b11111111111111111100011111001011;
assign LUT_4[55086] = 32'b00000000000000000010101101110111;
assign LUT_4[55087] = 32'b11111111111111111011111001101111;
assign LUT_4[55088] = 32'b00000000000000001010111000010000;
assign LUT_4[55089] = 32'b00000000000000000100000100001000;
assign LUT_4[55090] = 32'b00000000000000001010010010110100;
assign LUT_4[55091] = 32'b00000000000000000011011110101100;
assign LUT_4[55092] = 32'b00000000000000000111111000101100;
assign LUT_4[55093] = 32'b00000000000000000001000100100100;
assign LUT_4[55094] = 32'b00000000000000000111010011010000;
assign LUT_4[55095] = 32'b00000000000000000000011111001000;
assign LUT_4[55096] = 32'b00000000000000000100000100100101;
assign LUT_4[55097] = 32'b11111111111111111101010000011101;
assign LUT_4[55098] = 32'b00000000000000000011011111001001;
assign LUT_4[55099] = 32'b11111111111111111100101011000001;
assign LUT_4[55100] = 32'b00000000000000000001000101000001;
assign LUT_4[55101] = 32'b11111111111111111010010000111001;
assign LUT_4[55102] = 32'b00000000000000000000011111100101;
assign LUT_4[55103] = 32'b11111111111111111001101011011101;
assign LUT_4[55104] = 32'b00000000000000010000000010101111;
assign LUT_4[55105] = 32'b00000000000000001001001110100111;
assign LUT_4[55106] = 32'b00000000000000001111011101010011;
assign LUT_4[55107] = 32'b00000000000000001000101001001011;
assign LUT_4[55108] = 32'b00000000000000001101000011001011;
assign LUT_4[55109] = 32'b00000000000000000110001111000011;
assign LUT_4[55110] = 32'b00000000000000001100011101101111;
assign LUT_4[55111] = 32'b00000000000000000101101001100111;
assign LUT_4[55112] = 32'b00000000000000001001001111000100;
assign LUT_4[55113] = 32'b00000000000000000010011010111100;
assign LUT_4[55114] = 32'b00000000000000001000101001101000;
assign LUT_4[55115] = 32'b00000000000000000001110101100000;
assign LUT_4[55116] = 32'b00000000000000000110001111100000;
assign LUT_4[55117] = 32'b11111111111111111111011011011000;
assign LUT_4[55118] = 32'b00000000000000000101101010000100;
assign LUT_4[55119] = 32'b11111111111111111110110101111100;
assign LUT_4[55120] = 32'b00000000000000001101110100011101;
assign LUT_4[55121] = 32'b00000000000000000111000000010101;
assign LUT_4[55122] = 32'b00000000000000001101001111000001;
assign LUT_4[55123] = 32'b00000000000000000110011010111001;
assign LUT_4[55124] = 32'b00000000000000001010110100111001;
assign LUT_4[55125] = 32'b00000000000000000100000000110001;
assign LUT_4[55126] = 32'b00000000000000001010001111011101;
assign LUT_4[55127] = 32'b00000000000000000011011011010101;
assign LUT_4[55128] = 32'b00000000000000000111000000110010;
assign LUT_4[55129] = 32'b00000000000000000000001100101010;
assign LUT_4[55130] = 32'b00000000000000000110011011010110;
assign LUT_4[55131] = 32'b11111111111111111111100111001110;
assign LUT_4[55132] = 32'b00000000000000000100000001001110;
assign LUT_4[55133] = 32'b11111111111111111101001101000110;
assign LUT_4[55134] = 32'b00000000000000000011011011110010;
assign LUT_4[55135] = 32'b11111111111111111100100111101010;
assign LUT_4[55136] = 32'b00000000000000001110011101110110;
assign LUT_4[55137] = 32'b00000000000000000111101001101110;
assign LUT_4[55138] = 32'b00000000000000001101111000011010;
assign LUT_4[55139] = 32'b00000000000000000111000100010010;
assign LUT_4[55140] = 32'b00000000000000001011011110010010;
assign LUT_4[55141] = 32'b00000000000000000100101010001010;
assign LUT_4[55142] = 32'b00000000000000001010111000110110;
assign LUT_4[55143] = 32'b00000000000000000100000100101110;
assign LUT_4[55144] = 32'b00000000000000000111101010001011;
assign LUT_4[55145] = 32'b00000000000000000000110110000011;
assign LUT_4[55146] = 32'b00000000000000000111000100101111;
assign LUT_4[55147] = 32'b00000000000000000000010000100111;
assign LUT_4[55148] = 32'b00000000000000000100101010100111;
assign LUT_4[55149] = 32'b11111111111111111101110110011111;
assign LUT_4[55150] = 32'b00000000000000000100000101001011;
assign LUT_4[55151] = 32'b11111111111111111101010001000011;
assign LUT_4[55152] = 32'b00000000000000001100001111100100;
assign LUT_4[55153] = 32'b00000000000000000101011011011100;
assign LUT_4[55154] = 32'b00000000000000001011101010001000;
assign LUT_4[55155] = 32'b00000000000000000100110110000000;
assign LUT_4[55156] = 32'b00000000000000001001010000000000;
assign LUT_4[55157] = 32'b00000000000000000010011011111000;
assign LUT_4[55158] = 32'b00000000000000001000101010100100;
assign LUT_4[55159] = 32'b00000000000000000001110110011100;
assign LUT_4[55160] = 32'b00000000000000000101011011111001;
assign LUT_4[55161] = 32'b11111111111111111110100111110001;
assign LUT_4[55162] = 32'b00000000000000000100110110011101;
assign LUT_4[55163] = 32'b11111111111111111110000010010101;
assign LUT_4[55164] = 32'b00000000000000000010011100010101;
assign LUT_4[55165] = 32'b11111111111111111011101000001101;
assign LUT_4[55166] = 32'b00000000000000000001110110111001;
assign LUT_4[55167] = 32'b11111111111111111011000010110001;
assign LUT_4[55168] = 32'b00000000000000010001010001100011;
assign LUT_4[55169] = 32'b00000000000000001010011101011011;
assign LUT_4[55170] = 32'b00000000000000010000101100000111;
assign LUT_4[55171] = 32'b00000000000000001001110111111111;
assign LUT_4[55172] = 32'b00000000000000001110010001111111;
assign LUT_4[55173] = 32'b00000000000000000111011101110111;
assign LUT_4[55174] = 32'b00000000000000001101101100100011;
assign LUT_4[55175] = 32'b00000000000000000110111000011011;
assign LUT_4[55176] = 32'b00000000000000001010011101111000;
assign LUT_4[55177] = 32'b00000000000000000011101001110000;
assign LUT_4[55178] = 32'b00000000000000001001111000011100;
assign LUT_4[55179] = 32'b00000000000000000011000100010100;
assign LUT_4[55180] = 32'b00000000000000000111011110010100;
assign LUT_4[55181] = 32'b00000000000000000000101010001100;
assign LUT_4[55182] = 32'b00000000000000000110111000111000;
assign LUT_4[55183] = 32'b00000000000000000000000100110000;
assign LUT_4[55184] = 32'b00000000000000001111000011010001;
assign LUT_4[55185] = 32'b00000000000000001000001111001001;
assign LUT_4[55186] = 32'b00000000000000001110011101110101;
assign LUT_4[55187] = 32'b00000000000000000111101001101101;
assign LUT_4[55188] = 32'b00000000000000001100000011101101;
assign LUT_4[55189] = 32'b00000000000000000101001111100101;
assign LUT_4[55190] = 32'b00000000000000001011011110010001;
assign LUT_4[55191] = 32'b00000000000000000100101010001001;
assign LUT_4[55192] = 32'b00000000000000001000001111100110;
assign LUT_4[55193] = 32'b00000000000000000001011011011110;
assign LUT_4[55194] = 32'b00000000000000000111101010001010;
assign LUT_4[55195] = 32'b00000000000000000000110110000010;
assign LUT_4[55196] = 32'b00000000000000000101010000000010;
assign LUT_4[55197] = 32'b11111111111111111110011011111010;
assign LUT_4[55198] = 32'b00000000000000000100101010100110;
assign LUT_4[55199] = 32'b11111111111111111101110110011110;
assign LUT_4[55200] = 32'b00000000000000001111101100101010;
assign LUT_4[55201] = 32'b00000000000000001000111000100010;
assign LUT_4[55202] = 32'b00000000000000001111000111001110;
assign LUT_4[55203] = 32'b00000000000000001000010011000110;
assign LUT_4[55204] = 32'b00000000000000001100101101000110;
assign LUT_4[55205] = 32'b00000000000000000101111000111110;
assign LUT_4[55206] = 32'b00000000000000001100000111101010;
assign LUT_4[55207] = 32'b00000000000000000101010011100010;
assign LUT_4[55208] = 32'b00000000000000001000111000111111;
assign LUT_4[55209] = 32'b00000000000000000010000100110111;
assign LUT_4[55210] = 32'b00000000000000001000010011100011;
assign LUT_4[55211] = 32'b00000000000000000001011111011011;
assign LUT_4[55212] = 32'b00000000000000000101111001011011;
assign LUT_4[55213] = 32'b11111111111111111111000101010011;
assign LUT_4[55214] = 32'b00000000000000000101010011111111;
assign LUT_4[55215] = 32'b11111111111111111110011111110111;
assign LUT_4[55216] = 32'b00000000000000001101011110011000;
assign LUT_4[55217] = 32'b00000000000000000110101010010000;
assign LUT_4[55218] = 32'b00000000000000001100111000111100;
assign LUT_4[55219] = 32'b00000000000000000110000100110100;
assign LUT_4[55220] = 32'b00000000000000001010011110110100;
assign LUT_4[55221] = 32'b00000000000000000011101010101100;
assign LUT_4[55222] = 32'b00000000000000001001111001011000;
assign LUT_4[55223] = 32'b00000000000000000011000101010000;
assign LUT_4[55224] = 32'b00000000000000000110101010101101;
assign LUT_4[55225] = 32'b11111111111111111111110110100101;
assign LUT_4[55226] = 32'b00000000000000000110000101010001;
assign LUT_4[55227] = 32'b11111111111111111111010001001001;
assign LUT_4[55228] = 32'b00000000000000000011101011001001;
assign LUT_4[55229] = 32'b11111111111111111100110111000001;
assign LUT_4[55230] = 32'b00000000000000000011000101101101;
assign LUT_4[55231] = 32'b11111111111111111100010001100101;
assign LUT_4[55232] = 32'b00000000000000010010101000110111;
assign LUT_4[55233] = 32'b00000000000000001011110100101111;
assign LUT_4[55234] = 32'b00000000000000010010000011011011;
assign LUT_4[55235] = 32'b00000000000000001011001111010011;
assign LUT_4[55236] = 32'b00000000000000001111101001010011;
assign LUT_4[55237] = 32'b00000000000000001000110101001011;
assign LUT_4[55238] = 32'b00000000000000001111000011110111;
assign LUT_4[55239] = 32'b00000000000000001000001111101111;
assign LUT_4[55240] = 32'b00000000000000001011110101001100;
assign LUT_4[55241] = 32'b00000000000000000101000001000100;
assign LUT_4[55242] = 32'b00000000000000001011001111110000;
assign LUT_4[55243] = 32'b00000000000000000100011011101000;
assign LUT_4[55244] = 32'b00000000000000001000110101101000;
assign LUT_4[55245] = 32'b00000000000000000010000001100000;
assign LUT_4[55246] = 32'b00000000000000001000010000001100;
assign LUT_4[55247] = 32'b00000000000000000001011100000100;
assign LUT_4[55248] = 32'b00000000000000010000011010100101;
assign LUT_4[55249] = 32'b00000000000000001001100110011101;
assign LUT_4[55250] = 32'b00000000000000001111110101001001;
assign LUT_4[55251] = 32'b00000000000000001001000001000001;
assign LUT_4[55252] = 32'b00000000000000001101011011000001;
assign LUT_4[55253] = 32'b00000000000000000110100110111001;
assign LUT_4[55254] = 32'b00000000000000001100110101100101;
assign LUT_4[55255] = 32'b00000000000000000110000001011101;
assign LUT_4[55256] = 32'b00000000000000001001100110111010;
assign LUT_4[55257] = 32'b00000000000000000010110010110010;
assign LUT_4[55258] = 32'b00000000000000001001000001011110;
assign LUT_4[55259] = 32'b00000000000000000010001101010110;
assign LUT_4[55260] = 32'b00000000000000000110100111010110;
assign LUT_4[55261] = 32'b11111111111111111111110011001110;
assign LUT_4[55262] = 32'b00000000000000000110000001111010;
assign LUT_4[55263] = 32'b11111111111111111111001101110010;
assign LUT_4[55264] = 32'b00000000000000010001000011111110;
assign LUT_4[55265] = 32'b00000000000000001010001111110110;
assign LUT_4[55266] = 32'b00000000000000010000011110100010;
assign LUT_4[55267] = 32'b00000000000000001001101010011010;
assign LUT_4[55268] = 32'b00000000000000001110000100011010;
assign LUT_4[55269] = 32'b00000000000000000111010000010010;
assign LUT_4[55270] = 32'b00000000000000001101011110111110;
assign LUT_4[55271] = 32'b00000000000000000110101010110110;
assign LUT_4[55272] = 32'b00000000000000001010010000010011;
assign LUT_4[55273] = 32'b00000000000000000011011100001011;
assign LUT_4[55274] = 32'b00000000000000001001101010110111;
assign LUT_4[55275] = 32'b00000000000000000010110110101111;
assign LUT_4[55276] = 32'b00000000000000000111010000101111;
assign LUT_4[55277] = 32'b00000000000000000000011100100111;
assign LUT_4[55278] = 32'b00000000000000000110101011010011;
assign LUT_4[55279] = 32'b11111111111111111111110111001011;
assign LUT_4[55280] = 32'b00000000000000001110110101101100;
assign LUT_4[55281] = 32'b00000000000000001000000001100100;
assign LUT_4[55282] = 32'b00000000000000001110010000010000;
assign LUT_4[55283] = 32'b00000000000000000111011100001000;
assign LUT_4[55284] = 32'b00000000000000001011110110001000;
assign LUT_4[55285] = 32'b00000000000000000101000010000000;
assign LUT_4[55286] = 32'b00000000000000001011010000101100;
assign LUT_4[55287] = 32'b00000000000000000100011100100100;
assign LUT_4[55288] = 32'b00000000000000001000000010000001;
assign LUT_4[55289] = 32'b00000000000000000001001101111001;
assign LUT_4[55290] = 32'b00000000000000000111011100100101;
assign LUT_4[55291] = 32'b00000000000000000000101000011101;
assign LUT_4[55292] = 32'b00000000000000000101000010011101;
assign LUT_4[55293] = 32'b11111111111111111110001110010101;
assign LUT_4[55294] = 32'b00000000000000000100011101000001;
assign LUT_4[55295] = 32'b11111111111111111101101000111001;
assign LUT_4[55296] = 32'b00000000000000000100100000011011;
assign LUT_4[55297] = 32'b11111111111111111101101100010011;
assign LUT_4[55298] = 32'b00000000000000000011111010111111;
assign LUT_4[55299] = 32'b11111111111111111101000110110111;
assign LUT_4[55300] = 32'b00000000000000000001100000110111;
assign LUT_4[55301] = 32'b11111111111111111010101100101111;
assign LUT_4[55302] = 32'b00000000000000000000111011011011;
assign LUT_4[55303] = 32'b11111111111111111010000111010011;
assign LUT_4[55304] = 32'b11111111111111111101101100110000;
assign LUT_4[55305] = 32'b11111111111111110110111000101000;
assign LUT_4[55306] = 32'b11111111111111111101000111010100;
assign LUT_4[55307] = 32'b11111111111111110110010011001100;
assign LUT_4[55308] = 32'b11111111111111111010101101001100;
assign LUT_4[55309] = 32'b11111111111111110011111001000100;
assign LUT_4[55310] = 32'b11111111111111111010000111110000;
assign LUT_4[55311] = 32'b11111111111111110011010011101000;
assign LUT_4[55312] = 32'b00000000000000000010010010001001;
assign LUT_4[55313] = 32'b11111111111111111011011110000001;
assign LUT_4[55314] = 32'b00000000000000000001101100101101;
assign LUT_4[55315] = 32'b11111111111111111010111000100101;
assign LUT_4[55316] = 32'b11111111111111111111010010100101;
assign LUT_4[55317] = 32'b11111111111111111000011110011101;
assign LUT_4[55318] = 32'b11111111111111111110101101001001;
assign LUT_4[55319] = 32'b11111111111111110111111001000001;
assign LUT_4[55320] = 32'b11111111111111111011011110011110;
assign LUT_4[55321] = 32'b11111111111111110100101010010110;
assign LUT_4[55322] = 32'b11111111111111111010111001000010;
assign LUT_4[55323] = 32'b11111111111111110100000100111010;
assign LUT_4[55324] = 32'b11111111111111111000011110111010;
assign LUT_4[55325] = 32'b11111111111111110001101010110010;
assign LUT_4[55326] = 32'b11111111111111110111111001011110;
assign LUT_4[55327] = 32'b11111111111111110001000101010110;
assign LUT_4[55328] = 32'b00000000000000000010111011100010;
assign LUT_4[55329] = 32'b11111111111111111100000111011010;
assign LUT_4[55330] = 32'b00000000000000000010010110000110;
assign LUT_4[55331] = 32'b11111111111111111011100001111110;
assign LUT_4[55332] = 32'b11111111111111111111111011111110;
assign LUT_4[55333] = 32'b11111111111111111001000111110110;
assign LUT_4[55334] = 32'b11111111111111111111010110100010;
assign LUT_4[55335] = 32'b11111111111111111000100010011010;
assign LUT_4[55336] = 32'b11111111111111111100000111110111;
assign LUT_4[55337] = 32'b11111111111111110101010011101111;
assign LUT_4[55338] = 32'b11111111111111111011100010011011;
assign LUT_4[55339] = 32'b11111111111111110100101110010011;
assign LUT_4[55340] = 32'b11111111111111111001001000010011;
assign LUT_4[55341] = 32'b11111111111111110010010100001011;
assign LUT_4[55342] = 32'b11111111111111111000100010110111;
assign LUT_4[55343] = 32'b11111111111111110001101110101111;
assign LUT_4[55344] = 32'b00000000000000000000101101010000;
assign LUT_4[55345] = 32'b11111111111111111001111001001000;
assign LUT_4[55346] = 32'b00000000000000000000000111110100;
assign LUT_4[55347] = 32'b11111111111111111001010011101100;
assign LUT_4[55348] = 32'b11111111111111111101101101101100;
assign LUT_4[55349] = 32'b11111111111111110110111001100100;
assign LUT_4[55350] = 32'b11111111111111111101001000010000;
assign LUT_4[55351] = 32'b11111111111111110110010100001000;
assign LUT_4[55352] = 32'b11111111111111111001111001100101;
assign LUT_4[55353] = 32'b11111111111111110011000101011101;
assign LUT_4[55354] = 32'b11111111111111111001010100001001;
assign LUT_4[55355] = 32'b11111111111111110010100000000001;
assign LUT_4[55356] = 32'b11111111111111110110111010000001;
assign LUT_4[55357] = 32'b11111111111111110000000101111001;
assign LUT_4[55358] = 32'b11111111111111110110010100100101;
assign LUT_4[55359] = 32'b11111111111111101111100000011101;
assign LUT_4[55360] = 32'b00000000000000000101110111101111;
assign LUT_4[55361] = 32'b11111111111111111111000011100111;
assign LUT_4[55362] = 32'b00000000000000000101010010010011;
assign LUT_4[55363] = 32'b11111111111111111110011110001011;
assign LUT_4[55364] = 32'b00000000000000000010111000001011;
assign LUT_4[55365] = 32'b11111111111111111100000100000011;
assign LUT_4[55366] = 32'b00000000000000000010010010101111;
assign LUT_4[55367] = 32'b11111111111111111011011110100111;
assign LUT_4[55368] = 32'b11111111111111111111000100000100;
assign LUT_4[55369] = 32'b11111111111111111000001111111100;
assign LUT_4[55370] = 32'b11111111111111111110011110101000;
assign LUT_4[55371] = 32'b11111111111111110111101010100000;
assign LUT_4[55372] = 32'b11111111111111111100000100100000;
assign LUT_4[55373] = 32'b11111111111111110101010000011000;
assign LUT_4[55374] = 32'b11111111111111111011011111000100;
assign LUT_4[55375] = 32'b11111111111111110100101010111100;
assign LUT_4[55376] = 32'b00000000000000000011101001011101;
assign LUT_4[55377] = 32'b11111111111111111100110101010101;
assign LUT_4[55378] = 32'b00000000000000000011000100000001;
assign LUT_4[55379] = 32'b11111111111111111100001111111001;
assign LUT_4[55380] = 32'b00000000000000000000101001111001;
assign LUT_4[55381] = 32'b11111111111111111001110101110001;
assign LUT_4[55382] = 32'b00000000000000000000000100011101;
assign LUT_4[55383] = 32'b11111111111111111001010000010101;
assign LUT_4[55384] = 32'b11111111111111111100110101110010;
assign LUT_4[55385] = 32'b11111111111111110110000001101010;
assign LUT_4[55386] = 32'b11111111111111111100010000010110;
assign LUT_4[55387] = 32'b11111111111111110101011100001110;
assign LUT_4[55388] = 32'b11111111111111111001110110001110;
assign LUT_4[55389] = 32'b11111111111111110011000010000110;
assign LUT_4[55390] = 32'b11111111111111111001010000110010;
assign LUT_4[55391] = 32'b11111111111111110010011100101010;
assign LUT_4[55392] = 32'b00000000000000000100010010110110;
assign LUT_4[55393] = 32'b11111111111111111101011110101110;
assign LUT_4[55394] = 32'b00000000000000000011101101011010;
assign LUT_4[55395] = 32'b11111111111111111100111001010010;
assign LUT_4[55396] = 32'b00000000000000000001010011010010;
assign LUT_4[55397] = 32'b11111111111111111010011111001010;
assign LUT_4[55398] = 32'b00000000000000000000101101110110;
assign LUT_4[55399] = 32'b11111111111111111001111001101110;
assign LUT_4[55400] = 32'b11111111111111111101011111001011;
assign LUT_4[55401] = 32'b11111111111111110110101011000011;
assign LUT_4[55402] = 32'b11111111111111111100111001101111;
assign LUT_4[55403] = 32'b11111111111111110110000101100111;
assign LUT_4[55404] = 32'b11111111111111111010011111100111;
assign LUT_4[55405] = 32'b11111111111111110011101011011111;
assign LUT_4[55406] = 32'b11111111111111111001111010001011;
assign LUT_4[55407] = 32'b11111111111111110011000110000011;
assign LUT_4[55408] = 32'b00000000000000000010000100100100;
assign LUT_4[55409] = 32'b11111111111111111011010000011100;
assign LUT_4[55410] = 32'b00000000000000000001011111001000;
assign LUT_4[55411] = 32'b11111111111111111010101011000000;
assign LUT_4[55412] = 32'b11111111111111111111000101000000;
assign LUT_4[55413] = 32'b11111111111111111000010000111000;
assign LUT_4[55414] = 32'b11111111111111111110011111100100;
assign LUT_4[55415] = 32'b11111111111111110111101011011100;
assign LUT_4[55416] = 32'b11111111111111111011010000111001;
assign LUT_4[55417] = 32'b11111111111111110100011100110001;
assign LUT_4[55418] = 32'b11111111111111111010101011011101;
assign LUT_4[55419] = 32'b11111111111111110011110111010101;
assign LUT_4[55420] = 32'b11111111111111111000010001010101;
assign LUT_4[55421] = 32'b11111111111111110001011101001101;
assign LUT_4[55422] = 32'b11111111111111110111101011111001;
assign LUT_4[55423] = 32'b11111111111111110000110111110001;
assign LUT_4[55424] = 32'b00000000000000000111000110100011;
assign LUT_4[55425] = 32'b00000000000000000000010010011011;
assign LUT_4[55426] = 32'b00000000000000000110100001000111;
assign LUT_4[55427] = 32'b11111111111111111111101100111111;
assign LUT_4[55428] = 32'b00000000000000000100000110111111;
assign LUT_4[55429] = 32'b11111111111111111101010010110111;
assign LUT_4[55430] = 32'b00000000000000000011100001100011;
assign LUT_4[55431] = 32'b11111111111111111100101101011011;
assign LUT_4[55432] = 32'b00000000000000000000010010111000;
assign LUT_4[55433] = 32'b11111111111111111001011110110000;
assign LUT_4[55434] = 32'b11111111111111111111101101011100;
assign LUT_4[55435] = 32'b11111111111111111000111001010100;
assign LUT_4[55436] = 32'b11111111111111111101010011010100;
assign LUT_4[55437] = 32'b11111111111111110110011111001100;
assign LUT_4[55438] = 32'b11111111111111111100101101111000;
assign LUT_4[55439] = 32'b11111111111111110101111001110000;
assign LUT_4[55440] = 32'b00000000000000000100111000010001;
assign LUT_4[55441] = 32'b11111111111111111110000100001001;
assign LUT_4[55442] = 32'b00000000000000000100010010110101;
assign LUT_4[55443] = 32'b11111111111111111101011110101101;
assign LUT_4[55444] = 32'b00000000000000000001111000101101;
assign LUT_4[55445] = 32'b11111111111111111011000100100101;
assign LUT_4[55446] = 32'b00000000000000000001010011010001;
assign LUT_4[55447] = 32'b11111111111111111010011111001001;
assign LUT_4[55448] = 32'b11111111111111111110000100100110;
assign LUT_4[55449] = 32'b11111111111111110111010000011110;
assign LUT_4[55450] = 32'b11111111111111111101011111001010;
assign LUT_4[55451] = 32'b11111111111111110110101011000010;
assign LUT_4[55452] = 32'b11111111111111111011000101000010;
assign LUT_4[55453] = 32'b11111111111111110100010000111010;
assign LUT_4[55454] = 32'b11111111111111111010011111100110;
assign LUT_4[55455] = 32'b11111111111111110011101011011110;
assign LUT_4[55456] = 32'b00000000000000000101100001101010;
assign LUT_4[55457] = 32'b11111111111111111110101101100010;
assign LUT_4[55458] = 32'b00000000000000000100111100001110;
assign LUT_4[55459] = 32'b11111111111111111110001000000110;
assign LUT_4[55460] = 32'b00000000000000000010100010000110;
assign LUT_4[55461] = 32'b11111111111111111011101101111110;
assign LUT_4[55462] = 32'b00000000000000000001111100101010;
assign LUT_4[55463] = 32'b11111111111111111011001000100010;
assign LUT_4[55464] = 32'b11111111111111111110101101111111;
assign LUT_4[55465] = 32'b11111111111111110111111001110111;
assign LUT_4[55466] = 32'b11111111111111111110001000100011;
assign LUT_4[55467] = 32'b11111111111111110111010100011011;
assign LUT_4[55468] = 32'b11111111111111111011101110011011;
assign LUT_4[55469] = 32'b11111111111111110100111010010011;
assign LUT_4[55470] = 32'b11111111111111111011001000111111;
assign LUT_4[55471] = 32'b11111111111111110100010100110111;
assign LUT_4[55472] = 32'b00000000000000000011010011011000;
assign LUT_4[55473] = 32'b11111111111111111100011111010000;
assign LUT_4[55474] = 32'b00000000000000000010101101111100;
assign LUT_4[55475] = 32'b11111111111111111011111001110100;
assign LUT_4[55476] = 32'b00000000000000000000010011110100;
assign LUT_4[55477] = 32'b11111111111111111001011111101100;
assign LUT_4[55478] = 32'b11111111111111111111101110011000;
assign LUT_4[55479] = 32'b11111111111111111000111010010000;
assign LUT_4[55480] = 32'b11111111111111111100011111101101;
assign LUT_4[55481] = 32'b11111111111111110101101011100101;
assign LUT_4[55482] = 32'b11111111111111111011111010010001;
assign LUT_4[55483] = 32'b11111111111111110101000110001001;
assign LUT_4[55484] = 32'b11111111111111111001100000001001;
assign LUT_4[55485] = 32'b11111111111111110010101100000001;
assign LUT_4[55486] = 32'b11111111111111111000111010101101;
assign LUT_4[55487] = 32'b11111111111111110010000110100101;
assign LUT_4[55488] = 32'b00000000000000001000011101110111;
assign LUT_4[55489] = 32'b00000000000000000001101001101111;
assign LUT_4[55490] = 32'b00000000000000000111111000011011;
assign LUT_4[55491] = 32'b00000000000000000001000100010011;
assign LUT_4[55492] = 32'b00000000000000000101011110010011;
assign LUT_4[55493] = 32'b11111111111111111110101010001011;
assign LUT_4[55494] = 32'b00000000000000000100111000110111;
assign LUT_4[55495] = 32'b11111111111111111110000100101111;
assign LUT_4[55496] = 32'b00000000000000000001101010001100;
assign LUT_4[55497] = 32'b11111111111111111010110110000100;
assign LUT_4[55498] = 32'b00000000000000000001000100110000;
assign LUT_4[55499] = 32'b11111111111111111010010000101000;
assign LUT_4[55500] = 32'b11111111111111111110101010101000;
assign LUT_4[55501] = 32'b11111111111111110111110110100000;
assign LUT_4[55502] = 32'b11111111111111111110000101001100;
assign LUT_4[55503] = 32'b11111111111111110111010001000100;
assign LUT_4[55504] = 32'b00000000000000000110001111100101;
assign LUT_4[55505] = 32'b11111111111111111111011011011101;
assign LUT_4[55506] = 32'b00000000000000000101101010001001;
assign LUT_4[55507] = 32'b11111111111111111110110110000001;
assign LUT_4[55508] = 32'b00000000000000000011010000000001;
assign LUT_4[55509] = 32'b11111111111111111100011011111001;
assign LUT_4[55510] = 32'b00000000000000000010101010100101;
assign LUT_4[55511] = 32'b11111111111111111011110110011101;
assign LUT_4[55512] = 32'b11111111111111111111011011111010;
assign LUT_4[55513] = 32'b11111111111111111000100111110010;
assign LUT_4[55514] = 32'b11111111111111111110110110011110;
assign LUT_4[55515] = 32'b11111111111111111000000010010110;
assign LUT_4[55516] = 32'b11111111111111111100011100010110;
assign LUT_4[55517] = 32'b11111111111111110101101000001110;
assign LUT_4[55518] = 32'b11111111111111111011110110111010;
assign LUT_4[55519] = 32'b11111111111111110101000010110010;
assign LUT_4[55520] = 32'b00000000000000000110111000111110;
assign LUT_4[55521] = 32'b00000000000000000000000100110110;
assign LUT_4[55522] = 32'b00000000000000000110010011100010;
assign LUT_4[55523] = 32'b11111111111111111111011111011010;
assign LUT_4[55524] = 32'b00000000000000000011111001011010;
assign LUT_4[55525] = 32'b11111111111111111101000101010010;
assign LUT_4[55526] = 32'b00000000000000000011010011111110;
assign LUT_4[55527] = 32'b11111111111111111100011111110110;
assign LUT_4[55528] = 32'b00000000000000000000000101010011;
assign LUT_4[55529] = 32'b11111111111111111001010001001011;
assign LUT_4[55530] = 32'b11111111111111111111011111110111;
assign LUT_4[55531] = 32'b11111111111111111000101011101111;
assign LUT_4[55532] = 32'b11111111111111111101000101101111;
assign LUT_4[55533] = 32'b11111111111111110110010001100111;
assign LUT_4[55534] = 32'b11111111111111111100100000010011;
assign LUT_4[55535] = 32'b11111111111111110101101100001011;
assign LUT_4[55536] = 32'b00000000000000000100101010101100;
assign LUT_4[55537] = 32'b11111111111111111101110110100100;
assign LUT_4[55538] = 32'b00000000000000000100000101010000;
assign LUT_4[55539] = 32'b11111111111111111101010001001000;
assign LUT_4[55540] = 32'b00000000000000000001101011001000;
assign LUT_4[55541] = 32'b11111111111111111010110111000000;
assign LUT_4[55542] = 32'b00000000000000000001000101101100;
assign LUT_4[55543] = 32'b11111111111111111010010001100100;
assign LUT_4[55544] = 32'b11111111111111111101110111000001;
assign LUT_4[55545] = 32'b11111111111111110111000010111001;
assign LUT_4[55546] = 32'b11111111111111111101010001100101;
assign LUT_4[55547] = 32'b11111111111111110110011101011101;
assign LUT_4[55548] = 32'b11111111111111111010110111011101;
assign LUT_4[55549] = 32'b11111111111111110100000011010101;
assign LUT_4[55550] = 32'b11111111111111111010010010000001;
assign LUT_4[55551] = 32'b11111111111111110011011101111001;
assign LUT_4[55552] = 32'b00000000000000001001011011111110;
assign LUT_4[55553] = 32'b00000000000000000010100111110110;
assign LUT_4[55554] = 32'b00000000000000001000110110100010;
assign LUT_4[55555] = 32'b00000000000000000010000010011010;
assign LUT_4[55556] = 32'b00000000000000000110011100011010;
assign LUT_4[55557] = 32'b11111111111111111111101000010010;
assign LUT_4[55558] = 32'b00000000000000000101110110111110;
assign LUT_4[55559] = 32'b11111111111111111111000010110110;
assign LUT_4[55560] = 32'b00000000000000000010101000010011;
assign LUT_4[55561] = 32'b11111111111111111011110100001011;
assign LUT_4[55562] = 32'b00000000000000000010000010110111;
assign LUT_4[55563] = 32'b11111111111111111011001110101111;
assign LUT_4[55564] = 32'b11111111111111111111101000101111;
assign LUT_4[55565] = 32'b11111111111111111000110100100111;
assign LUT_4[55566] = 32'b11111111111111111111000011010011;
assign LUT_4[55567] = 32'b11111111111111111000001111001011;
assign LUT_4[55568] = 32'b00000000000000000111001101101100;
assign LUT_4[55569] = 32'b00000000000000000000011001100100;
assign LUT_4[55570] = 32'b00000000000000000110101000010000;
assign LUT_4[55571] = 32'b11111111111111111111110100001000;
assign LUT_4[55572] = 32'b00000000000000000100001110001000;
assign LUT_4[55573] = 32'b11111111111111111101011010000000;
assign LUT_4[55574] = 32'b00000000000000000011101000101100;
assign LUT_4[55575] = 32'b11111111111111111100110100100100;
assign LUT_4[55576] = 32'b00000000000000000000011010000001;
assign LUT_4[55577] = 32'b11111111111111111001100101111001;
assign LUT_4[55578] = 32'b11111111111111111111110100100101;
assign LUT_4[55579] = 32'b11111111111111111001000000011101;
assign LUT_4[55580] = 32'b11111111111111111101011010011101;
assign LUT_4[55581] = 32'b11111111111111110110100110010101;
assign LUT_4[55582] = 32'b11111111111111111100110101000001;
assign LUT_4[55583] = 32'b11111111111111110110000000111001;
assign LUT_4[55584] = 32'b00000000000000000111110111000101;
assign LUT_4[55585] = 32'b00000000000000000001000010111101;
assign LUT_4[55586] = 32'b00000000000000000111010001101001;
assign LUT_4[55587] = 32'b00000000000000000000011101100001;
assign LUT_4[55588] = 32'b00000000000000000100110111100001;
assign LUT_4[55589] = 32'b11111111111111111110000011011001;
assign LUT_4[55590] = 32'b00000000000000000100010010000101;
assign LUT_4[55591] = 32'b11111111111111111101011101111101;
assign LUT_4[55592] = 32'b00000000000000000001000011011010;
assign LUT_4[55593] = 32'b11111111111111111010001111010010;
assign LUT_4[55594] = 32'b00000000000000000000011101111110;
assign LUT_4[55595] = 32'b11111111111111111001101001110110;
assign LUT_4[55596] = 32'b11111111111111111110000011110110;
assign LUT_4[55597] = 32'b11111111111111110111001111101110;
assign LUT_4[55598] = 32'b11111111111111111101011110011010;
assign LUT_4[55599] = 32'b11111111111111110110101010010010;
assign LUT_4[55600] = 32'b00000000000000000101101000110011;
assign LUT_4[55601] = 32'b11111111111111111110110100101011;
assign LUT_4[55602] = 32'b00000000000000000101000011010111;
assign LUT_4[55603] = 32'b11111111111111111110001111001111;
assign LUT_4[55604] = 32'b00000000000000000010101001001111;
assign LUT_4[55605] = 32'b11111111111111111011110101000111;
assign LUT_4[55606] = 32'b00000000000000000010000011110011;
assign LUT_4[55607] = 32'b11111111111111111011001111101011;
assign LUT_4[55608] = 32'b11111111111111111110110101001000;
assign LUT_4[55609] = 32'b11111111111111111000000001000000;
assign LUT_4[55610] = 32'b11111111111111111110001111101100;
assign LUT_4[55611] = 32'b11111111111111110111011011100100;
assign LUT_4[55612] = 32'b11111111111111111011110101100100;
assign LUT_4[55613] = 32'b11111111111111110101000001011100;
assign LUT_4[55614] = 32'b11111111111111111011010000001000;
assign LUT_4[55615] = 32'b11111111111111110100011100000000;
assign LUT_4[55616] = 32'b00000000000000001010110011010010;
assign LUT_4[55617] = 32'b00000000000000000011111111001010;
assign LUT_4[55618] = 32'b00000000000000001010001101110110;
assign LUT_4[55619] = 32'b00000000000000000011011001101110;
assign LUT_4[55620] = 32'b00000000000000000111110011101110;
assign LUT_4[55621] = 32'b00000000000000000000111111100110;
assign LUT_4[55622] = 32'b00000000000000000111001110010010;
assign LUT_4[55623] = 32'b00000000000000000000011010001010;
assign LUT_4[55624] = 32'b00000000000000000011111111100111;
assign LUT_4[55625] = 32'b11111111111111111101001011011111;
assign LUT_4[55626] = 32'b00000000000000000011011010001011;
assign LUT_4[55627] = 32'b11111111111111111100100110000011;
assign LUT_4[55628] = 32'b00000000000000000001000000000011;
assign LUT_4[55629] = 32'b11111111111111111010001011111011;
assign LUT_4[55630] = 32'b00000000000000000000011010100111;
assign LUT_4[55631] = 32'b11111111111111111001100110011111;
assign LUT_4[55632] = 32'b00000000000000001000100101000000;
assign LUT_4[55633] = 32'b00000000000000000001110000111000;
assign LUT_4[55634] = 32'b00000000000000000111111111100100;
assign LUT_4[55635] = 32'b00000000000000000001001011011100;
assign LUT_4[55636] = 32'b00000000000000000101100101011100;
assign LUT_4[55637] = 32'b11111111111111111110110001010100;
assign LUT_4[55638] = 32'b00000000000000000101000000000000;
assign LUT_4[55639] = 32'b11111111111111111110001011111000;
assign LUT_4[55640] = 32'b00000000000000000001110001010101;
assign LUT_4[55641] = 32'b11111111111111111010111101001101;
assign LUT_4[55642] = 32'b00000000000000000001001011111001;
assign LUT_4[55643] = 32'b11111111111111111010010111110001;
assign LUT_4[55644] = 32'b11111111111111111110110001110001;
assign LUT_4[55645] = 32'b11111111111111110111111101101001;
assign LUT_4[55646] = 32'b11111111111111111110001100010101;
assign LUT_4[55647] = 32'b11111111111111110111011000001101;
assign LUT_4[55648] = 32'b00000000000000001001001110011001;
assign LUT_4[55649] = 32'b00000000000000000010011010010001;
assign LUT_4[55650] = 32'b00000000000000001000101000111101;
assign LUT_4[55651] = 32'b00000000000000000001110100110101;
assign LUT_4[55652] = 32'b00000000000000000110001110110101;
assign LUT_4[55653] = 32'b11111111111111111111011010101101;
assign LUT_4[55654] = 32'b00000000000000000101101001011001;
assign LUT_4[55655] = 32'b11111111111111111110110101010001;
assign LUT_4[55656] = 32'b00000000000000000010011010101110;
assign LUT_4[55657] = 32'b11111111111111111011100110100110;
assign LUT_4[55658] = 32'b00000000000000000001110101010010;
assign LUT_4[55659] = 32'b11111111111111111011000001001010;
assign LUT_4[55660] = 32'b11111111111111111111011011001010;
assign LUT_4[55661] = 32'b11111111111111111000100111000010;
assign LUT_4[55662] = 32'b11111111111111111110110101101110;
assign LUT_4[55663] = 32'b11111111111111111000000001100110;
assign LUT_4[55664] = 32'b00000000000000000111000000000111;
assign LUT_4[55665] = 32'b00000000000000000000001011111111;
assign LUT_4[55666] = 32'b00000000000000000110011010101011;
assign LUT_4[55667] = 32'b11111111111111111111100110100011;
assign LUT_4[55668] = 32'b00000000000000000100000000100011;
assign LUT_4[55669] = 32'b11111111111111111101001100011011;
assign LUT_4[55670] = 32'b00000000000000000011011011000111;
assign LUT_4[55671] = 32'b11111111111111111100100110111111;
assign LUT_4[55672] = 32'b00000000000000000000001100011100;
assign LUT_4[55673] = 32'b11111111111111111001011000010100;
assign LUT_4[55674] = 32'b11111111111111111111100111000000;
assign LUT_4[55675] = 32'b11111111111111111000110010111000;
assign LUT_4[55676] = 32'b11111111111111111101001100111000;
assign LUT_4[55677] = 32'b11111111111111110110011000110000;
assign LUT_4[55678] = 32'b11111111111111111100100111011100;
assign LUT_4[55679] = 32'b11111111111111110101110011010100;
assign LUT_4[55680] = 32'b00000000000000001100000010000110;
assign LUT_4[55681] = 32'b00000000000000000101001101111110;
assign LUT_4[55682] = 32'b00000000000000001011011100101010;
assign LUT_4[55683] = 32'b00000000000000000100101000100010;
assign LUT_4[55684] = 32'b00000000000000001001000010100010;
assign LUT_4[55685] = 32'b00000000000000000010001110011010;
assign LUT_4[55686] = 32'b00000000000000001000011101000110;
assign LUT_4[55687] = 32'b00000000000000000001101000111110;
assign LUT_4[55688] = 32'b00000000000000000101001110011011;
assign LUT_4[55689] = 32'b11111111111111111110011010010011;
assign LUT_4[55690] = 32'b00000000000000000100101000111111;
assign LUT_4[55691] = 32'b11111111111111111101110100110111;
assign LUT_4[55692] = 32'b00000000000000000010001110110111;
assign LUT_4[55693] = 32'b11111111111111111011011010101111;
assign LUT_4[55694] = 32'b00000000000000000001101001011011;
assign LUT_4[55695] = 32'b11111111111111111010110101010011;
assign LUT_4[55696] = 32'b00000000000000001001110011110100;
assign LUT_4[55697] = 32'b00000000000000000010111111101100;
assign LUT_4[55698] = 32'b00000000000000001001001110011000;
assign LUT_4[55699] = 32'b00000000000000000010011010010000;
assign LUT_4[55700] = 32'b00000000000000000110110100010000;
assign LUT_4[55701] = 32'b00000000000000000000000000001000;
assign LUT_4[55702] = 32'b00000000000000000110001110110100;
assign LUT_4[55703] = 32'b11111111111111111111011010101100;
assign LUT_4[55704] = 32'b00000000000000000011000000001001;
assign LUT_4[55705] = 32'b11111111111111111100001100000001;
assign LUT_4[55706] = 32'b00000000000000000010011010101101;
assign LUT_4[55707] = 32'b11111111111111111011100110100101;
assign LUT_4[55708] = 32'b00000000000000000000000000100101;
assign LUT_4[55709] = 32'b11111111111111111001001100011101;
assign LUT_4[55710] = 32'b11111111111111111111011011001001;
assign LUT_4[55711] = 32'b11111111111111111000100111000001;
assign LUT_4[55712] = 32'b00000000000000001010011101001101;
assign LUT_4[55713] = 32'b00000000000000000011101001000101;
assign LUT_4[55714] = 32'b00000000000000001001110111110001;
assign LUT_4[55715] = 32'b00000000000000000011000011101001;
assign LUT_4[55716] = 32'b00000000000000000111011101101001;
assign LUT_4[55717] = 32'b00000000000000000000101001100001;
assign LUT_4[55718] = 32'b00000000000000000110111000001101;
assign LUT_4[55719] = 32'b00000000000000000000000100000101;
assign LUT_4[55720] = 32'b00000000000000000011101001100010;
assign LUT_4[55721] = 32'b11111111111111111100110101011010;
assign LUT_4[55722] = 32'b00000000000000000011000100000110;
assign LUT_4[55723] = 32'b11111111111111111100001111111110;
assign LUT_4[55724] = 32'b00000000000000000000101001111110;
assign LUT_4[55725] = 32'b11111111111111111001110101110110;
assign LUT_4[55726] = 32'b00000000000000000000000100100010;
assign LUT_4[55727] = 32'b11111111111111111001010000011010;
assign LUT_4[55728] = 32'b00000000000000001000001110111011;
assign LUT_4[55729] = 32'b00000000000000000001011010110011;
assign LUT_4[55730] = 32'b00000000000000000111101001011111;
assign LUT_4[55731] = 32'b00000000000000000000110101010111;
assign LUT_4[55732] = 32'b00000000000000000101001111010111;
assign LUT_4[55733] = 32'b11111111111111111110011011001111;
assign LUT_4[55734] = 32'b00000000000000000100101001111011;
assign LUT_4[55735] = 32'b11111111111111111101110101110011;
assign LUT_4[55736] = 32'b00000000000000000001011011010000;
assign LUT_4[55737] = 32'b11111111111111111010100111001000;
assign LUT_4[55738] = 32'b00000000000000000000110101110100;
assign LUT_4[55739] = 32'b11111111111111111010000001101100;
assign LUT_4[55740] = 32'b11111111111111111110011011101100;
assign LUT_4[55741] = 32'b11111111111111110111100111100100;
assign LUT_4[55742] = 32'b11111111111111111101110110010000;
assign LUT_4[55743] = 32'b11111111111111110111000010001000;
assign LUT_4[55744] = 32'b00000000000000001101011001011010;
assign LUT_4[55745] = 32'b00000000000000000110100101010010;
assign LUT_4[55746] = 32'b00000000000000001100110011111110;
assign LUT_4[55747] = 32'b00000000000000000101111111110110;
assign LUT_4[55748] = 32'b00000000000000001010011001110110;
assign LUT_4[55749] = 32'b00000000000000000011100101101110;
assign LUT_4[55750] = 32'b00000000000000001001110100011010;
assign LUT_4[55751] = 32'b00000000000000000011000000010010;
assign LUT_4[55752] = 32'b00000000000000000110100101101111;
assign LUT_4[55753] = 32'b11111111111111111111110001100111;
assign LUT_4[55754] = 32'b00000000000000000110000000010011;
assign LUT_4[55755] = 32'b11111111111111111111001100001011;
assign LUT_4[55756] = 32'b00000000000000000011100110001011;
assign LUT_4[55757] = 32'b11111111111111111100110010000011;
assign LUT_4[55758] = 32'b00000000000000000011000000101111;
assign LUT_4[55759] = 32'b11111111111111111100001100100111;
assign LUT_4[55760] = 32'b00000000000000001011001011001000;
assign LUT_4[55761] = 32'b00000000000000000100010111000000;
assign LUT_4[55762] = 32'b00000000000000001010100101101100;
assign LUT_4[55763] = 32'b00000000000000000011110001100100;
assign LUT_4[55764] = 32'b00000000000000001000001011100100;
assign LUT_4[55765] = 32'b00000000000000000001010111011100;
assign LUT_4[55766] = 32'b00000000000000000111100110001000;
assign LUT_4[55767] = 32'b00000000000000000000110010000000;
assign LUT_4[55768] = 32'b00000000000000000100010111011101;
assign LUT_4[55769] = 32'b11111111111111111101100011010101;
assign LUT_4[55770] = 32'b00000000000000000011110010000001;
assign LUT_4[55771] = 32'b11111111111111111100111101111001;
assign LUT_4[55772] = 32'b00000000000000000001010111111001;
assign LUT_4[55773] = 32'b11111111111111111010100011110001;
assign LUT_4[55774] = 32'b00000000000000000000110010011101;
assign LUT_4[55775] = 32'b11111111111111111001111110010101;
assign LUT_4[55776] = 32'b00000000000000001011110100100001;
assign LUT_4[55777] = 32'b00000000000000000101000000011001;
assign LUT_4[55778] = 32'b00000000000000001011001111000101;
assign LUT_4[55779] = 32'b00000000000000000100011010111101;
assign LUT_4[55780] = 32'b00000000000000001000110100111101;
assign LUT_4[55781] = 32'b00000000000000000010000000110101;
assign LUT_4[55782] = 32'b00000000000000001000001111100001;
assign LUT_4[55783] = 32'b00000000000000000001011011011001;
assign LUT_4[55784] = 32'b00000000000000000101000000110110;
assign LUT_4[55785] = 32'b11111111111111111110001100101110;
assign LUT_4[55786] = 32'b00000000000000000100011011011010;
assign LUT_4[55787] = 32'b11111111111111111101100111010010;
assign LUT_4[55788] = 32'b00000000000000000010000001010010;
assign LUT_4[55789] = 32'b11111111111111111011001101001010;
assign LUT_4[55790] = 32'b00000000000000000001011011110110;
assign LUT_4[55791] = 32'b11111111111111111010100111101110;
assign LUT_4[55792] = 32'b00000000000000001001100110001111;
assign LUT_4[55793] = 32'b00000000000000000010110010000111;
assign LUT_4[55794] = 32'b00000000000000001001000000110011;
assign LUT_4[55795] = 32'b00000000000000000010001100101011;
assign LUT_4[55796] = 32'b00000000000000000110100110101011;
assign LUT_4[55797] = 32'b11111111111111111111110010100011;
assign LUT_4[55798] = 32'b00000000000000000110000001001111;
assign LUT_4[55799] = 32'b11111111111111111111001101000111;
assign LUT_4[55800] = 32'b00000000000000000010110010100100;
assign LUT_4[55801] = 32'b11111111111111111011111110011100;
assign LUT_4[55802] = 32'b00000000000000000010001101001000;
assign LUT_4[55803] = 32'b11111111111111111011011001000000;
assign LUT_4[55804] = 32'b11111111111111111111110011000000;
assign LUT_4[55805] = 32'b11111111111111111000111110111000;
assign LUT_4[55806] = 32'b11111111111111111111001101100100;
assign LUT_4[55807] = 32'b11111111111111111000011001011100;
assign LUT_4[55808] = 32'b00000000000000000011100100100011;
assign LUT_4[55809] = 32'b11111111111111111100110000011011;
assign LUT_4[55810] = 32'b00000000000000000010111111000111;
assign LUT_4[55811] = 32'b11111111111111111100001010111111;
assign LUT_4[55812] = 32'b00000000000000000000100100111111;
assign LUT_4[55813] = 32'b11111111111111111001110000110111;
assign LUT_4[55814] = 32'b11111111111111111111111111100011;
assign LUT_4[55815] = 32'b11111111111111111001001011011011;
assign LUT_4[55816] = 32'b11111111111111111100110000111000;
assign LUT_4[55817] = 32'b11111111111111110101111100110000;
assign LUT_4[55818] = 32'b11111111111111111100001011011100;
assign LUT_4[55819] = 32'b11111111111111110101010111010100;
assign LUT_4[55820] = 32'b11111111111111111001110001010100;
assign LUT_4[55821] = 32'b11111111111111110010111101001100;
assign LUT_4[55822] = 32'b11111111111111111001001011111000;
assign LUT_4[55823] = 32'b11111111111111110010010111110000;
assign LUT_4[55824] = 32'b00000000000000000001010110010001;
assign LUT_4[55825] = 32'b11111111111111111010100010001001;
assign LUT_4[55826] = 32'b00000000000000000000110000110101;
assign LUT_4[55827] = 32'b11111111111111111001111100101101;
assign LUT_4[55828] = 32'b11111111111111111110010110101101;
assign LUT_4[55829] = 32'b11111111111111110111100010100101;
assign LUT_4[55830] = 32'b11111111111111111101110001010001;
assign LUT_4[55831] = 32'b11111111111111110110111101001001;
assign LUT_4[55832] = 32'b11111111111111111010100010100110;
assign LUT_4[55833] = 32'b11111111111111110011101110011110;
assign LUT_4[55834] = 32'b11111111111111111001111101001010;
assign LUT_4[55835] = 32'b11111111111111110011001001000010;
assign LUT_4[55836] = 32'b11111111111111110111100011000010;
assign LUT_4[55837] = 32'b11111111111111110000101110111010;
assign LUT_4[55838] = 32'b11111111111111110110111101100110;
assign LUT_4[55839] = 32'b11111111111111110000001001011110;
assign LUT_4[55840] = 32'b00000000000000000001111111101010;
assign LUT_4[55841] = 32'b11111111111111111011001011100010;
assign LUT_4[55842] = 32'b00000000000000000001011010001110;
assign LUT_4[55843] = 32'b11111111111111111010100110000110;
assign LUT_4[55844] = 32'b11111111111111111111000000000110;
assign LUT_4[55845] = 32'b11111111111111111000001011111110;
assign LUT_4[55846] = 32'b11111111111111111110011010101010;
assign LUT_4[55847] = 32'b11111111111111110111100110100010;
assign LUT_4[55848] = 32'b11111111111111111011001011111111;
assign LUT_4[55849] = 32'b11111111111111110100010111110111;
assign LUT_4[55850] = 32'b11111111111111111010100110100011;
assign LUT_4[55851] = 32'b11111111111111110011110010011011;
assign LUT_4[55852] = 32'b11111111111111111000001100011011;
assign LUT_4[55853] = 32'b11111111111111110001011000010011;
assign LUT_4[55854] = 32'b11111111111111110111100110111111;
assign LUT_4[55855] = 32'b11111111111111110000110010110111;
assign LUT_4[55856] = 32'b11111111111111111111110001011000;
assign LUT_4[55857] = 32'b11111111111111111000111101010000;
assign LUT_4[55858] = 32'b11111111111111111111001011111100;
assign LUT_4[55859] = 32'b11111111111111111000010111110100;
assign LUT_4[55860] = 32'b11111111111111111100110001110100;
assign LUT_4[55861] = 32'b11111111111111110101111101101100;
assign LUT_4[55862] = 32'b11111111111111111100001100011000;
assign LUT_4[55863] = 32'b11111111111111110101011000010000;
assign LUT_4[55864] = 32'b11111111111111111000111101101101;
assign LUT_4[55865] = 32'b11111111111111110010001001100101;
assign LUT_4[55866] = 32'b11111111111111111000011000010001;
assign LUT_4[55867] = 32'b11111111111111110001100100001001;
assign LUT_4[55868] = 32'b11111111111111110101111110001001;
assign LUT_4[55869] = 32'b11111111111111101111001010000001;
assign LUT_4[55870] = 32'b11111111111111110101011000101101;
assign LUT_4[55871] = 32'b11111111111111101110100100100101;
assign LUT_4[55872] = 32'b00000000000000000100111011110111;
assign LUT_4[55873] = 32'b11111111111111111110000111101111;
assign LUT_4[55874] = 32'b00000000000000000100010110011011;
assign LUT_4[55875] = 32'b11111111111111111101100010010011;
assign LUT_4[55876] = 32'b00000000000000000001111100010011;
assign LUT_4[55877] = 32'b11111111111111111011001000001011;
assign LUT_4[55878] = 32'b00000000000000000001010110110111;
assign LUT_4[55879] = 32'b11111111111111111010100010101111;
assign LUT_4[55880] = 32'b11111111111111111110001000001100;
assign LUT_4[55881] = 32'b11111111111111110111010100000100;
assign LUT_4[55882] = 32'b11111111111111111101100010110000;
assign LUT_4[55883] = 32'b11111111111111110110101110101000;
assign LUT_4[55884] = 32'b11111111111111111011001000101000;
assign LUT_4[55885] = 32'b11111111111111110100010100100000;
assign LUT_4[55886] = 32'b11111111111111111010100011001100;
assign LUT_4[55887] = 32'b11111111111111110011101111000100;
assign LUT_4[55888] = 32'b00000000000000000010101101100101;
assign LUT_4[55889] = 32'b11111111111111111011111001011101;
assign LUT_4[55890] = 32'b00000000000000000010001000001001;
assign LUT_4[55891] = 32'b11111111111111111011010100000001;
assign LUT_4[55892] = 32'b11111111111111111111101110000001;
assign LUT_4[55893] = 32'b11111111111111111000111001111001;
assign LUT_4[55894] = 32'b11111111111111111111001000100101;
assign LUT_4[55895] = 32'b11111111111111111000010100011101;
assign LUT_4[55896] = 32'b11111111111111111011111001111010;
assign LUT_4[55897] = 32'b11111111111111110101000101110010;
assign LUT_4[55898] = 32'b11111111111111111011010100011110;
assign LUT_4[55899] = 32'b11111111111111110100100000010110;
assign LUT_4[55900] = 32'b11111111111111111000111010010110;
assign LUT_4[55901] = 32'b11111111111111110010000110001110;
assign LUT_4[55902] = 32'b11111111111111111000010100111010;
assign LUT_4[55903] = 32'b11111111111111110001100000110010;
assign LUT_4[55904] = 32'b00000000000000000011010110111110;
assign LUT_4[55905] = 32'b11111111111111111100100010110110;
assign LUT_4[55906] = 32'b00000000000000000010110001100010;
assign LUT_4[55907] = 32'b11111111111111111011111101011010;
assign LUT_4[55908] = 32'b00000000000000000000010111011010;
assign LUT_4[55909] = 32'b11111111111111111001100011010010;
assign LUT_4[55910] = 32'b11111111111111111111110001111110;
assign LUT_4[55911] = 32'b11111111111111111000111101110110;
assign LUT_4[55912] = 32'b11111111111111111100100011010011;
assign LUT_4[55913] = 32'b11111111111111110101101111001011;
assign LUT_4[55914] = 32'b11111111111111111011111101110111;
assign LUT_4[55915] = 32'b11111111111111110101001001101111;
assign LUT_4[55916] = 32'b11111111111111111001100011101111;
assign LUT_4[55917] = 32'b11111111111111110010101111100111;
assign LUT_4[55918] = 32'b11111111111111111000111110010011;
assign LUT_4[55919] = 32'b11111111111111110010001010001011;
assign LUT_4[55920] = 32'b00000000000000000001001000101100;
assign LUT_4[55921] = 32'b11111111111111111010010100100100;
assign LUT_4[55922] = 32'b00000000000000000000100011010000;
assign LUT_4[55923] = 32'b11111111111111111001101111001000;
assign LUT_4[55924] = 32'b11111111111111111110001001001000;
assign LUT_4[55925] = 32'b11111111111111110111010101000000;
assign LUT_4[55926] = 32'b11111111111111111101100011101100;
assign LUT_4[55927] = 32'b11111111111111110110101111100100;
assign LUT_4[55928] = 32'b11111111111111111010010101000001;
assign LUT_4[55929] = 32'b11111111111111110011100000111001;
assign LUT_4[55930] = 32'b11111111111111111001101111100101;
assign LUT_4[55931] = 32'b11111111111111110010111011011101;
assign LUT_4[55932] = 32'b11111111111111110111010101011101;
assign LUT_4[55933] = 32'b11111111111111110000100001010101;
assign LUT_4[55934] = 32'b11111111111111110110110000000001;
assign LUT_4[55935] = 32'b11111111111111101111111011111001;
assign LUT_4[55936] = 32'b00000000000000000110001010101011;
assign LUT_4[55937] = 32'b11111111111111111111010110100011;
assign LUT_4[55938] = 32'b00000000000000000101100101001111;
assign LUT_4[55939] = 32'b11111111111111111110110001000111;
assign LUT_4[55940] = 32'b00000000000000000011001011000111;
assign LUT_4[55941] = 32'b11111111111111111100010110111111;
assign LUT_4[55942] = 32'b00000000000000000010100101101011;
assign LUT_4[55943] = 32'b11111111111111111011110001100011;
assign LUT_4[55944] = 32'b11111111111111111111010111000000;
assign LUT_4[55945] = 32'b11111111111111111000100010111000;
assign LUT_4[55946] = 32'b11111111111111111110110001100100;
assign LUT_4[55947] = 32'b11111111111111110111111101011100;
assign LUT_4[55948] = 32'b11111111111111111100010111011100;
assign LUT_4[55949] = 32'b11111111111111110101100011010100;
assign LUT_4[55950] = 32'b11111111111111111011110010000000;
assign LUT_4[55951] = 32'b11111111111111110100111101111000;
assign LUT_4[55952] = 32'b00000000000000000011111100011001;
assign LUT_4[55953] = 32'b11111111111111111101001000010001;
assign LUT_4[55954] = 32'b00000000000000000011010110111101;
assign LUT_4[55955] = 32'b11111111111111111100100010110101;
assign LUT_4[55956] = 32'b00000000000000000000111100110101;
assign LUT_4[55957] = 32'b11111111111111111010001000101101;
assign LUT_4[55958] = 32'b00000000000000000000010111011001;
assign LUT_4[55959] = 32'b11111111111111111001100011010001;
assign LUT_4[55960] = 32'b11111111111111111101001000101110;
assign LUT_4[55961] = 32'b11111111111111110110010100100110;
assign LUT_4[55962] = 32'b11111111111111111100100011010010;
assign LUT_4[55963] = 32'b11111111111111110101101111001010;
assign LUT_4[55964] = 32'b11111111111111111010001001001010;
assign LUT_4[55965] = 32'b11111111111111110011010101000010;
assign LUT_4[55966] = 32'b11111111111111111001100011101110;
assign LUT_4[55967] = 32'b11111111111111110010101111100110;
assign LUT_4[55968] = 32'b00000000000000000100100101110010;
assign LUT_4[55969] = 32'b11111111111111111101110001101010;
assign LUT_4[55970] = 32'b00000000000000000100000000010110;
assign LUT_4[55971] = 32'b11111111111111111101001100001110;
assign LUT_4[55972] = 32'b00000000000000000001100110001110;
assign LUT_4[55973] = 32'b11111111111111111010110010000110;
assign LUT_4[55974] = 32'b00000000000000000001000000110010;
assign LUT_4[55975] = 32'b11111111111111111010001100101010;
assign LUT_4[55976] = 32'b11111111111111111101110010000111;
assign LUT_4[55977] = 32'b11111111111111110110111101111111;
assign LUT_4[55978] = 32'b11111111111111111101001100101011;
assign LUT_4[55979] = 32'b11111111111111110110011000100011;
assign LUT_4[55980] = 32'b11111111111111111010110010100011;
assign LUT_4[55981] = 32'b11111111111111110011111110011011;
assign LUT_4[55982] = 32'b11111111111111111010001101000111;
assign LUT_4[55983] = 32'b11111111111111110011011000111111;
assign LUT_4[55984] = 32'b00000000000000000010010111100000;
assign LUT_4[55985] = 32'b11111111111111111011100011011000;
assign LUT_4[55986] = 32'b00000000000000000001110010000100;
assign LUT_4[55987] = 32'b11111111111111111010111101111100;
assign LUT_4[55988] = 32'b11111111111111111111010111111100;
assign LUT_4[55989] = 32'b11111111111111111000100011110100;
assign LUT_4[55990] = 32'b11111111111111111110110010100000;
assign LUT_4[55991] = 32'b11111111111111110111111110011000;
assign LUT_4[55992] = 32'b11111111111111111011100011110101;
assign LUT_4[55993] = 32'b11111111111111110100101111101101;
assign LUT_4[55994] = 32'b11111111111111111010111110011001;
assign LUT_4[55995] = 32'b11111111111111110100001010010001;
assign LUT_4[55996] = 32'b11111111111111111000100100010001;
assign LUT_4[55997] = 32'b11111111111111110001110000001001;
assign LUT_4[55998] = 32'b11111111111111110111111110110101;
assign LUT_4[55999] = 32'b11111111111111110001001010101101;
assign LUT_4[56000] = 32'b00000000000000000111100001111111;
assign LUT_4[56001] = 32'b00000000000000000000101101110111;
assign LUT_4[56002] = 32'b00000000000000000110111100100011;
assign LUT_4[56003] = 32'b00000000000000000000001000011011;
assign LUT_4[56004] = 32'b00000000000000000100100010011011;
assign LUT_4[56005] = 32'b11111111111111111101101110010011;
assign LUT_4[56006] = 32'b00000000000000000011111100111111;
assign LUT_4[56007] = 32'b11111111111111111101001000110111;
assign LUT_4[56008] = 32'b00000000000000000000101110010100;
assign LUT_4[56009] = 32'b11111111111111111001111010001100;
assign LUT_4[56010] = 32'b00000000000000000000001000111000;
assign LUT_4[56011] = 32'b11111111111111111001010100110000;
assign LUT_4[56012] = 32'b11111111111111111101101110110000;
assign LUT_4[56013] = 32'b11111111111111110110111010101000;
assign LUT_4[56014] = 32'b11111111111111111101001001010100;
assign LUT_4[56015] = 32'b11111111111111110110010101001100;
assign LUT_4[56016] = 32'b00000000000000000101010011101101;
assign LUT_4[56017] = 32'b11111111111111111110011111100101;
assign LUT_4[56018] = 32'b00000000000000000100101110010001;
assign LUT_4[56019] = 32'b11111111111111111101111010001001;
assign LUT_4[56020] = 32'b00000000000000000010010100001001;
assign LUT_4[56021] = 32'b11111111111111111011100000000001;
assign LUT_4[56022] = 32'b00000000000000000001101110101101;
assign LUT_4[56023] = 32'b11111111111111111010111010100101;
assign LUT_4[56024] = 32'b11111111111111111110100000000010;
assign LUT_4[56025] = 32'b11111111111111110111101011111010;
assign LUT_4[56026] = 32'b11111111111111111101111010100110;
assign LUT_4[56027] = 32'b11111111111111110111000110011110;
assign LUT_4[56028] = 32'b11111111111111111011100000011110;
assign LUT_4[56029] = 32'b11111111111111110100101100010110;
assign LUT_4[56030] = 32'b11111111111111111010111011000010;
assign LUT_4[56031] = 32'b11111111111111110100000110111010;
assign LUT_4[56032] = 32'b00000000000000000101111101000110;
assign LUT_4[56033] = 32'b11111111111111111111001000111110;
assign LUT_4[56034] = 32'b00000000000000000101010111101010;
assign LUT_4[56035] = 32'b11111111111111111110100011100010;
assign LUT_4[56036] = 32'b00000000000000000010111101100010;
assign LUT_4[56037] = 32'b11111111111111111100001001011010;
assign LUT_4[56038] = 32'b00000000000000000010011000000110;
assign LUT_4[56039] = 32'b11111111111111111011100011111110;
assign LUT_4[56040] = 32'b11111111111111111111001001011011;
assign LUT_4[56041] = 32'b11111111111111111000010101010011;
assign LUT_4[56042] = 32'b11111111111111111110100011111111;
assign LUT_4[56043] = 32'b11111111111111110111101111110111;
assign LUT_4[56044] = 32'b11111111111111111100001001110111;
assign LUT_4[56045] = 32'b11111111111111110101010101101111;
assign LUT_4[56046] = 32'b11111111111111111011100100011011;
assign LUT_4[56047] = 32'b11111111111111110100110000010011;
assign LUT_4[56048] = 32'b00000000000000000011101110110100;
assign LUT_4[56049] = 32'b11111111111111111100111010101100;
assign LUT_4[56050] = 32'b00000000000000000011001001011000;
assign LUT_4[56051] = 32'b11111111111111111100010101010000;
assign LUT_4[56052] = 32'b00000000000000000000101111010000;
assign LUT_4[56053] = 32'b11111111111111111001111011001000;
assign LUT_4[56054] = 32'b00000000000000000000001001110100;
assign LUT_4[56055] = 32'b11111111111111111001010101101100;
assign LUT_4[56056] = 32'b11111111111111111100111011001001;
assign LUT_4[56057] = 32'b11111111111111110110000111000001;
assign LUT_4[56058] = 32'b11111111111111111100010101101101;
assign LUT_4[56059] = 32'b11111111111111110101100001100101;
assign LUT_4[56060] = 32'b11111111111111111001111011100101;
assign LUT_4[56061] = 32'b11111111111111110011000111011101;
assign LUT_4[56062] = 32'b11111111111111111001010110001001;
assign LUT_4[56063] = 32'b11111111111111110010100010000001;
assign LUT_4[56064] = 32'b00000000000000001000100000000110;
assign LUT_4[56065] = 32'b00000000000000000001101011111110;
assign LUT_4[56066] = 32'b00000000000000000111111010101010;
assign LUT_4[56067] = 32'b00000000000000000001000110100010;
assign LUT_4[56068] = 32'b00000000000000000101100000100010;
assign LUT_4[56069] = 32'b11111111111111111110101100011010;
assign LUT_4[56070] = 32'b00000000000000000100111011000110;
assign LUT_4[56071] = 32'b11111111111111111110000110111110;
assign LUT_4[56072] = 32'b00000000000000000001101100011011;
assign LUT_4[56073] = 32'b11111111111111111010111000010011;
assign LUT_4[56074] = 32'b00000000000000000001000110111111;
assign LUT_4[56075] = 32'b11111111111111111010010010110111;
assign LUT_4[56076] = 32'b11111111111111111110101100110111;
assign LUT_4[56077] = 32'b11111111111111110111111000101111;
assign LUT_4[56078] = 32'b11111111111111111110000111011011;
assign LUT_4[56079] = 32'b11111111111111110111010011010011;
assign LUT_4[56080] = 32'b00000000000000000110010001110100;
assign LUT_4[56081] = 32'b11111111111111111111011101101100;
assign LUT_4[56082] = 32'b00000000000000000101101100011000;
assign LUT_4[56083] = 32'b11111111111111111110111000010000;
assign LUT_4[56084] = 32'b00000000000000000011010010010000;
assign LUT_4[56085] = 32'b11111111111111111100011110001000;
assign LUT_4[56086] = 32'b00000000000000000010101100110100;
assign LUT_4[56087] = 32'b11111111111111111011111000101100;
assign LUT_4[56088] = 32'b11111111111111111111011110001001;
assign LUT_4[56089] = 32'b11111111111111111000101010000001;
assign LUT_4[56090] = 32'b11111111111111111110111000101101;
assign LUT_4[56091] = 32'b11111111111111111000000100100101;
assign LUT_4[56092] = 32'b11111111111111111100011110100101;
assign LUT_4[56093] = 32'b11111111111111110101101010011101;
assign LUT_4[56094] = 32'b11111111111111111011111001001001;
assign LUT_4[56095] = 32'b11111111111111110101000101000001;
assign LUT_4[56096] = 32'b00000000000000000110111011001101;
assign LUT_4[56097] = 32'b00000000000000000000000111000101;
assign LUT_4[56098] = 32'b00000000000000000110010101110001;
assign LUT_4[56099] = 32'b11111111111111111111100001101001;
assign LUT_4[56100] = 32'b00000000000000000011111011101001;
assign LUT_4[56101] = 32'b11111111111111111101000111100001;
assign LUT_4[56102] = 32'b00000000000000000011010110001101;
assign LUT_4[56103] = 32'b11111111111111111100100010000101;
assign LUT_4[56104] = 32'b00000000000000000000000111100010;
assign LUT_4[56105] = 32'b11111111111111111001010011011010;
assign LUT_4[56106] = 32'b11111111111111111111100010000110;
assign LUT_4[56107] = 32'b11111111111111111000101101111110;
assign LUT_4[56108] = 32'b11111111111111111101000111111110;
assign LUT_4[56109] = 32'b11111111111111110110010011110110;
assign LUT_4[56110] = 32'b11111111111111111100100010100010;
assign LUT_4[56111] = 32'b11111111111111110101101110011010;
assign LUT_4[56112] = 32'b00000000000000000100101100111011;
assign LUT_4[56113] = 32'b11111111111111111101111000110011;
assign LUT_4[56114] = 32'b00000000000000000100000111011111;
assign LUT_4[56115] = 32'b11111111111111111101010011010111;
assign LUT_4[56116] = 32'b00000000000000000001101101010111;
assign LUT_4[56117] = 32'b11111111111111111010111001001111;
assign LUT_4[56118] = 32'b00000000000000000001000111111011;
assign LUT_4[56119] = 32'b11111111111111111010010011110011;
assign LUT_4[56120] = 32'b11111111111111111101111001010000;
assign LUT_4[56121] = 32'b11111111111111110111000101001000;
assign LUT_4[56122] = 32'b11111111111111111101010011110100;
assign LUT_4[56123] = 32'b11111111111111110110011111101100;
assign LUT_4[56124] = 32'b11111111111111111010111001101100;
assign LUT_4[56125] = 32'b11111111111111110100000101100100;
assign LUT_4[56126] = 32'b11111111111111111010010100010000;
assign LUT_4[56127] = 32'b11111111111111110011100000001000;
assign LUT_4[56128] = 32'b00000000000000001001110111011010;
assign LUT_4[56129] = 32'b00000000000000000011000011010010;
assign LUT_4[56130] = 32'b00000000000000001001010001111110;
assign LUT_4[56131] = 32'b00000000000000000010011101110110;
assign LUT_4[56132] = 32'b00000000000000000110110111110110;
assign LUT_4[56133] = 32'b00000000000000000000000011101110;
assign LUT_4[56134] = 32'b00000000000000000110010010011010;
assign LUT_4[56135] = 32'b11111111111111111111011110010010;
assign LUT_4[56136] = 32'b00000000000000000011000011101111;
assign LUT_4[56137] = 32'b11111111111111111100001111100111;
assign LUT_4[56138] = 32'b00000000000000000010011110010011;
assign LUT_4[56139] = 32'b11111111111111111011101010001011;
assign LUT_4[56140] = 32'b00000000000000000000000100001011;
assign LUT_4[56141] = 32'b11111111111111111001010000000011;
assign LUT_4[56142] = 32'b11111111111111111111011110101111;
assign LUT_4[56143] = 32'b11111111111111111000101010100111;
assign LUT_4[56144] = 32'b00000000000000000111101001001000;
assign LUT_4[56145] = 32'b00000000000000000000110101000000;
assign LUT_4[56146] = 32'b00000000000000000111000011101100;
assign LUT_4[56147] = 32'b00000000000000000000001111100100;
assign LUT_4[56148] = 32'b00000000000000000100101001100100;
assign LUT_4[56149] = 32'b11111111111111111101110101011100;
assign LUT_4[56150] = 32'b00000000000000000100000100001000;
assign LUT_4[56151] = 32'b11111111111111111101010000000000;
assign LUT_4[56152] = 32'b00000000000000000000110101011101;
assign LUT_4[56153] = 32'b11111111111111111010000001010101;
assign LUT_4[56154] = 32'b00000000000000000000010000000001;
assign LUT_4[56155] = 32'b11111111111111111001011011111001;
assign LUT_4[56156] = 32'b11111111111111111101110101111001;
assign LUT_4[56157] = 32'b11111111111111110111000001110001;
assign LUT_4[56158] = 32'b11111111111111111101010000011101;
assign LUT_4[56159] = 32'b11111111111111110110011100010101;
assign LUT_4[56160] = 32'b00000000000000001000010010100001;
assign LUT_4[56161] = 32'b00000000000000000001011110011001;
assign LUT_4[56162] = 32'b00000000000000000111101101000101;
assign LUT_4[56163] = 32'b00000000000000000000111000111101;
assign LUT_4[56164] = 32'b00000000000000000101010010111101;
assign LUT_4[56165] = 32'b11111111111111111110011110110101;
assign LUT_4[56166] = 32'b00000000000000000100101101100001;
assign LUT_4[56167] = 32'b11111111111111111101111001011001;
assign LUT_4[56168] = 32'b00000000000000000001011110110110;
assign LUT_4[56169] = 32'b11111111111111111010101010101110;
assign LUT_4[56170] = 32'b00000000000000000000111001011010;
assign LUT_4[56171] = 32'b11111111111111111010000101010010;
assign LUT_4[56172] = 32'b11111111111111111110011111010010;
assign LUT_4[56173] = 32'b11111111111111110111101011001010;
assign LUT_4[56174] = 32'b11111111111111111101111001110110;
assign LUT_4[56175] = 32'b11111111111111110111000101101110;
assign LUT_4[56176] = 32'b00000000000000000110000100001111;
assign LUT_4[56177] = 32'b11111111111111111111010000000111;
assign LUT_4[56178] = 32'b00000000000000000101011110110011;
assign LUT_4[56179] = 32'b11111111111111111110101010101011;
assign LUT_4[56180] = 32'b00000000000000000011000100101011;
assign LUT_4[56181] = 32'b11111111111111111100010000100011;
assign LUT_4[56182] = 32'b00000000000000000010011111001111;
assign LUT_4[56183] = 32'b11111111111111111011101011000111;
assign LUT_4[56184] = 32'b11111111111111111111010000100100;
assign LUT_4[56185] = 32'b11111111111111111000011100011100;
assign LUT_4[56186] = 32'b11111111111111111110101011001000;
assign LUT_4[56187] = 32'b11111111111111110111110111000000;
assign LUT_4[56188] = 32'b11111111111111111100010001000000;
assign LUT_4[56189] = 32'b11111111111111110101011100111000;
assign LUT_4[56190] = 32'b11111111111111111011101011100100;
assign LUT_4[56191] = 32'b11111111111111110100110111011100;
assign LUT_4[56192] = 32'b00000000000000001011000110001110;
assign LUT_4[56193] = 32'b00000000000000000100010010000110;
assign LUT_4[56194] = 32'b00000000000000001010100000110010;
assign LUT_4[56195] = 32'b00000000000000000011101100101010;
assign LUT_4[56196] = 32'b00000000000000001000000110101010;
assign LUT_4[56197] = 32'b00000000000000000001010010100010;
assign LUT_4[56198] = 32'b00000000000000000111100001001110;
assign LUT_4[56199] = 32'b00000000000000000000101101000110;
assign LUT_4[56200] = 32'b00000000000000000100010010100011;
assign LUT_4[56201] = 32'b11111111111111111101011110011011;
assign LUT_4[56202] = 32'b00000000000000000011101101000111;
assign LUT_4[56203] = 32'b11111111111111111100111000111111;
assign LUT_4[56204] = 32'b00000000000000000001010010111111;
assign LUT_4[56205] = 32'b11111111111111111010011110110111;
assign LUT_4[56206] = 32'b00000000000000000000101101100011;
assign LUT_4[56207] = 32'b11111111111111111001111001011011;
assign LUT_4[56208] = 32'b00000000000000001000110111111100;
assign LUT_4[56209] = 32'b00000000000000000010000011110100;
assign LUT_4[56210] = 32'b00000000000000001000010010100000;
assign LUT_4[56211] = 32'b00000000000000000001011110011000;
assign LUT_4[56212] = 32'b00000000000000000101111000011000;
assign LUT_4[56213] = 32'b11111111111111111111000100010000;
assign LUT_4[56214] = 32'b00000000000000000101010010111100;
assign LUT_4[56215] = 32'b11111111111111111110011110110100;
assign LUT_4[56216] = 32'b00000000000000000010000100010001;
assign LUT_4[56217] = 32'b11111111111111111011010000001001;
assign LUT_4[56218] = 32'b00000000000000000001011110110101;
assign LUT_4[56219] = 32'b11111111111111111010101010101101;
assign LUT_4[56220] = 32'b11111111111111111111000100101101;
assign LUT_4[56221] = 32'b11111111111111111000010000100101;
assign LUT_4[56222] = 32'b11111111111111111110011111010001;
assign LUT_4[56223] = 32'b11111111111111110111101011001001;
assign LUT_4[56224] = 32'b00000000000000001001100001010101;
assign LUT_4[56225] = 32'b00000000000000000010101101001101;
assign LUT_4[56226] = 32'b00000000000000001000111011111001;
assign LUT_4[56227] = 32'b00000000000000000010000111110001;
assign LUT_4[56228] = 32'b00000000000000000110100001110001;
assign LUT_4[56229] = 32'b11111111111111111111101101101001;
assign LUT_4[56230] = 32'b00000000000000000101111100010101;
assign LUT_4[56231] = 32'b11111111111111111111001000001101;
assign LUT_4[56232] = 32'b00000000000000000010101101101010;
assign LUT_4[56233] = 32'b11111111111111111011111001100010;
assign LUT_4[56234] = 32'b00000000000000000010001000001110;
assign LUT_4[56235] = 32'b11111111111111111011010100000110;
assign LUT_4[56236] = 32'b11111111111111111111101110000110;
assign LUT_4[56237] = 32'b11111111111111111000111001111110;
assign LUT_4[56238] = 32'b11111111111111111111001000101010;
assign LUT_4[56239] = 32'b11111111111111111000010100100010;
assign LUT_4[56240] = 32'b00000000000000000111010011000011;
assign LUT_4[56241] = 32'b00000000000000000000011110111011;
assign LUT_4[56242] = 32'b00000000000000000110101101100111;
assign LUT_4[56243] = 32'b11111111111111111111111001011111;
assign LUT_4[56244] = 32'b00000000000000000100010011011111;
assign LUT_4[56245] = 32'b11111111111111111101011111010111;
assign LUT_4[56246] = 32'b00000000000000000011101110000011;
assign LUT_4[56247] = 32'b11111111111111111100111001111011;
assign LUT_4[56248] = 32'b00000000000000000000011111011000;
assign LUT_4[56249] = 32'b11111111111111111001101011010000;
assign LUT_4[56250] = 32'b11111111111111111111111001111100;
assign LUT_4[56251] = 32'b11111111111111111001000101110100;
assign LUT_4[56252] = 32'b11111111111111111101011111110100;
assign LUT_4[56253] = 32'b11111111111111110110101011101100;
assign LUT_4[56254] = 32'b11111111111111111100111010011000;
assign LUT_4[56255] = 32'b11111111111111110110000110010000;
assign LUT_4[56256] = 32'b00000000000000001100011101100010;
assign LUT_4[56257] = 32'b00000000000000000101101001011010;
assign LUT_4[56258] = 32'b00000000000000001011111000000110;
assign LUT_4[56259] = 32'b00000000000000000101000011111110;
assign LUT_4[56260] = 32'b00000000000000001001011101111110;
assign LUT_4[56261] = 32'b00000000000000000010101001110110;
assign LUT_4[56262] = 32'b00000000000000001000111000100010;
assign LUT_4[56263] = 32'b00000000000000000010000100011010;
assign LUT_4[56264] = 32'b00000000000000000101101001110111;
assign LUT_4[56265] = 32'b11111111111111111110110101101111;
assign LUT_4[56266] = 32'b00000000000000000101000100011011;
assign LUT_4[56267] = 32'b11111111111111111110010000010011;
assign LUT_4[56268] = 32'b00000000000000000010101010010011;
assign LUT_4[56269] = 32'b11111111111111111011110110001011;
assign LUT_4[56270] = 32'b00000000000000000010000100110111;
assign LUT_4[56271] = 32'b11111111111111111011010000101111;
assign LUT_4[56272] = 32'b00000000000000001010001111010000;
assign LUT_4[56273] = 32'b00000000000000000011011011001000;
assign LUT_4[56274] = 32'b00000000000000001001101001110100;
assign LUT_4[56275] = 32'b00000000000000000010110101101100;
assign LUT_4[56276] = 32'b00000000000000000111001111101100;
assign LUT_4[56277] = 32'b00000000000000000000011011100100;
assign LUT_4[56278] = 32'b00000000000000000110101010010000;
assign LUT_4[56279] = 32'b11111111111111111111110110001000;
assign LUT_4[56280] = 32'b00000000000000000011011011100101;
assign LUT_4[56281] = 32'b11111111111111111100100111011101;
assign LUT_4[56282] = 32'b00000000000000000010110110001001;
assign LUT_4[56283] = 32'b11111111111111111100000010000001;
assign LUT_4[56284] = 32'b00000000000000000000011100000001;
assign LUT_4[56285] = 32'b11111111111111111001100111111001;
assign LUT_4[56286] = 32'b11111111111111111111110110100101;
assign LUT_4[56287] = 32'b11111111111111111001000010011101;
assign LUT_4[56288] = 32'b00000000000000001010111000101001;
assign LUT_4[56289] = 32'b00000000000000000100000100100001;
assign LUT_4[56290] = 32'b00000000000000001010010011001101;
assign LUT_4[56291] = 32'b00000000000000000011011111000101;
assign LUT_4[56292] = 32'b00000000000000000111111001000101;
assign LUT_4[56293] = 32'b00000000000000000001000100111101;
assign LUT_4[56294] = 32'b00000000000000000111010011101001;
assign LUT_4[56295] = 32'b00000000000000000000011111100001;
assign LUT_4[56296] = 32'b00000000000000000100000100111110;
assign LUT_4[56297] = 32'b11111111111111111101010000110110;
assign LUT_4[56298] = 32'b00000000000000000011011111100010;
assign LUT_4[56299] = 32'b11111111111111111100101011011010;
assign LUT_4[56300] = 32'b00000000000000000001000101011010;
assign LUT_4[56301] = 32'b11111111111111111010010001010010;
assign LUT_4[56302] = 32'b00000000000000000000011111111110;
assign LUT_4[56303] = 32'b11111111111111111001101011110110;
assign LUT_4[56304] = 32'b00000000000000001000101010010111;
assign LUT_4[56305] = 32'b00000000000000000001110110001111;
assign LUT_4[56306] = 32'b00000000000000001000000100111011;
assign LUT_4[56307] = 32'b00000000000000000001010000110011;
assign LUT_4[56308] = 32'b00000000000000000101101010110011;
assign LUT_4[56309] = 32'b11111111111111111110110110101011;
assign LUT_4[56310] = 32'b00000000000000000101000101010111;
assign LUT_4[56311] = 32'b11111111111111111110010001001111;
assign LUT_4[56312] = 32'b00000000000000000001110110101100;
assign LUT_4[56313] = 32'b11111111111111111011000010100100;
assign LUT_4[56314] = 32'b00000000000000000001010001010000;
assign LUT_4[56315] = 32'b11111111111111111010011101001000;
assign LUT_4[56316] = 32'b11111111111111111110110111001000;
assign LUT_4[56317] = 32'b11111111111111111000000011000000;
assign LUT_4[56318] = 32'b11111111111111111110010001101100;
assign LUT_4[56319] = 32'b11111111111111110111011101100100;
assign LUT_4[56320] = 32'b00000000000000000110001010111010;
assign LUT_4[56321] = 32'b11111111111111111111010110110010;
assign LUT_4[56322] = 32'b00000000000000000101100101011110;
assign LUT_4[56323] = 32'b11111111111111111110110001010110;
assign LUT_4[56324] = 32'b00000000000000000011001011010110;
assign LUT_4[56325] = 32'b11111111111111111100010111001110;
assign LUT_4[56326] = 32'b00000000000000000010100101111010;
assign LUT_4[56327] = 32'b11111111111111111011110001110010;
assign LUT_4[56328] = 32'b11111111111111111111010111001111;
assign LUT_4[56329] = 32'b11111111111111111000100011000111;
assign LUT_4[56330] = 32'b11111111111111111110110001110011;
assign LUT_4[56331] = 32'b11111111111111110111111101101011;
assign LUT_4[56332] = 32'b11111111111111111100010111101011;
assign LUT_4[56333] = 32'b11111111111111110101100011100011;
assign LUT_4[56334] = 32'b11111111111111111011110010001111;
assign LUT_4[56335] = 32'b11111111111111110100111110000111;
assign LUT_4[56336] = 32'b00000000000000000011111100101000;
assign LUT_4[56337] = 32'b11111111111111111101001000100000;
assign LUT_4[56338] = 32'b00000000000000000011010111001100;
assign LUT_4[56339] = 32'b11111111111111111100100011000100;
assign LUT_4[56340] = 32'b00000000000000000000111101000100;
assign LUT_4[56341] = 32'b11111111111111111010001000111100;
assign LUT_4[56342] = 32'b00000000000000000000010111101000;
assign LUT_4[56343] = 32'b11111111111111111001100011100000;
assign LUT_4[56344] = 32'b11111111111111111101001000111101;
assign LUT_4[56345] = 32'b11111111111111110110010100110101;
assign LUT_4[56346] = 32'b11111111111111111100100011100001;
assign LUT_4[56347] = 32'b11111111111111110101101111011001;
assign LUT_4[56348] = 32'b11111111111111111010001001011001;
assign LUT_4[56349] = 32'b11111111111111110011010101010001;
assign LUT_4[56350] = 32'b11111111111111111001100011111101;
assign LUT_4[56351] = 32'b11111111111111110010101111110101;
assign LUT_4[56352] = 32'b00000000000000000100100110000001;
assign LUT_4[56353] = 32'b11111111111111111101110001111001;
assign LUT_4[56354] = 32'b00000000000000000100000000100101;
assign LUT_4[56355] = 32'b11111111111111111101001100011101;
assign LUT_4[56356] = 32'b00000000000000000001100110011101;
assign LUT_4[56357] = 32'b11111111111111111010110010010101;
assign LUT_4[56358] = 32'b00000000000000000001000001000001;
assign LUT_4[56359] = 32'b11111111111111111010001100111001;
assign LUT_4[56360] = 32'b11111111111111111101110010010110;
assign LUT_4[56361] = 32'b11111111111111110110111110001110;
assign LUT_4[56362] = 32'b11111111111111111101001100111010;
assign LUT_4[56363] = 32'b11111111111111110110011000110010;
assign LUT_4[56364] = 32'b11111111111111111010110010110010;
assign LUT_4[56365] = 32'b11111111111111110011111110101010;
assign LUT_4[56366] = 32'b11111111111111111010001101010110;
assign LUT_4[56367] = 32'b11111111111111110011011001001110;
assign LUT_4[56368] = 32'b00000000000000000010010111101111;
assign LUT_4[56369] = 32'b11111111111111111011100011100111;
assign LUT_4[56370] = 32'b00000000000000000001110010010011;
assign LUT_4[56371] = 32'b11111111111111111010111110001011;
assign LUT_4[56372] = 32'b11111111111111111111011000001011;
assign LUT_4[56373] = 32'b11111111111111111000100100000011;
assign LUT_4[56374] = 32'b11111111111111111110110010101111;
assign LUT_4[56375] = 32'b11111111111111110111111110100111;
assign LUT_4[56376] = 32'b11111111111111111011100100000100;
assign LUT_4[56377] = 32'b11111111111111110100101111111100;
assign LUT_4[56378] = 32'b11111111111111111010111110101000;
assign LUT_4[56379] = 32'b11111111111111110100001010100000;
assign LUT_4[56380] = 32'b11111111111111111000100100100000;
assign LUT_4[56381] = 32'b11111111111111110001110000011000;
assign LUT_4[56382] = 32'b11111111111111110111111111000100;
assign LUT_4[56383] = 32'b11111111111111110001001010111100;
assign LUT_4[56384] = 32'b00000000000000000111100010001110;
assign LUT_4[56385] = 32'b00000000000000000000101110000110;
assign LUT_4[56386] = 32'b00000000000000000110111100110010;
assign LUT_4[56387] = 32'b00000000000000000000001000101010;
assign LUT_4[56388] = 32'b00000000000000000100100010101010;
assign LUT_4[56389] = 32'b11111111111111111101101110100010;
assign LUT_4[56390] = 32'b00000000000000000011111101001110;
assign LUT_4[56391] = 32'b11111111111111111101001001000110;
assign LUT_4[56392] = 32'b00000000000000000000101110100011;
assign LUT_4[56393] = 32'b11111111111111111001111010011011;
assign LUT_4[56394] = 32'b00000000000000000000001001000111;
assign LUT_4[56395] = 32'b11111111111111111001010100111111;
assign LUT_4[56396] = 32'b11111111111111111101101110111111;
assign LUT_4[56397] = 32'b11111111111111110110111010110111;
assign LUT_4[56398] = 32'b11111111111111111101001001100011;
assign LUT_4[56399] = 32'b11111111111111110110010101011011;
assign LUT_4[56400] = 32'b00000000000000000101010011111100;
assign LUT_4[56401] = 32'b11111111111111111110011111110100;
assign LUT_4[56402] = 32'b00000000000000000100101110100000;
assign LUT_4[56403] = 32'b11111111111111111101111010011000;
assign LUT_4[56404] = 32'b00000000000000000010010100011000;
assign LUT_4[56405] = 32'b11111111111111111011100000010000;
assign LUT_4[56406] = 32'b00000000000000000001101110111100;
assign LUT_4[56407] = 32'b11111111111111111010111010110100;
assign LUT_4[56408] = 32'b11111111111111111110100000010001;
assign LUT_4[56409] = 32'b11111111111111110111101100001001;
assign LUT_4[56410] = 32'b11111111111111111101111010110101;
assign LUT_4[56411] = 32'b11111111111111110111000110101101;
assign LUT_4[56412] = 32'b11111111111111111011100000101101;
assign LUT_4[56413] = 32'b11111111111111110100101100100101;
assign LUT_4[56414] = 32'b11111111111111111010111011010001;
assign LUT_4[56415] = 32'b11111111111111110100000111001001;
assign LUT_4[56416] = 32'b00000000000000000101111101010101;
assign LUT_4[56417] = 32'b11111111111111111111001001001101;
assign LUT_4[56418] = 32'b00000000000000000101010111111001;
assign LUT_4[56419] = 32'b11111111111111111110100011110001;
assign LUT_4[56420] = 32'b00000000000000000010111101110001;
assign LUT_4[56421] = 32'b11111111111111111100001001101001;
assign LUT_4[56422] = 32'b00000000000000000010011000010101;
assign LUT_4[56423] = 32'b11111111111111111011100100001101;
assign LUT_4[56424] = 32'b11111111111111111111001001101010;
assign LUT_4[56425] = 32'b11111111111111111000010101100010;
assign LUT_4[56426] = 32'b11111111111111111110100100001110;
assign LUT_4[56427] = 32'b11111111111111110111110000000110;
assign LUT_4[56428] = 32'b11111111111111111100001010000110;
assign LUT_4[56429] = 32'b11111111111111110101010101111110;
assign LUT_4[56430] = 32'b11111111111111111011100100101010;
assign LUT_4[56431] = 32'b11111111111111110100110000100010;
assign LUT_4[56432] = 32'b00000000000000000011101111000011;
assign LUT_4[56433] = 32'b11111111111111111100111010111011;
assign LUT_4[56434] = 32'b00000000000000000011001001100111;
assign LUT_4[56435] = 32'b11111111111111111100010101011111;
assign LUT_4[56436] = 32'b00000000000000000000101111011111;
assign LUT_4[56437] = 32'b11111111111111111001111011010111;
assign LUT_4[56438] = 32'b00000000000000000000001010000011;
assign LUT_4[56439] = 32'b11111111111111111001010101111011;
assign LUT_4[56440] = 32'b11111111111111111100111011011000;
assign LUT_4[56441] = 32'b11111111111111110110000111010000;
assign LUT_4[56442] = 32'b11111111111111111100010101111100;
assign LUT_4[56443] = 32'b11111111111111110101100001110100;
assign LUT_4[56444] = 32'b11111111111111111001111011110100;
assign LUT_4[56445] = 32'b11111111111111110011000111101100;
assign LUT_4[56446] = 32'b11111111111111111001010110011000;
assign LUT_4[56447] = 32'b11111111111111110010100010010000;
assign LUT_4[56448] = 32'b00000000000000001000110001000010;
assign LUT_4[56449] = 32'b00000000000000000001111100111010;
assign LUT_4[56450] = 32'b00000000000000001000001011100110;
assign LUT_4[56451] = 32'b00000000000000000001010111011110;
assign LUT_4[56452] = 32'b00000000000000000101110001011110;
assign LUT_4[56453] = 32'b11111111111111111110111101010110;
assign LUT_4[56454] = 32'b00000000000000000101001100000010;
assign LUT_4[56455] = 32'b11111111111111111110010111111010;
assign LUT_4[56456] = 32'b00000000000000000001111101010111;
assign LUT_4[56457] = 32'b11111111111111111011001001001111;
assign LUT_4[56458] = 32'b00000000000000000001010111111011;
assign LUT_4[56459] = 32'b11111111111111111010100011110011;
assign LUT_4[56460] = 32'b11111111111111111110111101110011;
assign LUT_4[56461] = 32'b11111111111111111000001001101011;
assign LUT_4[56462] = 32'b11111111111111111110011000010111;
assign LUT_4[56463] = 32'b11111111111111110111100100001111;
assign LUT_4[56464] = 32'b00000000000000000110100010110000;
assign LUT_4[56465] = 32'b11111111111111111111101110101000;
assign LUT_4[56466] = 32'b00000000000000000101111101010100;
assign LUT_4[56467] = 32'b11111111111111111111001001001100;
assign LUT_4[56468] = 32'b00000000000000000011100011001100;
assign LUT_4[56469] = 32'b11111111111111111100101111000100;
assign LUT_4[56470] = 32'b00000000000000000010111101110000;
assign LUT_4[56471] = 32'b11111111111111111100001001101000;
assign LUT_4[56472] = 32'b11111111111111111111101111000101;
assign LUT_4[56473] = 32'b11111111111111111000111010111101;
assign LUT_4[56474] = 32'b11111111111111111111001001101001;
assign LUT_4[56475] = 32'b11111111111111111000010101100001;
assign LUT_4[56476] = 32'b11111111111111111100101111100001;
assign LUT_4[56477] = 32'b11111111111111110101111011011001;
assign LUT_4[56478] = 32'b11111111111111111100001010000101;
assign LUT_4[56479] = 32'b11111111111111110101010101111101;
assign LUT_4[56480] = 32'b00000000000000000111001100001001;
assign LUT_4[56481] = 32'b00000000000000000000011000000001;
assign LUT_4[56482] = 32'b00000000000000000110100110101101;
assign LUT_4[56483] = 32'b11111111111111111111110010100101;
assign LUT_4[56484] = 32'b00000000000000000100001100100101;
assign LUT_4[56485] = 32'b11111111111111111101011000011101;
assign LUT_4[56486] = 32'b00000000000000000011100111001001;
assign LUT_4[56487] = 32'b11111111111111111100110011000001;
assign LUT_4[56488] = 32'b00000000000000000000011000011110;
assign LUT_4[56489] = 32'b11111111111111111001100100010110;
assign LUT_4[56490] = 32'b11111111111111111111110011000010;
assign LUT_4[56491] = 32'b11111111111111111000111110111010;
assign LUT_4[56492] = 32'b11111111111111111101011000111010;
assign LUT_4[56493] = 32'b11111111111111110110100100110010;
assign LUT_4[56494] = 32'b11111111111111111100110011011110;
assign LUT_4[56495] = 32'b11111111111111110101111111010110;
assign LUT_4[56496] = 32'b00000000000000000100111101110111;
assign LUT_4[56497] = 32'b11111111111111111110001001101111;
assign LUT_4[56498] = 32'b00000000000000000100011000011011;
assign LUT_4[56499] = 32'b11111111111111111101100100010011;
assign LUT_4[56500] = 32'b00000000000000000001111110010011;
assign LUT_4[56501] = 32'b11111111111111111011001010001011;
assign LUT_4[56502] = 32'b00000000000000000001011000110111;
assign LUT_4[56503] = 32'b11111111111111111010100100101111;
assign LUT_4[56504] = 32'b11111111111111111110001010001100;
assign LUT_4[56505] = 32'b11111111111111110111010110000100;
assign LUT_4[56506] = 32'b11111111111111111101100100110000;
assign LUT_4[56507] = 32'b11111111111111110110110000101000;
assign LUT_4[56508] = 32'b11111111111111111011001010101000;
assign LUT_4[56509] = 32'b11111111111111110100010110100000;
assign LUT_4[56510] = 32'b11111111111111111010100101001100;
assign LUT_4[56511] = 32'b11111111111111110011110001000100;
assign LUT_4[56512] = 32'b00000000000000001010001000010110;
assign LUT_4[56513] = 32'b00000000000000000011010100001110;
assign LUT_4[56514] = 32'b00000000000000001001100010111010;
assign LUT_4[56515] = 32'b00000000000000000010101110110010;
assign LUT_4[56516] = 32'b00000000000000000111001000110010;
assign LUT_4[56517] = 32'b00000000000000000000010100101010;
assign LUT_4[56518] = 32'b00000000000000000110100011010110;
assign LUT_4[56519] = 32'b11111111111111111111101111001110;
assign LUT_4[56520] = 32'b00000000000000000011010100101011;
assign LUT_4[56521] = 32'b11111111111111111100100000100011;
assign LUT_4[56522] = 32'b00000000000000000010101111001111;
assign LUT_4[56523] = 32'b11111111111111111011111011000111;
assign LUT_4[56524] = 32'b00000000000000000000010101000111;
assign LUT_4[56525] = 32'b11111111111111111001100000111111;
assign LUT_4[56526] = 32'b11111111111111111111101111101011;
assign LUT_4[56527] = 32'b11111111111111111000111011100011;
assign LUT_4[56528] = 32'b00000000000000000111111010000100;
assign LUT_4[56529] = 32'b00000000000000000001000101111100;
assign LUT_4[56530] = 32'b00000000000000000111010100101000;
assign LUT_4[56531] = 32'b00000000000000000000100000100000;
assign LUT_4[56532] = 32'b00000000000000000100111010100000;
assign LUT_4[56533] = 32'b11111111111111111110000110011000;
assign LUT_4[56534] = 32'b00000000000000000100010101000100;
assign LUT_4[56535] = 32'b11111111111111111101100000111100;
assign LUT_4[56536] = 32'b00000000000000000001000110011001;
assign LUT_4[56537] = 32'b11111111111111111010010010010001;
assign LUT_4[56538] = 32'b00000000000000000000100000111101;
assign LUT_4[56539] = 32'b11111111111111111001101100110101;
assign LUT_4[56540] = 32'b11111111111111111110000110110101;
assign LUT_4[56541] = 32'b11111111111111110111010010101101;
assign LUT_4[56542] = 32'b11111111111111111101100001011001;
assign LUT_4[56543] = 32'b11111111111111110110101101010001;
assign LUT_4[56544] = 32'b00000000000000001000100011011101;
assign LUT_4[56545] = 32'b00000000000000000001101111010101;
assign LUT_4[56546] = 32'b00000000000000000111111110000001;
assign LUT_4[56547] = 32'b00000000000000000001001001111001;
assign LUT_4[56548] = 32'b00000000000000000101100011111001;
assign LUT_4[56549] = 32'b11111111111111111110101111110001;
assign LUT_4[56550] = 32'b00000000000000000100111110011101;
assign LUT_4[56551] = 32'b11111111111111111110001010010101;
assign LUT_4[56552] = 32'b00000000000000000001101111110010;
assign LUT_4[56553] = 32'b11111111111111111010111011101010;
assign LUT_4[56554] = 32'b00000000000000000001001010010110;
assign LUT_4[56555] = 32'b11111111111111111010010110001110;
assign LUT_4[56556] = 32'b11111111111111111110110000001110;
assign LUT_4[56557] = 32'b11111111111111110111111100000110;
assign LUT_4[56558] = 32'b11111111111111111110001010110010;
assign LUT_4[56559] = 32'b11111111111111110111010110101010;
assign LUT_4[56560] = 32'b00000000000000000110010101001011;
assign LUT_4[56561] = 32'b11111111111111111111100001000011;
assign LUT_4[56562] = 32'b00000000000000000101101111101111;
assign LUT_4[56563] = 32'b11111111111111111110111011100111;
assign LUT_4[56564] = 32'b00000000000000000011010101100111;
assign LUT_4[56565] = 32'b11111111111111111100100001011111;
assign LUT_4[56566] = 32'b00000000000000000010110000001011;
assign LUT_4[56567] = 32'b11111111111111111011111100000011;
assign LUT_4[56568] = 32'b11111111111111111111100001100000;
assign LUT_4[56569] = 32'b11111111111111111000101101011000;
assign LUT_4[56570] = 32'b11111111111111111110111100000100;
assign LUT_4[56571] = 32'b11111111111111111000000111111100;
assign LUT_4[56572] = 32'b11111111111111111100100001111100;
assign LUT_4[56573] = 32'b11111111111111110101101101110100;
assign LUT_4[56574] = 32'b11111111111111111011111100100000;
assign LUT_4[56575] = 32'b11111111111111110101001000011000;
assign LUT_4[56576] = 32'b00000000000000001011000110011101;
assign LUT_4[56577] = 32'b00000000000000000100010010010101;
assign LUT_4[56578] = 32'b00000000000000001010100001000001;
assign LUT_4[56579] = 32'b00000000000000000011101100111001;
assign LUT_4[56580] = 32'b00000000000000001000000110111001;
assign LUT_4[56581] = 32'b00000000000000000001010010110001;
assign LUT_4[56582] = 32'b00000000000000000111100001011101;
assign LUT_4[56583] = 32'b00000000000000000000101101010101;
assign LUT_4[56584] = 32'b00000000000000000100010010110010;
assign LUT_4[56585] = 32'b11111111111111111101011110101010;
assign LUT_4[56586] = 32'b00000000000000000011101101010110;
assign LUT_4[56587] = 32'b11111111111111111100111001001110;
assign LUT_4[56588] = 32'b00000000000000000001010011001110;
assign LUT_4[56589] = 32'b11111111111111111010011111000110;
assign LUT_4[56590] = 32'b00000000000000000000101101110010;
assign LUT_4[56591] = 32'b11111111111111111001111001101010;
assign LUT_4[56592] = 32'b00000000000000001000111000001011;
assign LUT_4[56593] = 32'b00000000000000000010000100000011;
assign LUT_4[56594] = 32'b00000000000000001000010010101111;
assign LUT_4[56595] = 32'b00000000000000000001011110100111;
assign LUT_4[56596] = 32'b00000000000000000101111000100111;
assign LUT_4[56597] = 32'b11111111111111111111000100011111;
assign LUT_4[56598] = 32'b00000000000000000101010011001011;
assign LUT_4[56599] = 32'b11111111111111111110011111000011;
assign LUT_4[56600] = 32'b00000000000000000010000100100000;
assign LUT_4[56601] = 32'b11111111111111111011010000011000;
assign LUT_4[56602] = 32'b00000000000000000001011111000100;
assign LUT_4[56603] = 32'b11111111111111111010101010111100;
assign LUT_4[56604] = 32'b11111111111111111111000100111100;
assign LUT_4[56605] = 32'b11111111111111111000010000110100;
assign LUT_4[56606] = 32'b11111111111111111110011111100000;
assign LUT_4[56607] = 32'b11111111111111110111101011011000;
assign LUT_4[56608] = 32'b00000000000000001001100001100100;
assign LUT_4[56609] = 32'b00000000000000000010101101011100;
assign LUT_4[56610] = 32'b00000000000000001000111100001000;
assign LUT_4[56611] = 32'b00000000000000000010001000000000;
assign LUT_4[56612] = 32'b00000000000000000110100010000000;
assign LUT_4[56613] = 32'b11111111111111111111101101111000;
assign LUT_4[56614] = 32'b00000000000000000101111100100100;
assign LUT_4[56615] = 32'b11111111111111111111001000011100;
assign LUT_4[56616] = 32'b00000000000000000010101101111001;
assign LUT_4[56617] = 32'b11111111111111111011111001110001;
assign LUT_4[56618] = 32'b00000000000000000010001000011101;
assign LUT_4[56619] = 32'b11111111111111111011010100010101;
assign LUT_4[56620] = 32'b11111111111111111111101110010101;
assign LUT_4[56621] = 32'b11111111111111111000111010001101;
assign LUT_4[56622] = 32'b11111111111111111111001000111001;
assign LUT_4[56623] = 32'b11111111111111111000010100110001;
assign LUT_4[56624] = 32'b00000000000000000111010011010010;
assign LUT_4[56625] = 32'b00000000000000000000011111001010;
assign LUT_4[56626] = 32'b00000000000000000110101101110110;
assign LUT_4[56627] = 32'b11111111111111111111111001101110;
assign LUT_4[56628] = 32'b00000000000000000100010011101110;
assign LUT_4[56629] = 32'b11111111111111111101011111100110;
assign LUT_4[56630] = 32'b00000000000000000011101110010010;
assign LUT_4[56631] = 32'b11111111111111111100111010001010;
assign LUT_4[56632] = 32'b00000000000000000000011111100111;
assign LUT_4[56633] = 32'b11111111111111111001101011011111;
assign LUT_4[56634] = 32'b11111111111111111111111010001011;
assign LUT_4[56635] = 32'b11111111111111111001000110000011;
assign LUT_4[56636] = 32'b11111111111111111101100000000011;
assign LUT_4[56637] = 32'b11111111111111110110101011111011;
assign LUT_4[56638] = 32'b11111111111111111100111010100111;
assign LUT_4[56639] = 32'b11111111111111110110000110011111;
assign LUT_4[56640] = 32'b00000000000000001100011101110001;
assign LUT_4[56641] = 32'b00000000000000000101101001101001;
assign LUT_4[56642] = 32'b00000000000000001011111000010101;
assign LUT_4[56643] = 32'b00000000000000000101000100001101;
assign LUT_4[56644] = 32'b00000000000000001001011110001101;
assign LUT_4[56645] = 32'b00000000000000000010101010000101;
assign LUT_4[56646] = 32'b00000000000000001000111000110001;
assign LUT_4[56647] = 32'b00000000000000000010000100101001;
assign LUT_4[56648] = 32'b00000000000000000101101010000110;
assign LUT_4[56649] = 32'b11111111111111111110110101111110;
assign LUT_4[56650] = 32'b00000000000000000101000100101010;
assign LUT_4[56651] = 32'b11111111111111111110010000100010;
assign LUT_4[56652] = 32'b00000000000000000010101010100010;
assign LUT_4[56653] = 32'b11111111111111111011110110011010;
assign LUT_4[56654] = 32'b00000000000000000010000101000110;
assign LUT_4[56655] = 32'b11111111111111111011010000111110;
assign LUT_4[56656] = 32'b00000000000000001010001111011111;
assign LUT_4[56657] = 32'b00000000000000000011011011010111;
assign LUT_4[56658] = 32'b00000000000000001001101010000011;
assign LUT_4[56659] = 32'b00000000000000000010110101111011;
assign LUT_4[56660] = 32'b00000000000000000111001111111011;
assign LUT_4[56661] = 32'b00000000000000000000011011110011;
assign LUT_4[56662] = 32'b00000000000000000110101010011111;
assign LUT_4[56663] = 32'b11111111111111111111110110010111;
assign LUT_4[56664] = 32'b00000000000000000011011011110100;
assign LUT_4[56665] = 32'b11111111111111111100100111101100;
assign LUT_4[56666] = 32'b00000000000000000010110110011000;
assign LUT_4[56667] = 32'b11111111111111111100000010010000;
assign LUT_4[56668] = 32'b00000000000000000000011100010000;
assign LUT_4[56669] = 32'b11111111111111111001101000001000;
assign LUT_4[56670] = 32'b11111111111111111111110110110100;
assign LUT_4[56671] = 32'b11111111111111111001000010101100;
assign LUT_4[56672] = 32'b00000000000000001010111000111000;
assign LUT_4[56673] = 32'b00000000000000000100000100110000;
assign LUT_4[56674] = 32'b00000000000000001010010011011100;
assign LUT_4[56675] = 32'b00000000000000000011011111010100;
assign LUT_4[56676] = 32'b00000000000000000111111001010100;
assign LUT_4[56677] = 32'b00000000000000000001000101001100;
assign LUT_4[56678] = 32'b00000000000000000111010011111000;
assign LUT_4[56679] = 32'b00000000000000000000011111110000;
assign LUT_4[56680] = 32'b00000000000000000100000101001101;
assign LUT_4[56681] = 32'b11111111111111111101010001000101;
assign LUT_4[56682] = 32'b00000000000000000011011111110001;
assign LUT_4[56683] = 32'b11111111111111111100101011101001;
assign LUT_4[56684] = 32'b00000000000000000001000101101001;
assign LUT_4[56685] = 32'b11111111111111111010010001100001;
assign LUT_4[56686] = 32'b00000000000000000000100000001101;
assign LUT_4[56687] = 32'b11111111111111111001101100000101;
assign LUT_4[56688] = 32'b00000000000000001000101010100110;
assign LUT_4[56689] = 32'b00000000000000000001110110011110;
assign LUT_4[56690] = 32'b00000000000000001000000101001010;
assign LUT_4[56691] = 32'b00000000000000000001010001000010;
assign LUT_4[56692] = 32'b00000000000000000101101011000010;
assign LUT_4[56693] = 32'b11111111111111111110110110111010;
assign LUT_4[56694] = 32'b00000000000000000101000101100110;
assign LUT_4[56695] = 32'b11111111111111111110010001011110;
assign LUT_4[56696] = 32'b00000000000000000001110110111011;
assign LUT_4[56697] = 32'b11111111111111111011000010110011;
assign LUT_4[56698] = 32'b00000000000000000001010001011111;
assign LUT_4[56699] = 32'b11111111111111111010011101010111;
assign LUT_4[56700] = 32'b11111111111111111110110111010111;
assign LUT_4[56701] = 32'b11111111111111111000000011001111;
assign LUT_4[56702] = 32'b11111111111111111110010001111011;
assign LUT_4[56703] = 32'b11111111111111110111011101110011;
assign LUT_4[56704] = 32'b00000000000000001101101100100101;
assign LUT_4[56705] = 32'b00000000000000000110111000011101;
assign LUT_4[56706] = 32'b00000000000000001101000111001001;
assign LUT_4[56707] = 32'b00000000000000000110010011000001;
assign LUT_4[56708] = 32'b00000000000000001010101101000001;
assign LUT_4[56709] = 32'b00000000000000000011111000111001;
assign LUT_4[56710] = 32'b00000000000000001010000111100101;
assign LUT_4[56711] = 32'b00000000000000000011010011011101;
assign LUT_4[56712] = 32'b00000000000000000110111000111010;
assign LUT_4[56713] = 32'b00000000000000000000000100110010;
assign LUT_4[56714] = 32'b00000000000000000110010011011110;
assign LUT_4[56715] = 32'b11111111111111111111011111010110;
assign LUT_4[56716] = 32'b00000000000000000011111001010110;
assign LUT_4[56717] = 32'b11111111111111111101000101001110;
assign LUT_4[56718] = 32'b00000000000000000011010011111010;
assign LUT_4[56719] = 32'b11111111111111111100011111110010;
assign LUT_4[56720] = 32'b00000000000000001011011110010011;
assign LUT_4[56721] = 32'b00000000000000000100101010001011;
assign LUT_4[56722] = 32'b00000000000000001010111000110111;
assign LUT_4[56723] = 32'b00000000000000000100000100101111;
assign LUT_4[56724] = 32'b00000000000000001000011110101111;
assign LUT_4[56725] = 32'b00000000000000000001101010100111;
assign LUT_4[56726] = 32'b00000000000000000111111001010011;
assign LUT_4[56727] = 32'b00000000000000000001000101001011;
assign LUT_4[56728] = 32'b00000000000000000100101010101000;
assign LUT_4[56729] = 32'b11111111111111111101110110100000;
assign LUT_4[56730] = 32'b00000000000000000100000101001100;
assign LUT_4[56731] = 32'b11111111111111111101010001000100;
assign LUT_4[56732] = 32'b00000000000000000001101011000100;
assign LUT_4[56733] = 32'b11111111111111111010110110111100;
assign LUT_4[56734] = 32'b00000000000000000001000101101000;
assign LUT_4[56735] = 32'b11111111111111111010010001100000;
assign LUT_4[56736] = 32'b00000000000000001100000111101100;
assign LUT_4[56737] = 32'b00000000000000000101010011100100;
assign LUT_4[56738] = 32'b00000000000000001011100010010000;
assign LUT_4[56739] = 32'b00000000000000000100101110001000;
assign LUT_4[56740] = 32'b00000000000000001001001000001000;
assign LUT_4[56741] = 32'b00000000000000000010010100000000;
assign LUT_4[56742] = 32'b00000000000000001000100010101100;
assign LUT_4[56743] = 32'b00000000000000000001101110100100;
assign LUT_4[56744] = 32'b00000000000000000101010100000001;
assign LUT_4[56745] = 32'b11111111111111111110011111111001;
assign LUT_4[56746] = 32'b00000000000000000100101110100101;
assign LUT_4[56747] = 32'b11111111111111111101111010011101;
assign LUT_4[56748] = 32'b00000000000000000010010100011101;
assign LUT_4[56749] = 32'b11111111111111111011100000010101;
assign LUT_4[56750] = 32'b00000000000000000001101111000001;
assign LUT_4[56751] = 32'b11111111111111111010111010111001;
assign LUT_4[56752] = 32'b00000000000000001001111001011010;
assign LUT_4[56753] = 32'b00000000000000000011000101010010;
assign LUT_4[56754] = 32'b00000000000000001001010011111110;
assign LUT_4[56755] = 32'b00000000000000000010011111110110;
assign LUT_4[56756] = 32'b00000000000000000110111001110110;
assign LUT_4[56757] = 32'b00000000000000000000000101101110;
assign LUT_4[56758] = 32'b00000000000000000110010100011010;
assign LUT_4[56759] = 32'b11111111111111111111100000010010;
assign LUT_4[56760] = 32'b00000000000000000011000101101111;
assign LUT_4[56761] = 32'b11111111111111111100010001100111;
assign LUT_4[56762] = 32'b00000000000000000010100000010011;
assign LUT_4[56763] = 32'b11111111111111111011101100001011;
assign LUT_4[56764] = 32'b00000000000000000000000110001011;
assign LUT_4[56765] = 32'b11111111111111111001010010000011;
assign LUT_4[56766] = 32'b11111111111111111111100000101111;
assign LUT_4[56767] = 32'b11111111111111111000101100100111;
assign LUT_4[56768] = 32'b00000000000000001111000011111001;
assign LUT_4[56769] = 32'b00000000000000001000001111110001;
assign LUT_4[56770] = 32'b00000000000000001110011110011101;
assign LUT_4[56771] = 32'b00000000000000000111101010010101;
assign LUT_4[56772] = 32'b00000000000000001100000100010101;
assign LUT_4[56773] = 32'b00000000000000000101010000001101;
assign LUT_4[56774] = 32'b00000000000000001011011110111001;
assign LUT_4[56775] = 32'b00000000000000000100101010110001;
assign LUT_4[56776] = 32'b00000000000000001000010000001110;
assign LUT_4[56777] = 32'b00000000000000000001011100000110;
assign LUT_4[56778] = 32'b00000000000000000111101010110010;
assign LUT_4[56779] = 32'b00000000000000000000110110101010;
assign LUT_4[56780] = 32'b00000000000000000101010000101010;
assign LUT_4[56781] = 32'b11111111111111111110011100100010;
assign LUT_4[56782] = 32'b00000000000000000100101011001110;
assign LUT_4[56783] = 32'b11111111111111111101110111000110;
assign LUT_4[56784] = 32'b00000000000000001100110101100111;
assign LUT_4[56785] = 32'b00000000000000000110000001011111;
assign LUT_4[56786] = 32'b00000000000000001100010000001011;
assign LUT_4[56787] = 32'b00000000000000000101011100000011;
assign LUT_4[56788] = 32'b00000000000000001001110110000011;
assign LUT_4[56789] = 32'b00000000000000000011000001111011;
assign LUT_4[56790] = 32'b00000000000000001001010000100111;
assign LUT_4[56791] = 32'b00000000000000000010011100011111;
assign LUT_4[56792] = 32'b00000000000000000110000001111100;
assign LUT_4[56793] = 32'b11111111111111111111001101110100;
assign LUT_4[56794] = 32'b00000000000000000101011100100000;
assign LUT_4[56795] = 32'b11111111111111111110101000011000;
assign LUT_4[56796] = 32'b00000000000000000011000010011000;
assign LUT_4[56797] = 32'b11111111111111111100001110010000;
assign LUT_4[56798] = 32'b00000000000000000010011100111100;
assign LUT_4[56799] = 32'b11111111111111111011101000110100;
assign LUT_4[56800] = 32'b00000000000000001101011111000000;
assign LUT_4[56801] = 32'b00000000000000000110101010111000;
assign LUT_4[56802] = 32'b00000000000000001100111001100100;
assign LUT_4[56803] = 32'b00000000000000000110000101011100;
assign LUT_4[56804] = 32'b00000000000000001010011111011100;
assign LUT_4[56805] = 32'b00000000000000000011101011010100;
assign LUT_4[56806] = 32'b00000000000000001001111010000000;
assign LUT_4[56807] = 32'b00000000000000000011000101111000;
assign LUT_4[56808] = 32'b00000000000000000110101011010101;
assign LUT_4[56809] = 32'b11111111111111111111110111001101;
assign LUT_4[56810] = 32'b00000000000000000110000101111001;
assign LUT_4[56811] = 32'b11111111111111111111010001110001;
assign LUT_4[56812] = 32'b00000000000000000011101011110001;
assign LUT_4[56813] = 32'b11111111111111111100110111101001;
assign LUT_4[56814] = 32'b00000000000000000011000110010101;
assign LUT_4[56815] = 32'b11111111111111111100010010001101;
assign LUT_4[56816] = 32'b00000000000000001011010000101110;
assign LUT_4[56817] = 32'b00000000000000000100011100100110;
assign LUT_4[56818] = 32'b00000000000000001010101011010010;
assign LUT_4[56819] = 32'b00000000000000000011110111001010;
assign LUT_4[56820] = 32'b00000000000000001000010001001010;
assign LUT_4[56821] = 32'b00000000000000000001011101000010;
assign LUT_4[56822] = 32'b00000000000000000111101011101110;
assign LUT_4[56823] = 32'b00000000000000000000110111100110;
assign LUT_4[56824] = 32'b00000000000000000100011101000011;
assign LUT_4[56825] = 32'b11111111111111111101101000111011;
assign LUT_4[56826] = 32'b00000000000000000011110111100111;
assign LUT_4[56827] = 32'b11111111111111111101000011011111;
assign LUT_4[56828] = 32'b00000000000000000001011101011111;
assign LUT_4[56829] = 32'b11111111111111111010101001010111;
assign LUT_4[56830] = 32'b00000000000000000000111000000011;
assign LUT_4[56831] = 32'b11111111111111111010000011111011;
assign LUT_4[56832] = 32'b00000000000000000101001111000010;
assign LUT_4[56833] = 32'b11111111111111111110011010111010;
assign LUT_4[56834] = 32'b00000000000000000100101001100110;
assign LUT_4[56835] = 32'b11111111111111111101110101011110;
assign LUT_4[56836] = 32'b00000000000000000010001111011110;
assign LUT_4[56837] = 32'b11111111111111111011011011010110;
assign LUT_4[56838] = 32'b00000000000000000001101010000010;
assign LUT_4[56839] = 32'b11111111111111111010110101111010;
assign LUT_4[56840] = 32'b11111111111111111110011011010111;
assign LUT_4[56841] = 32'b11111111111111110111100111001111;
assign LUT_4[56842] = 32'b11111111111111111101110101111011;
assign LUT_4[56843] = 32'b11111111111111110111000001110011;
assign LUT_4[56844] = 32'b11111111111111111011011011110011;
assign LUT_4[56845] = 32'b11111111111111110100100111101011;
assign LUT_4[56846] = 32'b11111111111111111010110110010111;
assign LUT_4[56847] = 32'b11111111111111110100000010001111;
assign LUT_4[56848] = 32'b00000000000000000011000000110000;
assign LUT_4[56849] = 32'b11111111111111111100001100101000;
assign LUT_4[56850] = 32'b00000000000000000010011011010100;
assign LUT_4[56851] = 32'b11111111111111111011100111001100;
assign LUT_4[56852] = 32'b00000000000000000000000001001100;
assign LUT_4[56853] = 32'b11111111111111111001001101000100;
assign LUT_4[56854] = 32'b11111111111111111111011011110000;
assign LUT_4[56855] = 32'b11111111111111111000100111101000;
assign LUT_4[56856] = 32'b11111111111111111100001101000101;
assign LUT_4[56857] = 32'b11111111111111110101011000111101;
assign LUT_4[56858] = 32'b11111111111111111011100111101001;
assign LUT_4[56859] = 32'b11111111111111110100110011100001;
assign LUT_4[56860] = 32'b11111111111111111001001101100001;
assign LUT_4[56861] = 32'b11111111111111110010011001011001;
assign LUT_4[56862] = 32'b11111111111111111000101000000101;
assign LUT_4[56863] = 32'b11111111111111110001110011111101;
assign LUT_4[56864] = 32'b00000000000000000011101010001001;
assign LUT_4[56865] = 32'b11111111111111111100110110000001;
assign LUT_4[56866] = 32'b00000000000000000011000100101101;
assign LUT_4[56867] = 32'b11111111111111111100010000100101;
assign LUT_4[56868] = 32'b00000000000000000000101010100101;
assign LUT_4[56869] = 32'b11111111111111111001110110011101;
assign LUT_4[56870] = 32'b00000000000000000000000101001001;
assign LUT_4[56871] = 32'b11111111111111111001010001000001;
assign LUT_4[56872] = 32'b11111111111111111100110110011110;
assign LUT_4[56873] = 32'b11111111111111110110000010010110;
assign LUT_4[56874] = 32'b11111111111111111100010001000010;
assign LUT_4[56875] = 32'b11111111111111110101011100111010;
assign LUT_4[56876] = 32'b11111111111111111001110110111010;
assign LUT_4[56877] = 32'b11111111111111110011000010110010;
assign LUT_4[56878] = 32'b11111111111111111001010001011110;
assign LUT_4[56879] = 32'b11111111111111110010011101010110;
assign LUT_4[56880] = 32'b00000000000000000001011011110111;
assign LUT_4[56881] = 32'b11111111111111111010100111101111;
assign LUT_4[56882] = 32'b00000000000000000000110110011011;
assign LUT_4[56883] = 32'b11111111111111111010000010010011;
assign LUT_4[56884] = 32'b11111111111111111110011100010011;
assign LUT_4[56885] = 32'b11111111111111110111101000001011;
assign LUT_4[56886] = 32'b11111111111111111101110110110111;
assign LUT_4[56887] = 32'b11111111111111110111000010101111;
assign LUT_4[56888] = 32'b11111111111111111010101000001100;
assign LUT_4[56889] = 32'b11111111111111110011110100000100;
assign LUT_4[56890] = 32'b11111111111111111010000010110000;
assign LUT_4[56891] = 32'b11111111111111110011001110101000;
assign LUT_4[56892] = 32'b11111111111111110111101000101000;
assign LUT_4[56893] = 32'b11111111111111110000110100100000;
assign LUT_4[56894] = 32'b11111111111111110111000011001100;
assign LUT_4[56895] = 32'b11111111111111110000001111000100;
assign LUT_4[56896] = 32'b00000000000000000110100110010110;
assign LUT_4[56897] = 32'b11111111111111111111110010001110;
assign LUT_4[56898] = 32'b00000000000000000110000000111010;
assign LUT_4[56899] = 32'b11111111111111111111001100110010;
assign LUT_4[56900] = 32'b00000000000000000011100110110010;
assign LUT_4[56901] = 32'b11111111111111111100110010101010;
assign LUT_4[56902] = 32'b00000000000000000011000001010110;
assign LUT_4[56903] = 32'b11111111111111111100001101001110;
assign LUT_4[56904] = 32'b11111111111111111111110010101011;
assign LUT_4[56905] = 32'b11111111111111111000111110100011;
assign LUT_4[56906] = 32'b11111111111111111111001101001111;
assign LUT_4[56907] = 32'b11111111111111111000011001000111;
assign LUT_4[56908] = 32'b11111111111111111100110011000111;
assign LUT_4[56909] = 32'b11111111111111110101111110111111;
assign LUT_4[56910] = 32'b11111111111111111100001101101011;
assign LUT_4[56911] = 32'b11111111111111110101011001100011;
assign LUT_4[56912] = 32'b00000000000000000100011000000100;
assign LUT_4[56913] = 32'b11111111111111111101100011111100;
assign LUT_4[56914] = 32'b00000000000000000011110010101000;
assign LUT_4[56915] = 32'b11111111111111111100111110100000;
assign LUT_4[56916] = 32'b00000000000000000001011000100000;
assign LUT_4[56917] = 32'b11111111111111111010100100011000;
assign LUT_4[56918] = 32'b00000000000000000000110011000100;
assign LUT_4[56919] = 32'b11111111111111111001111110111100;
assign LUT_4[56920] = 32'b11111111111111111101100100011001;
assign LUT_4[56921] = 32'b11111111111111110110110000010001;
assign LUT_4[56922] = 32'b11111111111111111100111110111101;
assign LUT_4[56923] = 32'b11111111111111110110001010110101;
assign LUT_4[56924] = 32'b11111111111111111010100100110101;
assign LUT_4[56925] = 32'b11111111111111110011110000101101;
assign LUT_4[56926] = 32'b11111111111111111001111111011001;
assign LUT_4[56927] = 32'b11111111111111110011001011010001;
assign LUT_4[56928] = 32'b00000000000000000101000001011101;
assign LUT_4[56929] = 32'b11111111111111111110001101010101;
assign LUT_4[56930] = 32'b00000000000000000100011100000001;
assign LUT_4[56931] = 32'b11111111111111111101100111111001;
assign LUT_4[56932] = 32'b00000000000000000010000001111001;
assign LUT_4[56933] = 32'b11111111111111111011001101110001;
assign LUT_4[56934] = 32'b00000000000000000001011100011101;
assign LUT_4[56935] = 32'b11111111111111111010101000010101;
assign LUT_4[56936] = 32'b11111111111111111110001101110010;
assign LUT_4[56937] = 32'b11111111111111110111011001101010;
assign LUT_4[56938] = 32'b11111111111111111101101000010110;
assign LUT_4[56939] = 32'b11111111111111110110110100001110;
assign LUT_4[56940] = 32'b11111111111111111011001110001110;
assign LUT_4[56941] = 32'b11111111111111110100011010000110;
assign LUT_4[56942] = 32'b11111111111111111010101000110010;
assign LUT_4[56943] = 32'b11111111111111110011110100101010;
assign LUT_4[56944] = 32'b00000000000000000010110011001011;
assign LUT_4[56945] = 32'b11111111111111111011111111000011;
assign LUT_4[56946] = 32'b00000000000000000010001101101111;
assign LUT_4[56947] = 32'b11111111111111111011011001100111;
assign LUT_4[56948] = 32'b11111111111111111111110011100111;
assign LUT_4[56949] = 32'b11111111111111111000111111011111;
assign LUT_4[56950] = 32'b11111111111111111111001110001011;
assign LUT_4[56951] = 32'b11111111111111111000011010000011;
assign LUT_4[56952] = 32'b11111111111111111011111111100000;
assign LUT_4[56953] = 32'b11111111111111110101001011011000;
assign LUT_4[56954] = 32'b11111111111111111011011010000100;
assign LUT_4[56955] = 32'b11111111111111110100100101111100;
assign LUT_4[56956] = 32'b11111111111111111000111111111100;
assign LUT_4[56957] = 32'b11111111111111110010001011110100;
assign LUT_4[56958] = 32'b11111111111111111000011010100000;
assign LUT_4[56959] = 32'b11111111111111110001100110011000;
assign LUT_4[56960] = 32'b00000000000000000111110101001010;
assign LUT_4[56961] = 32'b00000000000000000001000001000010;
assign LUT_4[56962] = 32'b00000000000000000111001111101110;
assign LUT_4[56963] = 32'b00000000000000000000011011100110;
assign LUT_4[56964] = 32'b00000000000000000100110101100110;
assign LUT_4[56965] = 32'b11111111111111111110000001011110;
assign LUT_4[56966] = 32'b00000000000000000100010000001010;
assign LUT_4[56967] = 32'b11111111111111111101011100000010;
assign LUT_4[56968] = 32'b00000000000000000001000001011111;
assign LUT_4[56969] = 32'b11111111111111111010001101010111;
assign LUT_4[56970] = 32'b00000000000000000000011100000011;
assign LUT_4[56971] = 32'b11111111111111111001100111111011;
assign LUT_4[56972] = 32'b11111111111111111110000001111011;
assign LUT_4[56973] = 32'b11111111111111110111001101110011;
assign LUT_4[56974] = 32'b11111111111111111101011100011111;
assign LUT_4[56975] = 32'b11111111111111110110101000010111;
assign LUT_4[56976] = 32'b00000000000000000101100110111000;
assign LUT_4[56977] = 32'b11111111111111111110110010110000;
assign LUT_4[56978] = 32'b00000000000000000101000001011100;
assign LUT_4[56979] = 32'b11111111111111111110001101010100;
assign LUT_4[56980] = 32'b00000000000000000010100111010100;
assign LUT_4[56981] = 32'b11111111111111111011110011001100;
assign LUT_4[56982] = 32'b00000000000000000010000001111000;
assign LUT_4[56983] = 32'b11111111111111111011001101110000;
assign LUT_4[56984] = 32'b11111111111111111110110011001101;
assign LUT_4[56985] = 32'b11111111111111110111111111000101;
assign LUT_4[56986] = 32'b11111111111111111110001101110001;
assign LUT_4[56987] = 32'b11111111111111110111011001101001;
assign LUT_4[56988] = 32'b11111111111111111011110011101001;
assign LUT_4[56989] = 32'b11111111111111110100111111100001;
assign LUT_4[56990] = 32'b11111111111111111011001110001101;
assign LUT_4[56991] = 32'b11111111111111110100011010000101;
assign LUT_4[56992] = 32'b00000000000000000110010000010001;
assign LUT_4[56993] = 32'b11111111111111111111011100001001;
assign LUT_4[56994] = 32'b00000000000000000101101010110101;
assign LUT_4[56995] = 32'b11111111111111111110110110101101;
assign LUT_4[56996] = 32'b00000000000000000011010000101101;
assign LUT_4[56997] = 32'b11111111111111111100011100100101;
assign LUT_4[56998] = 32'b00000000000000000010101011010001;
assign LUT_4[56999] = 32'b11111111111111111011110111001001;
assign LUT_4[57000] = 32'b11111111111111111111011100100110;
assign LUT_4[57001] = 32'b11111111111111111000101000011110;
assign LUT_4[57002] = 32'b11111111111111111110110111001010;
assign LUT_4[57003] = 32'b11111111111111111000000011000010;
assign LUT_4[57004] = 32'b11111111111111111100011101000010;
assign LUT_4[57005] = 32'b11111111111111110101101000111010;
assign LUT_4[57006] = 32'b11111111111111111011110111100110;
assign LUT_4[57007] = 32'b11111111111111110101000011011110;
assign LUT_4[57008] = 32'b00000000000000000100000001111111;
assign LUT_4[57009] = 32'b11111111111111111101001101110111;
assign LUT_4[57010] = 32'b00000000000000000011011100100011;
assign LUT_4[57011] = 32'b11111111111111111100101000011011;
assign LUT_4[57012] = 32'b00000000000000000001000010011011;
assign LUT_4[57013] = 32'b11111111111111111010001110010011;
assign LUT_4[57014] = 32'b00000000000000000000011100111111;
assign LUT_4[57015] = 32'b11111111111111111001101000110111;
assign LUT_4[57016] = 32'b11111111111111111101001110010100;
assign LUT_4[57017] = 32'b11111111111111110110011010001100;
assign LUT_4[57018] = 32'b11111111111111111100101000111000;
assign LUT_4[57019] = 32'b11111111111111110101110100110000;
assign LUT_4[57020] = 32'b11111111111111111010001110110000;
assign LUT_4[57021] = 32'b11111111111111110011011010101000;
assign LUT_4[57022] = 32'b11111111111111111001101001010100;
assign LUT_4[57023] = 32'b11111111111111110010110101001100;
assign LUT_4[57024] = 32'b00000000000000001001001100011110;
assign LUT_4[57025] = 32'b00000000000000000010011000010110;
assign LUT_4[57026] = 32'b00000000000000001000100111000010;
assign LUT_4[57027] = 32'b00000000000000000001110010111010;
assign LUT_4[57028] = 32'b00000000000000000110001100111010;
assign LUT_4[57029] = 32'b11111111111111111111011000110010;
assign LUT_4[57030] = 32'b00000000000000000101100111011110;
assign LUT_4[57031] = 32'b11111111111111111110110011010110;
assign LUT_4[57032] = 32'b00000000000000000010011000110011;
assign LUT_4[57033] = 32'b11111111111111111011100100101011;
assign LUT_4[57034] = 32'b00000000000000000001110011010111;
assign LUT_4[57035] = 32'b11111111111111111010111111001111;
assign LUT_4[57036] = 32'b11111111111111111111011001001111;
assign LUT_4[57037] = 32'b11111111111111111000100101000111;
assign LUT_4[57038] = 32'b11111111111111111110110011110011;
assign LUT_4[57039] = 32'b11111111111111110111111111101011;
assign LUT_4[57040] = 32'b00000000000000000110111110001100;
assign LUT_4[57041] = 32'b00000000000000000000001010000100;
assign LUT_4[57042] = 32'b00000000000000000110011000110000;
assign LUT_4[57043] = 32'b11111111111111111111100100101000;
assign LUT_4[57044] = 32'b00000000000000000011111110101000;
assign LUT_4[57045] = 32'b11111111111111111101001010100000;
assign LUT_4[57046] = 32'b00000000000000000011011001001100;
assign LUT_4[57047] = 32'b11111111111111111100100101000100;
assign LUT_4[57048] = 32'b00000000000000000000001010100001;
assign LUT_4[57049] = 32'b11111111111111111001010110011001;
assign LUT_4[57050] = 32'b11111111111111111111100101000101;
assign LUT_4[57051] = 32'b11111111111111111000110000111101;
assign LUT_4[57052] = 32'b11111111111111111101001010111101;
assign LUT_4[57053] = 32'b11111111111111110110010110110101;
assign LUT_4[57054] = 32'b11111111111111111100100101100001;
assign LUT_4[57055] = 32'b11111111111111110101110001011001;
assign LUT_4[57056] = 32'b00000000000000000111100111100101;
assign LUT_4[57057] = 32'b00000000000000000000110011011101;
assign LUT_4[57058] = 32'b00000000000000000111000010001001;
assign LUT_4[57059] = 32'b00000000000000000000001110000001;
assign LUT_4[57060] = 32'b00000000000000000100101000000001;
assign LUT_4[57061] = 32'b11111111111111111101110011111001;
assign LUT_4[57062] = 32'b00000000000000000100000010100101;
assign LUT_4[57063] = 32'b11111111111111111101001110011101;
assign LUT_4[57064] = 32'b00000000000000000000110011111010;
assign LUT_4[57065] = 32'b11111111111111111001111111110010;
assign LUT_4[57066] = 32'b00000000000000000000001110011110;
assign LUT_4[57067] = 32'b11111111111111111001011010010110;
assign LUT_4[57068] = 32'b11111111111111111101110100010110;
assign LUT_4[57069] = 32'b11111111111111110111000000001110;
assign LUT_4[57070] = 32'b11111111111111111101001110111010;
assign LUT_4[57071] = 32'b11111111111111110110011010110010;
assign LUT_4[57072] = 32'b00000000000000000101011001010011;
assign LUT_4[57073] = 32'b11111111111111111110100101001011;
assign LUT_4[57074] = 32'b00000000000000000100110011110111;
assign LUT_4[57075] = 32'b11111111111111111101111111101111;
assign LUT_4[57076] = 32'b00000000000000000010011001101111;
assign LUT_4[57077] = 32'b11111111111111111011100101100111;
assign LUT_4[57078] = 32'b00000000000000000001110100010011;
assign LUT_4[57079] = 32'b11111111111111111011000000001011;
assign LUT_4[57080] = 32'b11111111111111111110100101101000;
assign LUT_4[57081] = 32'b11111111111111110111110001100000;
assign LUT_4[57082] = 32'b11111111111111111110000000001100;
assign LUT_4[57083] = 32'b11111111111111110111001100000100;
assign LUT_4[57084] = 32'b11111111111111111011100110000100;
assign LUT_4[57085] = 32'b11111111111111110100110001111100;
assign LUT_4[57086] = 32'b11111111111111111011000000101000;
assign LUT_4[57087] = 32'b11111111111111110100001100100000;
assign LUT_4[57088] = 32'b00000000000000001010001010100101;
assign LUT_4[57089] = 32'b00000000000000000011010110011101;
assign LUT_4[57090] = 32'b00000000000000001001100101001001;
assign LUT_4[57091] = 32'b00000000000000000010110001000001;
assign LUT_4[57092] = 32'b00000000000000000111001011000001;
assign LUT_4[57093] = 32'b00000000000000000000010110111001;
assign LUT_4[57094] = 32'b00000000000000000110100101100101;
assign LUT_4[57095] = 32'b11111111111111111111110001011101;
assign LUT_4[57096] = 32'b00000000000000000011010110111010;
assign LUT_4[57097] = 32'b11111111111111111100100010110010;
assign LUT_4[57098] = 32'b00000000000000000010110001011110;
assign LUT_4[57099] = 32'b11111111111111111011111101010110;
assign LUT_4[57100] = 32'b00000000000000000000010111010110;
assign LUT_4[57101] = 32'b11111111111111111001100011001110;
assign LUT_4[57102] = 32'b11111111111111111111110001111010;
assign LUT_4[57103] = 32'b11111111111111111000111101110010;
assign LUT_4[57104] = 32'b00000000000000000111111100010011;
assign LUT_4[57105] = 32'b00000000000000000001001000001011;
assign LUT_4[57106] = 32'b00000000000000000111010110110111;
assign LUT_4[57107] = 32'b00000000000000000000100010101111;
assign LUT_4[57108] = 32'b00000000000000000100111100101111;
assign LUT_4[57109] = 32'b11111111111111111110001000100111;
assign LUT_4[57110] = 32'b00000000000000000100010111010011;
assign LUT_4[57111] = 32'b11111111111111111101100011001011;
assign LUT_4[57112] = 32'b00000000000000000001001000101000;
assign LUT_4[57113] = 32'b11111111111111111010010100100000;
assign LUT_4[57114] = 32'b00000000000000000000100011001100;
assign LUT_4[57115] = 32'b11111111111111111001101111000100;
assign LUT_4[57116] = 32'b11111111111111111110001001000100;
assign LUT_4[57117] = 32'b11111111111111110111010100111100;
assign LUT_4[57118] = 32'b11111111111111111101100011101000;
assign LUT_4[57119] = 32'b11111111111111110110101111100000;
assign LUT_4[57120] = 32'b00000000000000001000100101101100;
assign LUT_4[57121] = 32'b00000000000000000001110001100100;
assign LUT_4[57122] = 32'b00000000000000001000000000010000;
assign LUT_4[57123] = 32'b00000000000000000001001100001000;
assign LUT_4[57124] = 32'b00000000000000000101100110001000;
assign LUT_4[57125] = 32'b11111111111111111110110010000000;
assign LUT_4[57126] = 32'b00000000000000000101000000101100;
assign LUT_4[57127] = 32'b11111111111111111110001100100100;
assign LUT_4[57128] = 32'b00000000000000000001110010000001;
assign LUT_4[57129] = 32'b11111111111111111010111101111001;
assign LUT_4[57130] = 32'b00000000000000000001001100100101;
assign LUT_4[57131] = 32'b11111111111111111010011000011101;
assign LUT_4[57132] = 32'b11111111111111111110110010011101;
assign LUT_4[57133] = 32'b11111111111111110111111110010101;
assign LUT_4[57134] = 32'b11111111111111111110001101000001;
assign LUT_4[57135] = 32'b11111111111111110111011000111001;
assign LUT_4[57136] = 32'b00000000000000000110010111011010;
assign LUT_4[57137] = 32'b11111111111111111111100011010010;
assign LUT_4[57138] = 32'b00000000000000000101110001111110;
assign LUT_4[57139] = 32'b11111111111111111110111101110110;
assign LUT_4[57140] = 32'b00000000000000000011010111110110;
assign LUT_4[57141] = 32'b11111111111111111100100011101110;
assign LUT_4[57142] = 32'b00000000000000000010110010011010;
assign LUT_4[57143] = 32'b11111111111111111011111110010010;
assign LUT_4[57144] = 32'b11111111111111111111100011101111;
assign LUT_4[57145] = 32'b11111111111111111000101111100111;
assign LUT_4[57146] = 32'b11111111111111111110111110010011;
assign LUT_4[57147] = 32'b11111111111111111000001010001011;
assign LUT_4[57148] = 32'b11111111111111111100100100001011;
assign LUT_4[57149] = 32'b11111111111111110101110000000011;
assign LUT_4[57150] = 32'b11111111111111111011111110101111;
assign LUT_4[57151] = 32'b11111111111111110101001010100111;
assign LUT_4[57152] = 32'b00000000000000001011100001111001;
assign LUT_4[57153] = 32'b00000000000000000100101101110001;
assign LUT_4[57154] = 32'b00000000000000001010111100011101;
assign LUT_4[57155] = 32'b00000000000000000100001000010101;
assign LUT_4[57156] = 32'b00000000000000001000100010010101;
assign LUT_4[57157] = 32'b00000000000000000001101110001101;
assign LUT_4[57158] = 32'b00000000000000000111111100111001;
assign LUT_4[57159] = 32'b00000000000000000001001000110001;
assign LUT_4[57160] = 32'b00000000000000000100101110001110;
assign LUT_4[57161] = 32'b11111111111111111101111010000110;
assign LUT_4[57162] = 32'b00000000000000000100001000110010;
assign LUT_4[57163] = 32'b11111111111111111101010100101010;
assign LUT_4[57164] = 32'b00000000000000000001101110101010;
assign LUT_4[57165] = 32'b11111111111111111010111010100010;
assign LUT_4[57166] = 32'b00000000000000000001001001001110;
assign LUT_4[57167] = 32'b11111111111111111010010101000110;
assign LUT_4[57168] = 32'b00000000000000001001010011100111;
assign LUT_4[57169] = 32'b00000000000000000010011111011111;
assign LUT_4[57170] = 32'b00000000000000001000101110001011;
assign LUT_4[57171] = 32'b00000000000000000001111010000011;
assign LUT_4[57172] = 32'b00000000000000000110010100000011;
assign LUT_4[57173] = 32'b11111111111111111111011111111011;
assign LUT_4[57174] = 32'b00000000000000000101101110100111;
assign LUT_4[57175] = 32'b11111111111111111110111010011111;
assign LUT_4[57176] = 32'b00000000000000000010011111111100;
assign LUT_4[57177] = 32'b11111111111111111011101011110100;
assign LUT_4[57178] = 32'b00000000000000000001111010100000;
assign LUT_4[57179] = 32'b11111111111111111011000110011000;
assign LUT_4[57180] = 32'b11111111111111111111100000011000;
assign LUT_4[57181] = 32'b11111111111111111000101100010000;
assign LUT_4[57182] = 32'b11111111111111111110111010111100;
assign LUT_4[57183] = 32'b11111111111111111000000110110100;
assign LUT_4[57184] = 32'b00000000000000001001111101000000;
assign LUT_4[57185] = 32'b00000000000000000011001000111000;
assign LUT_4[57186] = 32'b00000000000000001001010111100100;
assign LUT_4[57187] = 32'b00000000000000000010100011011100;
assign LUT_4[57188] = 32'b00000000000000000110111101011100;
assign LUT_4[57189] = 32'b00000000000000000000001001010100;
assign LUT_4[57190] = 32'b00000000000000000110011000000000;
assign LUT_4[57191] = 32'b11111111111111111111100011111000;
assign LUT_4[57192] = 32'b00000000000000000011001001010101;
assign LUT_4[57193] = 32'b11111111111111111100010101001101;
assign LUT_4[57194] = 32'b00000000000000000010100011111001;
assign LUT_4[57195] = 32'b11111111111111111011101111110001;
assign LUT_4[57196] = 32'b00000000000000000000001001110001;
assign LUT_4[57197] = 32'b11111111111111111001010101101001;
assign LUT_4[57198] = 32'b11111111111111111111100100010101;
assign LUT_4[57199] = 32'b11111111111111111000110000001101;
assign LUT_4[57200] = 32'b00000000000000000111101110101110;
assign LUT_4[57201] = 32'b00000000000000000000111010100110;
assign LUT_4[57202] = 32'b00000000000000000111001001010010;
assign LUT_4[57203] = 32'b00000000000000000000010101001010;
assign LUT_4[57204] = 32'b00000000000000000100101111001010;
assign LUT_4[57205] = 32'b11111111111111111101111011000010;
assign LUT_4[57206] = 32'b00000000000000000100001001101110;
assign LUT_4[57207] = 32'b11111111111111111101010101100110;
assign LUT_4[57208] = 32'b00000000000000000000111011000011;
assign LUT_4[57209] = 32'b11111111111111111010000110111011;
assign LUT_4[57210] = 32'b00000000000000000000010101100111;
assign LUT_4[57211] = 32'b11111111111111111001100001011111;
assign LUT_4[57212] = 32'b11111111111111111101111011011111;
assign LUT_4[57213] = 32'b11111111111111110111000111010111;
assign LUT_4[57214] = 32'b11111111111111111101010110000011;
assign LUT_4[57215] = 32'b11111111111111110110100001111011;
assign LUT_4[57216] = 32'b00000000000000001100110000101101;
assign LUT_4[57217] = 32'b00000000000000000101111100100101;
assign LUT_4[57218] = 32'b00000000000000001100001011010001;
assign LUT_4[57219] = 32'b00000000000000000101010111001001;
assign LUT_4[57220] = 32'b00000000000000001001110001001001;
assign LUT_4[57221] = 32'b00000000000000000010111101000001;
assign LUT_4[57222] = 32'b00000000000000001001001011101101;
assign LUT_4[57223] = 32'b00000000000000000010010111100101;
assign LUT_4[57224] = 32'b00000000000000000101111101000010;
assign LUT_4[57225] = 32'b11111111111111111111001000111010;
assign LUT_4[57226] = 32'b00000000000000000101010111100110;
assign LUT_4[57227] = 32'b11111111111111111110100011011110;
assign LUT_4[57228] = 32'b00000000000000000010111101011110;
assign LUT_4[57229] = 32'b11111111111111111100001001010110;
assign LUT_4[57230] = 32'b00000000000000000010011000000010;
assign LUT_4[57231] = 32'b11111111111111111011100011111010;
assign LUT_4[57232] = 32'b00000000000000001010100010011011;
assign LUT_4[57233] = 32'b00000000000000000011101110010011;
assign LUT_4[57234] = 32'b00000000000000001001111100111111;
assign LUT_4[57235] = 32'b00000000000000000011001000110111;
assign LUT_4[57236] = 32'b00000000000000000111100010110111;
assign LUT_4[57237] = 32'b00000000000000000000101110101111;
assign LUT_4[57238] = 32'b00000000000000000110111101011011;
assign LUT_4[57239] = 32'b00000000000000000000001001010011;
assign LUT_4[57240] = 32'b00000000000000000011101110110000;
assign LUT_4[57241] = 32'b11111111111111111100111010101000;
assign LUT_4[57242] = 32'b00000000000000000011001001010100;
assign LUT_4[57243] = 32'b11111111111111111100010101001100;
assign LUT_4[57244] = 32'b00000000000000000000101111001100;
assign LUT_4[57245] = 32'b11111111111111111001111011000100;
assign LUT_4[57246] = 32'b00000000000000000000001001110000;
assign LUT_4[57247] = 32'b11111111111111111001010101101000;
assign LUT_4[57248] = 32'b00000000000000001011001011110100;
assign LUT_4[57249] = 32'b00000000000000000100010111101100;
assign LUT_4[57250] = 32'b00000000000000001010100110011000;
assign LUT_4[57251] = 32'b00000000000000000011110010010000;
assign LUT_4[57252] = 32'b00000000000000001000001100010000;
assign LUT_4[57253] = 32'b00000000000000000001011000001000;
assign LUT_4[57254] = 32'b00000000000000000111100110110100;
assign LUT_4[57255] = 32'b00000000000000000000110010101100;
assign LUT_4[57256] = 32'b00000000000000000100011000001001;
assign LUT_4[57257] = 32'b11111111111111111101100100000001;
assign LUT_4[57258] = 32'b00000000000000000011110010101101;
assign LUT_4[57259] = 32'b11111111111111111100111110100101;
assign LUT_4[57260] = 32'b00000000000000000001011000100101;
assign LUT_4[57261] = 32'b11111111111111111010100100011101;
assign LUT_4[57262] = 32'b00000000000000000000110011001001;
assign LUT_4[57263] = 32'b11111111111111111001111111000001;
assign LUT_4[57264] = 32'b00000000000000001000111101100010;
assign LUT_4[57265] = 32'b00000000000000000010001001011010;
assign LUT_4[57266] = 32'b00000000000000001000011000000110;
assign LUT_4[57267] = 32'b00000000000000000001100011111110;
assign LUT_4[57268] = 32'b00000000000000000101111101111110;
assign LUT_4[57269] = 32'b11111111111111111111001001110110;
assign LUT_4[57270] = 32'b00000000000000000101011000100010;
assign LUT_4[57271] = 32'b11111111111111111110100100011010;
assign LUT_4[57272] = 32'b00000000000000000010001001110111;
assign LUT_4[57273] = 32'b11111111111111111011010101101111;
assign LUT_4[57274] = 32'b00000000000000000001100100011011;
assign LUT_4[57275] = 32'b11111111111111111010110000010011;
assign LUT_4[57276] = 32'b11111111111111111111001010010011;
assign LUT_4[57277] = 32'b11111111111111111000010110001011;
assign LUT_4[57278] = 32'b11111111111111111110100100110111;
assign LUT_4[57279] = 32'b11111111111111110111110000101111;
assign LUT_4[57280] = 32'b00000000000000001110001000000001;
assign LUT_4[57281] = 32'b00000000000000000111010011111001;
assign LUT_4[57282] = 32'b00000000000000001101100010100101;
assign LUT_4[57283] = 32'b00000000000000000110101110011101;
assign LUT_4[57284] = 32'b00000000000000001011001000011101;
assign LUT_4[57285] = 32'b00000000000000000100010100010101;
assign LUT_4[57286] = 32'b00000000000000001010100011000001;
assign LUT_4[57287] = 32'b00000000000000000011101110111001;
assign LUT_4[57288] = 32'b00000000000000000111010100010110;
assign LUT_4[57289] = 32'b00000000000000000000100000001110;
assign LUT_4[57290] = 32'b00000000000000000110101110111010;
assign LUT_4[57291] = 32'b11111111111111111111111010110010;
assign LUT_4[57292] = 32'b00000000000000000100010100110010;
assign LUT_4[57293] = 32'b11111111111111111101100000101010;
assign LUT_4[57294] = 32'b00000000000000000011101111010110;
assign LUT_4[57295] = 32'b11111111111111111100111011001110;
assign LUT_4[57296] = 32'b00000000000000001011111001101111;
assign LUT_4[57297] = 32'b00000000000000000101000101100111;
assign LUT_4[57298] = 32'b00000000000000001011010100010011;
assign LUT_4[57299] = 32'b00000000000000000100100000001011;
assign LUT_4[57300] = 32'b00000000000000001000111010001011;
assign LUT_4[57301] = 32'b00000000000000000010000110000011;
assign LUT_4[57302] = 32'b00000000000000001000010100101111;
assign LUT_4[57303] = 32'b00000000000000000001100000100111;
assign LUT_4[57304] = 32'b00000000000000000101000110000100;
assign LUT_4[57305] = 32'b11111111111111111110010001111100;
assign LUT_4[57306] = 32'b00000000000000000100100000101000;
assign LUT_4[57307] = 32'b11111111111111111101101100100000;
assign LUT_4[57308] = 32'b00000000000000000010000110100000;
assign LUT_4[57309] = 32'b11111111111111111011010010011000;
assign LUT_4[57310] = 32'b00000000000000000001100001000100;
assign LUT_4[57311] = 32'b11111111111111111010101100111100;
assign LUT_4[57312] = 32'b00000000000000001100100011001000;
assign LUT_4[57313] = 32'b00000000000000000101101111000000;
assign LUT_4[57314] = 32'b00000000000000001011111101101100;
assign LUT_4[57315] = 32'b00000000000000000101001001100100;
assign LUT_4[57316] = 32'b00000000000000001001100011100100;
assign LUT_4[57317] = 32'b00000000000000000010101111011100;
assign LUT_4[57318] = 32'b00000000000000001000111110001000;
assign LUT_4[57319] = 32'b00000000000000000010001010000000;
assign LUT_4[57320] = 32'b00000000000000000101101111011101;
assign LUT_4[57321] = 32'b11111111111111111110111011010101;
assign LUT_4[57322] = 32'b00000000000000000101001010000001;
assign LUT_4[57323] = 32'b11111111111111111110010101111001;
assign LUT_4[57324] = 32'b00000000000000000010101111111001;
assign LUT_4[57325] = 32'b11111111111111111011111011110001;
assign LUT_4[57326] = 32'b00000000000000000010001010011101;
assign LUT_4[57327] = 32'b11111111111111111011010110010101;
assign LUT_4[57328] = 32'b00000000000000001010010100110110;
assign LUT_4[57329] = 32'b00000000000000000011100000101110;
assign LUT_4[57330] = 32'b00000000000000001001101111011010;
assign LUT_4[57331] = 32'b00000000000000000010111011010010;
assign LUT_4[57332] = 32'b00000000000000000111010101010010;
assign LUT_4[57333] = 32'b00000000000000000000100001001010;
assign LUT_4[57334] = 32'b00000000000000000110101111110110;
assign LUT_4[57335] = 32'b11111111111111111111111011101110;
assign LUT_4[57336] = 32'b00000000000000000011100001001011;
assign LUT_4[57337] = 32'b11111111111111111100101101000011;
assign LUT_4[57338] = 32'b00000000000000000010111011101111;
assign LUT_4[57339] = 32'b11111111111111111100000111100111;
assign LUT_4[57340] = 32'b00000000000000000000100001100111;
assign LUT_4[57341] = 32'b11111111111111111001101101011111;
assign LUT_4[57342] = 32'b11111111111111111111111100001011;
assign LUT_4[57343] = 32'b11111111111111111001001000000011;
assign LUT_4[57344] = 32'b00000000000000010011000000101100;
assign LUT_4[57345] = 32'b00000000000000001100001100100100;
assign LUT_4[57346] = 32'b00000000000000010010011011010000;
assign LUT_4[57347] = 32'b00000000000000001011100111001000;
assign LUT_4[57348] = 32'b00000000000000010000000001001000;
assign LUT_4[57349] = 32'b00000000000000001001001101000000;
assign LUT_4[57350] = 32'b00000000000000001111011011101100;
assign LUT_4[57351] = 32'b00000000000000001000100111100100;
assign LUT_4[57352] = 32'b00000000000000001100001101000001;
assign LUT_4[57353] = 32'b00000000000000000101011000111001;
assign LUT_4[57354] = 32'b00000000000000001011100111100101;
assign LUT_4[57355] = 32'b00000000000000000100110011011101;
assign LUT_4[57356] = 32'b00000000000000001001001101011101;
assign LUT_4[57357] = 32'b00000000000000000010011001010101;
assign LUT_4[57358] = 32'b00000000000000001000101000000001;
assign LUT_4[57359] = 32'b00000000000000000001110011111001;
assign LUT_4[57360] = 32'b00000000000000010000110010011010;
assign LUT_4[57361] = 32'b00000000000000001001111110010010;
assign LUT_4[57362] = 32'b00000000000000010000001100111110;
assign LUT_4[57363] = 32'b00000000000000001001011000110110;
assign LUT_4[57364] = 32'b00000000000000001101110010110110;
assign LUT_4[57365] = 32'b00000000000000000110111110101110;
assign LUT_4[57366] = 32'b00000000000000001101001101011010;
assign LUT_4[57367] = 32'b00000000000000000110011001010010;
assign LUT_4[57368] = 32'b00000000000000001001111110101111;
assign LUT_4[57369] = 32'b00000000000000000011001010100111;
assign LUT_4[57370] = 32'b00000000000000001001011001010011;
assign LUT_4[57371] = 32'b00000000000000000010100101001011;
assign LUT_4[57372] = 32'b00000000000000000110111111001011;
assign LUT_4[57373] = 32'b00000000000000000000001011000011;
assign LUT_4[57374] = 32'b00000000000000000110011001101111;
assign LUT_4[57375] = 32'b11111111111111111111100101100111;
assign LUT_4[57376] = 32'b00000000000000010001011011110011;
assign LUT_4[57377] = 32'b00000000000000001010100111101011;
assign LUT_4[57378] = 32'b00000000000000010000110110010111;
assign LUT_4[57379] = 32'b00000000000000001010000010001111;
assign LUT_4[57380] = 32'b00000000000000001110011100001111;
assign LUT_4[57381] = 32'b00000000000000000111101000000111;
assign LUT_4[57382] = 32'b00000000000000001101110110110011;
assign LUT_4[57383] = 32'b00000000000000000111000010101011;
assign LUT_4[57384] = 32'b00000000000000001010101000001000;
assign LUT_4[57385] = 32'b00000000000000000011110100000000;
assign LUT_4[57386] = 32'b00000000000000001010000010101100;
assign LUT_4[57387] = 32'b00000000000000000011001110100100;
assign LUT_4[57388] = 32'b00000000000000000111101000100100;
assign LUT_4[57389] = 32'b00000000000000000000110100011100;
assign LUT_4[57390] = 32'b00000000000000000111000011001000;
assign LUT_4[57391] = 32'b00000000000000000000001111000000;
assign LUT_4[57392] = 32'b00000000000000001111001101100001;
assign LUT_4[57393] = 32'b00000000000000001000011001011001;
assign LUT_4[57394] = 32'b00000000000000001110101000000101;
assign LUT_4[57395] = 32'b00000000000000000111110011111101;
assign LUT_4[57396] = 32'b00000000000000001100001101111101;
assign LUT_4[57397] = 32'b00000000000000000101011001110101;
assign LUT_4[57398] = 32'b00000000000000001011101000100001;
assign LUT_4[57399] = 32'b00000000000000000100110100011001;
assign LUT_4[57400] = 32'b00000000000000001000011001110110;
assign LUT_4[57401] = 32'b00000000000000000001100101101110;
assign LUT_4[57402] = 32'b00000000000000000111110100011010;
assign LUT_4[57403] = 32'b00000000000000000001000000010010;
assign LUT_4[57404] = 32'b00000000000000000101011010010010;
assign LUT_4[57405] = 32'b11111111111111111110100110001010;
assign LUT_4[57406] = 32'b00000000000000000100110100110110;
assign LUT_4[57407] = 32'b11111111111111111110000000101110;
assign LUT_4[57408] = 32'b00000000000000010100011000000000;
assign LUT_4[57409] = 32'b00000000000000001101100011111000;
assign LUT_4[57410] = 32'b00000000000000010011110010100100;
assign LUT_4[57411] = 32'b00000000000000001100111110011100;
assign LUT_4[57412] = 32'b00000000000000010001011000011100;
assign LUT_4[57413] = 32'b00000000000000001010100100010100;
assign LUT_4[57414] = 32'b00000000000000010000110011000000;
assign LUT_4[57415] = 32'b00000000000000001001111110111000;
assign LUT_4[57416] = 32'b00000000000000001101100100010101;
assign LUT_4[57417] = 32'b00000000000000000110110000001101;
assign LUT_4[57418] = 32'b00000000000000001100111110111001;
assign LUT_4[57419] = 32'b00000000000000000110001010110001;
assign LUT_4[57420] = 32'b00000000000000001010100100110001;
assign LUT_4[57421] = 32'b00000000000000000011110000101001;
assign LUT_4[57422] = 32'b00000000000000001001111111010101;
assign LUT_4[57423] = 32'b00000000000000000011001011001101;
assign LUT_4[57424] = 32'b00000000000000010010001001101110;
assign LUT_4[57425] = 32'b00000000000000001011010101100110;
assign LUT_4[57426] = 32'b00000000000000010001100100010010;
assign LUT_4[57427] = 32'b00000000000000001010110000001010;
assign LUT_4[57428] = 32'b00000000000000001111001010001010;
assign LUT_4[57429] = 32'b00000000000000001000010110000010;
assign LUT_4[57430] = 32'b00000000000000001110100100101110;
assign LUT_4[57431] = 32'b00000000000000000111110000100110;
assign LUT_4[57432] = 32'b00000000000000001011010110000011;
assign LUT_4[57433] = 32'b00000000000000000100100001111011;
assign LUT_4[57434] = 32'b00000000000000001010110000100111;
assign LUT_4[57435] = 32'b00000000000000000011111100011111;
assign LUT_4[57436] = 32'b00000000000000001000010110011111;
assign LUT_4[57437] = 32'b00000000000000000001100010010111;
assign LUT_4[57438] = 32'b00000000000000000111110001000011;
assign LUT_4[57439] = 32'b00000000000000000000111100111011;
assign LUT_4[57440] = 32'b00000000000000010010110011000111;
assign LUT_4[57441] = 32'b00000000000000001011111110111111;
assign LUT_4[57442] = 32'b00000000000000010010001101101011;
assign LUT_4[57443] = 32'b00000000000000001011011001100011;
assign LUT_4[57444] = 32'b00000000000000001111110011100011;
assign LUT_4[57445] = 32'b00000000000000001000111111011011;
assign LUT_4[57446] = 32'b00000000000000001111001110000111;
assign LUT_4[57447] = 32'b00000000000000001000011001111111;
assign LUT_4[57448] = 32'b00000000000000001011111111011100;
assign LUT_4[57449] = 32'b00000000000000000101001011010100;
assign LUT_4[57450] = 32'b00000000000000001011011010000000;
assign LUT_4[57451] = 32'b00000000000000000100100101111000;
assign LUT_4[57452] = 32'b00000000000000001000111111111000;
assign LUT_4[57453] = 32'b00000000000000000010001011110000;
assign LUT_4[57454] = 32'b00000000000000001000011010011100;
assign LUT_4[57455] = 32'b00000000000000000001100110010100;
assign LUT_4[57456] = 32'b00000000000000010000100100110101;
assign LUT_4[57457] = 32'b00000000000000001001110000101101;
assign LUT_4[57458] = 32'b00000000000000001111111111011001;
assign LUT_4[57459] = 32'b00000000000000001001001011010001;
assign LUT_4[57460] = 32'b00000000000000001101100101010001;
assign LUT_4[57461] = 32'b00000000000000000110110001001001;
assign LUT_4[57462] = 32'b00000000000000001100111111110101;
assign LUT_4[57463] = 32'b00000000000000000110001011101101;
assign LUT_4[57464] = 32'b00000000000000001001110001001010;
assign LUT_4[57465] = 32'b00000000000000000010111101000010;
assign LUT_4[57466] = 32'b00000000000000001001001011101110;
assign LUT_4[57467] = 32'b00000000000000000010010111100110;
assign LUT_4[57468] = 32'b00000000000000000110110001100110;
assign LUT_4[57469] = 32'b11111111111111111111111101011110;
assign LUT_4[57470] = 32'b00000000000000000110001100001010;
assign LUT_4[57471] = 32'b11111111111111111111011000000010;
assign LUT_4[57472] = 32'b00000000000000010101100110110100;
assign LUT_4[57473] = 32'b00000000000000001110110010101100;
assign LUT_4[57474] = 32'b00000000000000010101000001011000;
assign LUT_4[57475] = 32'b00000000000000001110001101010000;
assign LUT_4[57476] = 32'b00000000000000010010100111010000;
assign LUT_4[57477] = 32'b00000000000000001011110011001000;
assign LUT_4[57478] = 32'b00000000000000010010000001110100;
assign LUT_4[57479] = 32'b00000000000000001011001101101100;
assign LUT_4[57480] = 32'b00000000000000001110110011001001;
assign LUT_4[57481] = 32'b00000000000000000111111111000001;
assign LUT_4[57482] = 32'b00000000000000001110001101101101;
assign LUT_4[57483] = 32'b00000000000000000111011001100101;
assign LUT_4[57484] = 32'b00000000000000001011110011100101;
assign LUT_4[57485] = 32'b00000000000000000100111111011101;
assign LUT_4[57486] = 32'b00000000000000001011001110001001;
assign LUT_4[57487] = 32'b00000000000000000100011010000001;
assign LUT_4[57488] = 32'b00000000000000010011011000100010;
assign LUT_4[57489] = 32'b00000000000000001100100100011010;
assign LUT_4[57490] = 32'b00000000000000010010110011000110;
assign LUT_4[57491] = 32'b00000000000000001011111110111110;
assign LUT_4[57492] = 32'b00000000000000010000011000111110;
assign LUT_4[57493] = 32'b00000000000000001001100100110110;
assign LUT_4[57494] = 32'b00000000000000001111110011100010;
assign LUT_4[57495] = 32'b00000000000000001000111111011010;
assign LUT_4[57496] = 32'b00000000000000001100100100110111;
assign LUT_4[57497] = 32'b00000000000000000101110000101111;
assign LUT_4[57498] = 32'b00000000000000001011111111011011;
assign LUT_4[57499] = 32'b00000000000000000101001011010011;
assign LUT_4[57500] = 32'b00000000000000001001100101010011;
assign LUT_4[57501] = 32'b00000000000000000010110001001011;
assign LUT_4[57502] = 32'b00000000000000001000111111110111;
assign LUT_4[57503] = 32'b00000000000000000010001011101111;
assign LUT_4[57504] = 32'b00000000000000010100000001111011;
assign LUT_4[57505] = 32'b00000000000000001101001101110011;
assign LUT_4[57506] = 32'b00000000000000010011011100011111;
assign LUT_4[57507] = 32'b00000000000000001100101000010111;
assign LUT_4[57508] = 32'b00000000000000010001000010010111;
assign LUT_4[57509] = 32'b00000000000000001010001110001111;
assign LUT_4[57510] = 32'b00000000000000010000011100111011;
assign LUT_4[57511] = 32'b00000000000000001001101000110011;
assign LUT_4[57512] = 32'b00000000000000001101001110010000;
assign LUT_4[57513] = 32'b00000000000000000110011010001000;
assign LUT_4[57514] = 32'b00000000000000001100101000110100;
assign LUT_4[57515] = 32'b00000000000000000101110100101100;
assign LUT_4[57516] = 32'b00000000000000001010001110101100;
assign LUT_4[57517] = 32'b00000000000000000011011010100100;
assign LUT_4[57518] = 32'b00000000000000001001101001010000;
assign LUT_4[57519] = 32'b00000000000000000010110101001000;
assign LUT_4[57520] = 32'b00000000000000010001110011101001;
assign LUT_4[57521] = 32'b00000000000000001010111111100001;
assign LUT_4[57522] = 32'b00000000000000010001001110001101;
assign LUT_4[57523] = 32'b00000000000000001010011010000101;
assign LUT_4[57524] = 32'b00000000000000001110110100000101;
assign LUT_4[57525] = 32'b00000000000000000111111111111101;
assign LUT_4[57526] = 32'b00000000000000001110001110101001;
assign LUT_4[57527] = 32'b00000000000000000111011010100001;
assign LUT_4[57528] = 32'b00000000000000001010111111111110;
assign LUT_4[57529] = 32'b00000000000000000100001011110110;
assign LUT_4[57530] = 32'b00000000000000001010011010100010;
assign LUT_4[57531] = 32'b00000000000000000011100110011010;
assign LUT_4[57532] = 32'b00000000000000001000000000011010;
assign LUT_4[57533] = 32'b00000000000000000001001100010010;
assign LUT_4[57534] = 32'b00000000000000000111011010111110;
assign LUT_4[57535] = 32'b00000000000000000000100110110110;
assign LUT_4[57536] = 32'b00000000000000010110111110001000;
assign LUT_4[57537] = 32'b00000000000000010000001010000000;
assign LUT_4[57538] = 32'b00000000000000010110011000101100;
assign LUT_4[57539] = 32'b00000000000000001111100100100100;
assign LUT_4[57540] = 32'b00000000000000010011111110100100;
assign LUT_4[57541] = 32'b00000000000000001101001010011100;
assign LUT_4[57542] = 32'b00000000000000010011011001001000;
assign LUT_4[57543] = 32'b00000000000000001100100101000000;
assign LUT_4[57544] = 32'b00000000000000010000001010011101;
assign LUT_4[57545] = 32'b00000000000000001001010110010101;
assign LUT_4[57546] = 32'b00000000000000001111100101000001;
assign LUT_4[57547] = 32'b00000000000000001000110000111001;
assign LUT_4[57548] = 32'b00000000000000001101001010111001;
assign LUT_4[57549] = 32'b00000000000000000110010110110001;
assign LUT_4[57550] = 32'b00000000000000001100100101011101;
assign LUT_4[57551] = 32'b00000000000000000101110001010101;
assign LUT_4[57552] = 32'b00000000000000010100101111110110;
assign LUT_4[57553] = 32'b00000000000000001101111011101110;
assign LUT_4[57554] = 32'b00000000000000010100001010011010;
assign LUT_4[57555] = 32'b00000000000000001101010110010010;
assign LUT_4[57556] = 32'b00000000000000010001110000010010;
assign LUT_4[57557] = 32'b00000000000000001010111100001010;
assign LUT_4[57558] = 32'b00000000000000010001001010110110;
assign LUT_4[57559] = 32'b00000000000000001010010110101110;
assign LUT_4[57560] = 32'b00000000000000001101111100001011;
assign LUT_4[57561] = 32'b00000000000000000111001000000011;
assign LUT_4[57562] = 32'b00000000000000001101010110101111;
assign LUT_4[57563] = 32'b00000000000000000110100010100111;
assign LUT_4[57564] = 32'b00000000000000001010111100100111;
assign LUT_4[57565] = 32'b00000000000000000100001000011111;
assign LUT_4[57566] = 32'b00000000000000001010010111001011;
assign LUT_4[57567] = 32'b00000000000000000011100011000011;
assign LUT_4[57568] = 32'b00000000000000010101011001001111;
assign LUT_4[57569] = 32'b00000000000000001110100101000111;
assign LUT_4[57570] = 32'b00000000000000010100110011110011;
assign LUT_4[57571] = 32'b00000000000000001101111111101011;
assign LUT_4[57572] = 32'b00000000000000010010011001101011;
assign LUT_4[57573] = 32'b00000000000000001011100101100011;
assign LUT_4[57574] = 32'b00000000000000010001110100001111;
assign LUT_4[57575] = 32'b00000000000000001011000000000111;
assign LUT_4[57576] = 32'b00000000000000001110100101100100;
assign LUT_4[57577] = 32'b00000000000000000111110001011100;
assign LUT_4[57578] = 32'b00000000000000001110000000001000;
assign LUT_4[57579] = 32'b00000000000000000111001100000000;
assign LUT_4[57580] = 32'b00000000000000001011100110000000;
assign LUT_4[57581] = 32'b00000000000000000100110001111000;
assign LUT_4[57582] = 32'b00000000000000001011000000100100;
assign LUT_4[57583] = 32'b00000000000000000100001100011100;
assign LUT_4[57584] = 32'b00000000000000010011001010111101;
assign LUT_4[57585] = 32'b00000000000000001100010110110101;
assign LUT_4[57586] = 32'b00000000000000010010100101100001;
assign LUT_4[57587] = 32'b00000000000000001011110001011001;
assign LUT_4[57588] = 32'b00000000000000010000001011011001;
assign LUT_4[57589] = 32'b00000000000000001001010111010001;
assign LUT_4[57590] = 32'b00000000000000001111100101111101;
assign LUT_4[57591] = 32'b00000000000000001000110001110101;
assign LUT_4[57592] = 32'b00000000000000001100010111010010;
assign LUT_4[57593] = 32'b00000000000000000101100011001010;
assign LUT_4[57594] = 32'b00000000000000001011110001110110;
assign LUT_4[57595] = 32'b00000000000000000100111101101110;
assign LUT_4[57596] = 32'b00000000000000001001010111101110;
assign LUT_4[57597] = 32'b00000000000000000010100011100110;
assign LUT_4[57598] = 32'b00000000000000001000110010010010;
assign LUT_4[57599] = 32'b00000000000000000001111110001010;
assign LUT_4[57600] = 32'b00000000000000010111111100001111;
assign LUT_4[57601] = 32'b00000000000000010001001000000111;
assign LUT_4[57602] = 32'b00000000000000010111010110110011;
assign LUT_4[57603] = 32'b00000000000000010000100010101011;
assign LUT_4[57604] = 32'b00000000000000010100111100101011;
assign LUT_4[57605] = 32'b00000000000000001110001000100011;
assign LUT_4[57606] = 32'b00000000000000010100010111001111;
assign LUT_4[57607] = 32'b00000000000000001101100011000111;
assign LUT_4[57608] = 32'b00000000000000010001001000100100;
assign LUT_4[57609] = 32'b00000000000000001010010100011100;
assign LUT_4[57610] = 32'b00000000000000010000100011001000;
assign LUT_4[57611] = 32'b00000000000000001001101111000000;
assign LUT_4[57612] = 32'b00000000000000001110001001000000;
assign LUT_4[57613] = 32'b00000000000000000111010100111000;
assign LUT_4[57614] = 32'b00000000000000001101100011100100;
assign LUT_4[57615] = 32'b00000000000000000110101111011100;
assign LUT_4[57616] = 32'b00000000000000010101101101111101;
assign LUT_4[57617] = 32'b00000000000000001110111001110101;
assign LUT_4[57618] = 32'b00000000000000010101001000100001;
assign LUT_4[57619] = 32'b00000000000000001110010100011001;
assign LUT_4[57620] = 32'b00000000000000010010101110011001;
assign LUT_4[57621] = 32'b00000000000000001011111010010001;
assign LUT_4[57622] = 32'b00000000000000010010001000111101;
assign LUT_4[57623] = 32'b00000000000000001011010100110101;
assign LUT_4[57624] = 32'b00000000000000001110111010010010;
assign LUT_4[57625] = 32'b00000000000000001000000110001010;
assign LUT_4[57626] = 32'b00000000000000001110010100110110;
assign LUT_4[57627] = 32'b00000000000000000111100000101110;
assign LUT_4[57628] = 32'b00000000000000001011111010101110;
assign LUT_4[57629] = 32'b00000000000000000101000110100110;
assign LUT_4[57630] = 32'b00000000000000001011010101010010;
assign LUT_4[57631] = 32'b00000000000000000100100001001010;
assign LUT_4[57632] = 32'b00000000000000010110010111010110;
assign LUT_4[57633] = 32'b00000000000000001111100011001110;
assign LUT_4[57634] = 32'b00000000000000010101110001111010;
assign LUT_4[57635] = 32'b00000000000000001110111101110010;
assign LUT_4[57636] = 32'b00000000000000010011010111110010;
assign LUT_4[57637] = 32'b00000000000000001100100011101010;
assign LUT_4[57638] = 32'b00000000000000010010110010010110;
assign LUT_4[57639] = 32'b00000000000000001011111110001110;
assign LUT_4[57640] = 32'b00000000000000001111100011101011;
assign LUT_4[57641] = 32'b00000000000000001000101111100011;
assign LUT_4[57642] = 32'b00000000000000001110111110001111;
assign LUT_4[57643] = 32'b00000000000000001000001010000111;
assign LUT_4[57644] = 32'b00000000000000001100100100000111;
assign LUT_4[57645] = 32'b00000000000000000101101111111111;
assign LUT_4[57646] = 32'b00000000000000001011111110101011;
assign LUT_4[57647] = 32'b00000000000000000101001010100011;
assign LUT_4[57648] = 32'b00000000000000010100001001000100;
assign LUT_4[57649] = 32'b00000000000000001101010100111100;
assign LUT_4[57650] = 32'b00000000000000010011100011101000;
assign LUT_4[57651] = 32'b00000000000000001100101111100000;
assign LUT_4[57652] = 32'b00000000000000010001001001100000;
assign LUT_4[57653] = 32'b00000000000000001010010101011000;
assign LUT_4[57654] = 32'b00000000000000010000100100000100;
assign LUT_4[57655] = 32'b00000000000000001001101111111100;
assign LUT_4[57656] = 32'b00000000000000001101010101011001;
assign LUT_4[57657] = 32'b00000000000000000110100001010001;
assign LUT_4[57658] = 32'b00000000000000001100101111111101;
assign LUT_4[57659] = 32'b00000000000000000101111011110101;
assign LUT_4[57660] = 32'b00000000000000001010010101110101;
assign LUT_4[57661] = 32'b00000000000000000011100001101101;
assign LUT_4[57662] = 32'b00000000000000001001110000011001;
assign LUT_4[57663] = 32'b00000000000000000010111100010001;
assign LUT_4[57664] = 32'b00000000000000011001010011100011;
assign LUT_4[57665] = 32'b00000000000000010010011111011011;
assign LUT_4[57666] = 32'b00000000000000011000101110000111;
assign LUT_4[57667] = 32'b00000000000000010001111001111111;
assign LUT_4[57668] = 32'b00000000000000010110010011111111;
assign LUT_4[57669] = 32'b00000000000000001111011111110111;
assign LUT_4[57670] = 32'b00000000000000010101101110100011;
assign LUT_4[57671] = 32'b00000000000000001110111010011011;
assign LUT_4[57672] = 32'b00000000000000010010011111111000;
assign LUT_4[57673] = 32'b00000000000000001011101011110000;
assign LUT_4[57674] = 32'b00000000000000010001111010011100;
assign LUT_4[57675] = 32'b00000000000000001011000110010100;
assign LUT_4[57676] = 32'b00000000000000001111100000010100;
assign LUT_4[57677] = 32'b00000000000000001000101100001100;
assign LUT_4[57678] = 32'b00000000000000001110111010111000;
assign LUT_4[57679] = 32'b00000000000000001000000110110000;
assign LUT_4[57680] = 32'b00000000000000010111000101010001;
assign LUT_4[57681] = 32'b00000000000000010000010001001001;
assign LUT_4[57682] = 32'b00000000000000010110011111110101;
assign LUT_4[57683] = 32'b00000000000000001111101011101101;
assign LUT_4[57684] = 32'b00000000000000010100000101101101;
assign LUT_4[57685] = 32'b00000000000000001101010001100101;
assign LUT_4[57686] = 32'b00000000000000010011100000010001;
assign LUT_4[57687] = 32'b00000000000000001100101100001001;
assign LUT_4[57688] = 32'b00000000000000010000010001100110;
assign LUT_4[57689] = 32'b00000000000000001001011101011110;
assign LUT_4[57690] = 32'b00000000000000001111101100001010;
assign LUT_4[57691] = 32'b00000000000000001000111000000010;
assign LUT_4[57692] = 32'b00000000000000001101010010000010;
assign LUT_4[57693] = 32'b00000000000000000110011101111010;
assign LUT_4[57694] = 32'b00000000000000001100101100100110;
assign LUT_4[57695] = 32'b00000000000000000101111000011110;
assign LUT_4[57696] = 32'b00000000000000010111101110101010;
assign LUT_4[57697] = 32'b00000000000000010000111010100010;
assign LUT_4[57698] = 32'b00000000000000010111001001001110;
assign LUT_4[57699] = 32'b00000000000000010000010101000110;
assign LUT_4[57700] = 32'b00000000000000010100101111000110;
assign LUT_4[57701] = 32'b00000000000000001101111010111110;
assign LUT_4[57702] = 32'b00000000000000010100001001101010;
assign LUT_4[57703] = 32'b00000000000000001101010101100010;
assign LUT_4[57704] = 32'b00000000000000010000111010111111;
assign LUT_4[57705] = 32'b00000000000000001010000110110111;
assign LUT_4[57706] = 32'b00000000000000010000010101100011;
assign LUT_4[57707] = 32'b00000000000000001001100001011011;
assign LUT_4[57708] = 32'b00000000000000001101111011011011;
assign LUT_4[57709] = 32'b00000000000000000111000111010011;
assign LUT_4[57710] = 32'b00000000000000001101010101111111;
assign LUT_4[57711] = 32'b00000000000000000110100001110111;
assign LUT_4[57712] = 32'b00000000000000010101100000011000;
assign LUT_4[57713] = 32'b00000000000000001110101100010000;
assign LUT_4[57714] = 32'b00000000000000010100111010111100;
assign LUT_4[57715] = 32'b00000000000000001110000110110100;
assign LUT_4[57716] = 32'b00000000000000010010100000110100;
assign LUT_4[57717] = 32'b00000000000000001011101100101100;
assign LUT_4[57718] = 32'b00000000000000010001111011011000;
assign LUT_4[57719] = 32'b00000000000000001011000111010000;
assign LUT_4[57720] = 32'b00000000000000001110101100101101;
assign LUT_4[57721] = 32'b00000000000000000111111000100101;
assign LUT_4[57722] = 32'b00000000000000001110000111010001;
assign LUT_4[57723] = 32'b00000000000000000111010011001001;
assign LUT_4[57724] = 32'b00000000000000001011101101001001;
assign LUT_4[57725] = 32'b00000000000000000100111001000001;
assign LUT_4[57726] = 32'b00000000000000001011000111101101;
assign LUT_4[57727] = 32'b00000000000000000100010011100101;
assign LUT_4[57728] = 32'b00000000000000011010100010010111;
assign LUT_4[57729] = 32'b00000000000000010011101110001111;
assign LUT_4[57730] = 32'b00000000000000011001111100111011;
assign LUT_4[57731] = 32'b00000000000000010011001000110011;
assign LUT_4[57732] = 32'b00000000000000010111100010110011;
assign LUT_4[57733] = 32'b00000000000000010000101110101011;
assign LUT_4[57734] = 32'b00000000000000010110111101010111;
assign LUT_4[57735] = 32'b00000000000000010000001001001111;
assign LUT_4[57736] = 32'b00000000000000010011101110101100;
assign LUT_4[57737] = 32'b00000000000000001100111010100100;
assign LUT_4[57738] = 32'b00000000000000010011001001010000;
assign LUT_4[57739] = 32'b00000000000000001100010101001000;
assign LUT_4[57740] = 32'b00000000000000010000101111001000;
assign LUT_4[57741] = 32'b00000000000000001001111011000000;
assign LUT_4[57742] = 32'b00000000000000010000001001101100;
assign LUT_4[57743] = 32'b00000000000000001001010101100100;
assign LUT_4[57744] = 32'b00000000000000011000010100000101;
assign LUT_4[57745] = 32'b00000000000000010001011111111101;
assign LUT_4[57746] = 32'b00000000000000010111101110101001;
assign LUT_4[57747] = 32'b00000000000000010000111010100001;
assign LUT_4[57748] = 32'b00000000000000010101010100100001;
assign LUT_4[57749] = 32'b00000000000000001110100000011001;
assign LUT_4[57750] = 32'b00000000000000010100101111000101;
assign LUT_4[57751] = 32'b00000000000000001101111010111101;
assign LUT_4[57752] = 32'b00000000000000010001100000011010;
assign LUT_4[57753] = 32'b00000000000000001010101100010010;
assign LUT_4[57754] = 32'b00000000000000010000111010111110;
assign LUT_4[57755] = 32'b00000000000000001010000110110110;
assign LUT_4[57756] = 32'b00000000000000001110100000110110;
assign LUT_4[57757] = 32'b00000000000000000111101100101110;
assign LUT_4[57758] = 32'b00000000000000001101111011011010;
assign LUT_4[57759] = 32'b00000000000000000111000111010010;
assign LUT_4[57760] = 32'b00000000000000011000111101011110;
assign LUT_4[57761] = 32'b00000000000000010010001001010110;
assign LUT_4[57762] = 32'b00000000000000011000011000000010;
assign LUT_4[57763] = 32'b00000000000000010001100011111010;
assign LUT_4[57764] = 32'b00000000000000010101111101111010;
assign LUT_4[57765] = 32'b00000000000000001111001001110010;
assign LUT_4[57766] = 32'b00000000000000010101011000011110;
assign LUT_4[57767] = 32'b00000000000000001110100100010110;
assign LUT_4[57768] = 32'b00000000000000010010001001110011;
assign LUT_4[57769] = 32'b00000000000000001011010101101011;
assign LUT_4[57770] = 32'b00000000000000010001100100010111;
assign LUT_4[57771] = 32'b00000000000000001010110000001111;
assign LUT_4[57772] = 32'b00000000000000001111001010001111;
assign LUT_4[57773] = 32'b00000000000000001000010110000111;
assign LUT_4[57774] = 32'b00000000000000001110100100110011;
assign LUT_4[57775] = 32'b00000000000000000111110000101011;
assign LUT_4[57776] = 32'b00000000000000010110101111001100;
assign LUT_4[57777] = 32'b00000000000000001111111011000100;
assign LUT_4[57778] = 32'b00000000000000010110001001110000;
assign LUT_4[57779] = 32'b00000000000000001111010101101000;
assign LUT_4[57780] = 32'b00000000000000010011101111101000;
assign LUT_4[57781] = 32'b00000000000000001100111011100000;
assign LUT_4[57782] = 32'b00000000000000010011001010001100;
assign LUT_4[57783] = 32'b00000000000000001100010110000100;
assign LUT_4[57784] = 32'b00000000000000001111111011100001;
assign LUT_4[57785] = 32'b00000000000000001001000111011001;
assign LUT_4[57786] = 32'b00000000000000001111010110000101;
assign LUT_4[57787] = 32'b00000000000000001000100001111101;
assign LUT_4[57788] = 32'b00000000000000001100111011111101;
assign LUT_4[57789] = 32'b00000000000000000110000111110101;
assign LUT_4[57790] = 32'b00000000000000001100010110100001;
assign LUT_4[57791] = 32'b00000000000000000101100010011001;
assign LUT_4[57792] = 32'b00000000000000011011111001101011;
assign LUT_4[57793] = 32'b00000000000000010101000101100011;
assign LUT_4[57794] = 32'b00000000000000011011010100001111;
assign LUT_4[57795] = 32'b00000000000000010100100000000111;
assign LUT_4[57796] = 32'b00000000000000011000111010000111;
assign LUT_4[57797] = 32'b00000000000000010010000101111111;
assign LUT_4[57798] = 32'b00000000000000011000010100101011;
assign LUT_4[57799] = 32'b00000000000000010001100000100011;
assign LUT_4[57800] = 32'b00000000000000010101000110000000;
assign LUT_4[57801] = 32'b00000000000000001110010001111000;
assign LUT_4[57802] = 32'b00000000000000010100100000100100;
assign LUT_4[57803] = 32'b00000000000000001101101100011100;
assign LUT_4[57804] = 32'b00000000000000010010000110011100;
assign LUT_4[57805] = 32'b00000000000000001011010010010100;
assign LUT_4[57806] = 32'b00000000000000010001100001000000;
assign LUT_4[57807] = 32'b00000000000000001010101100111000;
assign LUT_4[57808] = 32'b00000000000000011001101011011001;
assign LUT_4[57809] = 32'b00000000000000010010110111010001;
assign LUT_4[57810] = 32'b00000000000000011001000101111101;
assign LUT_4[57811] = 32'b00000000000000010010010001110101;
assign LUT_4[57812] = 32'b00000000000000010110101011110101;
assign LUT_4[57813] = 32'b00000000000000001111110111101101;
assign LUT_4[57814] = 32'b00000000000000010110000110011001;
assign LUT_4[57815] = 32'b00000000000000001111010010010001;
assign LUT_4[57816] = 32'b00000000000000010010110111101110;
assign LUT_4[57817] = 32'b00000000000000001100000011100110;
assign LUT_4[57818] = 32'b00000000000000010010010010010010;
assign LUT_4[57819] = 32'b00000000000000001011011110001010;
assign LUT_4[57820] = 32'b00000000000000001111111000001010;
assign LUT_4[57821] = 32'b00000000000000001001000100000010;
assign LUT_4[57822] = 32'b00000000000000001111010010101110;
assign LUT_4[57823] = 32'b00000000000000001000011110100110;
assign LUT_4[57824] = 32'b00000000000000011010010100110010;
assign LUT_4[57825] = 32'b00000000000000010011100000101010;
assign LUT_4[57826] = 32'b00000000000000011001101111010110;
assign LUT_4[57827] = 32'b00000000000000010010111011001110;
assign LUT_4[57828] = 32'b00000000000000010111010101001110;
assign LUT_4[57829] = 32'b00000000000000010000100001000110;
assign LUT_4[57830] = 32'b00000000000000010110101111110010;
assign LUT_4[57831] = 32'b00000000000000001111111011101010;
assign LUT_4[57832] = 32'b00000000000000010011100001000111;
assign LUT_4[57833] = 32'b00000000000000001100101100111111;
assign LUT_4[57834] = 32'b00000000000000010010111011101011;
assign LUT_4[57835] = 32'b00000000000000001100000111100011;
assign LUT_4[57836] = 32'b00000000000000010000100001100011;
assign LUT_4[57837] = 32'b00000000000000001001101101011011;
assign LUT_4[57838] = 32'b00000000000000001111111100000111;
assign LUT_4[57839] = 32'b00000000000000001001000111111111;
assign LUT_4[57840] = 32'b00000000000000011000000110100000;
assign LUT_4[57841] = 32'b00000000000000010001010010011000;
assign LUT_4[57842] = 32'b00000000000000010111100001000100;
assign LUT_4[57843] = 32'b00000000000000010000101100111100;
assign LUT_4[57844] = 32'b00000000000000010101000110111100;
assign LUT_4[57845] = 32'b00000000000000001110010010110100;
assign LUT_4[57846] = 32'b00000000000000010100100001100000;
assign LUT_4[57847] = 32'b00000000000000001101101101011000;
assign LUT_4[57848] = 32'b00000000000000010001010010110101;
assign LUT_4[57849] = 32'b00000000000000001010011110101101;
assign LUT_4[57850] = 32'b00000000000000010000101101011001;
assign LUT_4[57851] = 32'b00000000000000001001111001010001;
assign LUT_4[57852] = 32'b00000000000000001110010011010001;
assign LUT_4[57853] = 32'b00000000000000000111011111001001;
assign LUT_4[57854] = 32'b00000000000000001101101101110101;
assign LUT_4[57855] = 32'b00000000000000000110111001101101;
assign LUT_4[57856] = 32'b00000000000000010010000100110100;
assign LUT_4[57857] = 32'b00000000000000001011010000101100;
assign LUT_4[57858] = 32'b00000000000000010001011111011000;
assign LUT_4[57859] = 32'b00000000000000001010101011010000;
assign LUT_4[57860] = 32'b00000000000000001111000101010000;
assign LUT_4[57861] = 32'b00000000000000001000010001001000;
assign LUT_4[57862] = 32'b00000000000000001110011111110100;
assign LUT_4[57863] = 32'b00000000000000000111101011101100;
assign LUT_4[57864] = 32'b00000000000000001011010001001001;
assign LUT_4[57865] = 32'b00000000000000000100011101000001;
assign LUT_4[57866] = 32'b00000000000000001010101011101101;
assign LUT_4[57867] = 32'b00000000000000000011110111100101;
assign LUT_4[57868] = 32'b00000000000000001000010001100101;
assign LUT_4[57869] = 32'b00000000000000000001011101011101;
assign LUT_4[57870] = 32'b00000000000000000111101100001001;
assign LUT_4[57871] = 32'b00000000000000000000111000000001;
assign LUT_4[57872] = 32'b00000000000000001111110110100010;
assign LUT_4[57873] = 32'b00000000000000001001000010011010;
assign LUT_4[57874] = 32'b00000000000000001111010001000110;
assign LUT_4[57875] = 32'b00000000000000001000011100111110;
assign LUT_4[57876] = 32'b00000000000000001100110110111110;
assign LUT_4[57877] = 32'b00000000000000000110000010110110;
assign LUT_4[57878] = 32'b00000000000000001100010001100010;
assign LUT_4[57879] = 32'b00000000000000000101011101011010;
assign LUT_4[57880] = 32'b00000000000000001001000010110111;
assign LUT_4[57881] = 32'b00000000000000000010001110101111;
assign LUT_4[57882] = 32'b00000000000000001000011101011011;
assign LUT_4[57883] = 32'b00000000000000000001101001010011;
assign LUT_4[57884] = 32'b00000000000000000110000011010011;
assign LUT_4[57885] = 32'b11111111111111111111001111001011;
assign LUT_4[57886] = 32'b00000000000000000101011101110111;
assign LUT_4[57887] = 32'b11111111111111111110101001101111;
assign LUT_4[57888] = 32'b00000000000000010000011111111011;
assign LUT_4[57889] = 32'b00000000000000001001101011110011;
assign LUT_4[57890] = 32'b00000000000000001111111010011111;
assign LUT_4[57891] = 32'b00000000000000001001000110010111;
assign LUT_4[57892] = 32'b00000000000000001101100000010111;
assign LUT_4[57893] = 32'b00000000000000000110101100001111;
assign LUT_4[57894] = 32'b00000000000000001100111010111011;
assign LUT_4[57895] = 32'b00000000000000000110000110110011;
assign LUT_4[57896] = 32'b00000000000000001001101100010000;
assign LUT_4[57897] = 32'b00000000000000000010111000001000;
assign LUT_4[57898] = 32'b00000000000000001001000110110100;
assign LUT_4[57899] = 32'b00000000000000000010010010101100;
assign LUT_4[57900] = 32'b00000000000000000110101100101100;
assign LUT_4[57901] = 32'b11111111111111111111111000100100;
assign LUT_4[57902] = 32'b00000000000000000110000111010000;
assign LUT_4[57903] = 32'b11111111111111111111010011001000;
assign LUT_4[57904] = 32'b00000000000000001110010001101001;
assign LUT_4[57905] = 32'b00000000000000000111011101100001;
assign LUT_4[57906] = 32'b00000000000000001101101100001101;
assign LUT_4[57907] = 32'b00000000000000000110111000000101;
assign LUT_4[57908] = 32'b00000000000000001011010010000101;
assign LUT_4[57909] = 32'b00000000000000000100011101111101;
assign LUT_4[57910] = 32'b00000000000000001010101100101001;
assign LUT_4[57911] = 32'b00000000000000000011111000100001;
assign LUT_4[57912] = 32'b00000000000000000111011101111110;
assign LUT_4[57913] = 32'b00000000000000000000101001110110;
assign LUT_4[57914] = 32'b00000000000000000110111000100010;
assign LUT_4[57915] = 32'b00000000000000000000000100011010;
assign LUT_4[57916] = 32'b00000000000000000100011110011010;
assign LUT_4[57917] = 32'b11111111111111111101101010010010;
assign LUT_4[57918] = 32'b00000000000000000011111000111110;
assign LUT_4[57919] = 32'b11111111111111111101000100110110;
assign LUT_4[57920] = 32'b00000000000000010011011100001000;
assign LUT_4[57921] = 32'b00000000000000001100101000000000;
assign LUT_4[57922] = 32'b00000000000000010010110110101100;
assign LUT_4[57923] = 32'b00000000000000001100000010100100;
assign LUT_4[57924] = 32'b00000000000000010000011100100100;
assign LUT_4[57925] = 32'b00000000000000001001101000011100;
assign LUT_4[57926] = 32'b00000000000000001111110111001000;
assign LUT_4[57927] = 32'b00000000000000001001000011000000;
assign LUT_4[57928] = 32'b00000000000000001100101000011101;
assign LUT_4[57929] = 32'b00000000000000000101110100010101;
assign LUT_4[57930] = 32'b00000000000000001100000011000001;
assign LUT_4[57931] = 32'b00000000000000000101001110111001;
assign LUT_4[57932] = 32'b00000000000000001001101000111001;
assign LUT_4[57933] = 32'b00000000000000000010110100110001;
assign LUT_4[57934] = 32'b00000000000000001001000011011101;
assign LUT_4[57935] = 32'b00000000000000000010001111010101;
assign LUT_4[57936] = 32'b00000000000000010001001101110110;
assign LUT_4[57937] = 32'b00000000000000001010011001101110;
assign LUT_4[57938] = 32'b00000000000000010000101000011010;
assign LUT_4[57939] = 32'b00000000000000001001110100010010;
assign LUT_4[57940] = 32'b00000000000000001110001110010010;
assign LUT_4[57941] = 32'b00000000000000000111011010001010;
assign LUT_4[57942] = 32'b00000000000000001101101000110110;
assign LUT_4[57943] = 32'b00000000000000000110110100101110;
assign LUT_4[57944] = 32'b00000000000000001010011010001011;
assign LUT_4[57945] = 32'b00000000000000000011100110000011;
assign LUT_4[57946] = 32'b00000000000000001001110100101111;
assign LUT_4[57947] = 32'b00000000000000000011000000100111;
assign LUT_4[57948] = 32'b00000000000000000111011010100111;
assign LUT_4[57949] = 32'b00000000000000000000100110011111;
assign LUT_4[57950] = 32'b00000000000000000110110101001011;
assign LUT_4[57951] = 32'b00000000000000000000000001000011;
assign LUT_4[57952] = 32'b00000000000000010001110111001111;
assign LUT_4[57953] = 32'b00000000000000001011000011000111;
assign LUT_4[57954] = 32'b00000000000000010001010001110011;
assign LUT_4[57955] = 32'b00000000000000001010011101101011;
assign LUT_4[57956] = 32'b00000000000000001110110111101011;
assign LUT_4[57957] = 32'b00000000000000001000000011100011;
assign LUT_4[57958] = 32'b00000000000000001110010010001111;
assign LUT_4[57959] = 32'b00000000000000000111011110000111;
assign LUT_4[57960] = 32'b00000000000000001011000011100100;
assign LUT_4[57961] = 32'b00000000000000000100001111011100;
assign LUT_4[57962] = 32'b00000000000000001010011110001000;
assign LUT_4[57963] = 32'b00000000000000000011101010000000;
assign LUT_4[57964] = 32'b00000000000000001000000100000000;
assign LUT_4[57965] = 32'b00000000000000000001001111111000;
assign LUT_4[57966] = 32'b00000000000000000111011110100100;
assign LUT_4[57967] = 32'b00000000000000000000101010011100;
assign LUT_4[57968] = 32'b00000000000000001111101000111101;
assign LUT_4[57969] = 32'b00000000000000001000110100110101;
assign LUT_4[57970] = 32'b00000000000000001111000011100001;
assign LUT_4[57971] = 32'b00000000000000001000001111011001;
assign LUT_4[57972] = 32'b00000000000000001100101001011001;
assign LUT_4[57973] = 32'b00000000000000000101110101010001;
assign LUT_4[57974] = 32'b00000000000000001100000011111101;
assign LUT_4[57975] = 32'b00000000000000000101001111110101;
assign LUT_4[57976] = 32'b00000000000000001000110101010010;
assign LUT_4[57977] = 32'b00000000000000000010000001001010;
assign LUT_4[57978] = 32'b00000000000000001000001111110110;
assign LUT_4[57979] = 32'b00000000000000000001011011101110;
assign LUT_4[57980] = 32'b00000000000000000101110101101110;
assign LUT_4[57981] = 32'b11111111111111111111000001100110;
assign LUT_4[57982] = 32'b00000000000000000101010000010010;
assign LUT_4[57983] = 32'b11111111111111111110011100001010;
assign LUT_4[57984] = 32'b00000000000000010100101010111100;
assign LUT_4[57985] = 32'b00000000000000001101110110110100;
assign LUT_4[57986] = 32'b00000000000000010100000101100000;
assign LUT_4[57987] = 32'b00000000000000001101010001011000;
assign LUT_4[57988] = 32'b00000000000000010001101011011000;
assign LUT_4[57989] = 32'b00000000000000001010110111010000;
assign LUT_4[57990] = 32'b00000000000000010001000101111100;
assign LUT_4[57991] = 32'b00000000000000001010010001110100;
assign LUT_4[57992] = 32'b00000000000000001101110111010001;
assign LUT_4[57993] = 32'b00000000000000000111000011001001;
assign LUT_4[57994] = 32'b00000000000000001101010001110101;
assign LUT_4[57995] = 32'b00000000000000000110011101101101;
assign LUT_4[57996] = 32'b00000000000000001010110111101101;
assign LUT_4[57997] = 32'b00000000000000000100000011100101;
assign LUT_4[57998] = 32'b00000000000000001010010010010001;
assign LUT_4[57999] = 32'b00000000000000000011011110001001;
assign LUT_4[58000] = 32'b00000000000000010010011100101010;
assign LUT_4[58001] = 32'b00000000000000001011101000100010;
assign LUT_4[58002] = 32'b00000000000000010001110111001110;
assign LUT_4[58003] = 32'b00000000000000001011000011000110;
assign LUT_4[58004] = 32'b00000000000000001111011101000110;
assign LUT_4[58005] = 32'b00000000000000001000101000111110;
assign LUT_4[58006] = 32'b00000000000000001110110111101010;
assign LUT_4[58007] = 32'b00000000000000001000000011100010;
assign LUT_4[58008] = 32'b00000000000000001011101000111111;
assign LUT_4[58009] = 32'b00000000000000000100110100110111;
assign LUT_4[58010] = 32'b00000000000000001011000011100011;
assign LUT_4[58011] = 32'b00000000000000000100001111011011;
assign LUT_4[58012] = 32'b00000000000000001000101001011011;
assign LUT_4[58013] = 32'b00000000000000000001110101010011;
assign LUT_4[58014] = 32'b00000000000000001000000011111111;
assign LUT_4[58015] = 32'b00000000000000000001001111110111;
assign LUT_4[58016] = 32'b00000000000000010011000110000011;
assign LUT_4[58017] = 32'b00000000000000001100010001111011;
assign LUT_4[58018] = 32'b00000000000000010010100000100111;
assign LUT_4[58019] = 32'b00000000000000001011101100011111;
assign LUT_4[58020] = 32'b00000000000000010000000110011111;
assign LUT_4[58021] = 32'b00000000000000001001010010010111;
assign LUT_4[58022] = 32'b00000000000000001111100001000011;
assign LUT_4[58023] = 32'b00000000000000001000101100111011;
assign LUT_4[58024] = 32'b00000000000000001100010010011000;
assign LUT_4[58025] = 32'b00000000000000000101011110010000;
assign LUT_4[58026] = 32'b00000000000000001011101100111100;
assign LUT_4[58027] = 32'b00000000000000000100111000110100;
assign LUT_4[58028] = 32'b00000000000000001001010010110100;
assign LUT_4[58029] = 32'b00000000000000000010011110101100;
assign LUT_4[58030] = 32'b00000000000000001000101101011000;
assign LUT_4[58031] = 32'b00000000000000000001111001010000;
assign LUT_4[58032] = 32'b00000000000000010000110111110001;
assign LUT_4[58033] = 32'b00000000000000001010000011101001;
assign LUT_4[58034] = 32'b00000000000000010000010010010101;
assign LUT_4[58035] = 32'b00000000000000001001011110001101;
assign LUT_4[58036] = 32'b00000000000000001101111000001101;
assign LUT_4[58037] = 32'b00000000000000000111000100000101;
assign LUT_4[58038] = 32'b00000000000000001101010010110001;
assign LUT_4[58039] = 32'b00000000000000000110011110101001;
assign LUT_4[58040] = 32'b00000000000000001010000100000110;
assign LUT_4[58041] = 32'b00000000000000000011001111111110;
assign LUT_4[58042] = 32'b00000000000000001001011110101010;
assign LUT_4[58043] = 32'b00000000000000000010101010100010;
assign LUT_4[58044] = 32'b00000000000000000111000100100010;
assign LUT_4[58045] = 32'b00000000000000000000010000011010;
assign LUT_4[58046] = 32'b00000000000000000110011111000110;
assign LUT_4[58047] = 32'b11111111111111111111101010111110;
assign LUT_4[58048] = 32'b00000000000000010110000010010000;
assign LUT_4[58049] = 32'b00000000000000001111001110001000;
assign LUT_4[58050] = 32'b00000000000000010101011100110100;
assign LUT_4[58051] = 32'b00000000000000001110101000101100;
assign LUT_4[58052] = 32'b00000000000000010011000010101100;
assign LUT_4[58053] = 32'b00000000000000001100001110100100;
assign LUT_4[58054] = 32'b00000000000000010010011101010000;
assign LUT_4[58055] = 32'b00000000000000001011101001001000;
assign LUT_4[58056] = 32'b00000000000000001111001110100101;
assign LUT_4[58057] = 32'b00000000000000001000011010011101;
assign LUT_4[58058] = 32'b00000000000000001110101001001001;
assign LUT_4[58059] = 32'b00000000000000000111110101000001;
assign LUT_4[58060] = 32'b00000000000000001100001111000001;
assign LUT_4[58061] = 32'b00000000000000000101011010111001;
assign LUT_4[58062] = 32'b00000000000000001011101001100101;
assign LUT_4[58063] = 32'b00000000000000000100110101011101;
assign LUT_4[58064] = 32'b00000000000000010011110011111110;
assign LUT_4[58065] = 32'b00000000000000001100111111110110;
assign LUT_4[58066] = 32'b00000000000000010011001110100010;
assign LUT_4[58067] = 32'b00000000000000001100011010011010;
assign LUT_4[58068] = 32'b00000000000000010000110100011010;
assign LUT_4[58069] = 32'b00000000000000001010000000010010;
assign LUT_4[58070] = 32'b00000000000000010000001110111110;
assign LUT_4[58071] = 32'b00000000000000001001011010110110;
assign LUT_4[58072] = 32'b00000000000000001101000000010011;
assign LUT_4[58073] = 32'b00000000000000000110001100001011;
assign LUT_4[58074] = 32'b00000000000000001100011010110111;
assign LUT_4[58075] = 32'b00000000000000000101100110101111;
assign LUT_4[58076] = 32'b00000000000000001010000000101111;
assign LUT_4[58077] = 32'b00000000000000000011001100100111;
assign LUT_4[58078] = 32'b00000000000000001001011011010011;
assign LUT_4[58079] = 32'b00000000000000000010100111001011;
assign LUT_4[58080] = 32'b00000000000000010100011101010111;
assign LUT_4[58081] = 32'b00000000000000001101101001001111;
assign LUT_4[58082] = 32'b00000000000000010011110111111011;
assign LUT_4[58083] = 32'b00000000000000001101000011110011;
assign LUT_4[58084] = 32'b00000000000000010001011101110011;
assign LUT_4[58085] = 32'b00000000000000001010101001101011;
assign LUT_4[58086] = 32'b00000000000000010000111000010111;
assign LUT_4[58087] = 32'b00000000000000001010000100001111;
assign LUT_4[58088] = 32'b00000000000000001101101001101100;
assign LUT_4[58089] = 32'b00000000000000000110110101100100;
assign LUT_4[58090] = 32'b00000000000000001101000100010000;
assign LUT_4[58091] = 32'b00000000000000000110010000001000;
assign LUT_4[58092] = 32'b00000000000000001010101010001000;
assign LUT_4[58093] = 32'b00000000000000000011110110000000;
assign LUT_4[58094] = 32'b00000000000000001010000100101100;
assign LUT_4[58095] = 32'b00000000000000000011010000100100;
assign LUT_4[58096] = 32'b00000000000000010010001111000101;
assign LUT_4[58097] = 32'b00000000000000001011011010111101;
assign LUT_4[58098] = 32'b00000000000000010001101001101001;
assign LUT_4[58099] = 32'b00000000000000001010110101100001;
assign LUT_4[58100] = 32'b00000000000000001111001111100001;
assign LUT_4[58101] = 32'b00000000000000001000011011011001;
assign LUT_4[58102] = 32'b00000000000000001110101010000101;
assign LUT_4[58103] = 32'b00000000000000000111110101111101;
assign LUT_4[58104] = 32'b00000000000000001011011011011010;
assign LUT_4[58105] = 32'b00000000000000000100100111010010;
assign LUT_4[58106] = 32'b00000000000000001010110101111110;
assign LUT_4[58107] = 32'b00000000000000000100000001110110;
assign LUT_4[58108] = 32'b00000000000000001000011011110110;
assign LUT_4[58109] = 32'b00000000000000000001100111101110;
assign LUT_4[58110] = 32'b00000000000000000111110110011010;
assign LUT_4[58111] = 32'b00000000000000000001000010010010;
assign LUT_4[58112] = 32'b00000000000000010111000000010111;
assign LUT_4[58113] = 32'b00000000000000010000001100001111;
assign LUT_4[58114] = 32'b00000000000000010110011010111011;
assign LUT_4[58115] = 32'b00000000000000001111100110110011;
assign LUT_4[58116] = 32'b00000000000000010100000000110011;
assign LUT_4[58117] = 32'b00000000000000001101001100101011;
assign LUT_4[58118] = 32'b00000000000000010011011011010111;
assign LUT_4[58119] = 32'b00000000000000001100100111001111;
assign LUT_4[58120] = 32'b00000000000000010000001100101100;
assign LUT_4[58121] = 32'b00000000000000001001011000100100;
assign LUT_4[58122] = 32'b00000000000000001111100111010000;
assign LUT_4[58123] = 32'b00000000000000001000110011001000;
assign LUT_4[58124] = 32'b00000000000000001101001101001000;
assign LUT_4[58125] = 32'b00000000000000000110011001000000;
assign LUT_4[58126] = 32'b00000000000000001100100111101100;
assign LUT_4[58127] = 32'b00000000000000000101110011100100;
assign LUT_4[58128] = 32'b00000000000000010100110010000101;
assign LUT_4[58129] = 32'b00000000000000001101111101111101;
assign LUT_4[58130] = 32'b00000000000000010100001100101001;
assign LUT_4[58131] = 32'b00000000000000001101011000100001;
assign LUT_4[58132] = 32'b00000000000000010001110010100001;
assign LUT_4[58133] = 32'b00000000000000001010111110011001;
assign LUT_4[58134] = 32'b00000000000000010001001101000101;
assign LUT_4[58135] = 32'b00000000000000001010011000111101;
assign LUT_4[58136] = 32'b00000000000000001101111110011010;
assign LUT_4[58137] = 32'b00000000000000000111001010010010;
assign LUT_4[58138] = 32'b00000000000000001101011000111110;
assign LUT_4[58139] = 32'b00000000000000000110100100110110;
assign LUT_4[58140] = 32'b00000000000000001010111110110110;
assign LUT_4[58141] = 32'b00000000000000000100001010101110;
assign LUT_4[58142] = 32'b00000000000000001010011001011010;
assign LUT_4[58143] = 32'b00000000000000000011100101010010;
assign LUT_4[58144] = 32'b00000000000000010101011011011110;
assign LUT_4[58145] = 32'b00000000000000001110100111010110;
assign LUT_4[58146] = 32'b00000000000000010100110110000010;
assign LUT_4[58147] = 32'b00000000000000001110000001111010;
assign LUT_4[58148] = 32'b00000000000000010010011011111010;
assign LUT_4[58149] = 32'b00000000000000001011100111110010;
assign LUT_4[58150] = 32'b00000000000000010001110110011110;
assign LUT_4[58151] = 32'b00000000000000001011000010010110;
assign LUT_4[58152] = 32'b00000000000000001110100111110011;
assign LUT_4[58153] = 32'b00000000000000000111110011101011;
assign LUT_4[58154] = 32'b00000000000000001110000010010111;
assign LUT_4[58155] = 32'b00000000000000000111001110001111;
assign LUT_4[58156] = 32'b00000000000000001011101000001111;
assign LUT_4[58157] = 32'b00000000000000000100110100000111;
assign LUT_4[58158] = 32'b00000000000000001011000010110011;
assign LUT_4[58159] = 32'b00000000000000000100001110101011;
assign LUT_4[58160] = 32'b00000000000000010011001101001100;
assign LUT_4[58161] = 32'b00000000000000001100011001000100;
assign LUT_4[58162] = 32'b00000000000000010010100111110000;
assign LUT_4[58163] = 32'b00000000000000001011110011101000;
assign LUT_4[58164] = 32'b00000000000000010000001101101000;
assign LUT_4[58165] = 32'b00000000000000001001011001100000;
assign LUT_4[58166] = 32'b00000000000000001111101000001100;
assign LUT_4[58167] = 32'b00000000000000001000110100000100;
assign LUT_4[58168] = 32'b00000000000000001100011001100001;
assign LUT_4[58169] = 32'b00000000000000000101100101011001;
assign LUT_4[58170] = 32'b00000000000000001011110100000101;
assign LUT_4[58171] = 32'b00000000000000000100111111111101;
assign LUT_4[58172] = 32'b00000000000000001001011001111101;
assign LUT_4[58173] = 32'b00000000000000000010100101110101;
assign LUT_4[58174] = 32'b00000000000000001000110100100001;
assign LUT_4[58175] = 32'b00000000000000000010000000011001;
assign LUT_4[58176] = 32'b00000000000000011000010111101011;
assign LUT_4[58177] = 32'b00000000000000010001100011100011;
assign LUT_4[58178] = 32'b00000000000000010111110010001111;
assign LUT_4[58179] = 32'b00000000000000010000111110000111;
assign LUT_4[58180] = 32'b00000000000000010101011000000111;
assign LUT_4[58181] = 32'b00000000000000001110100011111111;
assign LUT_4[58182] = 32'b00000000000000010100110010101011;
assign LUT_4[58183] = 32'b00000000000000001101111110100011;
assign LUT_4[58184] = 32'b00000000000000010001100100000000;
assign LUT_4[58185] = 32'b00000000000000001010101111111000;
assign LUT_4[58186] = 32'b00000000000000010000111110100100;
assign LUT_4[58187] = 32'b00000000000000001010001010011100;
assign LUT_4[58188] = 32'b00000000000000001110100100011100;
assign LUT_4[58189] = 32'b00000000000000000111110000010100;
assign LUT_4[58190] = 32'b00000000000000001101111111000000;
assign LUT_4[58191] = 32'b00000000000000000111001010111000;
assign LUT_4[58192] = 32'b00000000000000010110001001011001;
assign LUT_4[58193] = 32'b00000000000000001111010101010001;
assign LUT_4[58194] = 32'b00000000000000010101100011111101;
assign LUT_4[58195] = 32'b00000000000000001110101111110101;
assign LUT_4[58196] = 32'b00000000000000010011001001110101;
assign LUT_4[58197] = 32'b00000000000000001100010101101101;
assign LUT_4[58198] = 32'b00000000000000010010100100011001;
assign LUT_4[58199] = 32'b00000000000000001011110000010001;
assign LUT_4[58200] = 32'b00000000000000001111010101101110;
assign LUT_4[58201] = 32'b00000000000000001000100001100110;
assign LUT_4[58202] = 32'b00000000000000001110110000010010;
assign LUT_4[58203] = 32'b00000000000000000111111100001010;
assign LUT_4[58204] = 32'b00000000000000001100010110001010;
assign LUT_4[58205] = 32'b00000000000000000101100010000010;
assign LUT_4[58206] = 32'b00000000000000001011110000101110;
assign LUT_4[58207] = 32'b00000000000000000100111100100110;
assign LUT_4[58208] = 32'b00000000000000010110110010110010;
assign LUT_4[58209] = 32'b00000000000000001111111110101010;
assign LUT_4[58210] = 32'b00000000000000010110001101010110;
assign LUT_4[58211] = 32'b00000000000000001111011001001110;
assign LUT_4[58212] = 32'b00000000000000010011110011001110;
assign LUT_4[58213] = 32'b00000000000000001100111111000110;
assign LUT_4[58214] = 32'b00000000000000010011001101110010;
assign LUT_4[58215] = 32'b00000000000000001100011001101010;
assign LUT_4[58216] = 32'b00000000000000001111111111000111;
assign LUT_4[58217] = 32'b00000000000000001001001010111111;
assign LUT_4[58218] = 32'b00000000000000001111011001101011;
assign LUT_4[58219] = 32'b00000000000000001000100101100011;
assign LUT_4[58220] = 32'b00000000000000001100111111100011;
assign LUT_4[58221] = 32'b00000000000000000110001011011011;
assign LUT_4[58222] = 32'b00000000000000001100011010000111;
assign LUT_4[58223] = 32'b00000000000000000101100101111111;
assign LUT_4[58224] = 32'b00000000000000010100100100100000;
assign LUT_4[58225] = 32'b00000000000000001101110000011000;
assign LUT_4[58226] = 32'b00000000000000010011111111000100;
assign LUT_4[58227] = 32'b00000000000000001101001010111100;
assign LUT_4[58228] = 32'b00000000000000010001100100111100;
assign LUT_4[58229] = 32'b00000000000000001010110000110100;
assign LUT_4[58230] = 32'b00000000000000010000111111100000;
assign LUT_4[58231] = 32'b00000000000000001010001011011000;
assign LUT_4[58232] = 32'b00000000000000001101110000110101;
assign LUT_4[58233] = 32'b00000000000000000110111100101101;
assign LUT_4[58234] = 32'b00000000000000001101001011011001;
assign LUT_4[58235] = 32'b00000000000000000110010111010001;
assign LUT_4[58236] = 32'b00000000000000001010110001010001;
assign LUT_4[58237] = 32'b00000000000000000011111101001001;
assign LUT_4[58238] = 32'b00000000000000001010001011110101;
assign LUT_4[58239] = 32'b00000000000000000011010111101101;
assign LUT_4[58240] = 32'b00000000000000011001100110011111;
assign LUT_4[58241] = 32'b00000000000000010010110010010111;
assign LUT_4[58242] = 32'b00000000000000011001000001000011;
assign LUT_4[58243] = 32'b00000000000000010010001100111011;
assign LUT_4[58244] = 32'b00000000000000010110100110111011;
assign LUT_4[58245] = 32'b00000000000000001111110010110011;
assign LUT_4[58246] = 32'b00000000000000010110000001011111;
assign LUT_4[58247] = 32'b00000000000000001111001101010111;
assign LUT_4[58248] = 32'b00000000000000010010110010110100;
assign LUT_4[58249] = 32'b00000000000000001011111110101100;
assign LUT_4[58250] = 32'b00000000000000010010001101011000;
assign LUT_4[58251] = 32'b00000000000000001011011001010000;
assign LUT_4[58252] = 32'b00000000000000001111110011010000;
assign LUT_4[58253] = 32'b00000000000000001000111111001000;
assign LUT_4[58254] = 32'b00000000000000001111001101110100;
assign LUT_4[58255] = 32'b00000000000000001000011001101100;
assign LUT_4[58256] = 32'b00000000000000010111011000001101;
assign LUT_4[58257] = 32'b00000000000000010000100100000101;
assign LUT_4[58258] = 32'b00000000000000010110110010110001;
assign LUT_4[58259] = 32'b00000000000000001111111110101001;
assign LUT_4[58260] = 32'b00000000000000010100011000101001;
assign LUT_4[58261] = 32'b00000000000000001101100100100001;
assign LUT_4[58262] = 32'b00000000000000010011110011001101;
assign LUT_4[58263] = 32'b00000000000000001100111111000101;
assign LUT_4[58264] = 32'b00000000000000010000100100100010;
assign LUT_4[58265] = 32'b00000000000000001001110000011010;
assign LUT_4[58266] = 32'b00000000000000001111111111000110;
assign LUT_4[58267] = 32'b00000000000000001001001010111110;
assign LUT_4[58268] = 32'b00000000000000001101100100111110;
assign LUT_4[58269] = 32'b00000000000000000110110000110110;
assign LUT_4[58270] = 32'b00000000000000001100111111100010;
assign LUT_4[58271] = 32'b00000000000000000110001011011010;
assign LUT_4[58272] = 32'b00000000000000011000000001100110;
assign LUT_4[58273] = 32'b00000000000000010001001101011110;
assign LUT_4[58274] = 32'b00000000000000010111011100001010;
assign LUT_4[58275] = 32'b00000000000000010000101000000010;
assign LUT_4[58276] = 32'b00000000000000010101000010000010;
assign LUT_4[58277] = 32'b00000000000000001110001101111010;
assign LUT_4[58278] = 32'b00000000000000010100011100100110;
assign LUT_4[58279] = 32'b00000000000000001101101000011110;
assign LUT_4[58280] = 32'b00000000000000010001001101111011;
assign LUT_4[58281] = 32'b00000000000000001010011001110011;
assign LUT_4[58282] = 32'b00000000000000010000101000011111;
assign LUT_4[58283] = 32'b00000000000000001001110100010111;
assign LUT_4[58284] = 32'b00000000000000001110001110010111;
assign LUT_4[58285] = 32'b00000000000000000111011010001111;
assign LUT_4[58286] = 32'b00000000000000001101101000111011;
assign LUT_4[58287] = 32'b00000000000000000110110100110011;
assign LUT_4[58288] = 32'b00000000000000010101110011010100;
assign LUT_4[58289] = 32'b00000000000000001110111111001100;
assign LUT_4[58290] = 32'b00000000000000010101001101111000;
assign LUT_4[58291] = 32'b00000000000000001110011001110000;
assign LUT_4[58292] = 32'b00000000000000010010110011110000;
assign LUT_4[58293] = 32'b00000000000000001011111111101000;
assign LUT_4[58294] = 32'b00000000000000010010001110010100;
assign LUT_4[58295] = 32'b00000000000000001011011010001100;
assign LUT_4[58296] = 32'b00000000000000001110111111101001;
assign LUT_4[58297] = 32'b00000000000000001000001011100001;
assign LUT_4[58298] = 32'b00000000000000001110011010001101;
assign LUT_4[58299] = 32'b00000000000000000111100110000101;
assign LUT_4[58300] = 32'b00000000000000001100000000000101;
assign LUT_4[58301] = 32'b00000000000000000101001011111101;
assign LUT_4[58302] = 32'b00000000000000001011011010101001;
assign LUT_4[58303] = 32'b00000000000000000100100110100001;
assign LUT_4[58304] = 32'b00000000000000011010111101110011;
assign LUT_4[58305] = 32'b00000000000000010100001001101011;
assign LUT_4[58306] = 32'b00000000000000011010011000010111;
assign LUT_4[58307] = 32'b00000000000000010011100100001111;
assign LUT_4[58308] = 32'b00000000000000010111111110001111;
assign LUT_4[58309] = 32'b00000000000000010001001010000111;
assign LUT_4[58310] = 32'b00000000000000010111011000110011;
assign LUT_4[58311] = 32'b00000000000000010000100100101011;
assign LUT_4[58312] = 32'b00000000000000010100001010001000;
assign LUT_4[58313] = 32'b00000000000000001101010110000000;
assign LUT_4[58314] = 32'b00000000000000010011100100101100;
assign LUT_4[58315] = 32'b00000000000000001100110000100100;
assign LUT_4[58316] = 32'b00000000000000010001001010100100;
assign LUT_4[58317] = 32'b00000000000000001010010110011100;
assign LUT_4[58318] = 32'b00000000000000010000100101001000;
assign LUT_4[58319] = 32'b00000000000000001001110001000000;
assign LUT_4[58320] = 32'b00000000000000011000101111100001;
assign LUT_4[58321] = 32'b00000000000000010001111011011001;
assign LUT_4[58322] = 32'b00000000000000011000001010000101;
assign LUT_4[58323] = 32'b00000000000000010001010101111101;
assign LUT_4[58324] = 32'b00000000000000010101101111111101;
assign LUT_4[58325] = 32'b00000000000000001110111011110101;
assign LUT_4[58326] = 32'b00000000000000010101001010100001;
assign LUT_4[58327] = 32'b00000000000000001110010110011001;
assign LUT_4[58328] = 32'b00000000000000010001111011110110;
assign LUT_4[58329] = 32'b00000000000000001011000111101110;
assign LUT_4[58330] = 32'b00000000000000010001010110011010;
assign LUT_4[58331] = 32'b00000000000000001010100010010010;
assign LUT_4[58332] = 32'b00000000000000001110111100010010;
assign LUT_4[58333] = 32'b00000000000000001000001000001010;
assign LUT_4[58334] = 32'b00000000000000001110010110110110;
assign LUT_4[58335] = 32'b00000000000000000111100010101110;
assign LUT_4[58336] = 32'b00000000000000011001011000111010;
assign LUT_4[58337] = 32'b00000000000000010010100100110010;
assign LUT_4[58338] = 32'b00000000000000011000110011011110;
assign LUT_4[58339] = 32'b00000000000000010001111111010110;
assign LUT_4[58340] = 32'b00000000000000010110011001010110;
assign LUT_4[58341] = 32'b00000000000000001111100101001110;
assign LUT_4[58342] = 32'b00000000000000010101110011111010;
assign LUT_4[58343] = 32'b00000000000000001110111111110010;
assign LUT_4[58344] = 32'b00000000000000010010100101001111;
assign LUT_4[58345] = 32'b00000000000000001011110001000111;
assign LUT_4[58346] = 32'b00000000000000010001111111110011;
assign LUT_4[58347] = 32'b00000000000000001011001011101011;
assign LUT_4[58348] = 32'b00000000000000001111100101101011;
assign LUT_4[58349] = 32'b00000000000000001000110001100011;
assign LUT_4[58350] = 32'b00000000000000001111000000001111;
assign LUT_4[58351] = 32'b00000000000000001000001100000111;
assign LUT_4[58352] = 32'b00000000000000010111001010101000;
assign LUT_4[58353] = 32'b00000000000000010000010110100000;
assign LUT_4[58354] = 32'b00000000000000010110100101001100;
assign LUT_4[58355] = 32'b00000000000000001111110001000100;
assign LUT_4[58356] = 32'b00000000000000010100001011000100;
assign LUT_4[58357] = 32'b00000000000000001101010110111100;
assign LUT_4[58358] = 32'b00000000000000010011100101101000;
assign LUT_4[58359] = 32'b00000000000000001100110001100000;
assign LUT_4[58360] = 32'b00000000000000010000010110111101;
assign LUT_4[58361] = 32'b00000000000000001001100010110101;
assign LUT_4[58362] = 32'b00000000000000001111110001100001;
assign LUT_4[58363] = 32'b00000000000000001000111101011001;
assign LUT_4[58364] = 32'b00000000000000001101010111011001;
assign LUT_4[58365] = 32'b00000000000000000110100011010001;
assign LUT_4[58366] = 32'b00000000000000001100110001111101;
assign LUT_4[58367] = 32'b00000000000000000101111101110101;
assign LUT_4[58368] = 32'b00000000000000010100101011001011;
assign LUT_4[58369] = 32'b00000000000000001101110111000011;
assign LUT_4[58370] = 32'b00000000000000010100000101101111;
assign LUT_4[58371] = 32'b00000000000000001101010001100111;
assign LUT_4[58372] = 32'b00000000000000010001101011100111;
assign LUT_4[58373] = 32'b00000000000000001010110111011111;
assign LUT_4[58374] = 32'b00000000000000010001000110001011;
assign LUT_4[58375] = 32'b00000000000000001010010010000011;
assign LUT_4[58376] = 32'b00000000000000001101110111100000;
assign LUT_4[58377] = 32'b00000000000000000111000011011000;
assign LUT_4[58378] = 32'b00000000000000001101010010000100;
assign LUT_4[58379] = 32'b00000000000000000110011101111100;
assign LUT_4[58380] = 32'b00000000000000001010110111111100;
assign LUT_4[58381] = 32'b00000000000000000100000011110100;
assign LUT_4[58382] = 32'b00000000000000001010010010100000;
assign LUT_4[58383] = 32'b00000000000000000011011110011000;
assign LUT_4[58384] = 32'b00000000000000010010011100111001;
assign LUT_4[58385] = 32'b00000000000000001011101000110001;
assign LUT_4[58386] = 32'b00000000000000010001110111011101;
assign LUT_4[58387] = 32'b00000000000000001011000011010101;
assign LUT_4[58388] = 32'b00000000000000001111011101010101;
assign LUT_4[58389] = 32'b00000000000000001000101001001101;
assign LUT_4[58390] = 32'b00000000000000001110110111111001;
assign LUT_4[58391] = 32'b00000000000000001000000011110001;
assign LUT_4[58392] = 32'b00000000000000001011101001001110;
assign LUT_4[58393] = 32'b00000000000000000100110101000110;
assign LUT_4[58394] = 32'b00000000000000001011000011110010;
assign LUT_4[58395] = 32'b00000000000000000100001111101010;
assign LUT_4[58396] = 32'b00000000000000001000101001101010;
assign LUT_4[58397] = 32'b00000000000000000001110101100010;
assign LUT_4[58398] = 32'b00000000000000001000000100001110;
assign LUT_4[58399] = 32'b00000000000000000001010000000110;
assign LUT_4[58400] = 32'b00000000000000010011000110010010;
assign LUT_4[58401] = 32'b00000000000000001100010010001010;
assign LUT_4[58402] = 32'b00000000000000010010100000110110;
assign LUT_4[58403] = 32'b00000000000000001011101100101110;
assign LUT_4[58404] = 32'b00000000000000010000000110101110;
assign LUT_4[58405] = 32'b00000000000000001001010010100110;
assign LUT_4[58406] = 32'b00000000000000001111100001010010;
assign LUT_4[58407] = 32'b00000000000000001000101101001010;
assign LUT_4[58408] = 32'b00000000000000001100010010100111;
assign LUT_4[58409] = 32'b00000000000000000101011110011111;
assign LUT_4[58410] = 32'b00000000000000001011101101001011;
assign LUT_4[58411] = 32'b00000000000000000100111001000011;
assign LUT_4[58412] = 32'b00000000000000001001010011000011;
assign LUT_4[58413] = 32'b00000000000000000010011110111011;
assign LUT_4[58414] = 32'b00000000000000001000101101100111;
assign LUT_4[58415] = 32'b00000000000000000001111001011111;
assign LUT_4[58416] = 32'b00000000000000010000111000000000;
assign LUT_4[58417] = 32'b00000000000000001010000011111000;
assign LUT_4[58418] = 32'b00000000000000010000010010100100;
assign LUT_4[58419] = 32'b00000000000000001001011110011100;
assign LUT_4[58420] = 32'b00000000000000001101111000011100;
assign LUT_4[58421] = 32'b00000000000000000111000100010100;
assign LUT_4[58422] = 32'b00000000000000001101010011000000;
assign LUT_4[58423] = 32'b00000000000000000110011110111000;
assign LUT_4[58424] = 32'b00000000000000001010000100010101;
assign LUT_4[58425] = 32'b00000000000000000011010000001101;
assign LUT_4[58426] = 32'b00000000000000001001011110111001;
assign LUT_4[58427] = 32'b00000000000000000010101010110001;
assign LUT_4[58428] = 32'b00000000000000000111000100110001;
assign LUT_4[58429] = 32'b00000000000000000000010000101001;
assign LUT_4[58430] = 32'b00000000000000000110011111010101;
assign LUT_4[58431] = 32'b11111111111111111111101011001101;
assign LUT_4[58432] = 32'b00000000000000010110000010011111;
assign LUT_4[58433] = 32'b00000000000000001111001110010111;
assign LUT_4[58434] = 32'b00000000000000010101011101000011;
assign LUT_4[58435] = 32'b00000000000000001110101000111011;
assign LUT_4[58436] = 32'b00000000000000010011000010111011;
assign LUT_4[58437] = 32'b00000000000000001100001110110011;
assign LUT_4[58438] = 32'b00000000000000010010011101011111;
assign LUT_4[58439] = 32'b00000000000000001011101001010111;
assign LUT_4[58440] = 32'b00000000000000001111001110110100;
assign LUT_4[58441] = 32'b00000000000000001000011010101100;
assign LUT_4[58442] = 32'b00000000000000001110101001011000;
assign LUT_4[58443] = 32'b00000000000000000111110101010000;
assign LUT_4[58444] = 32'b00000000000000001100001111010000;
assign LUT_4[58445] = 32'b00000000000000000101011011001000;
assign LUT_4[58446] = 32'b00000000000000001011101001110100;
assign LUT_4[58447] = 32'b00000000000000000100110101101100;
assign LUT_4[58448] = 32'b00000000000000010011110100001101;
assign LUT_4[58449] = 32'b00000000000000001101000000000101;
assign LUT_4[58450] = 32'b00000000000000010011001110110001;
assign LUT_4[58451] = 32'b00000000000000001100011010101001;
assign LUT_4[58452] = 32'b00000000000000010000110100101001;
assign LUT_4[58453] = 32'b00000000000000001010000000100001;
assign LUT_4[58454] = 32'b00000000000000010000001111001101;
assign LUT_4[58455] = 32'b00000000000000001001011011000101;
assign LUT_4[58456] = 32'b00000000000000001101000000100010;
assign LUT_4[58457] = 32'b00000000000000000110001100011010;
assign LUT_4[58458] = 32'b00000000000000001100011011000110;
assign LUT_4[58459] = 32'b00000000000000000101100110111110;
assign LUT_4[58460] = 32'b00000000000000001010000000111110;
assign LUT_4[58461] = 32'b00000000000000000011001100110110;
assign LUT_4[58462] = 32'b00000000000000001001011011100010;
assign LUT_4[58463] = 32'b00000000000000000010100111011010;
assign LUT_4[58464] = 32'b00000000000000010100011101100110;
assign LUT_4[58465] = 32'b00000000000000001101101001011110;
assign LUT_4[58466] = 32'b00000000000000010011111000001010;
assign LUT_4[58467] = 32'b00000000000000001101000100000010;
assign LUT_4[58468] = 32'b00000000000000010001011110000010;
assign LUT_4[58469] = 32'b00000000000000001010101001111010;
assign LUT_4[58470] = 32'b00000000000000010000111000100110;
assign LUT_4[58471] = 32'b00000000000000001010000100011110;
assign LUT_4[58472] = 32'b00000000000000001101101001111011;
assign LUT_4[58473] = 32'b00000000000000000110110101110011;
assign LUT_4[58474] = 32'b00000000000000001101000100011111;
assign LUT_4[58475] = 32'b00000000000000000110010000010111;
assign LUT_4[58476] = 32'b00000000000000001010101010010111;
assign LUT_4[58477] = 32'b00000000000000000011110110001111;
assign LUT_4[58478] = 32'b00000000000000001010000100111011;
assign LUT_4[58479] = 32'b00000000000000000011010000110011;
assign LUT_4[58480] = 32'b00000000000000010010001111010100;
assign LUT_4[58481] = 32'b00000000000000001011011011001100;
assign LUT_4[58482] = 32'b00000000000000010001101001111000;
assign LUT_4[58483] = 32'b00000000000000001010110101110000;
assign LUT_4[58484] = 32'b00000000000000001111001111110000;
assign LUT_4[58485] = 32'b00000000000000001000011011101000;
assign LUT_4[58486] = 32'b00000000000000001110101010010100;
assign LUT_4[58487] = 32'b00000000000000000111110110001100;
assign LUT_4[58488] = 32'b00000000000000001011011011101001;
assign LUT_4[58489] = 32'b00000000000000000100100111100001;
assign LUT_4[58490] = 32'b00000000000000001010110110001101;
assign LUT_4[58491] = 32'b00000000000000000100000010000101;
assign LUT_4[58492] = 32'b00000000000000001000011100000101;
assign LUT_4[58493] = 32'b00000000000000000001100111111101;
assign LUT_4[58494] = 32'b00000000000000000111110110101001;
assign LUT_4[58495] = 32'b00000000000000000001000010100001;
assign LUT_4[58496] = 32'b00000000000000010111010001010011;
assign LUT_4[58497] = 32'b00000000000000010000011101001011;
assign LUT_4[58498] = 32'b00000000000000010110101011110111;
assign LUT_4[58499] = 32'b00000000000000001111110111101111;
assign LUT_4[58500] = 32'b00000000000000010100010001101111;
assign LUT_4[58501] = 32'b00000000000000001101011101100111;
assign LUT_4[58502] = 32'b00000000000000010011101100010011;
assign LUT_4[58503] = 32'b00000000000000001100111000001011;
assign LUT_4[58504] = 32'b00000000000000010000011101101000;
assign LUT_4[58505] = 32'b00000000000000001001101001100000;
assign LUT_4[58506] = 32'b00000000000000001111111000001100;
assign LUT_4[58507] = 32'b00000000000000001001000100000100;
assign LUT_4[58508] = 32'b00000000000000001101011110000100;
assign LUT_4[58509] = 32'b00000000000000000110101001111100;
assign LUT_4[58510] = 32'b00000000000000001100111000101000;
assign LUT_4[58511] = 32'b00000000000000000110000100100000;
assign LUT_4[58512] = 32'b00000000000000010101000011000001;
assign LUT_4[58513] = 32'b00000000000000001110001110111001;
assign LUT_4[58514] = 32'b00000000000000010100011101100101;
assign LUT_4[58515] = 32'b00000000000000001101101001011101;
assign LUT_4[58516] = 32'b00000000000000010010000011011101;
assign LUT_4[58517] = 32'b00000000000000001011001111010101;
assign LUT_4[58518] = 32'b00000000000000010001011110000001;
assign LUT_4[58519] = 32'b00000000000000001010101001111001;
assign LUT_4[58520] = 32'b00000000000000001110001111010110;
assign LUT_4[58521] = 32'b00000000000000000111011011001110;
assign LUT_4[58522] = 32'b00000000000000001101101001111010;
assign LUT_4[58523] = 32'b00000000000000000110110101110010;
assign LUT_4[58524] = 32'b00000000000000001011001111110010;
assign LUT_4[58525] = 32'b00000000000000000100011011101010;
assign LUT_4[58526] = 32'b00000000000000001010101010010110;
assign LUT_4[58527] = 32'b00000000000000000011110110001110;
assign LUT_4[58528] = 32'b00000000000000010101101100011010;
assign LUT_4[58529] = 32'b00000000000000001110111000010010;
assign LUT_4[58530] = 32'b00000000000000010101000110111110;
assign LUT_4[58531] = 32'b00000000000000001110010010110110;
assign LUT_4[58532] = 32'b00000000000000010010101100110110;
assign LUT_4[58533] = 32'b00000000000000001011111000101110;
assign LUT_4[58534] = 32'b00000000000000010010000111011010;
assign LUT_4[58535] = 32'b00000000000000001011010011010010;
assign LUT_4[58536] = 32'b00000000000000001110111000101111;
assign LUT_4[58537] = 32'b00000000000000001000000100100111;
assign LUT_4[58538] = 32'b00000000000000001110010011010011;
assign LUT_4[58539] = 32'b00000000000000000111011111001011;
assign LUT_4[58540] = 32'b00000000000000001011111001001011;
assign LUT_4[58541] = 32'b00000000000000000101000101000011;
assign LUT_4[58542] = 32'b00000000000000001011010011101111;
assign LUT_4[58543] = 32'b00000000000000000100011111100111;
assign LUT_4[58544] = 32'b00000000000000010011011110001000;
assign LUT_4[58545] = 32'b00000000000000001100101010000000;
assign LUT_4[58546] = 32'b00000000000000010010111000101100;
assign LUT_4[58547] = 32'b00000000000000001100000100100100;
assign LUT_4[58548] = 32'b00000000000000010000011110100100;
assign LUT_4[58549] = 32'b00000000000000001001101010011100;
assign LUT_4[58550] = 32'b00000000000000001111111001001000;
assign LUT_4[58551] = 32'b00000000000000001001000101000000;
assign LUT_4[58552] = 32'b00000000000000001100101010011101;
assign LUT_4[58553] = 32'b00000000000000000101110110010101;
assign LUT_4[58554] = 32'b00000000000000001100000101000001;
assign LUT_4[58555] = 32'b00000000000000000101010000111001;
assign LUT_4[58556] = 32'b00000000000000001001101010111001;
assign LUT_4[58557] = 32'b00000000000000000010110110110001;
assign LUT_4[58558] = 32'b00000000000000001001000101011101;
assign LUT_4[58559] = 32'b00000000000000000010010001010101;
assign LUT_4[58560] = 32'b00000000000000011000101000100111;
assign LUT_4[58561] = 32'b00000000000000010001110100011111;
assign LUT_4[58562] = 32'b00000000000000011000000011001011;
assign LUT_4[58563] = 32'b00000000000000010001001111000011;
assign LUT_4[58564] = 32'b00000000000000010101101001000011;
assign LUT_4[58565] = 32'b00000000000000001110110100111011;
assign LUT_4[58566] = 32'b00000000000000010101000011100111;
assign LUT_4[58567] = 32'b00000000000000001110001111011111;
assign LUT_4[58568] = 32'b00000000000000010001110100111100;
assign LUT_4[58569] = 32'b00000000000000001011000000110100;
assign LUT_4[58570] = 32'b00000000000000010001001111100000;
assign LUT_4[58571] = 32'b00000000000000001010011011011000;
assign LUT_4[58572] = 32'b00000000000000001110110101011000;
assign LUT_4[58573] = 32'b00000000000000001000000001010000;
assign LUT_4[58574] = 32'b00000000000000001110001111111100;
assign LUT_4[58575] = 32'b00000000000000000111011011110100;
assign LUT_4[58576] = 32'b00000000000000010110011010010101;
assign LUT_4[58577] = 32'b00000000000000001111100110001101;
assign LUT_4[58578] = 32'b00000000000000010101110100111001;
assign LUT_4[58579] = 32'b00000000000000001111000000110001;
assign LUT_4[58580] = 32'b00000000000000010011011010110001;
assign LUT_4[58581] = 32'b00000000000000001100100110101001;
assign LUT_4[58582] = 32'b00000000000000010010110101010101;
assign LUT_4[58583] = 32'b00000000000000001100000001001101;
assign LUT_4[58584] = 32'b00000000000000001111100110101010;
assign LUT_4[58585] = 32'b00000000000000001000110010100010;
assign LUT_4[58586] = 32'b00000000000000001111000001001110;
assign LUT_4[58587] = 32'b00000000000000001000001101000110;
assign LUT_4[58588] = 32'b00000000000000001100100111000110;
assign LUT_4[58589] = 32'b00000000000000000101110010111110;
assign LUT_4[58590] = 32'b00000000000000001100000001101010;
assign LUT_4[58591] = 32'b00000000000000000101001101100010;
assign LUT_4[58592] = 32'b00000000000000010111000011101110;
assign LUT_4[58593] = 32'b00000000000000010000001111100110;
assign LUT_4[58594] = 32'b00000000000000010110011110010010;
assign LUT_4[58595] = 32'b00000000000000001111101010001010;
assign LUT_4[58596] = 32'b00000000000000010100000100001010;
assign LUT_4[58597] = 32'b00000000000000001101010000000010;
assign LUT_4[58598] = 32'b00000000000000010011011110101110;
assign LUT_4[58599] = 32'b00000000000000001100101010100110;
assign LUT_4[58600] = 32'b00000000000000010000010000000011;
assign LUT_4[58601] = 32'b00000000000000001001011011111011;
assign LUT_4[58602] = 32'b00000000000000001111101010100111;
assign LUT_4[58603] = 32'b00000000000000001000110110011111;
assign LUT_4[58604] = 32'b00000000000000001101010000011111;
assign LUT_4[58605] = 32'b00000000000000000110011100010111;
assign LUT_4[58606] = 32'b00000000000000001100101011000011;
assign LUT_4[58607] = 32'b00000000000000000101110110111011;
assign LUT_4[58608] = 32'b00000000000000010100110101011100;
assign LUT_4[58609] = 32'b00000000000000001110000001010100;
assign LUT_4[58610] = 32'b00000000000000010100010000000000;
assign LUT_4[58611] = 32'b00000000000000001101011011111000;
assign LUT_4[58612] = 32'b00000000000000010001110101111000;
assign LUT_4[58613] = 32'b00000000000000001011000001110000;
assign LUT_4[58614] = 32'b00000000000000010001010000011100;
assign LUT_4[58615] = 32'b00000000000000001010011100010100;
assign LUT_4[58616] = 32'b00000000000000001110000001110001;
assign LUT_4[58617] = 32'b00000000000000000111001101101001;
assign LUT_4[58618] = 32'b00000000000000001101011100010101;
assign LUT_4[58619] = 32'b00000000000000000110101000001101;
assign LUT_4[58620] = 32'b00000000000000001011000010001101;
assign LUT_4[58621] = 32'b00000000000000000100001110000101;
assign LUT_4[58622] = 32'b00000000000000001010011100110001;
assign LUT_4[58623] = 32'b00000000000000000011101000101001;
assign LUT_4[58624] = 32'b00000000000000011001100110101110;
assign LUT_4[58625] = 32'b00000000000000010010110010100110;
assign LUT_4[58626] = 32'b00000000000000011001000001010010;
assign LUT_4[58627] = 32'b00000000000000010010001101001010;
assign LUT_4[58628] = 32'b00000000000000010110100111001010;
assign LUT_4[58629] = 32'b00000000000000001111110011000010;
assign LUT_4[58630] = 32'b00000000000000010110000001101110;
assign LUT_4[58631] = 32'b00000000000000001111001101100110;
assign LUT_4[58632] = 32'b00000000000000010010110011000011;
assign LUT_4[58633] = 32'b00000000000000001011111110111011;
assign LUT_4[58634] = 32'b00000000000000010010001101100111;
assign LUT_4[58635] = 32'b00000000000000001011011001011111;
assign LUT_4[58636] = 32'b00000000000000001111110011011111;
assign LUT_4[58637] = 32'b00000000000000001000111111010111;
assign LUT_4[58638] = 32'b00000000000000001111001110000011;
assign LUT_4[58639] = 32'b00000000000000001000011001111011;
assign LUT_4[58640] = 32'b00000000000000010111011000011100;
assign LUT_4[58641] = 32'b00000000000000010000100100010100;
assign LUT_4[58642] = 32'b00000000000000010110110011000000;
assign LUT_4[58643] = 32'b00000000000000001111111110111000;
assign LUT_4[58644] = 32'b00000000000000010100011000111000;
assign LUT_4[58645] = 32'b00000000000000001101100100110000;
assign LUT_4[58646] = 32'b00000000000000010011110011011100;
assign LUT_4[58647] = 32'b00000000000000001100111111010100;
assign LUT_4[58648] = 32'b00000000000000010000100100110001;
assign LUT_4[58649] = 32'b00000000000000001001110000101001;
assign LUT_4[58650] = 32'b00000000000000001111111111010101;
assign LUT_4[58651] = 32'b00000000000000001001001011001101;
assign LUT_4[58652] = 32'b00000000000000001101100101001101;
assign LUT_4[58653] = 32'b00000000000000000110110001000101;
assign LUT_4[58654] = 32'b00000000000000001100111111110001;
assign LUT_4[58655] = 32'b00000000000000000110001011101001;
assign LUT_4[58656] = 32'b00000000000000011000000001110101;
assign LUT_4[58657] = 32'b00000000000000010001001101101101;
assign LUT_4[58658] = 32'b00000000000000010111011100011001;
assign LUT_4[58659] = 32'b00000000000000010000101000010001;
assign LUT_4[58660] = 32'b00000000000000010101000010010001;
assign LUT_4[58661] = 32'b00000000000000001110001110001001;
assign LUT_4[58662] = 32'b00000000000000010100011100110101;
assign LUT_4[58663] = 32'b00000000000000001101101000101101;
assign LUT_4[58664] = 32'b00000000000000010001001110001010;
assign LUT_4[58665] = 32'b00000000000000001010011010000010;
assign LUT_4[58666] = 32'b00000000000000010000101000101110;
assign LUT_4[58667] = 32'b00000000000000001001110100100110;
assign LUT_4[58668] = 32'b00000000000000001110001110100110;
assign LUT_4[58669] = 32'b00000000000000000111011010011110;
assign LUT_4[58670] = 32'b00000000000000001101101001001010;
assign LUT_4[58671] = 32'b00000000000000000110110101000010;
assign LUT_4[58672] = 32'b00000000000000010101110011100011;
assign LUT_4[58673] = 32'b00000000000000001110111111011011;
assign LUT_4[58674] = 32'b00000000000000010101001110000111;
assign LUT_4[58675] = 32'b00000000000000001110011001111111;
assign LUT_4[58676] = 32'b00000000000000010010110011111111;
assign LUT_4[58677] = 32'b00000000000000001011111111110111;
assign LUT_4[58678] = 32'b00000000000000010010001110100011;
assign LUT_4[58679] = 32'b00000000000000001011011010011011;
assign LUT_4[58680] = 32'b00000000000000001110111111111000;
assign LUT_4[58681] = 32'b00000000000000001000001011110000;
assign LUT_4[58682] = 32'b00000000000000001110011010011100;
assign LUT_4[58683] = 32'b00000000000000000111100110010100;
assign LUT_4[58684] = 32'b00000000000000001100000000010100;
assign LUT_4[58685] = 32'b00000000000000000101001100001100;
assign LUT_4[58686] = 32'b00000000000000001011011010111000;
assign LUT_4[58687] = 32'b00000000000000000100100110110000;
assign LUT_4[58688] = 32'b00000000000000011010111110000010;
assign LUT_4[58689] = 32'b00000000000000010100001001111010;
assign LUT_4[58690] = 32'b00000000000000011010011000100110;
assign LUT_4[58691] = 32'b00000000000000010011100100011110;
assign LUT_4[58692] = 32'b00000000000000010111111110011110;
assign LUT_4[58693] = 32'b00000000000000010001001010010110;
assign LUT_4[58694] = 32'b00000000000000010111011001000010;
assign LUT_4[58695] = 32'b00000000000000010000100100111010;
assign LUT_4[58696] = 32'b00000000000000010100001010010111;
assign LUT_4[58697] = 32'b00000000000000001101010110001111;
assign LUT_4[58698] = 32'b00000000000000010011100100111011;
assign LUT_4[58699] = 32'b00000000000000001100110000110011;
assign LUT_4[58700] = 32'b00000000000000010001001010110011;
assign LUT_4[58701] = 32'b00000000000000001010010110101011;
assign LUT_4[58702] = 32'b00000000000000010000100101010111;
assign LUT_4[58703] = 32'b00000000000000001001110001001111;
assign LUT_4[58704] = 32'b00000000000000011000101111110000;
assign LUT_4[58705] = 32'b00000000000000010001111011101000;
assign LUT_4[58706] = 32'b00000000000000011000001010010100;
assign LUT_4[58707] = 32'b00000000000000010001010110001100;
assign LUT_4[58708] = 32'b00000000000000010101110000001100;
assign LUT_4[58709] = 32'b00000000000000001110111100000100;
assign LUT_4[58710] = 32'b00000000000000010101001010110000;
assign LUT_4[58711] = 32'b00000000000000001110010110101000;
assign LUT_4[58712] = 32'b00000000000000010001111100000101;
assign LUT_4[58713] = 32'b00000000000000001011000111111101;
assign LUT_4[58714] = 32'b00000000000000010001010110101001;
assign LUT_4[58715] = 32'b00000000000000001010100010100001;
assign LUT_4[58716] = 32'b00000000000000001110111100100001;
assign LUT_4[58717] = 32'b00000000000000001000001000011001;
assign LUT_4[58718] = 32'b00000000000000001110010111000101;
assign LUT_4[58719] = 32'b00000000000000000111100010111101;
assign LUT_4[58720] = 32'b00000000000000011001011001001001;
assign LUT_4[58721] = 32'b00000000000000010010100101000001;
assign LUT_4[58722] = 32'b00000000000000011000110011101101;
assign LUT_4[58723] = 32'b00000000000000010001111111100101;
assign LUT_4[58724] = 32'b00000000000000010110011001100101;
assign LUT_4[58725] = 32'b00000000000000001111100101011101;
assign LUT_4[58726] = 32'b00000000000000010101110100001001;
assign LUT_4[58727] = 32'b00000000000000001111000000000001;
assign LUT_4[58728] = 32'b00000000000000010010100101011110;
assign LUT_4[58729] = 32'b00000000000000001011110001010110;
assign LUT_4[58730] = 32'b00000000000000010010000000000010;
assign LUT_4[58731] = 32'b00000000000000001011001011111010;
assign LUT_4[58732] = 32'b00000000000000001111100101111010;
assign LUT_4[58733] = 32'b00000000000000001000110001110010;
assign LUT_4[58734] = 32'b00000000000000001111000000011110;
assign LUT_4[58735] = 32'b00000000000000001000001100010110;
assign LUT_4[58736] = 32'b00000000000000010111001010110111;
assign LUT_4[58737] = 32'b00000000000000010000010110101111;
assign LUT_4[58738] = 32'b00000000000000010110100101011011;
assign LUT_4[58739] = 32'b00000000000000001111110001010011;
assign LUT_4[58740] = 32'b00000000000000010100001011010011;
assign LUT_4[58741] = 32'b00000000000000001101010111001011;
assign LUT_4[58742] = 32'b00000000000000010011100101110111;
assign LUT_4[58743] = 32'b00000000000000001100110001101111;
assign LUT_4[58744] = 32'b00000000000000010000010111001100;
assign LUT_4[58745] = 32'b00000000000000001001100011000100;
assign LUT_4[58746] = 32'b00000000000000001111110001110000;
assign LUT_4[58747] = 32'b00000000000000001000111101101000;
assign LUT_4[58748] = 32'b00000000000000001101010111101000;
assign LUT_4[58749] = 32'b00000000000000000110100011100000;
assign LUT_4[58750] = 32'b00000000000000001100110010001100;
assign LUT_4[58751] = 32'b00000000000000000101111110000100;
assign LUT_4[58752] = 32'b00000000000000011100001100110110;
assign LUT_4[58753] = 32'b00000000000000010101011000101110;
assign LUT_4[58754] = 32'b00000000000000011011100111011010;
assign LUT_4[58755] = 32'b00000000000000010100110011010010;
assign LUT_4[58756] = 32'b00000000000000011001001101010010;
assign LUT_4[58757] = 32'b00000000000000010010011001001010;
assign LUT_4[58758] = 32'b00000000000000011000100111110110;
assign LUT_4[58759] = 32'b00000000000000010001110011101110;
assign LUT_4[58760] = 32'b00000000000000010101011001001011;
assign LUT_4[58761] = 32'b00000000000000001110100101000011;
assign LUT_4[58762] = 32'b00000000000000010100110011101111;
assign LUT_4[58763] = 32'b00000000000000001101111111100111;
assign LUT_4[58764] = 32'b00000000000000010010011001100111;
assign LUT_4[58765] = 32'b00000000000000001011100101011111;
assign LUT_4[58766] = 32'b00000000000000010001110100001011;
assign LUT_4[58767] = 32'b00000000000000001011000000000011;
assign LUT_4[58768] = 32'b00000000000000011001111110100100;
assign LUT_4[58769] = 32'b00000000000000010011001010011100;
assign LUT_4[58770] = 32'b00000000000000011001011001001000;
assign LUT_4[58771] = 32'b00000000000000010010100101000000;
assign LUT_4[58772] = 32'b00000000000000010110111111000000;
assign LUT_4[58773] = 32'b00000000000000010000001010111000;
assign LUT_4[58774] = 32'b00000000000000010110011001100100;
assign LUT_4[58775] = 32'b00000000000000001111100101011100;
assign LUT_4[58776] = 32'b00000000000000010011001010111001;
assign LUT_4[58777] = 32'b00000000000000001100010110110001;
assign LUT_4[58778] = 32'b00000000000000010010100101011101;
assign LUT_4[58779] = 32'b00000000000000001011110001010101;
assign LUT_4[58780] = 32'b00000000000000010000001011010101;
assign LUT_4[58781] = 32'b00000000000000001001010111001101;
assign LUT_4[58782] = 32'b00000000000000001111100101111001;
assign LUT_4[58783] = 32'b00000000000000001000110001110001;
assign LUT_4[58784] = 32'b00000000000000011010100111111101;
assign LUT_4[58785] = 32'b00000000000000010011110011110101;
assign LUT_4[58786] = 32'b00000000000000011010000010100001;
assign LUT_4[58787] = 32'b00000000000000010011001110011001;
assign LUT_4[58788] = 32'b00000000000000010111101000011001;
assign LUT_4[58789] = 32'b00000000000000010000110100010001;
assign LUT_4[58790] = 32'b00000000000000010111000010111101;
assign LUT_4[58791] = 32'b00000000000000010000001110110101;
assign LUT_4[58792] = 32'b00000000000000010011110100010010;
assign LUT_4[58793] = 32'b00000000000000001101000000001010;
assign LUT_4[58794] = 32'b00000000000000010011001110110110;
assign LUT_4[58795] = 32'b00000000000000001100011010101110;
assign LUT_4[58796] = 32'b00000000000000010000110100101110;
assign LUT_4[58797] = 32'b00000000000000001010000000100110;
assign LUT_4[58798] = 32'b00000000000000010000001111010010;
assign LUT_4[58799] = 32'b00000000000000001001011011001010;
assign LUT_4[58800] = 32'b00000000000000011000011001101011;
assign LUT_4[58801] = 32'b00000000000000010001100101100011;
assign LUT_4[58802] = 32'b00000000000000010111110100001111;
assign LUT_4[58803] = 32'b00000000000000010001000000000111;
assign LUT_4[58804] = 32'b00000000000000010101011010000111;
assign LUT_4[58805] = 32'b00000000000000001110100101111111;
assign LUT_4[58806] = 32'b00000000000000010100110100101011;
assign LUT_4[58807] = 32'b00000000000000001110000000100011;
assign LUT_4[58808] = 32'b00000000000000010001100110000000;
assign LUT_4[58809] = 32'b00000000000000001010110001111000;
assign LUT_4[58810] = 32'b00000000000000010001000000100100;
assign LUT_4[58811] = 32'b00000000000000001010001100011100;
assign LUT_4[58812] = 32'b00000000000000001110100110011100;
assign LUT_4[58813] = 32'b00000000000000000111110010010100;
assign LUT_4[58814] = 32'b00000000000000001110000001000000;
assign LUT_4[58815] = 32'b00000000000000000111001100111000;
assign LUT_4[58816] = 32'b00000000000000011101100100001010;
assign LUT_4[58817] = 32'b00000000000000010110110000000010;
assign LUT_4[58818] = 32'b00000000000000011100111110101110;
assign LUT_4[58819] = 32'b00000000000000010110001010100110;
assign LUT_4[58820] = 32'b00000000000000011010100100100110;
assign LUT_4[58821] = 32'b00000000000000010011110000011110;
assign LUT_4[58822] = 32'b00000000000000011001111111001010;
assign LUT_4[58823] = 32'b00000000000000010011001011000010;
assign LUT_4[58824] = 32'b00000000000000010110110000011111;
assign LUT_4[58825] = 32'b00000000000000001111111100010111;
assign LUT_4[58826] = 32'b00000000000000010110001011000011;
assign LUT_4[58827] = 32'b00000000000000001111010110111011;
assign LUT_4[58828] = 32'b00000000000000010011110000111011;
assign LUT_4[58829] = 32'b00000000000000001100111100110011;
assign LUT_4[58830] = 32'b00000000000000010011001011011111;
assign LUT_4[58831] = 32'b00000000000000001100010111010111;
assign LUT_4[58832] = 32'b00000000000000011011010101111000;
assign LUT_4[58833] = 32'b00000000000000010100100001110000;
assign LUT_4[58834] = 32'b00000000000000011010110000011100;
assign LUT_4[58835] = 32'b00000000000000010011111100010100;
assign LUT_4[58836] = 32'b00000000000000011000010110010100;
assign LUT_4[58837] = 32'b00000000000000010001100010001100;
assign LUT_4[58838] = 32'b00000000000000010111110000111000;
assign LUT_4[58839] = 32'b00000000000000010000111100110000;
assign LUT_4[58840] = 32'b00000000000000010100100010001101;
assign LUT_4[58841] = 32'b00000000000000001101101110000101;
assign LUT_4[58842] = 32'b00000000000000010011111100110001;
assign LUT_4[58843] = 32'b00000000000000001101001000101001;
assign LUT_4[58844] = 32'b00000000000000010001100010101001;
assign LUT_4[58845] = 32'b00000000000000001010101110100001;
assign LUT_4[58846] = 32'b00000000000000010000111101001101;
assign LUT_4[58847] = 32'b00000000000000001010001001000101;
assign LUT_4[58848] = 32'b00000000000000011011111111010001;
assign LUT_4[58849] = 32'b00000000000000010101001011001001;
assign LUT_4[58850] = 32'b00000000000000011011011001110101;
assign LUT_4[58851] = 32'b00000000000000010100100101101101;
assign LUT_4[58852] = 32'b00000000000000011000111111101101;
assign LUT_4[58853] = 32'b00000000000000010010001011100101;
assign LUT_4[58854] = 32'b00000000000000011000011010010001;
assign LUT_4[58855] = 32'b00000000000000010001100110001001;
assign LUT_4[58856] = 32'b00000000000000010101001011100110;
assign LUT_4[58857] = 32'b00000000000000001110010111011110;
assign LUT_4[58858] = 32'b00000000000000010100100110001010;
assign LUT_4[58859] = 32'b00000000000000001101110010000010;
assign LUT_4[58860] = 32'b00000000000000010010001100000010;
assign LUT_4[58861] = 32'b00000000000000001011010111111010;
assign LUT_4[58862] = 32'b00000000000000010001100110100110;
assign LUT_4[58863] = 32'b00000000000000001010110010011110;
assign LUT_4[58864] = 32'b00000000000000011001110000111111;
assign LUT_4[58865] = 32'b00000000000000010010111100110111;
assign LUT_4[58866] = 32'b00000000000000011001001011100011;
assign LUT_4[58867] = 32'b00000000000000010010010111011011;
assign LUT_4[58868] = 32'b00000000000000010110110001011011;
assign LUT_4[58869] = 32'b00000000000000001111111101010011;
assign LUT_4[58870] = 32'b00000000000000010110001011111111;
assign LUT_4[58871] = 32'b00000000000000001111010111110111;
assign LUT_4[58872] = 32'b00000000000000010010111101010100;
assign LUT_4[58873] = 32'b00000000000000001100001001001100;
assign LUT_4[58874] = 32'b00000000000000010010010111111000;
assign LUT_4[58875] = 32'b00000000000000001011100011110000;
assign LUT_4[58876] = 32'b00000000000000001111111101110000;
assign LUT_4[58877] = 32'b00000000000000001001001001101000;
assign LUT_4[58878] = 32'b00000000000000001111011000010100;
assign LUT_4[58879] = 32'b00000000000000001000100100001100;
assign LUT_4[58880] = 32'b00000000000000010011101111010011;
assign LUT_4[58881] = 32'b00000000000000001100111011001011;
assign LUT_4[58882] = 32'b00000000000000010011001001110111;
assign LUT_4[58883] = 32'b00000000000000001100010101101111;
assign LUT_4[58884] = 32'b00000000000000010000101111101111;
assign LUT_4[58885] = 32'b00000000000000001001111011100111;
assign LUT_4[58886] = 32'b00000000000000010000001010010011;
assign LUT_4[58887] = 32'b00000000000000001001010110001011;
assign LUT_4[58888] = 32'b00000000000000001100111011101000;
assign LUT_4[58889] = 32'b00000000000000000110000111100000;
assign LUT_4[58890] = 32'b00000000000000001100010110001100;
assign LUT_4[58891] = 32'b00000000000000000101100010000100;
assign LUT_4[58892] = 32'b00000000000000001001111100000100;
assign LUT_4[58893] = 32'b00000000000000000011000111111100;
assign LUT_4[58894] = 32'b00000000000000001001010110101000;
assign LUT_4[58895] = 32'b00000000000000000010100010100000;
assign LUT_4[58896] = 32'b00000000000000010001100001000001;
assign LUT_4[58897] = 32'b00000000000000001010101100111001;
assign LUT_4[58898] = 32'b00000000000000010000111011100101;
assign LUT_4[58899] = 32'b00000000000000001010000111011101;
assign LUT_4[58900] = 32'b00000000000000001110100001011101;
assign LUT_4[58901] = 32'b00000000000000000111101101010101;
assign LUT_4[58902] = 32'b00000000000000001101111100000001;
assign LUT_4[58903] = 32'b00000000000000000111000111111001;
assign LUT_4[58904] = 32'b00000000000000001010101101010110;
assign LUT_4[58905] = 32'b00000000000000000011111001001110;
assign LUT_4[58906] = 32'b00000000000000001010000111111010;
assign LUT_4[58907] = 32'b00000000000000000011010011110010;
assign LUT_4[58908] = 32'b00000000000000000111101101110010;
assign LUT_4[58909] = 32'b00000000000000000000111001101010;
assign LUT_4[58910] = 32'b00000000000000000111001000010110;
assign LUT_4[58911] = 32'b00000000000000000000010100001110;
assign LUT_4[58912] = 32'b00000000000000010010001010011010;
assign LUT_4[58913] = 32'b00000000000000001011010110010010;
assign LUT_4[58914] = 32'b00000000000000010001100100111110;
assign LUT_4[58915] = 32'b00000000000000001010110000110110;
assign LUT_4[58916] = 32'b00000000000000001111001010110110;
assign LUT_4[58917] = 32'b00000000000000001000010110101110;
assign LUT_4[58918] = 32'b00000000000000001110100101011010;
assign LUT_4[58919] = 32'b00000000000000000111110001010010;
assign LUT_4[58920] = 32'b00000000000000001011010110101111;
assign LUT_4[58921] = 32'b00000000000000000100100010100111;
assign LUT_4[58922] = 32'b00000000000000001010110001010011;
assign LUT_4[58923] = 32'b00000000000000000011111101001011;
assign LUT_4[58924] = 32'b00000000000000001000010111001011;
assign LUT_4[58925] = 32'b00000000000000000001100011000011;
assign LUT_4[58926] = 32'b00000000000000000111110001101111;
assign LUT_4[58927] = 32'b00000000000000000000111101100111;
assign LUT_4[58928] = 32'b00000000000000001111111100001000;
assign LUT_4[58929] = 32'b00000000000000001001001000000000;
assign LUT_4[58930] = 32'b00000000000000001111010110101100;
assign LUT_4[58931] = 32'b00000000000000001000100010100100;
assign LUT_4[58932] = 32'b00000000000000001100111100100100;
assign LUT_4[58933] = 32'b00000000000000000110001000011100;
assign LUT_4[58934] = 32'b00000000000000001100010111001000;
assign LUT_4[58935] = 32'b00000000000000000101100011000000;
assign LUT_4[58936] = 32'b00000000000000001001001000011101;
assign LUT_4[58937] = 32'b00000000000000000010010100010101;
assign LUT_4[58938] = 32'b00000000000000001000100011000001;
assign LUT_4[58939] = 32'b00000000000000000001101110111001;
assign LUT_4[58940] = 32'b00000000000000000110001000111001;
assign LUT_4[58941] = 32'b11111111111111111111010100110001;
assign LUT_4[58942] = 32'b00000000000000000101100011011101;
assign LUT_4[58943] = 32'b11111111111111111110101111010101;
assign LUT_4[58944] = 32'b00000000000000010101000110100111;
assign LUT_4[58945] = 32'b00000000000000001110010010011111;
assign LUT_4[58946] = 32'b00000000000000010100100001001011;
assign LUT_4[58947] = 32'b00000000000000001101101101000011;
assign LUT_4[58948] = 32'b00000000000000010010000111000011;
assign LUT_4[58949] = 32'b00000000000000001011010010111011;
assign LUT_4[58950] = 32'b00000000000000010001100001100111;
assign LUT_4[58951] = 32'b00000000000000001010101101011111;
assign LUT_4[58952] = 32'b00000000000000001110010010111100;
assign LUT_4[58953] = 32'b00000000000000000111011110110100;
assign LUT_4[58954] = 32'b00000000000000001101101101100000;
assign LUT_4[58955] = 32'b00000000000000000110111001011000;
assign LUT_4[58956] = 32'b00000000000000001011010011011000;
assign LUT_4[58957] = 32'b00000000000000000100011111010000;
assign LUT_4[58958] = 32'b00000000000000001010101101111100;
assign LUT_4[58959] = 32'b00000000000000000011111001110100;
assign LUT_4[58960] = 32'b00000000000000010010111000010101;
assign LUT_4[58961] = 32'b00000000000000001100000100001101;
assign LUT_4[58962] = 32'b00000000000000010010010010111001;
assign LUT_4[58963] = 32'b00000000000000001011011110110001;
assign LUT_4[58964] = 32'b00000000000000001111111000110001;
assign LUT_4[58965] = 32'b00000000000000001001000100101001;
assign LUT_4[58966] = 32'b00000000000000001111010011010101;
assign LUT_4[58967] = 32'b00000000000000001000011111001101;
assign LUT_4[58968] = 32'b00000000000000001100000100101010;
assign LUT_4[58969] = 32'b00000000000000000101010000100010;
assign LUT_4[58970] = 32'b00000000000000001011011111001110;
assign LUT_4[58971] = 32'b00000000000000000100101011000110;
assign LUT_4[58972] = 32'b00000000000000001001000101000110;
assign LUT_4[58973] = 32'b00000000000000000010010000111110;
assign LUT_4[58974] = 32'b00000000000000001000011111101010;
assign LUT_4[58975] = 32'b00000000000000000001101011100010;
assign LUT_4[58976] = 32'b00000000000000010011100001101110;
assign LUT_4[58977] = 32'b00000000000000001100101101100110;
assign LUT_4[58978] = 32'b00000000000000010010111100010010;
assign LUT_4[58979] = 32'b00000000000000001100001000001010;
assign LUT_4[58980] = 32'b00000000000000010000100010001010;
assign LUT_4[58981] = 32'b00000000000000001001101110000010;
assign LUT_4[58982] = 32'b00000000000000001111111100101110;
assign LUT_4[58983] = 32'b00000000000000001001001000100110;
assign LUT_4[58984] = 32'b00000000000000001100101110000011;
assign LUT_4[58985] = 32'b00000000000000000101111001111011;
assign LUT_4[58986] = 32'b00000000000000001100001000100111;
assign LUT_4[58987] = 32'b00000000000000000101010100011111;
assign LUT_4[58988] = 32'b00000000000000001001101110011111;
assign LUT_4[58989] = 32'b00000000000000000010111010010111;
assign LUT_4[58990] = 32'b00000000000000001001001001000011;
assign LUT_4[58991] = 32'b00000000000000000010010100111011;
assign LUT_4[58992] = 32'b00000000000000010001010011011100;
assign LUT_4[58993] = 32'b00000000000000001010011111010100;
assign LUT_4[58994] = 32'b00000000000000010000101110000000;
assign LUT_4[58995] = 32'b00000000000000001001111001111000;
assign LUT_4[58996] = 32'b00000000000000001110010011111000;
assign LUT_4[58997] = 32'b00000000000000000111011111110000;
assign LUT_4[58998] = 32'b00000000000000001101101110011100;
assign LUT_4[58999] = 32'b00000000000000000110111010010100;
assign LUT_4[59000] = 32'b00000000000000001010011111110001;
assign LUT_4[59001] = 32'b00000000000000000011101011101001;
assign LUT_4[59002] = 32'b00000000000000001001111010010101;
assign LUT_4[59003] = 32'b00000000000000000011000110001101;
assign LUT_4[59004] = 32'b00000000000000000111100000001101;
assign LUT_4[59005] = 32'b00000000000000000000101100000101;
assign LUT_4[59006] = 32'b00000000000000000110111010110001;
assign LUT_4[59007] = 32'b00000000000000000000000110101001;
assign LUT_4[59008] = 32'b00000000000000010110010101011011;
assign LUT_4[59009] = 32'b00000000000000001111100001010011;
assign LUT_4[59010] = 32'b00000000000000010101101111111111;
assign LUT_4[59011] = 32'b00000000000000001110111011110111;
assign LUT_4[59012] = 32'b00000000000000010011010101110111;
assign LUT_4[59013] = 32'b00000000000000001100100001101111;
assign LUT_4[59014] = 32'b00000000000000010010110000011011;
assign LUT_4[59015] = 32'b00000000000000001011111100010011;
assign LUT_4[59016] = 32'b00000000000000001111100001110000;
assign LUT_4[59017] = 32'b00000000000000001000101101101000;
assign LUT_4[59018] = 32'b00000000000000001110111100010100;
assign LUT_4[59019] = 32'b00000000000000001000001000001100;
assign LUT_4[59020] = 32'b00000000000000001100100010001100;
assign LUT_4[59021] = 32'b00000000000000000101101110000100;
assign LUT_4[59022] = 32'b00000000000000001011111100110000;
assign LUT_4[59023] = 32'b00000000000000000101001000101000;
assign LUT_4[59024] = 32'b00000000000000010100000111001001;
assign LUT_4[59025] = 32'b00000000000000001101010011000001;
assign LUT_4[59026] = 32'b00000000000000010011100001101101;
assign LUT_4[59027] = 32'b00000000000000001100101101100101;
assign LUT_4[59028] = 32'b00000000000000010001000111100101;
assign LUT_4[59029] = 32'b00000000000000001010010011011101;
assign LUT_4[59030] = 32'b00000000000000010000100010001001;
assign LUT_4[59031] = 32'b00000000000000001001101110000001;
assign LUT_4[59032] = 32'b00000000000000001101010011011110;
assign LUT_4[59033] = 32'b00000000000000000110011111010110;
assign LUT_4[59034] = 32'b00000000000000001100101110000010;
assign LUT_4[59035] = 32'b00000000000000000101111001111010;
assign LUT_4[59036] = 32'b00000000000000001010010011111010;
assign LUT_4[59037] = 32'b00000000000000000011011111110010;
assign LUT_4[59038] = 32'b00000000000000001001101110011110;
assign LUT_4[59039] = 32'b00000000000000000010111010010110;
assign LUT_4[59040] = 32'b00000000000000010100110000100010;
assign LUT_4[59041] = 32'b00000000000000001101111100011010;
assign LUT_4[59042] = 32'b00000000000000010100001011000110;
assign LUT_4[59043] = 32'b00000000000000001101010110111110;
assign LUT_4[59044] = 32'b00000000000000010001110000111110;
assign LUT_4[59045] = 32'b00000000000000001010111100110110;
assign LUT_4[59046] = 32'b00000000000000010001001011100010;
assign LUT_4[59047] = 32'b00000000000000001010010111011010;
assign LUT_4[59048] = 32'b00000000000000001101111100110111;
assign LUT_4[59049] = 32'b00000000000000000111001000101111;
assign LUT_4[59050] = 32'b00000000000000001101010111011011;
assign LUT_4[59051] = 32'b00000000000000000110100011010011;
assign LUT_4[59052] = 32'b00000000000000001010111101010011;
assign LUT_4[59053] = 32'b00000000000000000100001001001011;
assign LUT_4[59054] = 32'b00000000000000001010010111110111;
assign LUT_4[59055] = 32'b00000000000000000011100011101111;
assign LUT_4[59056] = 32'b00000000000000010010100010010000;
assign LUT_4[59057] = 32'b00000000000000001011101110001000;
assign LUT_4[59058] = 32'b00000000000000010001111100110100;
assign LUT_4[59059] = 32'b00000000000000001011001000101100;
assign LUT_4[59060] = 32'b00000000000000001111100010101100;
assign LUT_4[59061] = 32'b00000000000000001000101110100100;
assign LUT_4[59062] = 32'b00000000000000001110111101010000;
assign LUT_4[59063] = 32'b00000000000000001000001001001000;
assign LUT_4[59064] = 32'b00000000000000001011101110100101;
assign LUT_4[59065] = 32'b00000000000000000100111010011101;
assign LUT_4[59066] = 32'b00000000000000001011001001001001;
assign LUT_4[59067] = 32'b00000000000000000100010101000001;
assign LUT_4[59068] = 32'b00000000000000001000101111000001;
assign LUT_4[59069] = 32'b00000000000000000001111010111001;
assign LUT_4[59070] = 32'b00000000000000001000001001100101;
assign LUT_4[59071] = 32'b00000000000000000001010101011101;
assign LUT_4[59072] = 32'b00000000000000010111101100101111;
assign LUT_4[59073] = 32'b00000000000000010000111000100111;
assign LUT_4[59074] = 32'b00000000000000010111000111010011;
assign LUT_4[59075] = 32'b00000000000000010000010011001011;
assign LUT_4[59076] = 32'b00000000000000010100101101001011;
assign LUT_4[59077] = 32'b00000000000000001101111001000011;
assign LUT_4[59078] = 32'b00000000000000010100000111101111;
assign LUT_4[59079] = 32'b00000000000000001101010011100111;
assign LUT_4[59080] = 32'b00000000000000010000111001000100;
assign LUT_4[59081] = 32'b00000000000000001010000100111100;
assign LUT_4[59082] = 32'b00000000000000010000010011101000;
assign LUT_4[59083] = 32'b00000000000000001001011111100000;
assign LUT_4[59084] = 32'b00000000000000001101111001100000;
assign LUT_4[59085] = 32'b00000000000000000111000101011000;
assign LUT_4[59086] = 32'b00000000000000001101010100000100;
assign LUT_4[59087] = 32'b00000000000000000110011111111100;
assign LUT_4[59088] = 32'b00000000000000010101011110011101;
assign LUT_4[59089] = 32'b00000000000000001110101010010101;
assign LUT_4[59090] = 32'b00000000000000010100111001000001;
assign LUT_4[59091] = 32'b00000000000000001110000100111001;
assign LUT_4[59092] = 32'b00000000000000010010011110111001;
assign LUT_4[59093] = 32'b00000000000000001011101010110001;
assign LUT_4[59094] = 32'b00000000000000010001111001011101;
assign LUT_4[59095] = 32'b00000000000000001011000101010101;
assign LUT_4[59096] = 32'b00000000000000001110101010110010;
assign LUT_4[59097] = 32'b00000000000000000111110110101010;
assign LUT_4[59098] = 32'b00000000000000001110000101010110;
assign LUT_4[59099] = 32'b00000000000000000111010001001110;
assign LUT_4[59100] = 32'b00000000000000001011101011001110;
assign LUT_4[59101] = 32'b00000000000000000100110111000110;
assign LUT_4[59102] = 32'b00000000000000001011000101110010;
assign LUT_4[59103] = 32'b00000000000000000100010001101010;
assign LUT_4[59104] = 32'b00000000000000010110000111110110;
assign LUT_4[59105] = 32'b00000000000000001111010011101110;
assign LUT_4[59106] = 32'b00000000000000010101100010011010;
assign LUT_4[59107] = 32'b00000000000000001110101110010010;
assign LUT_4[59108] = 32'b00000000000000010011001000010010;
assign LUT_4[59109] = 32'b00000000000000001100010100001010;
assign LUT_4[59110] = 32'b00000000000000010010100010110110;
assign LUT_4[59111] = 32'b00000000000000001011101110101110;
assign LUT_4[59112] = 32'b00000000000000001111010100001011;
assign LUT_4[59113] = 32'b00000000000000001000100000000011;
assign LUT_4[59114] = 32'b00000000000000001110101110101111;
assign LUT_4[59115] = 32'b00000000000000000111111010100111;
assign LUT_4[59116] = 32'b00000000000000001100010100100111;
assign LUT_4[59117] = 32'b00000000000000000101100000011111;
assign LUT_4[59118] = 32'b00000000000000001011101111001011;
assign LUT_4[59119] = 32'b00000000000000000100111011000011;
assign LUT_4[59120] = 32'b00000000000000010011111001100100;
assign LUT_4[59121] = 32'b00000000000000001101000101011100;
assign LUT_4[59122] = 32'b00000000000000010011010100001000;
assign LUT_4[59123] = 32'b00000000000000001100100000000000;
assign LUT_4[59124] = 32'b00000000000000010000111010000000;
assign LUT_4[59125] = 32'b00000000000000001010000101111000;
assign LUT_4[59126] = 32'b00000000000000010000010100100100;
assign LUT_4[59127] = 32'b00000000000000001001100000011100;
assign LUT_4[59128] = 32'b00000000000000001101000101111001;
assign LUT_4[59129] = 32'b00000000000000000110010001110001;
assign LUT_4[59130] = 32'b00000000000000001100100000011101;
assign LUT_4[59131] = 32'b00000000000000000101101100010101;
assign LUT_4[59132] = 32'b00000000000000001010000110010101;
assign LUT_4[59133] = 32'b00000000000000000011010010001101;
assign LUT_4[59134] = 32'b00000000000000001001100000111001;
assign LUT_4[59135] = 32'b00000000000000000010101100110001;
assign LUT_4[59136] = 32'b00000000000000011000101010110110;
assign LUT_4[59137] = 32'b00000000000000010001110110101110;
assign LUT_4[59138] = 32'b00000000000000011000000101011010;
assign LUT_4[59139] = 32'b00000000000000010001010001010010;
assign LUT_4[59140] = 32'b00000000000000010101101011010010;
assign LUT_4[59141] = 32'b00000000000000001110110111001010;
assign LUT_4[59142] = 32'b00000000000000010101000101110110;
assign LUT_4[59143] = 32'b00000000000000001110010001101110;
assign LUT_4[59144] = 32'b00000000000000010001110111001011;
assign LUT_4[59145] = 32'b00000000000000001011000011000011;
assign LUT_4[59146] = 32'b00000000000000010001010001101111;
assign LUT_4[59147] = 32'b00000000000000001010011101100111;
assign LUT_4[59148] = 32'b00000000000000001110110111100111;
assign LUT_4[59149] = 32'b00000000000000001000000011011111;
assign LUT_4[59150] = 32'b00000000000000001110010010001011;
assign LUT_4[59151] = 32'b00000000000000000111011110000011;
assign LUT_4[59152] = 32'b00000000000000010110011100100100;
assign LUT_4[59153] = 32'b00000000000000001111101000011100;
assign LUT_4[59154] = 32'b00000000000000010101110111001000;
assign LUT_4[59155] = 32'b00000000000000001111000011000000;
assign LUT_4[59156] = 32'b00000000000000010011011101000000;
assign LUT_4[59157] = 32'b00000000000000001100101000111000;
assign LUT_4[59158] = 32'b00000000000000010010110111100100;
assign LUT_4[59159] = 32'b00000000000000001100000011011100;
assign LUT_4[59160] = 32'b00000000000000001111101000111001;
assign LUT_4[59161] = 32'b00000000000000001000110100110001;
assign LUT_4[59162] = 32'b00000000000000001111000011011101;
assign LUT_4[59163] = 32'b00000000000000001000001111010101;
assign LUT_4[59164] = 32'b00000000000000001100101001010101;
assign LUT_4[59165] = 32'b00000000000000000101110101001101;
assign LUT_4[59166] = 32'b00000000000000001100000011111001;
assign LUT_4[59167] = 32'b00000000000000000101001111110001;
assign LUT_4[59168] = 32'b00000000000000010111000101111101;
assign LUT_4[59169] = 32'b00000000000000010000010001110101;
assign LUT_4[59170] = 32'b00000000000000010110100000100001;
assign LUT_4[59171] = 32'b00000000000000001111101100011001;
assign LUT_4[59172] = 32'b00000000000000010100000110011001;
assign LUT_4[59173] = 32'b00000000000000001101010010010001;
assign LUT_4[59174] = 32'b00000000000000010011100000111101;
assign LUT_4[59175] = 32'b00000000000000001100101100110101;
assign LUT_4[59176] = 32'b00000000000000010000010010010010;
assign LUT_4[59177] = 32'b00000000000000001001011110001010;
assign LUT_4[59178] = 32'b00000000000000001111101100110110;
assign LUT_4[59179] = 32'b00000000000000001000111000101110;
assign LUT_4[59180] = 32'b00000000000000001101010010101110;
assign LUT_4[59181] = 32'b00000000000000000110011110100110;
assign LUT_4[59182] = 32'b00000000000000001100101101010010;
assign LUT_4[59183] = 32'b00000000000000000101111001001010;
assign LUT_4[59184] = 32'b00000000000000010100110111101011;
assign LUT_4[59185] = 32'b00000000000000001110000011100011;
assign LUT_4[59186] = 32'b00000000000000010100010010001111;
assign LUT_4[59187] = 32'b00000000000000001101011110000111;
assign LUT_4[59188] = 32'b00000000000000010001111000000111;
assign LUT_4[59189] = 32'b00000000000000001011000011111111;
assign LUT_4[59190] = 32'b00000000000000010001010010101011;
assign LUT_4[59191] = 32'b00000000000000001010011110100011;
assign LUT_4[59192] = 32'b00000000000000001110000100000000;
assign LUT_4[59193] = 32'b00000000000000000111001111111000;
assign LUT_4[59194] = 32'b00000000000000001101011110100100;
assign LUT_4[59195] = 32'b00000000000000000110101010011100;
assign LUT_4[59196] = 32'b00000000000000001011000100011100;
assign LUT_4[59197] = 32'b00000000000000000100010000010100;
assign LUT_4[59198] = 32'b00000000000000001010011111000000;
assign LUT_4[59199] = 32'b00000000000000000011101010111000;
assign LUT_4[59200] = 32'b00000000000000011010000010001010;
assign LUT_4[59201] = 32'b00000000000000010011001110000010;
assign LUT_4[59202] = 32'b00000000000000011001011100101110;
assign LUT_4[59203] = 32'b00000000000000010010101000100110;
assign LUT_4[59204] = 32'b00000000000000010111000010100110;
assign LUT_4[59205] = 32'b00000000000000010000001110011110;
assign LUT_4[59206] = 32'b00000000000000010110011101001010;
assign LUT_4[59207] = 32'b00000000000000001111101001000010;
assign LUT_4[59208] = 32'b00000000000000010011001110011111;
assign LUT_4[59209] = 32'b00000000000000001100011010010111;
assign LUT_4[59210] = 32'b00000000000000010010101001000011;
assign LUT_4[59211] = 32'b00000000000000001011110100111011;
assign LUT_4[59212] = 32'b00000000000000010000001110111011;
assign LUT_4[59213] = 32'b00000000000000001001011010110011;
assign LUT_4[59214] = 32'b00000000000000001111101001011111;
assign LUT_4[59215] = 32'b00000000000000001000110101010111;
assign LUT_4[59216] = 32'b00000000000000010111110011111000;
assign LUT_4[59217] = 32'b00000000000000010000111111110000;
assign LUT_4[59218] = 32'b00000000000000010111001110011100;
assign LUT_4[59219] = 32'b00000000000000010000011010010100;
assign LUT_4[59220] = 32'b00000000000000010100110100010100;
assign LUT_4[59221] = 32'b00000000000000001110000000001100;
assign LUT_4[59222] = 32'b00000000000000010100001110111000;
assign LUT_4[59223] = 32'b00000000000000001101011010110000;
assign LUT_4[59224] = 32'b00000000000000010001000000001101;
assign LUT_4[59225] = 32'b00000000000000001010001100000101;
assign LUT_4[59226] = 32'b00000000000000010000011010110001;
assign LUT_4[59227] = 32'b00000000000000001001100110101001;
assign LUT_4[59228] = 32'b00000000000000001110000000101001;
assign LUT_4[59229] = 32'b00000000000000000111001100100001;
assign LUT_4[59230] = 32'b00000000000000001101011011001101;
assign LUT_4[59231] = 32'b00000000000000000110100111000101;
assign LUT_4[59232] = 32'b00000000000000011000011101010001;
assign LUT_4[59233] = 32'b00000000000000010001101001001001;
assign LUT_4[59234] = 32'b00000000000000010111110111110101;
assign LUT_4[59235] = 32'b00000000000000010001000011101101;
assign LUT_4[59236] = 32'b00000000000000010101011101101101;
assign LUT_4[59237] = 32'b00000000000000001110101001100101;
assign LUT_4[59238] = 32'b00000000000000010100111000010001;
assign LUT_4[59239] = 32'b00000000000000001110000100001001;
assign LUT_4[59240] = 32'b00000000000000010001101001100110;
assign LUT_4[59241] = 32'b00000000000000001010110101011110;
assign LUT_4[59242] = 32'b00000000000000010001000100001010;
assign LUT_4[59243] = 32'b00000000000000001010010000000010;
assign LUT_4[59244] = 32'b00000000000000001110101010000010;
assign LUT_4[59245] = 32'b00000000000000000111110101111010;
assign LUT_4[59246] = 32'b00000000000000001110000100100110;
assign LUT_4[59247] = 32'b00000000000000000111010000011110;
assign LUT_4[59248] = 32'b00000000000000010110001110111111;
assign LUT_4[59249] = 32'b00000000000000001111011010110111;
assign LUT_4[59250] = 32'b00000000000000010101101001100011;
assign LUT_4[59251] = 32'b00000000000000001110110101011011;
assign LUT_4[59252] = 32'b00000000000000010011001111011011;
assign LUT_4[59253] = 32'b00000000000000001100011011010011;
assign LUT_4[59254] = 32'b00000000000000010010101001111111;
assign LUT_4[59255] = 32'b00000000000000001011110101110111;
assign LUT_4[59256] = 32'b00000000000000001111011011010100;
assign LUT_4[59257] = 32'b00000000000000001000100111001100;
assign LUT_4[59258] = 32'b00000000000000001110110101111000;
assign LUT_4[59259] = 32'b00000000000000001000000001110000;
assign LUT_4[59260] = 32'b00000000000000001100011011110000;
assign LUT_4[59261] = 32'b00000000000000000101100111101000;
assign LUT_4[59262] = 32'b00000000000000001011110110010100;
assign LUT_4[59263] = 32'b00000000000000000101000010001100;
assign LUT_4[59264] = 32'b00000000000000011011010000111110;
assign LUT_4[59265] = 32'b00000000000000010100011100110110;
assign LUT_4[59266] = 32'b00000000000000011010101011100010;
assign LUT_4[59267] = 32'b00000000000000010011110111011010;
assign LUT_4[59268] = 32'b00000000000000011000010001011010;
assign LUT_4[59269] = 32'b00000000000000010001011101010010;
assign LUT_4[59270] = 32'b00000000000000010111101011111110;
assign LUT_4[59271] = 32'b00000000000000010000110111110110;
assign LUT_4[59272] = 32'b00000000000000010100011101010011;
assign LUT_4[59273] = 32'b00000000000000001101101001001011;
assign LUT_4[59274] = 32'b00000000000000010011110111110111;
assign LUT_4[59275] = 32'b00000000000000001101000011101111;
assign LUT_4[59276] = 32'b00000000000000010001011101101111;
assign LUT_4[59277] = 32'b00000000000000001010101001100111;
assign LUT_4[59278] = 32'b00000000000000010000111000010011;
assign LUT_4[59279] = 32'b00000000000000001010000100001011;
assign LUT_4[59280] = 32'b00000000000000011001000010101100;
assign LUT_4[59281] = 32'b00000000000000010010001110100100;
assign LUT_4[59282] = 32'b00000000000000011000011101010000;
assign LUT_4[59283] = 32'b00000000000000010001101001001000;
assign LUT_4[59284] = 32'b00000000000000010110000011001000;
assign LUT_4[59285] = 32'b00000000000000001111001111000000;
assign LUT_4[59286] = 32'b00000000000000010101011101101100;
assign LUT_4[59287] = 32'b00000000000000001110101001100100;
assign LUT_4[59288] = 32'b00000000000000010010001111000001;
assign LUT_4[59289] = 32'b00000000000000001011011010111001;
assign LUT_4[59290] = 32'b00000000000000010001101001100101;
assign LUT_4[59291] = 32'b00000000000000001010110101011101;
assign LUT_4[59292] = 32'b00000000000000001111001111011101;
assign LUT_4[59293] = 32'b00000000000000001000011011010101;
assign LUT_4[59294] = 32'b00000000000000001110101010000001;
assign LUT_4[59295] = 32'b00000000000000000111110101111001;
assign LUT_4[59296] = 32'b00000000000000011001101100000101;
assign LUT_4[59297] = 32'b00000000000000010010110111111101;
assign LUT_4[59298] = 32'b00000000000000011001000110101001;
assign LUT_4[59299] = 32'b00000000000000010010010010100001;
assign LUT_4[59300] = 32'b00000000000000010110101100100001;
assign LUT_4[59301] = 32'b00000000000000001111111000011001;
assign LUT_4[59302] = 32'b00000000000000010110000111000101;
assign LUT_4[59303] = 32'b00000000000000001111010010111101;
assign LUT_4[59304] = 32'b00000000000000010010111000011010;
assign LUT_4[59305] = 32'b00000000000000001100000100010010;
assign LUT_4[59306] = 32'b00000000000000010010010010111110;
assign LUT_4[59307] = 32'b00000000000000001011011110110110;
assign LUT_4[59308] = 32'b00000000000000001111111000110110;
assign LUT_4[59309] = 32'b00000000000000001001000100101110;
assign LUT_4[59310] = 32'b00000000000000001111010011011010;
assign LUT_4[59311] = 32'b00000000000000001000011111010010;
assign LUT_4[59312] = 32'b00000000000000010111011101110011;
assign LUT_4[59313] = 32'b00000000000000010000101001101011;
assign LUT_4[59314] = 32'b00000000000000010110111000010111;
assign LUT_4[59315] = 32'b00000000000000010000000100001111;
assign LUT_4[59316] = 32'b00000000000000010100011110001111;
assign LUT_4[59317] = 32'b00000000000000001101101010000111;
assign LUT_4[59318] = 32'b00000000000000010011111000110011;
assign LUT_4[59319] = 32'b00000000000000001101000100101011;
assign LUT_4[59320] = 32'b00000000000000010000101010001000;
assign LUT_4[59321] = 32'b00000000000000001001110110000000;
assign LUT_4[59322] = 32'b00000000000000010000000100101100;
assign LUT_4[59323] = 32'b00000000000000001001010000100100;
assign LUT_4[59324] = 32'b00000000000000001101101010100100;
assign LUT_4[59325] = 32'b00000000000000000110110110011100;
assign LUT_4[59326] = 32'b00000000000000001101000101001000;
assign LUT_4[59327] = 32'b00000000000000000110010001000000;
assign LUT_4[59328] = 32'b00000000000000011100101000010010;
assign LUT_4[59329] = 32'b00000000000000010101110100001010;
assign LUT_4[59330] = 32'b00000000000000011100000010110110;
assign LUT_4[59331] = 32'b00000000000000010101001110101110;
assign LUT_4[59332] = 32'b00000000000000011001101000101110;
assign LUT_4[59333] = 32'b00000000000000010010110100100110;
assign LUT_4[59334] = 32'b00000000000000011001000011010010;
assign LUT_4[59335] = 32'b00000000000000010010001111001010;
assign LUT_4[59336] = 32'b00000000000000010101110100100111;
assign LUT_4[59337] = 32'b00000000000000001111000000011111;
assign LUT_4[59338] = 32'b00000000000000010101001111001011;
assign LUT_4[59339] = 32'b00000000000000001110011011000011;
assign LUT_4[59340] = 32'b00000000000000010010110101000011;
assign LUT_4[59341] = 32'b00000000000000001100000000111011;
assign LUT_4[59342] = 32'b00000000000000010010001111100111;
assign LUT_4[59343] = 32'b00000000000000001011011011011111;
assign LUT_4[59344] = 32'b00000000000000011010011010000000;
assign LUT_4[59345] = 32'b00000000000000010011100101111000;
assign LUT_4[59346] = 32'b00000000000000011001110100100100;
assign LUT_4[59347] = 32'b00000000000000010011000000011100;
assign LUT_4[59348] = 32'b00000000000000010111011010011100;
assign LUT_4[59349] = 32'b00000000000000010000100110010100;
assign LUT_4[59350] = 32'b00000000000000010110110101000000;
assign LUT_4[59351] = 32'b00000000000000010000000000111000;
assign LUT_4[59352] = 32'b00000000000000010011100110010101;
assign LUT_4[59353] = 32'b00000000000000001100110010001101;
assign LUT_4[59354] = 32'b00000000000000010011000000111001;
assign LUT_4[59355] = 32'b00000000000000001100001100110001;
assign LUT_4[59356] = 32'b00000000000000010000100110110001;
assign LUT_4[59357] = 32'b00000000000000001001110010101001;
assign LUT_4[59358] = 32'b00000000000000010000000001010101;
assign LUT_4[59359] = 32'b00000000000000001001001101001101;
assign LUT_4[59360] = 32'b00000000000000011011000011011001;
assign LUT_4[59361] = 32'b00000000000000010100001111010001;
assign LUT_4[59362] = 32'b00000000000000011010011101111101;
assign LUT_4[59363] = 32'b00000000000000010011101001110101;
assign LUT_4[59364] = 32'b00000000000000011000000011110101;
assign LUT_4[59365] = 32'b00000000000000010001001111101101;
assign LUT_4[59366] = 32'b00000000000000010111011110011001;
assign LUT_4[59367] = 32'b00000000000000010000101010010001;
assign LUT_4[59368] = 32'b00000000000000010100001111101110;
assign LUT_4[59369] = 32'b00000000000000001101011011100110;
assign LUT_4[59370] = 32'b00000000000000010011101010010010;
assign LUT_4[59371] = 32'b00000000000000001100110110001010;
assign LUT_4[59372] = 32'b00000000000000010001010000001010;
assign LUT_4[59373] = 32'b00000000000000001010011100000010;
assign LUT_4[59374] = 32'b00000000000000010000101010101110;
assign LUT_4[59375] = 32'b00000000000000001001110110100110;
assign LUT_4[59376] = 32'b00000000000000011000110101000111;
assign LUT_4[59377] = 32'b00000000000000010010000000111111;
assign LUT_4[59378] = 32'b00000000000000011000001111101011;
assign LUT_4[59379] = 32'b00000000000000010001011011100011;
assign LUT_4[59380] = 32'b00000000000000010101110101100011;
assign LUT_4[59381] = 32'b00000000000000001111000001011011;
assign LUT_4[59382] = 32'b00000000000000010101010000000111;
assign LUT_4[59383] = 32'b00000000000000001110011011111111;
assign LUT_4[59384] = 32'b00000000000000010010000001011100;
assign LUT_4[59385] = 32'b00000000000000001011001101010100;
assign LUT_4[59386] = 32'b00000000000000010001011100000000;
assign LUT_4[59387] = 32'b00000000000000001010100111111000;
assign LUT_4[59388] = 32'b00000000000000001111000001111000;
assign LUT_4[59389] = 32'b00000000000000001000001101110000;
assign LUT_4[59390] = 32'b00000000000000001110011100011100;
assign LUT_4[59391] = 32'b00000000000000000111101000010100;
assign LUT_4[59392] = 32'b00000000000000001110011111110110;
assign LUT_4[59393] = 32'b00000000000000000111101011101110;
assign LUT_4[59394] = 32'b00000000000000001101111010011010;
assign LUT_4[59395] = 32'b00000000000000000111000110010010;
assign LUT_4[59396] = 32'b00000000000000001011100000010010;
assign LUT_4[59397] = 32'b00000000000000000100101100001010;
assign LUT_4[59398] = 32'b00000000000000001010111010110110;
assign LUT_4[59399] = 32'b00000000000000000100000110101110;
assign LUT_4[59400] = 32'b00000000000000000111101100001011;
assign LUT_4[59401] = 32'b00000000000000000000111000000011;
assign LUT_4[59402] = 32'b00000000000000000111000110101111;
assign LUT_4[59403] = 32'b00000000000000000000010010100111;
assign LUT_4[59404] = 32'b00000000000000000100101100100111;
assign LUT_4[59405] = 32'b11111111111111111101111000011111;
assign LUT_4[59406] = 32'b00000000000000000100000111001011;
assign LUT_4[59407] = 32'b11111111111111111101010011000011;
assign LUT_4[59408] = 32'b00000000000000001100010001100100;
assign LUT_4[59409] = 32'b00000000000000000101011101011100;
assign LUT_4[59410] = 32'b00000000000000001011101100001000;
assign LUT_4[59411] = 32'b00000000000000000100111000000000;
assign LUT_4[59412] = 32'b00000000000000001001010010000000;
assign LUT_4[59413] = 32'b00000000000000000010011101111000;
assign LUT_4[59414] = 32'b00000000000000001000101100100100;
assign LUT_4[59415] = 32'b00000000000000000001111000011100;
assign LUT_4[59416] = 32'b00000000000000000101011101111001;
assign LUT_4[59417] = 32'b11111111111111111110101001110001;
assign LUT_4[59418] = 32'b00000000000000000100111000011101;
assign LUT_4[59419] = 32'b11111111111111111110000100010101;
assign LUT_4[59420] = 32'b00000000000000000010011110010101;
assign LUT_4[59421] = 32'b11111111111111111011101010001101;
assign LUT_4[59422] = 32'b00000000000000000001111000111001;
assign LUT_4[59423] = 32'b11111111111111111011000100110001;
assign LUT_4[59424] = 32'b00000000000000001100111010111101;
assign LUT_4[59425] = 32'b00000000000000000110000110110101;
assign LUT_4[59426] = 32'b00000000000000001100010101100001;
assign LUT_4[59427] = 32'b00000000000000000101100001011001;
assign LUT_4[59428] = 32'b00000000000000001001111011011001;
assign LUT_4[59429] = 32'b00000000000000000011000111010001;
assign LUT_4[59430] = 32'b00000000000000001001010101111101;
assign LUT_4[59431] = 32'b00000000000000000010100001110101;
assign LUT_4[59432] = 32'b00000000000000000110000111010010;
assign LUT_4[59433] = 32'b11111111111111111111010011001010;
assign LUT_4[59434] = 32'b00000000000000000101100001110110;
assign LUT_4[59435] = 32'b11111111111111111110101101101110;
assign LUT_4[59436] = 32'b00000000000000000011000111101110;
assign LUT_4[59437] = 32'b11111111111111111100010011100110;
assign LUT_4[59438] = 32'b00000000000000000010100010010010;
assign LUT_4[59439] = 32'b11111111111111111011101110001010;
assign LUT_4[59440] = 32'b00000000000000001010101100101011;
assign LUT_4[59441] = 32'b00000000000000000011111000100011;
assign LUT_4[59442] = 32'b00000000000000001010000111001111;
assign LUT_4[59443] = 32'b00000000000000000011010011000111;
assign LUT_4[59444] = 32'b00000000000000000111101101000111;
assign LUT_4[59445] = 32'b00000000000000000000111000111111;
assign LUT_4[59446] = 32'b00000000000000000111000111101011;
assign LUT_4[59447] = 32'b00000000000000000000010011100011;
assign LUT_4[59448] = 32'b00000000000000000011111001000000;
assign LUT_4[59449] = 32'b11111111111111111101000100111000;
assign LUT_4[59450] = 32'b00000000000000000011010011100100;
assign LUT_4[59451] = 32'b11111111111111111100011111011100;
assign LUT_4[59452] = 32'b00000000000000000000111001011100;
assign LUT_4[59453] = 32'b11111111111111111010000101010100;
assign LUT_4[59454] = 32'b00000000000000000000010100000000;
assign LUT_4[59455] = 32'b11111111111111111001011111111000;
assign LUT_4[59456] = 32'b00000000000000001111110111001010;
assign LUT_4[59457] = 32'b00000000000000001001000011000010;
assign LUT_4[59458] = 32'b00000000000000001111010001101110;
assign LUT_4[59459] = 32'b00000000000000001000011101100110;
assign LUT_4[59460] = 32'b00000000000000001100110111100110;
assign LUT_4[59461] = 32'b00000000000000000110000011011110;
assign LUT_4[59462] = 32'b00000000000000001100010010001010;
assign LUT_4[59463] = 32'b00000000000000000101011110000010;
assign LUT_4[59464] = 32'b00000000000000001001000011011111;
assign LUT_4[59465] = 32'b00000000000000000010001111010111;
assign LUT_4[59466] = 32'b00000000000000001000011110000011;
assign LUT_4[59467] = 32'b00000000000000000001101001111011;
assign LUT_4[59468] = 32'b00000000000000000110000011111011;
assign LUT_4[59469] = 32'b11111111111111111111001111110011;
assign LUT_4[59470] = 32'b00000000000000000101011110011111;
assign LUT_4[59471] = 32'b11111111111111111110101010010111;
assign LUT_4[59472] = 32'b00000000000000001101101000111000;
assign LUT_4[59473] = 32'b00000000000000000110110100110000;
assign LUT_4[59474] = 32'b00000000000000001101000011011100;
assign LUT_4[59475] = 32'b00000000000000000110001111010100;
assign LUT_4[59476] = 32'b00000000000000001010101001010100;
assign LUT_4[59477] = 32'b00000000000000000011110101001100;
assign LUT_4[59478] = 32'b00000000000000001010000011111000;
assign LUT_4[59479] = 32'b00000000000000000011001111110000;
assign LUT_4[59480] = 32'b00000000000000000110110101001101;
assign LUT_4[59481] = 32'b00000000000000000000000001000101;
assign LUT_4[59482] = 32'b00000000000000000110001111110001;
assign LUT_4[59483] = 32'b11111111111111111111011011101001;
assign LUT_4[59484] = 32'b00000000000000000011110101101001;
assign LUT_4[59485] = 32'b11111111111111111101000001100001;
assign LUT_4[59486] = 32'b00000000000000000011010000001101;
assign LUT_4[59487] = 32'b11111111111111111100011100000101;
assign LUT_4[59488] = 32'b00000000000000001110010010010001;
assign LUT_4[59489] = 32'b00000000000000000111011110001001;
assign LUT_4[59490] = 32'b00000000000000001101101100110101;
assign LUT_4[59491] = 32'b00000000000000000110111000101101;
assign LUT_4[59492] = 32'b00000000000000001011010010101101;
assign LUT_4[59493] = 32'b00000000000000000100011110100101;
assign LUT_4[59494] = 32'b00000000000000001010101101010001;
assign LUT_4[59495] = 32'b00000000000000000011111001001001;
assign LUT_4[59496] = 32'b00000000000000000111011110100110;
assign LUT_4[59497] = 32'b00000000000000000000101010011110;
assign LUT_4[59498] = 32'b00000000000000000110111001001010;
assign LUT_4[59499] = 32'b00000000000000000000000101000010;
assign LUT_4[59500] = 32'b00000000000000000100011111000010;
assign LUT_4[59501] = 32'b11111111111111111101101010111010;
assign LUT_4[59502] = 32'b00000000000000000011111001100110;
assign LUT_4[59503] = 32'b11111111111111111101000101011110;
assign LUT_4[59504] = 32'b00000000000000001100000011111111;
assign LUT_4[59505] = 32'b00000000000000000101001111110111;
assign LUT_4[59506] = 32'b00000000000000001011011110100011;
assign LUT_4[59507] = 32'b00000000000000000100101010011011;
assign LUT_4[59508] = 32'b00000000000000001001000100011011;
assign LUT_4[59509] = 32'b00000000000000000010010000010011;
assign LUT_4[59510] = 32'b00000000000000001000011110111111;
assign LUT_4[59511] = 32'b00000000000000000001101010110111;
assign LUT_4[59512] = 32'b00000000000000000101010000010100;
assign LUT_4[59513] = 32'b11111111111111111110011100001100;
assign LUT_4[59514] = 32'b00000000000000000100101010111000;
assign LUT_4[59515] = 32'b11111111111111111101110110110000;
assign LUT_4[59516] = 32'b00000000000000000010010000110000;
assign LUT_4[59517] = 32'b11111111111111111011011100101000;
assign LUT_4[59518] = 32'b00000000000000000001101011010100;
assign LUT_4[59519] = 32'b11111111111111111010110111001100;
assign LUT_4[59520] = 32'b00000000000000010001000101111110;
assign LUT_4[59521] = 32'b00000000000000001010010001110110;
assign LUT_4[59522] = 32'b00000000000000010000100000100010;
assign LUT_4[59523] = 32'b00000000000000001001101100011010;
assign LUT_4[59524] = 32'b00000000000000001110000110011010;
assign LUT_4[59525] = 32'b00000000000000000111010010010010;
assign LUT_4[59526] = 32'b00000000000000001101100000111110;
assign LUT_4[59527] = 32'b00000000000000000110101100110110;
assign LUT_4[59528] = 32'b00000000000000001010010010010011;
assign LUT_4[59529] = 32'b00000000000000000011011110001011;
assign LUT_4[59530] = 32'b00000000000000001001101100110111;
assign LUT_4[59531] = 32'b00000000000000000010111000101111;
assign LUT_4[59532] = 32'b00000000000000000111010010101111;
assign LUT_4[59533] = 32'b00000000000000000000011110100111;
assign LUT_4[59534] = 32'b00000000000000000110101101010011;
assign LUT_4[59535] = 32'b11111111111111111111111001001011;
assign LUT_4[59536] = 32'b00000000000000001110110111101100;
assign LUT_4[59537] = 32'b00000000000000001000000011100100;
assign LUT_4[59538] = 32'b00000000000000001110010010010000;
assign LUT_4[59539] = 32'b00000000000000000111011110001000;
assign LUT_4[59540] = 32'b00000000000000001011111000001000;
assign LUT_4[59541] = 32'b00000000000000000101000100000000;
assign LUT_4[59542] = 32'b00000000000000001011010010101100;
assign LUT_4[59543] = 32'b00000000000000000100011110100100;
assign LUT_4[59544] = 32'b00000000000000001000000100000001;
assign LUT_4[59545] = 32'b00000000000000000001001111111001;
assign LUT_4[59546] = 32'b00000000000000000111011110100101;
assign LUT_4[59547] = 32'b00000000000000000000101010011101;
assign LUT_4[59548] = 32'b00000000000000000101000100011101;
assign LUT_4[59549] = 32'b11111111111111111110010000010101;
assign LUT_4[59550] = 32'b00000000000000000100011111000001;
assign LUT_4[59551] = 32'b11111111111111111101101010111001;
assign LUT_4[59552] = 32'b00000000000000001111100001000101;
assign LUT_4[59553] = 32'b00000000000000001000101100111101;
assign LUT_4[59554] = 32'b00000000000000001110111011101001;
assign LUT_4[59555] = 32'b00000000000000001000000111100001;
assign LUT_4[59556] = 32'b00000000000000001100100001100001;
assign LUT_4[59557] = 32'b00000000000000000101101101011001;
assign LUT_4[59558] = 32'b00000000000000001011111100000101;
assign LUT_4[59559] = 32'b00000000000000000101000111111101;
assign LUT_4[59560] = 32'b00000000000000001000101101011010;
assign LUT_4[59561] = 32'b00000000000000000001111001010010;
assign LUT_4[59562] = 32'b00000000000000001000000111111110;
assign LUT_4[59563] = 32'b00000000000000000001010011110110;
assign LUT_4[59564] = 32'b00000000000000000101101101110110;
assign LUT_4[59565] = 32'b11111111111111111110111001101110;
assign LUT_4[59566] = 32'b00000000000000000101001000011010;
assign LUT_4[59567] = 32'b11111111111111111110010100010010;
assign LUT_4[59568] = 32'b00000000000000001101010010110011;
assign LUT_4[59569] = 32'b00000000000000000110011110101011;
assign LUT_4[59570] = 32'b00000000000000001100101101010111;
assign LUT_4[59571] = 32'b00000000000000000101111001001111;
assign LUT_4[59572] = 32'b00000000000000001010010011001111;
assign LUT_4[59573] = 32'b00000000000000000011011111000111;
assign LUT_4[59574] = 32'b00000000000000001001101101110011;
assign LUT_4[59575] = 32'b00000000000000000010111001101011;
assign LUT_4[59576] = 32'b00000000000000000110011111001000;
assign LUT_4[59577] = 32'b11111111111111111111101011000000;
assign LUT_4[59578] = 32'b00000000000000000101111001101100;
assign LUT_4[59579] = 32'b11111111111111111111000101100100;
assign LUT_4[59580] = 32'b00000000000000000011011111100100;
assign LUT_4[59581] = 32'b11111111111111111100101011011100;
assign LUT_4[59582] = 32'b00000000000000000010111010001000;
assign LUT_4[59583] = 32'b11111111111111111100000110000000;
assign LUT_4[59584] = 32'b00000000000000010010011101010010;
assign LUT_4[59585] = 32'b00000000000000001011101001001010;
assign LUT_4[59586] = 32'b00000000000000010001110111110110;
assign LUT_4[59587] = 32'b00000000000000001011000011101110;
assign LUT_4[59588] = 32'b00000000000000001111011101101110;
assign LUT_4[59589] = 32'b00000000000000001000101001100110;
assign LUT_4[59590] = 32'b00000000000000001110111000010010;
assign LUT_4[59591] = 32'b00000000000000001000000100001010;
assign LUT_4[59592] = 32'b00000000000000001011101001100111;
assign LUT_4[59593] = 32'b00000000000000000100110101011111;
assign LUT_4[59594] = 32'b00000000000000001011000100001011;
assign LUT_4[59595] = 32'b00000000000000000100010000000011;
assign LUT_4[59596] = 32'b00000000000000001000101010000011;
assign LUT_4[59597] = 32'b00000000000000000001110101111011;
assign LUT_4[59598] = 32'b00000000000000001000000100100111;
assign LUT_4[59599] = 32'b00000000000000000001010000011111;
assign LUT_4[59600] = 32'b00000000000000010000001111000000;
assign LUT_4[59601] = 32'b00000000000000001001011010111000;
assign LUT_4[59602] = 32'b00000000000000001111101001100100;
assign LUT_4[59603] = 32'b00000000000000001000110101011100;
assign LUT_4[59604] = 32'b00000000000000001101001111011100;
assign LUT_4[59605] = 32'b00000000000000000110011011010100;
assign LUT_4[59606] = 32'b00000000000000001100101010000000;
assign LUT_4[59607] = 32'b00000000000000000101110101111000;
assign LUT_4[59608] = 32'b00000000000000001001011011010101;
assign LUT_4[59609] = 32'b00000000000000000010100111001101;
assign LUT_4[59610] = 32'b00000000000000001000110101111001;
assign LUT_4[59611] = 32'b00000000000000000010000001110001;
assign LUT_4[59612] = 32'b00000000000000000110011011110001;
assign LUT_4[59613] = 32'b11111111111111111111100111101001;
assign LUT_4[59614] = 32'b00000000000000000101110110010101;
assign LUT_4[59615] = 32'b11111111111111111111000010001101;
assign LUT_4[59616] = 32'b00000000000000010000111000011001;
assign LUT_4[59617] = 32'b00000000000000001010000100010001;
assign LUT_4[59618] = 32'b00000000000000010000010010111101;
assign LUT_4[59619] = 32'b00000000000000001001011110110101;
assign LUT_4[59620] = 32'b00000000000000001101111000110101;
assign LUT_4[59621] = 32'b00000000000000000111000100101101;
assign LUT_4[59622] = 32'b00000000000000001101010011011001;
assign LUT_4[59623] = 32'b00000000000000000110011111010001;
assign LUT_4[59624] = 32'b00000000000000001010000100101110;
assign LUT_4[59625] = 32'b00000000000000000011010000100110;
assign LUT_4[59626] = 32'b00000000000000001001011111010010;
assign LUT_4[59627] = 32'b00000000000000000010101011001010;
assign LUT_4[59628] = 32'b00000000000000000111000101001010;
assign LUT_4[59629] = 32'b00000000000000000000010001000010;
assign LUT_4[59630] = 32'b00000000000000000110011111101110;
assign LUT_4[59631] = 32'b11111111111111111111101011100110;
assign LUT_4[59632] = 32'b00000000000000001110101010000111;
assign LUT_4[59633] = 32'b00000000000000000111110101111111;
assign LUT_4[59634] = 32'b00000000000000001110000100101011;
assign LUT_4[59635] = 32'b00000000000000000111010000100011;
assign LUT_4[59636] = 32'b00000000000000001011101010100011;
assign LUT_4[59637] = 32'b00000000000000000100110110011011;
assign LUT_4[59638] = 32'b00000000000000001011000101000111;
assign LUT_4[59639] = 32'b00000000000000000100010000111111;
assign LUT_4[59640] = 32'b00000000000000000111110110011100;
assign LUT_4[59641] = 32'b00000000000000000001000010010100;
assign LUT_4[59642] = 32'b00000000000000000111010001000000;
assign LUT_4[59643] = 32'b00000000000000000000011100111000;
assign LUT_4[59644] = 32'b00000000000000000100110110111000;
assign LUT_4[59645] = 32'b11111111111111111110000010110000;
assign LUT_4[59646] = 32'b00000000000000000100010001011100;
assign LUT_4[59647] = 32'b11111111111111111101011101010100;
assign LUT_4[59648] = 32'b00000000000000010011011011011001;
assign LUT_4[59649] = 32'b00000000000000001100100111010001;
assign LUT_4[59650] = 32'b00000000000000010010110101111101;
assign LUT_4[59651] = 32'b00000000000000001100000001110101;
assign LUT_4[59652] = 32'b00000000000000010000011011110101;
assign LUT_4[59653] = 32'b00000000000000001001100111101101;
assign LUT_4[59654] = 32'b00000000000000001111110110011001;
assign LUT_4[59655] = 32'b00000000000000001001000010010001;
assign LUT_4[59656] = 32'b00000000000000001100100111101110;
assign LUT_4[59657] = 32'b00000000000000000101110011100110;
assign LUT_4[59658] = 32'b00000000000000001100000010010010;
assign LUT_4[59659] = 32'b00000000000000000101001110001010;
assign LUT_4[59660] = 32'b00000000000000001001101000001010;
assign LUT_4[59661] = 32'b00000000000000000010110100000010;
assign LUT_4[59662] = 32'b00000000000000001001000010101110;
assign LUT_4[59663] = 32'b00000000000000000010001110100110;
assign LUT_4[59664] = 32'b00000000000000010001001101000111;
assign LUT_4[59665] = 32'b00000000000000001010011000111111;
assign LUT_4[59666] = 32'b00000000000000010000100111101011;
assign LUT_4[59667] = 32'b00000000000000001001110011100011;
assign LUT_4[59668] = 32'b00000000000000001110001101100011;
assign LUT_4[59669] = 32'b00000000000000000111011001011011;
assign LUT_4[59670] = 32'b00000000000000001101101000000111;
assign LUT_4[59671] = 32'b00000000000000000110110011111111;
assign LUT_4[59672] = 32'b00000000000000001010011001011100;
assign LUT_4[59673] = 32'b00000000000000000011100101010100;
assign LUT_4[59674] = 32'b00000000000000001001110100000000;
assign LUT_4[59675] = 32'b00000000000000000010111111111000;
assign LUT_4[59676] = 32'b00000000000000000111011001111000;
assign LUT_4[59677] = 32'b00000000000000000000100101110000;
assign LUT_4[59678] = 32'b00000000000000000110110100011100;
assign LUT_4[59679] = 32'b00000000000000000000000000010100;
assign LUT_4[59680] = 32'b00000000000000010001110110100000;
assign LUT_4[59681] = 32'b00000000000000001011000010011000;
assign LUT_4[59682] = 32'b00000000000000010001010001000100;
assign LUT_4[59683] = 32'b00000000000000001010011100111100;
assign LUT_4[59684] = 32'b00000000000000001110110110111100;
assign LUT_4[59685] = 32'b00000000000000001000000010110100;
assign LUT_4[59686] = 32'b00000000000000001110010001100000;
assign LUT_4[59687] = 32'b00000000000000000111011101011000;
assign LUT_4[59688] = 32'b00000000000000001011000010110101;
assign LUT_4[59689] = 32'b00000000000000000100001110101101;
assign LUT_4[59690] = 32'b00000000000000001010011101011001;
assign LUT_4[59691] = 32'b00000000000000000011101001010001;
assign LUT_4[59692] = 32'b00000000000000001000000011010001;
assign LUT_4[59693] = 32'b00000000000000000001001111001001;
assign LUT_4[59694] = 32'b00000000000000000111011101110101;
assign LUT_4[59695] = 32'b00000000000000000000101001101101;
assign LUT_4[59696] = 32'b00000000000000001111101000001110;
assign LUT_4[59697] = 32'b00000000000000001000110100000110;
assign LUT_4[59698] = 32'b00000000000000001111000010110010;
assign LUT_4[59699] = 32'b00000000000000001000001110101010;
assign LUT_4[59700] = 32'b00000000000000001100101000101010;
assign LUT_4[59701] = 32'b00000000000000000101110100100010;
assign LUT_4[59702] = 32'b00000000000000001100000011001110;
assign LUT_4[59703] = 32'b00000000000000000101001111000110;
assign LUT_4[59704] = 32'b00000000000000001000110100100011;
assign LUT_4[59705] = 32'b00000000000000000010000000011011;
assign LUT_4[59706] = 32'b00000000000000001000001111000111;
assign LUT_4[59707] = 32'b00000000000000000001011010111111;
assign LUT_4[59708] = 32'b00000000000000000101110100111111;
assign LUT_4[59709] = 32'b11111111111111111111000000110111;
assign LUT_4[59710] = 32'b00000000000000000101001111100011;
assign LUT_4[59711] = 32'b11111111111111111110011011011011;
assign LUT_4[59712] = 32'b00000000000000010100110010101101;
assign LUT_4[59713] = 32'b00000000000000001101111110100101;
assign LUT_4[59714] = 32'b00000000000000010100001101010001;
assign LUT_4[59715] = 32'b00000000000000001101011001001001;
assign LUT_4[59716] = 32'b00000000000000010001110011001001;
assign LUT_4[59717] = 32'b00000000000000001010111111000001;
assign LUT_4[59718] = 32'b00000000000000010001001101101101;
assign LUT_4[59719] = 32'b00000000000000001010011001100101;
assign LUT_4[59720] = 32'b00000000000000001101111111000010;
assign LUT_4[59721] = 32'b00000000000000000111001010111010;
assign LUT_4[59722] = 32'b00000000000000001101011001100110;
assign LUT_4[59723] = 32'b00000000000000000110100101011110;
assign LUT_4[59724] = 32'b00000000000000001010111111011110;
assign LUT_4[59725] = 32'b00000000000000000100001011010110;
assign LUT_4[59726] = 32'b00000000000000001010011010000010;
assign LUT_4[59727] = 32'b00000000000000000011100101111010;
assign LUT_4[59728] = 32'b00000000000000010010100100011011;
assign LUT_4[59729] = 32'b00000000000000001011110000010011;
assign LUT_4[59730] = 32'b00000000000000010001111110111111;
assign LUT_4[59731] = 32'b00000000000000001011001010110111;
assign LUT_4[59732] = 32'b00000000000000001111100100110111;
assign LUT_4[59733] = 32'b00000000000000001000110000101111;
assign LUT_4[59734] = 32'b00000000000000001110111111011011;
assign LUT_4[59735] = 32'b00000000000000001000001011010011;
assign LUT_4[59736] = 32'b00000000000000001011110000110000;
assign LUT_4[59737] = 32'b00000000000000000100111100101000;
assign LUT_4[59738] = 32'b00000000000000001011001011010100;
assign LUT_4[59739] = 32'b00000000000000000100010111001100;
assign LUT_4[59740] = 32'b00000000000000001000110001001100;
assign LUT_4[59741] = 32'b00000000000000000001111101000100;
assign LUT_4[59742] = 32'b00000000000000001000001011110000;
assign LUT_4[59743] = 32'b00000000000000000001010111101000;
assign LUT_4[59744] = 32'b00000000000000010011001101110100;
assign LUT_4[59745] = 32'b00000000000000001100011001101100;
assign LUT_4[59746] = 32'b00000000000000010010101000011000;
assign LUT_4[59747] = 32'b00000000000000001011110100010000;
assign LUT_4[59748] = 32'b00000000000000010000001110010000;
assign LUT_4[59749] = 32'b00000000000000001001011010001000;
assign LUT_4[59750] = 32'b00000000000000001111101000110100;
assign LUT_4[59751] = 32'b00000000000000001000110100101100;
assign LUT_4[59752] = 32'b00000000000000001100011010001001;
assign LUT_4[59753] = 32'b00000000000000000101100110000001;
assign LUT_4[59754] = 32'b00000000000000001011110100101101;
assign LUT_4[59755] = 32'b00000000000000000101000000100101;
assign LUT_4[59756] = 32'b00000000000000001001011010100101;
assign LUT_4[59757] = 32'b00000000000000000010100110011101;
assign LUT_4[59758] = 32'b00000000000000001000110101001001;
assign LUT_4[59759] = 32'b00000000000000000010000001000001;
assign LUT_4[59760] = 32'b00000000000000010000111111100010;
assign LUT_4[59761] = 32'b00000000000000001010001011011010;
assign LUT_4[59762] = 32'b00000000000000010000011010000110;
assign LUT_4[59763] = 32'b00000000000000001001100101111110;
assign LUT_4[59764] = 32'b00000000000000001101111111111110;
assign LUT_4[59765] = 32'b00000000000000000111001011110110;
assign LUT_4[59766] = 32'b00000000000000001101011010100010;
assign LUT_4[59767] = 32'b00000000000000000110100110011010;
assign LUT_4[59768] = 32'b00000000000000001010001011110111;
assign LUT_4[59769] = 32'b00000000000000000011010111101111;
assign LUT_4[59770] = 32'b00000000000000001001100110011011;
assign LUT_4[59771] = 32'b00000000000000000010110010010011;
assign LUT_4[59772] = 32'b00000000000000000111001100010011;
assign LUT_4[59773] = 32'b00000000000000000000011000001011;
assign LUT_4[59774] = 32'b00000000000000000110100110110111;
assign LUT_4[59775] = 32'b11111111111111111111110010101111;
assign LUT_4[59776] = 32'b00000000000000010110000001100001;
assign LUT_4[59777] = 32'b00000000000000001111001101011001;
assign LUT_4[59778] = 32'b00000000000000010101011100000101;
assign LUT_4[59779] = 32'b00000000000000001110100111111101;
assign LUT_4[59780] = 32'b00000000000000010011000001111101;
assign LUT_4[59781] = 32'b00000000000000001100001101110101;
assign LUT_4[59782] = 32'b00000000000000010010011100100001;
assign LUT_4[59783] = 32'b00000000000000001011101000011001;
assign LUT_4[59784] = 32'b00000000000000001111001101110110;
assign LUT_4[59785] = 32'b00000000000000001000011001101110;
assign LUT_4[59786] = 32'b00000000000000001110101000011010;
assign LUT_4[59787] = 32'b00000000000000000111110100010010;
assign LUT_4[59788] = 32'b00000000000000001100001110010010;
assign LUT_4[59789] = 32'b00000000000000000101011010001010;
assign LUT_4[59790] = 32'b00000000000000001011101000110110;
assign LUT_4[59791] = 32'b00000000000000000100110100101110;
assign LUT_4[59792] = 32'b00000000000000010011110011001111;
assign LUT_4[59793] = 32'b00000000000000001100111111000111;
assign LUT_4[59794] = 32'b00000000000000010011001101110011;
assign LUT_4[59795] = 32'b00000000000000001100011001101011;
assign LUT_4[59796] = 32'b00000000000000010000110011101011;
assign LUT_4[59797] = 32'b00000000000000001001111111100011;
assign LUT_4[59798] = 32'b00000000000000010000001110001111;
assign LUT_4[59799] = 32'b00000000000000001001011010000111;
assign LUT_4[59800] = 32'b00000000000000001100111111100100;
assign LUT_4[59801] = 32'b00000000000000000110001011011100;
assign LUT_4[59802] = 32'b00000000000000001100011010001000;
assign LUT_4[59803] = 32'b00000000000000000101100110000000;
assign LUT_4[59804] = 32'b00000000000000001010000000000000;
assign LUT_4[59805] = 32'b00000000000000000011001011111000;
assign LUT_4[59806] = 32'b00000000000000001001011010100100;
assign LUT_4[59807] = 32'b00000000000000000010100110011100;
assign LUT_4[59808] = 32'b00000000000000010100011100101000;
assign LUT_4[59809] = 32'b00000000000000001101101000100000;
assign LUT_4[59810] = 32'b00000000000000010011110111001100;
assign LUT_4[59811] = 32'b00000000000000001101000011000100;
assign LUT_4[59812] = 32'b00000000000000010001011101000100;
assign LUT_4[59813] = 32'b00000000000000001010101000111100;
assign LUT_4[59814] = 32'b00000000000000010000110111101000;
assign LUT_4[59815] = 32'b00000000000000001010000011100000;
assign LUT_4[59816] = 32'b00000000000000001101101000111101;
assign LUT_4[59817] = 32'b00000000000000000110110100110101;
assign LUT_4[59818] = 32'b00000000000000001101000011100001;
assign LUT_4[59819] = 32'b00000000000000000110001111011001;
assign LUT_4[59820] = 32'b00000000000000001010101001011001;
assign LUT_4[59821] = 32'b00000000000000000011110101010001;
assign LUT_4[59822] = 32'b00000000000000001010000011111101;
assign LUT_4[59823] = 32'b00000000000000000011001111110101;
assign LUT_4[59824] = 32'b00000000000000010010001110010110;
assign LUT_4[59825] = 32'b00000000000000001011011010001110;
assign LUT_4[59826] = 32'b00000000000000010001101000111010;
assign LUT_4[59827] = 32'b00000000000000001010110100110010;
assign LUT_4[59828] = 32'b00000000000000001111001110110010;
assign LUT_4[59829] = 32'b00000000000000001000011010101010;
assign LUT_4[59830] = 32'b00000000000000001110101001010110;
assign LUT_4[59831] = 32'b00000000000000000111110101001110;
assign LUT_4[59832] = 32'b00000000000000001011011010101011;
assign LUT_4[59833] = 32'b00000000000000000100100110100011;
assign LUT_4[59834] = 32'b00000000000000001010110101001111;
assign LUT_4[59835] = 32'b00000000000000000100000001000111;
assign LUT_4[59836] = 32'b00000000000000001000011011000111;
assign LUT_4[59837] = 32'b00000000000000000001100110111111;
assign LUT_4[59838] = 32'b00000000000000000111110101101011;
assign LUT_4[59839] = 32'b00000000000000000001000001100011;
assign LUT_4[59840] = 32'b00000000000000010111011000110101;
assign LUT_4[59841] = 32'b00000000000000010000100100101101;
assign LUT_4[59842] = 32'b00000000000000010110110011011001;
assign LUT_4[59843] = 32'b00000000000000001111111111010001;
assign LUT_4[59844] = 32'b00000000000000010100011001010001;
assign LUT_4[59845] = 32'b00000000000000001101100101001001;
assign LUT_4[59846] = 32'b00000000000000010011110011110101;
assign LUT_4[59847] = 32'b00000000000000001100111111101101;
assign LUT_4[59848] = 32'b00000000000000010000100101001010;
assign LUT_4[59849] = 32'b00000000000000001001110001000010;
assign LUT_4[59850] = 32'b00000000000000001111111111101110;
assign LUT_4[59851] = 32'b00000000000000001001001011100110;
assign LUT_4[59852] = 32'b00000000000000001101100101100110;
assign LUT_4[59853] = 32'b00000000000000000110110001011110;
assign LUT_4[59854] = 32'b00000000000000001101000000001010;
assign LUT_4[59855] = 32'b00000000000000000110001100000010;
assign LUT_4[59856] = 32'b00000000000000010101001010100011;
assign LUT_4[59857] = 32'b00000000000000001110010110011011;
assign LUT_4[59858] = 32'b00000000000000010100100101000111;
assign LUT_4[59859] = 32'b00000000000000001101110000111111;
assign LUT_4[59860] = 32'b00000000000000010010001010111111;
assign LUT_4[59861] = 32'b00000000000000001011010110110111;
assign LUT_4[59862] = 32'b00000000000000010001100101100011;
assign LUT_4[59863] = 32'b00000000000000001010110001011011;
assign LUT_4[59864] = 32'b00000000000000001110010110111000;
assign LUT_4[59865] = 32'b00000000000000000111100010110000;
assign LUT_4[59866] = 32'b00000000000000001101110001011100;
assign LUT_4[59867] = 32'b00000000000000000110111101010100;
assign LUT_4[59868] = 32'b00000000000000001011010111010100;
assign LUT_4[59869] = 32'b00000000000000000100100011001100;
assign LUT_4[59870] = 32'b00000000000000001010110001111000;
assign LUT_4[59871] = 32'b00000000000000000011111101110000;
assign LUT_4[59872] = 32'b00000000000000010101110011111100;
assign LUT_4[59873] = 32'b00000000000000001110111111110100;
assign LUT_4[59874] = 32'b00000000000000010101001110100000;
assign LUT_4[59875] = 32'b00000000000000001110011010011000;
assign LUT_4[59876] = 32'b00000000000000010010110100011000;
assign LUT_4[59877] = 32'b00000000000000001100000000010000;
assign LUT_4[59878] = 32'b00000000000000010010001110111100;
assign LUT_4[59879] = 32'b00000000000000001011011010110100;
assign LUT_4[59880] = 32'b00000000000000001111000000010001;
assign LUT_4[59881] = 32'b00000000000000001000001100001001;
assign LUT_4[59882] = 32'b00000000000000001110011010110101;
assign LUT_4[59883] = 32'b00000000000000000111100110101101;
assign LUT_4[59884] = 32'b00000000000000001100000000101101;
assign LUT_4[59885] = 32'b00000000000000000101001100100101;
assign LUT_4[59886] = 32'b00000000000000001011011011010001;
assign LUT_4[59887] = 32'b00000000000000000100100111001001;
assign LUT_4[59888] = 32'b00000000000000010011100101101010;
assign LUT_4[59889] = 32'b00000000000000001100110001100010;
assign LUT_4[59890] = 32'b00000000000000010011000000001110;
assign LUT_4[59891] = 32'b00000000000000001100001100000110;
assign LUT_4[59892] = 32'b00000000000000010000100110000110;
assign LUT_4[59893] = 32'b00000000000000001001110001111110;
assign LUT_4[59894] = 32'b00000000000000010000000000101010;
assign LUT_4[59895] = 32'b00000000000000001001001100100010;
assign LUT_4[59896] = 32'b00000000000000001100110001111111;
assign LUT_4[59897] = 32'b00000000000000000101111101110111;
assign LUT_4[59898] = 32'b00000000000000001100001100100011;
assign LUT_4[59899] = 32'b00000000000000000101011000011011;
assign LUT_4[59900] = 32'b00000000000000001001110010011011;
assign LUT_4[59901] = 32'b00000000000000000010111110010011;
assign LUT_4[59902] = 32'b00000000000000001001001100111111;
assign LUT_4[59903] = 32'b00000000000000000010011000110111;
assign LUT_4[59904] = 32'b00000000000000001101100011111110;
assign LUT_4[59905] = 32'b00000000000000000110101111110110;
assign LUT_4[59906] = 32'b00000000000000001100111110100010;
assign LUT_4[59907] = 32'b00000000000000000110001010011010;
assign LUT_4[59908] = 32'b00000000000000001010100100011010;
assign LUT_4[59909] = 32'b00000000000000000011110000010010;
assign LUT_4[59910] = 32'b00000000000000001001111110111110;
assign LUT_4[59911] = 32'b00000000000000000011001010110110;
assign LUT_4[59912] = 32'b00000000000000000110110000010011;
assign LUT_4[59913] = 32'b11111111111111111111111100001011;
assign LUT_4[59914] = 32'b00000000000000000110001010110111;
assign LUT_4[59915] = 32'b11111111111111111111010110101111;
assign LUT_4[59916] = 32'b00000000000000000011110000101111;
assign LUT_4[59917] = 32'b11111111111111111100111100100111;
assign LUT_4[59918] = 32'b00000000000000000011001011010011;
assign LUT_4[59919] = 32'b11111111111111111100010111001011;
assign LUT_4[59920] = 32'b00000000000000001011010101101100;
assign LUT_4[59921] = 32'b00000000000000000100100001100100;
assign LUT_4[59922] = 32'b00000000000000001010110000010000;
assign LUT_4[59923] = 32'b00000000000000000011111100001000;
assign LUT_4[59924] = 32'b00000000000000001000010110001000;
assign LUT_4[59925] = 32'b00000000000000000001100010000000;
assign LUT_4[59926] = 32'b00000000000000000111110000101100;
assign LUT_4[59927] = 32'b00000000000000000000111100100100;
assign LUT_4[59928] = 32'b00000000000000000100100010000001;
assign LUT_4[59929] = 32'b11111111111111111101101101111001;
assign LUT_4[59930] = 32'b00000000000000000011111100100101;
assign LUT_4[59931] = 32'b11111111111111111101001000011101;
assign LUT_4[59932] = 32'b00000000000000000001100010011101;
assign LUT_4[59933] = 32'b11111111111111111010101110010101;
assign LUT_4[59934] = 32'b00000000000000000000111101000001;
assign LUT_4[59935] = 32'b11111111111111111010001000111001;
assign LUT_4[59936] = 32'b00000000000000001011111111000101;
assign LUT_4[59937] = 32'b00000000000000000101001010111101;
assign LUT_4[59938] = 32'b00000000000000001011011001101001;
assign LUT_4[59939] = 32'b00000000000000000100100101100001;
assign LUT_4[59940] = 32'b00000000000000001000111111100001;
assign LUT_4[59941] = 32'b00000000000000000010001011011001;
assign LUT_4[59942] = 32'b00000000000000001000011010000101;
assign LUT_4[59943] = 32'b00000000000000000001100101111101;
assign LUT_4[59944] = 32'b00000000000000000101001011011010;
assign LUT_4[59945] = 32'b11111111111111111110010111010010;
assign LUT_4[59946] = 32'b00000000000000000100100101111110;
assign LUT_4[59947] = 32'b11111111111111111101110001110110;
assign LUT_4[59948] = 32'b00000000000000000010001011110110;
assign LUT_4[59949] = 32'b11111111111111111011010111101110;
assign LUT_4[59950] = 32'b00000000000000000001100110011010;
assign LUT_4[59951] = 32'b11111111111111111010110010010010;
assign LUT_4[59952] = 32'b00000000000000001001110000110011;
assign LUT_4[59953] = 32'b00000000000000000010111100101011;
assign LUT_4[59954] = 32'b00000000000000001001001011010111;
assign LUT_4[59955] = 32'b00000000000000000010010111001111;
assign LUT_4[59956] = 32'b00000000000000000110110001001111;
assign LUT_4[59957] = 32'b11111111111111111111111101000111;
assign LUT_4[59958] = 32'b00000000000000000110001011110011;
assign LUT_4[59959] = 32'b11111111111111111111010111101011;
assign LUT_4[59960] = 32'b00000000000000000010111101001000;
assign LUT_4[59961] = 32'b11111111111111111100001001000000;
assign LUT_4[59962] = 32'b00000000000000000010010111101100;
assign LUT_4[59963] = 32'b11111111111111111011100011100100;
assign LUT_4[59964] = 32'b11111111111111111111111101100100;
assign LUT_4[59965] = 32'b11111111111111111001001001011100;
assign LUT_4[59966] = 32'b11111111111111111111011000001000;
assign LUT_4[59967] = 32'b11111111111111111000100100000000;
assign LUT_4[59968] = 32'b00000000000000001110111011010010;
assign LUT_4[59969] = 32'b00000000000000001000000111001010;
assign LUT_4[59970] = 32'b00000000000000001110010101110110;
assign LUT_4[59971] = 32'b00000000000000000111100001101110;
assign LUT_4[59972] = 32'b00000000000000001011111011101110;
assign LUT_4[59973] = 32'b00000000000000000101000111100110;
assign LUT_4[59974] = 32'b00000000000000001011010110010010;
assign LUT_4[59975] = 32'b00000000000000000100100010001010;
assign LUT_4[59976] = 32'b00000000000000001000000111100111;
assign LUT_4[59977] = 32'b00000000000000000001010011011111;
assign LUT_4[59978] = 32'b00000000000000000111100010001011;
assign LUT_4[59979] = 32'b00000000000000000000101110000011;
assign LUT_4[59980] = 32'b00000000000000000101001000000011;
assign LUT_4[59981] = 32'b11111111111111111110010011111011;
assign LUT_4[59982] = 32'b00000000000000000100100010100111;
assign LUT_4[59983] = 32'b11111111111111111101101110011111;
assign LUT_4[59984] = 32'b00000000000000001100101101000000;
assign LUT_4[59985] = 32'b00000000000000000101111000111000;
assign LUT_4[59986] = 32'b00000000000000001100000111100100;
assign LUT_4[59987] = 32'b00000000000000000101010011011100;
assign LUT_4[59988] = 32'b00000000000000001001101101011100;
assign LUT_4[59989] = 32'b00000000000000000010111001010100;
assign LUT_4[59990] = 32'b00000000000000001001001000000000;
assign LUT_4[59991] = 32'b00000000000000000010010011111000;
assign LUT_4[59992] = 32'b00000000000000000101111001010101;
assign LUT_4[59993] = 32'b11111111111111111111000101001101;
assign LUT_4[59994] = 32'b00000000000000000101010011111001;
assign LUT_4[59995] = 32'b11111111111111111110011111110001;
assign LUT_4[59996] = 32'b00000000000000000010111001110001;
assign LUT_4[59997] = 32'b11111111111111111100000101101001;
assign LUT_4[59998] = 32'b00000000000000000010010100010101;
assign LUT_4[59999] = 32'b11111111111111111011100000001101;
assign LUT_4[60000] = 32'b00000000000000001101010110011001;
assign LUT_4[60001] = 32'b00000000000000000110100010010001;
assign LUT_4[60002] = 32'b00000000000000001100110000111101;
assign LUT_4[60003] = 32'b00000000000000000101111100110101;
assign LUT_4[60004] = 32'b00000000000000001010010110110101;
assign LUT_4[60005] = 32'b00000000000000000011100010101101;
assign LUT_4[60006] = 32'b00000000000000001001110001011001;
assign LUT_4[60007] = 32'b00000000000000000010111101010001;
assign LUT_4[60008] = 32'b00000000000000000110100010101110;
assign LUT_4[60009] = 32'b11111111111111111111101110100110;
assign LUT_4[60010] = 32'b00000000000000000101111101010010;
assign LUT_4[60011] = 32'b11111111111111111111001001001010;
assign LUT_4[60012] = 32'b00000000000000000011100011001010;
assign LUT_4[60013] = 32'b11111111111111111100101111000010;
assign LUT_4[60014] = 32'b00000000000000000010111101101110;
assign LUT_4[60015] = 32'b11111111111111111100001001100110;
assign LUT_4[60016] = 32'b00000000000000001011001000000111;
assign LUT_4[60017] = 32'b00000000000000000100010011111111;
assign LUT_4[60018] = 32'b00000000000000001010100010101011;
assign LUT_4[60019] = 32'b00000000000000000011101110100011;
assign LUT_4[60020] = 32'b00000000000000001000001000100011;
assign LUT_4[60021] = 32'b00000000000000000001010100011011;
assign LUT_4[60022] = 32'b00000000000000000111100011000111;
assign LUT_4[60023] = 32'b00000000000000000000101110111111;
assign LUT_4[60024] = 32'b00000000000000000100010100011100;
assign LUT_4[60025] = 32'b11111111111111111101100000010100;
assign LUT_4[60026] = 32'b00000000000000000011101111000000;
assign LUT_4[60027] = 32'b11111111111111111100111010111000;
assign LUT_4[60028] = 32'b00000000000000000001010100111000;
assign LUT_4[60029] = 32'b11111111111111111010100000110000;
assign LUT_4[60030] = 32'b00000000000000000000101111011100;
assign LUT_4[60031] = 32'b11111111111111111001111011010100;
assign LUT_4[60032] = 32'b00000000000000010000001010000110;
assign LUT_4[60033] = 32'b00000000000000001001010101111110;
assign LUT_4[60034] = 32'b00000000000000001111100100101010;
assign LUT_4[60035] = 32'b00000000000000001000110000100010;
assign LUT_4[60036] = 32'b00000000000000001101001010100010;
assign LUT_4[60037] = 32'b00000000000000000110010110011010;
assign LUT_4[60038] = 32'b00000000000000001100100101000110;
assign LUT_4[60039] = 32'b00000000000000000101110000111110;
assign LUT_4[60040] = 32'b00000000000000001001010110011011;
assign LUT_4[60041] = 32'b00000000000000000010100010010011;
assign LUT_4[60042] = 32'b00000000000000001000110000111111;
assign LUT_4[60043] = 32'b00000000000000000001111100110111;
assign LUT_4[60044] = 32'b00000000000000000110010110110111;
assign LUT_4[60045] = 32'b11111111111111111111100010101111;
assign LUT_4[60046] = 32'b00000000000000000101110001011011;
assign LUT_4[60047] = 32'b11111111111111111110111101010011;
assign LUT_4[60048] = 32'b00000000000000001101111011110100;
assign LUT_4[60049] = 32'b00000000000000000111000111101100;
assign LUT_4[60050] = 32'b00000000000000001101010110011000;
assign LUT_4[60051] = 32'b00000000000000000110100010010000;
assign LUT_4[60052] = 32'b00000000000000001010111100010000;
assign LUT_4[60053] = 32'b00000000000000000100001000001000;
assign LUT_4[60054] = 32'b00000000000000001010010110110100;
assign LUT_4[60055] = 32'b00000000000000000011100010101100;
assign LUT_4[60056] = 32'b00000000000000000111001000001001;
assign LUT_4[60057] = 32'b00000000000000000000010100000001;
assign LUT_4[60058] = 32'b00000000000000000110100010101101;
assign LUT_4[60059] = 32'b11111111111111111111101110100101;
assign LUT_4[60060] = 32'b00000000000000000100001000100101;
assign LUT_4[60061] = 32'b11111111111111111101010100011101;
assign LUT_4[60062] = 32'b00000000000000000011100011001001;
assign LUT_4[60063] = 32'b11111111111111111100101111000001;
assign LUT_4[60064] = 32'b00000000000000001110100101001101;
assign LUT_4[60065] = 32'b00000000000000000111110001000101;
assign LUT_4[60066] = 32'b00000000000000001101111111110001;
assign LUT_4[60067] = 32'b00000000000000000111001011101001;
assign LUT_4[60068] = 32'b00000000000000001011100101101001;
assign LUT_4[60069] = 32'b00000000000000000100110001100001;
assign LUT_4[60070] = 32'b00000000000000001011000000001101;
assign LUT_4[60071] = 32'b00000000000000000100001100000101;
assign LUT_4[60072] = 32'b00000000000000000111110001100010;
assign LUT_4[60073] = 32'b00000000000000000000111101011010;
assign LUT_4[60074] = 32'b00000000000000000111001100000110;
assign LUT_4[60075] = 32'b00000000000000000000010111111110;
assign LUT_4[60076] = 32'b00000000000000000100110001111110;
assign LUT_4[60077] = 32'b11111111111111111101111101110110;
assign LUT_4[60078] = 32'b00000000000000000100001100100010;
assign LUT_4[60079] = 32'b11111111111111111101011000011010;
assign LUT_4[60080] = 32'b00000000000000001100010110111011;
assign LUT_4[60081] = 32'b00000000000000000101100010110011;
assign LUT_4[60082] = 32'b00000000000000001011110001011111;
assign LUT_4[60083] = 32'b00000000000000000100111101010111;
assign LUT_4[60084] = 32'b00000000000000001001010111010111;
assign LUT_4[60085] = 32'b00000000000000000010100011001111;
assign LUT_4[60086] = 32'b00000000000000001000110001111011;
assign LUT_4[60087] = 32'b00000000000000000001111101110011;
assign LUT_4[60088] = 32'b00000000000000000101100011010000;
assign LUT_4[60089] = 32'b11111111111111111110101111001000;
assign LUT_4[60090] = 32'b00000000000000000100111101110100;
assign LUT_4[60091] = 32'b11111111111111111110001001101100;
assign LUT_4[60092] = 32'b00000000000000000010100011101100;
assign LUT_4[60093] = 32'b11111111111111111011101111100100;
assign LUT_4[60094] = 32'b00000000000000000001111110010000;
assign LUT_4[60095] = 32'b11111111111111111011001010001000;
assign LUT_4[60096] = 32'b00000000000000010001100001011010;
assign LUT_4[60097] = 32'b00000000000000001010101101010010;
assign LUT_4[60098] = 32'b00000000000000010000111011111110;
assign LUT_4[60099] = 32'b00000000000000001010000111110110;
assign LUT_4[60100] = 32'b00000000000000001110100001110110;
assign LUT_4[60101] = 32'b00000000000000000111101101101110;
assign LUT_4[60102] = 32'b00000000000000001101111100011010;
assign LUT_4[60103] = 32'b00000000000000000111001000010010;
assign LUT_4[60104] = 32'b00000000000000001010101101101111;
assign LUT_4[60105] = 32'b00000000000000000011111001100111;
assign LUT_4[60106] = 32'b00000000000000001010001000010011;
assign LUT_4[60107] = 32'b00000000000000000011010100001011;
assign LUT_4[60108] = 32'b00000000000000000111101110001011;
assign LUT_4[60109] = 32'b00000000000000000000111010000011;
assign LUT_4[60110] = 32'b00000000000000000111001000101111;
assign LUT_4[60111] = 32'b00000000000000000000010100100111;
assign LUT_4[60112] = 32'b00000000000000001111010011001000;
assign LUT_4[60113] = 32'b00000000000000001000011111000000;
assign LUT_4[60114] = 32'b00000000000000001110101101101100;
assign LUT_4[60115] = 32'b00000000000000000111111001100100;
assign LUT_4[60116] = 32'b00000000000000001100010011100100;
assign LUT_4[60117] = 32'b00000000000000000101011111011100;
assign LUT_4[60118] = 32'b00000000000000001011101110001000;
assign LUT_4[60119] = 32'b00000000000000000100111010000000;
assign LUT_4[60120] = 32'b00000000000000001000011111011101;
assign LUT_4[60121] = 32'b00000000000000000001101011010101;
assign LUT_4[60122] = 32'b00000000000000000111111010000001;
assign LUT_4[60123] = 32'b00000000000000000001000101111001;
assign LUT_4[60124] = 32'b00000000000000000101011111111001;
assign LUT_4[60125] = 32'b11111111111111111110101011110001;
assign LUT_4[60126] = 32'b00000000000000000100111010011101;
assign LUT_4[60127] = 32'b11111111111111111110000110010101;
assign LUT_4[60128] = 32'b00000000000000001111111100100001;
assign LUT_4[60129] = 32'b00000000000000001001001000011001;
assign LUT_4[60130] = 32'b00000000000000001111010111000101;
assign LUT_4[60131] = 32'b00000000000000001000100010111101;
assign LUT_4[60132] = 32'b00000000000000001100111100111101;
assign LUT_4[60133] = 32'b00000000000000000110001000110101;
assign LUT_4[60134] = 32'b00000000000000001100010111100001;
assign LUT_4[60135] = 32'b00000000000000000101100011011001;
assign LUT_4[60136] = 32'b00000000000000001001001000110110;
assign LUT_4[60137] = 32'b00000000000000000010010100101110;
assign LUT_4[60138] = 32'b00000000000000001000100011011010;
assign LUT_4[60139] = 32'b00000000000000000001101111010010;
assign LUT_4[60140] = 32'b00000000000000000110001001010010;
assign LUT_4[60141] = 32'b11111111111111111111010101001010;
assign LUT_4[60142] = 32'b00000000000000000101100011110110;
assign LUT_4[60143] = 32'b11111111111111111110101111101110;
assign LUT_4[60144] = 32'b00000000000000001101101110001111;
assign LUT_4[60145] = 32'b00000000000000000110111010000111;
assign LUT_4[60146] = 32'b00000000000000001101001000110011;
assign LUT_4[60147] = 32'b00000000000000000110010100101011;
assign LUT_4[60148] = 32'b00000000000000001010101110101011;
assign LUT_4[60149] = 32'b00000000000000000011111010100011;
assign LUT_4[60150] = 32'b00000000000000001010001001001111;
assign LUT_4[60151] = 32'b00000000000000000011010101000111;
assign LUT_4[60152] = 32'b00000000000000000110111010100100;
assign LUT_4[60153] = 32'b00000000000000000000000110011100;
assign LUT_4[60154] = 32'b00000000000000000110010101001000;
assign LUT_4[60155] = 32'b11111111111111111111100001000000;
assign LUT_4[60156] = 32'b00000000000000000011111011000000;
assign LUT_4[60157] = 32'b11111111111111111101000110111000;
assign LUT_4[60158] = 32'b00000000000000000011010101100100;
assign LUT_4[60159] = 32'b11111111111111111100100001011100;
assign LUT_4[60160] = 32'b00000000000000010010011111100001;
assign LUT_4[60161] = 32'b00000000000000001011101011011001;
assign LUT_4[60162] = 32'b00000000000000010001111010000101;
assign LUT_4[60163] = 32'b00000000000000001011000101111101;
assign LUT_4[60164] = 32'b00000000000000001111011111111101;
assign LUT_4[60165] = 32'b00000000000000001000101011110101;
assign LUT_4[60166] = 32'b00000000000000001110111010100001;
assign LUT_4[60167] = 32'b00000000000000001000000110011001;
assign LUT_4[60168] = 32'b00000000000000001011101011110110;
assign LUT_4[60169] = 32'b00000000000000000100110111101110;
assign LUT_4[60170] = 32'b00000000000000001011000110011010;
assign LUT_4[60171] = 32'b00000000000000000100010010010010;
assign LUT_4[60172] = 32'b00000000000000001000101100010010;
assign LUT_4[60173] = 32'b00000000000000000001111000001010;
assign LUT_4[60174] = 32'b00000000000000001000000110110110;
assign LUT_4[60175] = 32'b00000000000000000001010010101110;
assign LUT_4[60176] = 32'b00000000000000010000010001001111;
assign LUT_4[60177] = 32'b00000000000000001001011101000111;
assign LUT_4[60178] = 32'b00000000000000001111101011110011;
assign LUT_4[60179] = 32'b00000000000000001000110111101011;
assign LUT_4[60180] = 32'b00000000000000001101010001101011;
assign LUT_4[60181] = 32'b00000000000000000110011101100011;
assign LUT_4[60182] = 32'b00000000000000001100101100001111;
assign LUT_4[60183] = 32'b00000000000000000101111000000111;
assign LUT_4[60184] = 32'b00000000000000001001011101100100;
assign LUT_4[60185] = 32'b00000000000000000010101001011100;
assign LUT_4[60186] = 32'b00000000000000001000111000001000;
assign LUT_4[60187] = 32'b00000000000000000010000100000000;
assign LUT_4[60188] = 32'b00000000000000000110011110000000;
assign LUT_4[60189] = 32'b11111111111111111111101001111000;
assign LUT_4[60190] = 32'b00000000000000000101111000100100;
assign LUT_4[60191] = 32'b11111111111111111111000100011100;
assign LUT_4[60192] = 32'b00000000000000010000111010101000;
assign LUT_4[60193] = 32'b00000000000000001010000110100000;
assign LUT_4[60194] = 32'b00000000000000010000010101001100;
assign LUT_4[60195] = 32'b00000000000000001001100001000100;
assign LUT_4[60196] = 32'b00000000000000001101111011000100;
assign LUT_4[60197] = 32'b00000000000000000111000110111100;
assign LUT_4[60198] = 32'b00000000000000001101010101101000;
assign LUT_4[60199] = 32'b00000000000000000110100001100000;
assign LUT_4[60200] = 32'b00000000000000001010000110111101;
assign LUT_4[60201] = 32'b00000000000000000011010010110101;
assign LUT_4[60202] = 32'b00000000000000001001100001100001;
assign LUT_4[60203] = 32'b00000000000000000010101101011001;
assign LUT_4[60204] = 32'b00000000000000000111000111011001;
assign LUT_4[60205] = 32'b00000000000000000000010011010001;
assign LUT_4[60206] = 32'b00000000000000000110100001111101;
assign LUT_4[60207] = 32'b11111111111111111111101101110101;
assign LUT_4[60208] = 32'b00000000000000001110101100010110;
assign LUT_4[60209] = 32'b00000000000000000111111000001110;
assign LUT_4[60210] = 32'b00000000000000001110000110111010;
assign LUT_4[60211] = 32'b00000000000000000111010010110010;
assign LUT_4[60212] = 32'b00000000000000001011101100110010;
assign LUT_4[60213] = 32'b00000000000000000100111000101010;
assign LUT_4[60214] = 32'b00000000000000001011000111010110;
assign LUT_4[60215] = 32'b00000000000000000100010011001110;
assign LUT_4[60216] = 32'b00000000000000000111111000101011;
assign LUT_4[60217] = 32'b00000000000000000001000100100011;
assign LUT_4[60218] = 32'b00000000000000000111010011001111;
assign LUT_4[60219] = 32'b00000000000000000000011111000111;
assign LUT_4[60220] = 32'b00000000000000000100111001000111;
assign LUT_4[60221] = 32'b11111111111111111110000100111111;
assign LUT_4[60222] = 32'b00000000000000000100010011101011;
assign LUT_4[60223] = 32'b11111111111111111101011111100011;
assign LUT_4[60224] = 32'b00000000000000010011110110110101;
assign LUT_4[60225] = 32'b00000000000000001101000010101101;
assign LUT_4[60226] = 32'b00000000000000010011010001011001;
assign LUT_4[60227] = 32'b00000000000000001100011101010001;
assign LUT_4[60228] = 32'b00000000000000010000110111010001;
assign LUT_4[60229] = 32'b00000000000000001010000011001001;
assign LUT_4[60230] = 32'b00000000000000010000010001110101;
assign LUT_4[60231] = 32'b00000000000000001001011101101101;
assign LUT_4[60232] = 32'b00000000000000001101000011001010;
assign LUT_4[60233] = 32'b00000000000000000110001111000010;
assign LUT_4[60234] = 32'b00000000000000001100011101101110;
assign LUT_4[60235] = 32'b00000000000000000101101001100110;
assign LUT_4[60236] = 32'b00000000000000001010000011100110;
assign LUT_4[60237] = 32'b00000000000000000011001111011110;
assign LUT_4[60238] = 32'b00000000000000001001011110001010;
assign LUT_4[60239] = 32'b00000000000000000010101010000010;
assign LUT_4[60240] = 32'b00000000000000010001101000100011;
assign LUT_4[60241] = 32'b00000000000000001010110100011011;
assign LUT_4[60242] = 32'b00000000000000010001000011000111;
assign LUT_4[60243] = 32'b00000000000000001010001110111111;
assign LUT_4[60244] = 32'b00000000000000001110101000111111;
assign LUT_4[60245] = 32'b00000000000000000111110100110111;
assign LUT_4[60246] = 32'b00000000000000001110000011100011;
assign LUT_4[60247] = 32'b00000000000000000111001111011011;
assign LUT_4[60248] = 32'b00000000000000001010110100111000;
assign LUT_4[60249] = 32'b00000000000000000100000000110000;
assign LUT_4[60250] = 32'b00000000000000001010001111011100;
assign LUT_4[60251] = 32'b00000000000000000011011011010100;
assign LUT_4[60252] = 32'b00000000000000000111110101010100;
assign LUT_4[60253] = 32'b00000000000000000001000001001100;
assign LUT_4[60254] = 32'b00000000000000000111001111111000;
assign LUT_4[60255] = 32'b00000000000000000000011011110000;
assign LUT_4[60256] = 32'b00000000000000010010010001111100;
assign LUT_4[60257] = 32'b00000000000000001011011101110100;
assign LUT_4[60258] = 32'b00000000000000010001101100100000;
assign LUT_4[60259] = 32'b00000000000000001010111000011000;
assign LUT_4[60260] = 32'b00000000000000001111010010011000;
assign LUT_4[60261] = 32'b00000000000000001000011110010000;
assign LUT_4[60262] = 32'b00000000000000001110101100111100;
assign LUT_4[60263] = 32'b00000000000000000111111000110100;
assign LUT_4[60264] = 32'b00000000000000001011011110010001;
assign LUT_4[60265] = 32'b00000000000000000100101010001001;
assign LUT_4[60266] = 32'b00000000000000001010111000110101;
assign LUT_4[60267] = 32'b00000000000000000100000100101101;
assign LUT_4[60268] = 32'b00000000000000001000011110101101;
assign LUT_4[60269] = 32'b00000000000000000001101010100101;
assign LUT_4[60270] = 32'b00000000000000000111111001010001;
assign LUT_4[60271] = 32'b00000000000000000001000101001001;
assign LUT_4[60272] = 32'b00000000000000010000000011101010;
assign LUT_4[60273] = 32'b00000000000000001001001111100010;
assign LUT_4[60274] = 32'b00000000000000001111011110001110;
assign LUT_4[60275] = 32'b00000000000000001000101010000110;
assign LUT_4[60276] = 32'b00000000000000001101000100000110;
assign LUT_4[60277] = 32'b00000000000000000110001111111110;
assign LUT_4[60278] = 32'b00000000000000001100011110101010;
assign LUT_4[60279] = 32'b00000000000000000101101010100010;
assign LUT_4[60280] = 32'b00000000000000001001001111111111;
assign LUT_4[60281] = 32'b00000000000000000010011011110111;
assign LUT_4[60282] = 32'b00000000000000001000101010100011;
assign LUT_4[60283] = 32'b00000000000000000001110110011011;
assign LUT_4[60284] = 32'b00000000000000000110010000011011;
assign LUT_4[60285] = 32'b11111111111111111111011100010011;
assign LUT_4[60286] = 32'b00000000000000000101101010111111;
assign LUT_4[60287] = 32'b11111111111111111110110110110111;
assign LUT_4[60288] = 32'b00000000000000010101000101101001;
assign LUT_4[60289] = 32'b00000000000000001110010001100001;
assign LUT_4[60290] = 32'b00000000000000010100100000001101;
assign LUT_4[60291] = 32'b00000000000000001101101100000101;
assign LUT_4[60292] = 32'b00000000000000010010000110000101;
assign LUT_4[60293] = 32'b00000000000000001011010001111101;
assign LUT_4[60294] = 32'b00000000000000010001100000101001;
assign LUT_4[60295] = 32'b00000000000000001010101100100001;
assign LUT_4[60296] = 32'b00000000000000001110010001111110;
assign LUT_4[60297] = 32'b00000000000000000111011101110110;
assign LUT_4[60298] = 32'b00000000000000001101101100100010;
assign LUT_4[60299] = 32'b00000000000000000110111000011010;
assign LUT_4[60300] = 32'b00000000000000001011010010011010;
assign LUT_4[60301] = 32'b00000000000000000100011110010010;
assign LUT_4[60302] = 32'b00000000000000001010101100111110;
assign LUT_4[60303] = 32'b00000000000000000011111000110110;
assign LUT_4[60304] = 32'b00000000000000010010110111010111;
assign LUT_4[60305] = 32'b00000000000000001100000011001111;
assign LUT_4[60306] = 32'b00000000000000010010010001111011;
assign LUT_4[60307] = 32'b00000000000000001011011101110011;
assign LUT_4[60308] = 32'b00000000000000001111110111110011;
assign LUT_4[60309] = 32'b00000000000000001001000011101011;
assign LUT_4[60310] = 32'b00000000000000001111010010010111;
assign LUT_4[60311] = 32'b00000000000000001000011110001111;
assign LUT_4[60312] = 32'b00000000000000001100000011101100;
assign LUT_4[60313] = 32'b00000000000000000101001111100100;
assign LUT_4[60314] = 32'b00000000000000001011011110010000;
assign LUT_4[60315] = 32'b00000000000000000100101010001000;
assign LUT_4[60316] = 32'b00000000000000001001000100001000;
assign LUT_4[60317] = 32'b00000000000000000010010000000000;
assign LUT_4[60318] = 32'b00000000000000001000011110101100;
assign LUT_4[60319] = 32'b00000000000000000001101010100100;
assign LUT_4[60320] = 32'b00000000000000010011100000110000;
assign LUT_4[60321] = 32'b00000000000000001100101100101000;
assign LUT_4[60322] = 32'b00000000000000010010111011010100;
assign LUT_4[60323] = 32'b00000000000000001100000111001100;
assign LUT_4[60324] = 32'b00000000000000010000100001001100;
assign LUT_4[60325] = 32'b00000000000000001001101101000100;
assign LUT_4[60326] = 32'b00000000000000001111111011110000;
assign LUT_4[60327] = 32'b00000000000000001001000111101000;
assign LUT_4[60328] = 32'b00000000000000001100101101000101;
assign LUT_4[60329] = 32'b00000000000000000101111000111101;
assign LUT_4[60330] = 32'b00000000000000001100000111101001;
assign LUT_4[60331] = 32'b00000000000000000101010011100001;
assign LUT_4[60332] = 32'b00000000000000001001101101100001;
assign LUT_4[60333] = 32'b00000000000000000010111001011001;
assign LUT_4[60334] = 32'b00000000000000001001001000000101;
assign LUT_4[60335] = 32'b00000000000000000010010011111101;
assign LUT_4[60336] = 32'b00000000000000010001010010011110;
assign LUT_4[60337] = 32'b00000000000000001010011110010110;
assign LUT_4[60338] = 32'b00000000000000010000101101000010;
assign LUT_4[60339] = 32'b00000000000000001001111000111010;
assign LUT_4[60340] = 32'b00000000000000001110010010111010;
assign LUT_4[60341] = 32'b00000000000000000111011110110010;
assign LUT_4[60342] = 32'b00000000000000001101101101011110;
assign LUT_4[60343] = 32'b00000000000000000110111001010110;
assign LUT_4[60344] = 32'b00000000000000001010011110110011;
assign LUT_4[60345] = 32'b00000000000000000011101010101011;
assign LUT_4[60346] = 32'b00000000000000001001111001010111;
assign LUT_4[60347] = 32'b00000000000000000011000101001111;
assign LUT_4[60348] = 32'b00000000000000000111011111001111;
assign LUT_4[60349] = 32'b00000000000000000000101011000111;
assign LUT_4[60350] = 32'b00000000000000000110111001110011;
assign LUT_4[60351] = 32'b00000000000000000000000101101011;
assign LUT_4[60352] = 32'b00000000000000010110011100111101;
assign LUT_4[60353] = 32'b00000000000000001111101000110101;
assign LUT_4[60354] = 32'b00000000000000010101110111100001;
assign LUT_4[60355] = 32'b00000000000000001111000011011001;
assign LUT_4[60356] = 32'b00000000000000010011011101011001;
assign LUT_4[60357] = 32'b00000000000000001100101001010001;
assign LUT_4[60358] = 32'b00000000000000010010110111111101;
assign LUT_4[60359] = 32'b00000000000000001100000011110101;
assign LUT_4[60360] = 32'b00000000000000001111101001010010;
assign LUT_4[60361] = 32'b00000000000000001000110101001010;
assign LUT_4[60362] = 32'b00000000000000001111000011110110;
assign LUT_4[60363] = 32'b00000000000000001000001111101110;
assign LUT_4[60364] = 32'b00000000000000001100101001101110;
assign LUT_4[60365] = 32'b00000000000000000101110101100110;
assign LUT_4[60366] = 32'b00000000000000001100000100010010;
assign LUT_4[60367] = 32'b00000000000000000101010000001010;
assign LUT_4[60368] = 32'b00000000000000010100001110101011;
assign LUT_4[60369] = 32'b00000000000000001101011010100011;
assign LUT_4[60370] = 32'b00000000000000010011101001001111;
assign LUT_4[60371] = 32'b00000000000000001100110101000111;
assign LUT_4[60372] = 32'b00000000000000010001001111000111;
assign LUT_4[60373] = 32'b00000000000000001010011010111111;
assign LUT_4[60374] = 32'b00000000000000010000101001101011;
assign LUT_4[60375] = 32'b00000000000000001001110101100011;
assign LUT_4[60376] = 32'b00000000000000001101011011000000;
assign LUT_4[60377] = 32'b00000000000000000110100110111000;
assign LUT_4[60378] = 32'b00000000000000001100110101100100;
assign LUT_4[60379] = 32'b00000000000000000110000001011100;
assign LUT_4[60380] = 32'b00000000000000001010011011011100;
assign LUT_4[60381] = 32'b00000000000000000011100111010100;
assign LUT_4[60382] = 32'b00000000000000001001110110000000;
assign LUT_4[60383] = 32'b00000000000000000011000001111000;
assign LUT_4[60384] = 32'b00000000000000010100111000000100;
assign LUT_4[60385] = 32'b00000000000000001110000011111100;
assign LUT_4[60386] = 32'b00000000000000010100010010101000;
assign LUT_4[60387] = 32'b00000000000000001101011110100000;
assign LUT_4[60388] = 32'b00000000000000010001111000100000;
assign LUT_4[60389] = 32'b00000000000000001011000100011000;
assign LUT_4[60390] = 32'b00000000000000010001010011000100;
assign LUT_4[60391] = 32'b00000000000000001010011110111100;
assign LUT_4[60392] = 32'b00000000000000001110000100011001;
assign LUT_4[60393] = 32'b00000000000000000111010000010001;
assign LUT_4[60394] = 32'b00000000000000001101011110111101;
assign LUT_4[60395] = 32'b00000000000000000110101010110101;
assign LUT_4[60396] = 32'b00000000000000001011000100110101;
assign LUT_4[60397] = 32'b00000000000000000100010000101101;
assign LUT_4[60398] = 32'b00000000000000001010011111011001;
assign LUT_4[60399] = 32'b00000000000000000011101011010001;
assign LUT_4[60400] = 32'b00000000000000010010101001110010;
assign LUT_4[60401] = 32'b00000000000000001011110101101010;
assign LUT_4[60402] = 32'b00000000000000010010000100010110;
assign LUT_4[60403] = 32'b00000000000000001011010000001110;
assign LUT_4[60404] = 32'b00000000000000001111101010001110;
assign LUT_4[60405] = 32'b00000000000000001000110110000110;
assign LUT_4[60406] = 32'b00000000000000001111000100110010;
assign LUT_4[60407] = 32'b00000000000000001000010000101010;
assign LUT_4[60408] = 32'b00000000000000001011110110000111;
assign LUT_4[60409] = 32'b00000000000000000101000001111111;
assign LUT_4[60410] = 32'b00000000000000001011010000101011;
assign LUT_4[60411] = 32'b00000000000000000100011100100011;
assign LUT_4[60412] = 32'b00000000000000001000110110100011;
assign LUT_4[60413] = 32'b00000000000000000010000010011011;
assign LUT_4[60414] = 32'b00000000000000001000010001000111;
assign LUT_4[60415] = 32'b00000000000000000001011100111111;
assign LUT_4[60416] = 32'b00000000000000010000001010010101;
assign LUT_4[60417] = 32'b00000000000000001001010110001101;
assign LUT_4[60418] = 32'b00000000000000001111100100111001;
assign LUT_4[60419] = 32'b00000000000000001000110000110001;
assign LUT_4[60420] = 32'b00000000000000001101001010110001;
assign LUT_4[60421] = 32'b00000000000000000110010110101001;
assign LUT_4[60422] = 32'b00000000000000001100100101010101;
assign LUT_4[60423] = 32'b00000000000000000101110001001101;
assign LUT_4[60424] = 32'b00000000000000001001010110101010;
assign LUT_4[60425] = 32'b00000000000000000010100010100010;
assign LUT_4[60426] = 32'b00000000000000001000110001001110;
assign LUT_4[60427] = 32'b00000000000000000001111101000110;
assign LUT_4[60428] = 32'b00000000000000000110010111000110;
assign LUT_4[60429] = 32'b11111111111111111111100010111110;
assign LUT_4[60430] = 32'b00000000000000000101110001101010;
assign LUT_4[60431] = 32'b11111111111111111110111101100010;
assign LUT_4[60432] = 32'b00000000000000001101111100000011;
assign LUT_4[60433] = 32'b00000000000000000111000111111011;
assign LUT_4[60434] = 32'b00000000000000001101010110100111;
assign LUT_4[60435] = 32'b00000000000000000110100010011111;
assign LUT_4[60436] = 32'b00000000000000001010111100011111;
assign LUT_4[60437] = 32'b00000000000000000100001000010111;
assign LUT_4[60438] = 32'b00000000000000001010010111000011;
assign LUT_4[60439] = 32'b00000000000000000011100010111011;
assign LUT_4[60440] = 32'b00000000000000000111001000011000;
assign LUT_4[60441] = 32'b00000000000000000000010100010000;
assign LUT_4[60442] = 32'b00000000000000000110100010111100;
assign LUT_4[60443] = 32'b11111111111111111111101110110100;
assign LUT_4[60444] = 32'b00000000000000000100001000110100;
assign LUT_4[60445] = 32'b11111111111111111101010100101100;
assign LUT_4[60446] = 32'b00000000000000000011100011011000;
assign LUT_4[60447] = 32'b11111111111111111100101111010000;
assign LUT_4[60448] = 32'b00000000000000001110100101011100;
assign LUT_4[60449] = 32'b00000000000000000111110001010100;
assign LUT_4[60450] = 32'b00000000000000001110000000000000;
assign LUT_4[60451] = 32'b00000000000000000111001011111000;
assign LUT_4[60452] = 32'b00000000000000001011100101111000;
assign LUT_4[60453] = 32'b00000000000000000100110001110000;
assign LUT_4[60454] = 32'b00000000000000001011000000011100;
assign LUT_4[60455] = 32'b00000000000000000100001100010100;
assign LUT_4[60456] = 32'b00000000000000000111110001110001;
assign LUT_4[60457] = 32'b00000000000000000000111101101001;
assign LUT_4[60458] = 32'b00000000000000000111001100010101;
assign LUT_4[60459] = 32'b00000000000000000000011000001101;
assign LUT_4[60460] = 32'b00000000000000000100110010001101;
assign LUT_4[60461] = 32'b11111111111111111101111110000101;
assign LUT_4[60462] = 32'b00000000000000000100001100110001;
assign LUT_4[60463] = 32'b11111111111111111101011000101001;
assign LUT_4[60464] = 32'b00000000000000001100010111001010;
assign LUT_4[60465] = 32'b00000000000000000101100011000010;
assign LUT_4[60466] = 32'b00000000000000001011110001101110;
assign LUT_4[60467] = 32'b00000000000000000100111101100110;
assign LUT_4[60468] = 32'b00000000000000001001010111100110;
assign LUT_4[60469] = 32'b00000000000000000010100011011110;
assign LUT_4[60470] = 32'b00000000000000001000110010001010;
assign LUT_4[60471] = 32'b00000000000000000001111110000010;
assign LUT_4[60472] = 32'b00000000000000000101100011011111;
assign LUT_4[60473] = 32'b11111111111111111110101111010111;
assign LUT_4[60474] = 32'b00000000000000000100111110000011;
assign LUT_4[60475] = 32'b11111111111111111110001001111011;
assign LUT_4[60476] = 32'b00000000000000000010100011111011;
assign LUT_4[60477] = 32'b11111111111111111011101111110011;
assign LUT_4[60478] = 32'b00000000000000000001111110011111;
assign LUT_4[60479] = 32'b11111111111111111011001010010111;
assign LUT_4[60480] = 32'b00000000000000010001100001101001;
assign LUT_4[60481] = 32'b00000000000000001010101101100001;
assign LUT_4[60482] = 32'b00000000000000010000111100001101;
assign LUT_4[60483] = 32'b00000000000000001010001000000101;
assign LUT_4[60484] = 32'b00000000000000001110100010000101;
assign LUT_4[60485] = 32'b00000000000000000111101101111101;
assign LUT_4[60486] = 32'b00000000000000001101111100101001;
assign LUT_4[60487] = 32'b00000000000000000111001000100001;
assign LUT_4[60488] = 32'b00000000000000001010101101111110;
assign LUT_4[60489] = 32'b00000000000000000011111001110110;
assign LUT_4[60490] = 32'b00000000000000001010001000100010;
assign LUT_4[60491] = 32'b00000000000000000011010100011010;
assign LUT_4[60492] = 32'b00000000000000000111101110011010;
assign LUT_4[60493] = 32'b00000000000000000000111010010010;
assign LUT_4[60494] = 32'b00000000000000000111001000111110;
assign LUT_4[60495] = 32'b00000000000000000000010100110110;
assign LUT_4[60496] = 32'b00000000000000001111010011010111;
assign LUT_4[60497] = 32'b00000000000000001000011111001111;
assign LUT_4[60498] = 32'b00000000000000001110101101111011;
assign LUT_4[60499] = 32'b00000000000000000111111001110011;
assign LUT_4[60500] = 32'b00000000000000001100010011110011;
assign LUT_4[60501] = 32'b00000000000000000101011111101011;
assign LUT_4[60502] = 32'b00000000000000001011101110010111;
assign LUT_4[60503] = 32'b00000000000000000100111010001111;
assign LUT_4[60504] = 32'b00000000000000001000011111101100;
assign LUT_4[60505] = 32'b00000000000000000001101011100100;
assign LUT_4[60506] = 32'b00000000000000000111111010010000;
assign LUT_4[60507] = 32'b00000000000000000001000110001000;
assign LUT_4[60508] = 32'b00000000000000000101100000001000;
assign LUT_4[60509] = 32'b11111111111111111110101100000000;
assign LUT_4[60510] = 32'b00000000000000000100111010101100;
assign LUT_4[60511] = 32'b11111111111111111110000110100100;
assign LUT_4[60512] = 32'b00000000000000001111111100110000;
assign LUT_4[60513] = 32'b00000000000000001001001000101000;
assign LUT_4[60514] = 32'b00000000000000001111010111010100;
assign LUT_4[60515] = 32'b00000000000000001000100011001100;
assign LUT_4[60516] = 32'b00000000000000001100111101001100;
assign LUT_4[60517] = 32'b00000000000000000110001001000100;
assign LUT_4[60518] = 32'b00000000000000001100010111110000;
assign LUT_4[60519] = 32'b00000000000000000101100011101000;
assign LUT_4[60520] = 32'b00000000000000001001001001000101;
assign LUT_4[60521] = 32'b00000000000000000010010100111101;
assign LUT_4[60522] = 32'b00000000000000001000100011101001;
assign LUT_4[60523] = 32'b00000000000000000001101111100001;
assign LUT_4[60524] = 32'b00000000000000000110001001100001;
assign LUT_4[60525] = 32'b11111111111111111111010101011001;
assign LUT_4[60526] = 32'b00000000000000000101100100000101;
assign LUT_4[60527] = 32'b11111111111111111110101111111101;
assign LUT_4[60528] = 32'b00000000000000001101101110011110;
assign LUT_4[60529] = 32'b00000000000000000110111010010110;
assign LUT_4[60530] = 32'b00000000000000001101001001000010;
assign LUT_4[60531] = 32'b00000000000000000110010100111010;
assign LUT_4[60532] = 32'b00000000000000001010101110111010;
assign LUT_4[60533] = 32'b00000000000000000011111010110010;
assign LUT_4[60534] = 32'b00000000000000001010001001011110;
assign LUT_4[60535] = 32'b00000000000000000011010101010110;
assign LUT_4[60536] = 32'b00000000000000000110111010110011;
assign LUT_4[60537] = 32'b00000000000000000000000110101011;
assign LUT_4[60538] = 32'b00000000000000000110010101010111;
assign LUT_4[60539] = 32'b11111111111111111111100001001111;
assign LUT_4[60540] = 32'b00000000000000000011111011001111;
assign LUT_4[60541] = 32'b11111111111111111101000111000111;
assign LUT_4[60542] = 32'b00000000000000000011010101110011;
assign LUT_4[60543] = 32'b11111111111111111100100001101011;
assign LUT_4[60544] = 32'b00000000000000010010110000011101;
assign LUT_4[60545] = 32'b00000000000000001011111100010101;
assign LUT_4[60546] = 32'b00000000000000010010001011000001;
assign LUT_4[60547] = 32'b00000000000000001011010110111001;
assign LUT_4[60548] = 32'b00000000000000001111110000111001;
assign LUT_4[60549] = 32'b00000000000000001000111100110001;
assign LUT_4[60550] = 32'b00000000000000001111001011011101;
assign LUT_4[60551] = 32'b00000000000000001000010111010101;
assign LUT_4[60552] = 32'b00000000000000001011111100110010;
assign LUT_4[60553] = 32'b00000000000000000101001000101010;
assign LUT_4[60554] = 32'b00000000000000001011010111010110;
assign LUT_4[60555] = 32'b00000000000000000100100011001110;
assign LUT_4[60556] = 32'b00000000000000001000111101001110;
assign LUT_4[60557] = 32'b00000000000000000010001001000110;
assign LUT_4[60558] = 32'b00000000000000001000010111110010;
assign LUT_4[60559] = 32'b00000000000000000001100011101010;
assign LUT_4[60560] = 32'b00000000000000010000100010001011;
assign LUT_4[60561] = 32'b00000000000000001001101110000011;
assign LUT_4[60562] = 32'b00000000000000001111111100101111;
assign LUT_4[60563] = 32'b00000000000000001001001000100111;
assign LUT_4[60564] = 32'b00000000000000001101100010100111;
assign LUT_4[60565] = 32'b00000000000000000110101110011111;
assign LUT_4[60566] = 32'b00000000000000001100111101001011;
assign LUT_4[60567] = 32'b00000000000000000110001001000011;
assign LUT_4[60568] = 32'b00000000000000001001101110100000;
assign LUT_4[60569] = 32'b00000000000000000010111010011000;
assign LUT_4[60570] = 32'b00000000000000001001001001000100;
assign LUT_4[60571] = 32'b00000000000000000010010100111100;
assign LUT_4[60572] = 32'b00000000000000000110101110111100;
assign LUT_4[60573] = 32'b11111111111111111111111010110100;
assign LUT_4[60574] = 32'b00000000000000000110001001100000;
assign LUT_4[60575] = 32'b11111111111111111111010101011000;
assign LUT_4[60576] = 32'b00000000000000010001001011100100;
assign LUT_4[60577] = 32'b00000000000000001010010111011100;
assign LUT_4[60578] = 32'b00000000000000010000100110001000;
assign LUT_4[60579] = 32'b00000000000000001001110010000000;
assign LUT_4[60580] = 32'b00000000000000001110001100000000;
assign LUT_4[60581] = 32'b00000000000000000111010111111000;
assign LUT_4[60582] = 32'b00000000000000001101100110100100;
assign LUT_4[60583] = 32'b00000000000000000110110010011100;
assign LUT_4[60584] = 32'b00000000000000001010010111111001;
assign LUT_4[60585] = 32'b00000000000000000011100011110001;
assign LUT_4[60586] = 32'b00000000000000001001110010011101;
assign LUT_4[60587] = 32'b00000000000000000010111110010101;
assign LUT_4[60588] = 32'b00000000000000000111011000010101;
assign LUT_4[60589] = 32'b00000000000000000000100100001101;
assign LUT_4[60590] = 32'b00000000000000000110110010111001;
assign LUT_4[60591] = 32'b11111111111111111111111110110001;
assign LUT_4[60592] = 32'b00000000000000001110111101010010;
assign LUT_4[60593] = 32'b00000000000000001000001001001010;
assign LUT_4[60594] = 32'b00000000000000001110010111110110;
assign LUT_4[60595] = 32'b00000000000000000111100011101110;
assign LUT_4[60596] = 32'b00000000000000001011111101101110;
assign LUT_4[60597] = 32'b00000000000000000101001001100110;
assign LUT_4[60598] = 32'b00000000000000001011011000010010;
assign LUT_4[60599] = 32'b00000000000000000100100100001010;
assign LUT_4[60600] = 32'b00000000000000001000001001100111;
assign LUT_4[60601] = 32'b00000000000000000001010101011111;
assign LUT_4[60602] = 32'b00000000000000000111100100001011;
assign LUT_4[60603] = 32'b00000000000000000000110000000011;
assign LUT_4[60604] = 32'b00000000000000000101001010000011;
assign LUT_4[60605] = 32'b11111111111111111110010101111011;
assign LUT_4[60606] = 32'b00000000000000000100100100100111;
assign LUT_4[60607] = 32'b11111111111111111101110000011111;
assign LUT_4[60608] = 32'b00000000000000010100000111110001;
assign LUT_4[60609] = 32'b00000000000000001101010011101001;
assign LUT_4[60610] = 32'b00000000000000010011100010010101;
assign LUT_4[60611] = 32'b00000000000000001100101110001101;
assign LUT_4[60612] = 32'b00000000000000010001001000001101;
assign LUT_4[60613] = 32'b00000000000000001010010100000101;
assign LUT_4[60614] = 32'b00000000000000010000100010110001;
assign LUT_4[60615] = 32'b00000000000000001001101110101001;
assign LUT_4[60616] = 32'b00000000000000001101010100000110;
assign LUT_4[60617] = 32'b00000000000000000110011111111110;
assign LUT_4[60618] = 32'b00000000000000001100101110101010;
assign LUT_4[60619] = 32'b00000000000000000101111010100010;
assign LUT_4[60620] = 32'b00000000000000001010010100100010;
assign LUT_4[60621] = 32'b00000000000000000011100000011010;
assign LUT_4[60622] = 32'b00000000000000001001101111000110;
assign LUT_4[60623] = 32'b00000000000000000010111010111110;
assign LUT_4[60624] = 32'b00000000000000010001111001011111;
assign LUT_4[60625] = 32'b00000000000000001011000101010111;
assign LUT_4[60626] = 32'b00000000000000010001010100000011;
assign LUT_4[60627] = 32'b00000000000000001010011111111011;
assign LUT_4[60628] = 32'b00000000000000001110111001111011;
assign LUT_4[60629] = 32'b00000000000000001000000101110011;
assign LUT_4[60630] = 32'b00000000000000001110010100011111;
assign LUT_4[60631] = 32'b00000000000000000111100000010111;
assign LUT_4[60632] = 32'b00000000000000001011000101110100;
assign LUT_4[60633] = 32'b00000000000000000100010001101100;
assign LUT_4[60634] = 32'b00000000000000001010100000011000;
assign LUT_4[60635] = 32'b00000000000000000011101100010000;
assign LUT_4[60636] = 32'b00000000000000001000000110010000;
assign LUT_4[60637] = 32'b00000000000000000001010010001000;
assign LUT_4[60638] = 32'b00000000000000000111100000110100;
assign LUT_4[60639] = 32'b00000000000000000000101100101100;
assign LUT_4[60640] = 32'b00000000000000010010100010111000;
assign LUT_4[60641] = 32'b00000000000000001011101110110000;
assign LUT_4[60642] = 32'b00000000000000010001111101011100;
assign LUT_4[60643] = 32'b00000000000000001011001001010100;
assign LUT_4[60644] = 32'b00000000000000001111100011010100;
assign LUT_4[60645] = 32'b00000000000000001000101111001100;
assign LUT_4[60646] = 32'b00000000000000001110111101111000;
assign LUT_4[60647] = 32'b00000000000000001000001001110000;
assign LUT_4[60648] = 32'b00000000000000001011101111001101;
assign LUT_4[60649] = 32'b00000000000000000100111011000101;
assign LUT_4[60650] = 32'b00000000000000001011001001110001;
assign LUT_4[60651] = 32'b00000000000000000100010101101001;
assign LUT_4[60652] = 32'b00000000000000001000101111101001;
assign LUT_4[60653] = 32'b00000000000000000001111011100001;
assign LUT_4[60654] = 32'b00000000000000001000001010001101;
assign LUT_4[60655] = 32'b00000000000000000001010110000101;
assign LUT_4[60656] = 32'b00000000000000010000010100100110;
assign LUT_4[60657] = 32'b00000000000000001001100000011110;
assign LUT_4[60658] = 32'b00000000000000001111101111001010;
assign LUT_4[60659] = 32'b00000000000000001000111011000010;
assign LUT_4[60660] = 32'b00000000000000001101010101000010;
assign LUT_4[60661] = 32'b00000000000000000110100000111010;
assign LUT_4[60662] = 32'b00000000000000001100101111100110;
assign LUT_4[60663] = 32'b00000000000000000101111011011110;
assign LUT_4[60664] = 32'b00000000000000001001100000111011;
assign LUT_4[60665] = 32'b00000000000000000010101100110011;
assign LUT_4[60666] = 32'b00000000000000001000111011011111;
assign LUT_4[60667] = 32'b00000000000000000010000111010111;
assign LUT_4[60668] = 32'b00000000000000000110100001010111;
assign LUT_4[60669] = 32'b11111111111111111111101101001111;
assign LUT_4[60670] = 32'b00000000000000000101111011111011;
assign LUT_4[60671] = 32'b11111111111111111111000111110011;
assign LUT_4[60672] = 32'b00000000000000010101000101111000;
assign LUT_4[60673] = 32'b00000000000000001110010001110000;
assign LUT_4[60674] = 32'b00000000000000010100100000011100;
assign LUT_4[60675] = 32'b00000000000000001101101100010100;
assign LUT_4[60676] = 32'b00000000000000010010000110010100;
assign LUT_4[60677] = 32'b00000000000000001011010010001100;
assign LUT_4[60678] = 32'b00000000000000010001100000111000;
assign LUT_4[60679] = 32'b00000000000000001010101100110000;
assign LUT_4[60680] = 32'b00000000000000001110010010001101;
assign LUT_4[60681] = 32'b00000000000000000111011110000101;
assign LUT_4[60682] = 32'b00000000000000001101101100110001;
assign LUT_4[60683] = 32'b00000000000000000110111000101001;
assign LUT_4[60684] = 32'b00000000000000001011010010101001;
assign LUT_4[60685] = 32'b00000000000000000100011110100001;
assign LUT_4[60686] = 32'b00000000000000001010101101001101;
assign LUT_4[60687] = 32'b00000000000000000011111001000101;
assign LUT_4[60688] = 32'b00000000000000010010110111100110;
assign LUT_4[60689] = 32'b00000000000000001100000011011110;
assign LUT_4[60690] = 32'b00000000000000010010010010001010;
assign LUT_4[60691] = 32'b00000000000000001011011110000010;
assign LUT_4[60692] = 32'b00000000000000001111111000000010;
assign LUT_4[60693] = 32'b00000000000000001001000011111010;
assign LUT_4[60694] = 32'b00000000000000001111010010100110;
assign LUT_4[60695] = 32'b00000000000000001000011110011110;
assign LUT_4[60696] = 32'b00000000000000001100000011111011;
assign LUT_4[60697] = 32'b00000000000000000101001111110011;
assign LUT_4[60698] = 32'b00000000000000001011011110011111;
assign LUT_4[60699] = 32'b00000000000000000100101010010111;
assign LUT_4[60700] = 32'b00000000000000001001000100010111;
assign LUT_4[60701] = 32'b00000000000000000010010000001111;
assign LUT_4[60702] = 32'b00000000000000001000011110111011;
assign LUT_4[60703] = 32'b00000000000000000001101010110011;
assign LUT_4[60704] = 32'b00000000000000010011100000111111;
assign LUT_4[60705] = 32'b00000000000000001100101100110111;
assign LUT_4[60706] = 32'b00000000000000010010111011100011;
assign LUT_4[60707] = 32'b00000000000000001100000111011011;
assign LUT_4[60708] = 32'b00000000000000010000100001011011;
assign LUT_4[60709] = 32'b00000000000000001001101101010011;
assign LUT_4[60710] = 32'b00000000000000001111111011111111;
assign LUT_4[60711] = 32'b00000000000000001001000111110111;
assign LUT_4[60712] = 32'b00000000000000001100101101010100;
assign LUT_4[60713] = 32'b00000000000000000101111001001100;
assign LUT_4[60714] = 32'b00000000000000001100000111111000;
assign LUT_4[60715] = 32'b00000000000000000101010011110000;
assign LUT_4[60716] = 32'b00000000000000001001101101110000;
assign LUT_4[60717] = 32'b00000000000000000010111001101000;
assign LUT_4[60718] = 32'b00000000000000001001001000010100;
assign LUT_4[60719] = 32'b00000000000000000010010100001100;
assign LUT_4[60720] = 32'b00000000000000010001010010101101;
assign LUT_4[60721] = 32'b00000000000000001010011110100101;
assign LUT_4[60722] = 32'b00000000000000010000101101010001;
assign LUT_4[60723] = 32'b00000000000000001001111001001001;
assign LUT_4[60724] = 32'b00000000000000001110010011001001;
assign LUT_4[60725] = 32'b00000000000000000111011111000001;
assign LUT_4[60726] = 32'b00000000000000001101101101101101;
assign LUT_4[60727] = 32'b00000000000000000110111001100101;
assign LUT_4[60728] = 32'b00000000000000001010011111000010;
assign LUT_4[60729] = 32'b00000000000000000011101010111010;
assign LUT_4[60730] = 32'b00000000000000001001111001100110;
assign LUT_4[60731] = 32'b00000000000000000011000101011110;
assign LUT_4[60732] = 32'b00000000000000000111011111011110;
assign LUT_4[60733] = 32'b00000000000000000000101011010110;
assign LUT_4[60734] = 32'b00000000000000000110111010000010;
assign LUT_4[60735] = 32'b00000000000000000000000101111010;
assign LUT_4[60736] = 32'b00000000000000010110011101001100;
assign LUT_4[60737] = 32'b00000000000000001111101001000100;
assign LUT_4[60738] = 32'b00000000000000010101110111110000;
assign LUT_4[60739] = 32'b00000000000000001111000011101000;
assign LUT_4[60740] = 32'b00000000000000010011011101101000;
assign LUT_4[60741] = 32'b00000000000000001100101001100000;
assign LUT_4[60742] = 32'b00000000000000010010111000001100;
assign LUT_4[60743] = 32'b00000000000000001100000100000100;
assign LUT_4[60744] = 32'b00000000000000001111101001100001;
assign LUT_4[60745] = 32'b00000000000000001000110101011001;
assign LUT_4[60746] = 32'b00000000000000001111000100000101;
assign LUT_4[60747] = 32'b00000000000000001000001111111101;
assign LUT_4[60748] = 32'b00000000000000001100101001111101;
assign LUT_4[60749] = 32'b00000000000000000101110101110101;
assign LUT_4[60750] = 32'b00000000000000001100000100100001;
assign LUT_4[60751] = 32'b00000000000000000101010000011001;
assign LUT_4[60752] = 32'b00000000000000010100001110111010;
assign LUT_4[60753] = 32'b00000000000000001101011010110010;
assign LUT_4[60754] = 32'b00000000000000010011101001011110;
assign LUT_4[60755] = 32'b00000000000000001100110101010110;
assign LUT_4[60756] = 32'b00000000000000010001001111010110;
assign LUT_4[60757] = 32'b00000000000000001010011011001110;
assign LUT_4[60758] = 32'b00000000000000010000101001111010;
assign LUT_4[60759] = 32'b00000000000000001001110101110010;
assign LUT_4[60760] = 32'b00000000000000001101011011001111;
assign LUT_4[60761] = 32'b00000000000000000110100111000111;
assign LUT_4[60762] = 32'b00000000000000001100110101110011;
assign LUT_4[60763] = 32'b00000000000000000110000001101011;
assign LUT_4[60764] = 32'b00000000000000001010011011101011;
assign LUT_4[60765] = 32'b00000000000000000011100111100011;
assign LUT_4[60766] = 32'b00000000000000001001110110001111;
assign LUT_4[60767] = 32'b00000000000000000011000010000111;
assign LUT_4[60768] = 32'b00000000000000010100111000010011;
assign LUT_4[60769] = 32'b00000000000000001110000100001011;
assign LUT_4[60770] = 32'b00000000000000010100010010110111;
assign LUT_4[60771] = 32'b00000000000000001101011110101111;
assign LUT_4[60772] = 32'b00000000000000010001111000101111;
assign LUT_4[60773] = 32'b00000000000000001011000100100111;
assign LUT_4[60774] = 32'b00000000000000010001010011010011;
assign LUT_4[60775] = 32'b00000000000000001010011111001011;
assign LUT_4[60776] = 32'b00000000000000001110000100101000;
assign LUT_4[60777] = 32'b00000000000000000111010000100000;
assign LUT_4[60778] = 32'b00000000000000001101011111001100;
assign LUT_4[60779] = 32'b00000000000000000110101011000100;
assign LUT_4[60780] = 32'b00000000000000001011000101000100;
assign LUT_4[60781] = 32'b00000000000000000100010000111100;
assign LUT_4[60782] = 32'b00000000000000001010011111101000;
assign LUT_4[60783] = 32'b00000000000000000011101011100000;
assign LUT_4[60784] = 32'b00000000000000010010101010000001;
assign LUT_4[60785] = 32'b00000000000000001011110101111001;
assign LUT_4[60786] = 32'b00000000000000010010000100100101;
assign LUT_4[60787] = 32'b00000000000000001011010000011101;
assign LUT_4[60788] = 32'b00000000000000001111101010011101;
assign LUT_4[60789] = 32'b00000000000000001000110110010101;
assign LUT_4[60790] = 32'b00000000000000001111000101000001;
assign LUT_4[60791] = 32'b00000000000000001000010000111001;
assign LUT_4[60792] = 32'b00000000000000001011110110010110;
assign LUT_4[60793] = 32'b00000000000000000101000010001110;
assign LUT_4[60794] = 32'b00000000000000001011010000111010;
assign LUT_4[60795] = 32'b00000000000000000100011100110010;
assign LUT_4[60796] = 32'b00000000000000001000110110110010;
assign LUT_4[60797] = 32'b00000000000000000010000010101010;
assign LUT_4[60798] = 32'b00000000000000001000010001010110;
assign LUT_4[60799] = 32'b00000000000000000001011101001110;
assign LUT_4[60800] = 32'b00000000000000010111101100000000;
assign LUT_4[60801] = 32'b00000000000000010000110111111000;
assign LUT_4[60802] = 32'b00000000000000010111000110100100;
assign LUT_4[60803] = 32'b00000000000000010000010010011100;
assign LUT_4[60804] = 32'b00000000000000010100101100011100;
assign LUT_4[60805] = 32'b00000000000000001101111000010100;
assign LUT_4[60806] = 32'b00000000000000010100000111000000;
assign LUT_4[60807] = 32'b00000000000000001101010010111000;
assign LUT_4[60808] = 32'b00000000000000010000111000010101;
assign LUT_4[60809] = 32'b00000000000000001010000100001101;
assign LUT_4[60810] = 32'b00000000000000010000010010111001;
assign LUT_4[60811] = 32'b00000000000000001001011110110001;
assign LUT_4[60812] = 32'b00000000000000001101111000110001;
assign LUT_4[60813] = 32'b00000000000000000111000100101001;
assign LUT_4[60814] = 32'b00000000000000001101010011010101;
assign LUT_4[60815] = 32'b00000000000000000110011111001101;
assign LUT_4[60816] = 32'b00000000000000010101011101101110;
assign LUT_4[60817] = 32'b00000000000000001110101001100110;
assign LUT_4[60818] = 32'b00000000000000010100111000010010;
assign LUT_4[60819] = 32'b00000000000000001110000100001010;
assign LUT_4[60820] = 32'b00000000000000010010011110001010;
assign LUT_4[60821] = 32'b00000000000000001011101010000010;
assign LUT_4[60822] = 32'b00000000000000010001111000101110;
assign LUT_4[60823] = 32'b00000000000000001011000100100110;
assign LUT_4[60824] = 32'b00000000000000001110101010000011;
assign LUT_4[60825] = 32'b00000000000000000111110101111011;
assign LUT_4[60826] = 32'b00000000000000001110000100100111;
assign LUT_4[60827] = 32'b00000000000000000111010000011111;
assign LUT_4[60828] = 32'b00000000000000001011101010011111;
assign LUT_4[60829] = 32'b00000000000000000100110110010111;
assign LUT_4[60830] = 32'b00000000000000001011000101000011;
assign LUT_4[60831] = 32'b00000000000000000100010000111011;
assign LUT_4[60832] = 32'b00000000000000010110000111000111;
assign LUT_4[60833] = 32'b00000000000000001111010010111111;
assign LUT_4[60834] = 32'b00000000000000010101100001101011;
assign LUT_4[60835] = 32'b00000000000000001110101101100011;
assign LUT_4[60836] = 32'b00000000000000010011000111100011;
assign LUT_4[60837] = 32'b00000000000000001100010011011011;
assign LUT_4[60838] = 32'b00000000000000010010100010000111;
assign LUT_4[60839] = 32'b00000000000000001011101101111111;
assign LUT_4[60840] = 32'b00000000000000001111010011011100;
assign LUT_4[60841] = 32'b00000000000000001000011111010100;
assign LUT_4[60842] = 32'b00000000000000001110101110000000;
assign LUT_4[60843] = 32'b00000000000000000111111001111000;
assign LUT_4[60844] = 32'b00000000000000001100010011111000;
assign LUT_4[60845] = 32'b00000000000000000101011111110000;
assign LUT_4[60846] = 32'b00000000000000001011101110011100;
assign LUT_4[60847] = 32'b00000000000000000100111010010100;
assign LUT_4[60848] = 32'b00000000000000010011111000110101;
assign LUT_4[60849] = 32'b00000000000000001101000100101101;
assign LUT_4[60850] = 32'b00000000000000010011010011011001;
assign LUT_4[60851] = 32'b00000000000000001100011111010001;
assign LUT_4[60852] = 32'b00000000000000010000111001010001;
assign LUT_4[60853] = 32'b00000000000000001010000101001001;
assign LUT_4[60854] = 32'b00000000000000010000010011110101;
assign LUT_4[60855] = 32'b00000000000000001001011111101101;
assign LUT_4[60856] = 32'b00000000000000001101000101001010;
assign LUT_4[60857] = 32'b00000000000000000110010001000010;
assign LUT_4[60858] = 32'b00000000000000001100011111101110;
assign LUT_4[60859] = 32'b00000000000000000101101011100110;
assign LUT_4[60860] = 32'b00000000000000001010000101100110;
assign LUT_4[60861] = 32'b00000000000000000011010001011110;
assign LUT_4[60862] = 32'b00000000000000001001100000001010;
assign LUT_4[60863] = 32'b00000000000000000010101100000010;
assign LUT_4[60864] = 32'b00000000000000011001000011010100;
assign LUT_4[60865] = 32'b00000000000000010010001111001100;
assign LUT_4[60866] = 32'b00000000000000011000011101111000;
assign LUT_4[60867] = 32'b00000000000000010001101001110000;
assign LUT_4[60868] = 32'b00000000000000010110000011110000;
assign LUT_4[60869] = 32'b00000000000000001111001111101000;
assign LUT_4[60870] = 32'b00000000000000010101011110010100;
assign LUT_4[60871] = 32'b00000000000000001110101010001100;
assign LUT_4[60872] = 32'b00000000000000010010001111101001;
assign LUT_4[60873] = 32'b00000000000000001011011011100001;
assign LUT_4[60874] = 32'b00000000000000010001101010001101;
assign LUT_4[60875] = 32'b00000000000000001010110110000101;
assign LUT_4[60876] = 32'b00000000000000001111010000000101;
assign LUT_4[60877] = 32'b00000000000000001000011011111101;
assign LUT_4[60878] = 32'b00000000000000001110101010101001;
assign LUT_4[60879] = 32'b00000000000000000111110110100001;
assign LUT_4[60880] = 32'b00000000000000010110110101000010;
assign LUT_4[60881] = 32'b00000000000000010000000000111010;
assign LUT_4[60882] = 32'b00000000000000010110001111100110;
assign LUT_4[60883] = 32'b00000000000000001111011011011110;
assign LUT_4[60884] = 32'b00000000000000010011110101011110;
assign LUT_4[60885] = 32'b00000000000000001101000001010110;
assign LUT_4[60886] = 32'b00000000000000010011010000000010;
assign LUT_4[60887] = 32'b00000000000000001100011011111010;
assign LUT_4[60888] = 32'b00000000000000010000000001010111;
assign LUT_4[60889] = 32'b00000000000000001001001101001111;
assign LUT_4[60890] = 32'b00000000000000001111011011111011;
assign LUT_4[60891] = 32'b00000000000000001000100111110011;
assign LUT_4[60892] = 32'b00000000000000001101000001110011;
assign LUT_4[60893] = 32'b00000000000000000110001101101011;
assign LUT_4[60894] = 32'b00000000000000001100011100010111;
assign LUT_4[60895] = 32'b00000000000000000101101000001111;
assign LUT_4[60896] = 32'b00000000000000010111011110011011;
assign LUT_4[60897] = 32'b00000000000000010000101010010011;
assign LUT_4[60898] = 32'b00000000000000010110111000111111;
assign LUT_4[60899] = 32'b00000000000000010000000100110111;
assign LUT_4[60900] = 32'b00000000000000010100011110110111;
assign LUT_4[60901] = 32'b00000000000000001101101010101111;
assign LUT_4[60902] = 32'b00000000000000010011111001011011;
assign LUT_4[60903] = 32'b00000000000000001101000101010011;
assign LUT_4[60904] = 32'b00000000000000010000101010110000;
assign LUT_4[60905] = 32'b00000000000000001001110110101000;
assign LUT_4[60906] = 32'b00000000000000010000000101010100;
assign LUT_4[60907] = 32'b00000000000000001001010001001100;
assign LUT_4[60908] = 32'b00000000000000001101101011001100;
assign LUT_4[60909] = 32'b00000000000000000110110111000100;
assign LUT_4[60910] = 32'b00000000000000001101000101110000;
assign LUT_4[60911] = 32'b00000000000000000110010001101000;
assign LUT_4[60912] = 32'b00000000000000010101010000001001;
assign LUT_4[60913] = 32'b00000000000000001110011100000001;
assign LUT_4[60914] = 32'b00000000000000010100101010101101;
assign LUT_4[60915] = 32'b00000000000000001101110110100101;
assign LUT_4[60916] = 32'b00000000000000010010010000100101;
assign LUT_4[60917] = 32'b00000000000000001011011100011101;
assign LUT_4[60918] = 32'b00000000000000010001101011001001;
assign LUT_4[60919] = 32'b00000000000000001010110111000001;
assign LUT_4[60920] = 32'b00000000000000001110011100011110;
assign LUT_4[60921] = 32'b00000000000000000111101000010110;
assign LUT_4[60922] = 32'b00000000000000001101110111000010;
assign LUT_4[60923] = 32'b00000000000000000111000010111010;
assign LUT_4[60924] = 32'b00000000000000001011011100111010;
assign LUT_4[60925] = 32'b00000000000000000100101000110010;
assign LUT_4[60926] = 32'b00000000000000001010110111011110;
assign LUT_4[60927] = 32'b00000000000000000100000011010110;
assign LUT_4[60928] = 32'b00000000000000001111001110011101;
assign LUT_4[60929] = 32'b00000000000000001000011010010101;
assign LUT_4[60930] = 32'b00000000000000001110101001000001;
assign LUT_4[60931] = 32'b00000000000000000111110100111001;
assign LUT_4[60932] = 32'b00000000000000001100001110111001;
assign LUT_4[60933] = 32'b00000000000000000101011010110001;
assign LUT_4[60934] = 32'b00000000000000001011101001011101;
assign LUT_4[60935] = 32'b00000000000000000100110101010101;
assign LUT_4[60936] = 32'b00000000000000001000011010110010;
assign LUT_4[60937] = 32'b00000000000000000001100110101010;
assign LUT_4[60938] = 32'b00000000000000000111110101010110;
assign LUT_4[60939] = 32'b00000000000000000001000001001110;
assign LUT_4[60940] = 32'b00000000000000000101011011001110;
assign LUT_4[60941] = 32'b11111111111111111110100111000110;
assign LUT_4[60942] = 32'b00000000000000000100110101110010;
assign LUT_4[60943] = 32'b11111111111111111110000001101010;
assign LUT_4[60944] = 32'b00000000000000001101000000001011;
assign LUT_4[60945] = 32'b00000000000000000110001100000011;
assign LUT_4[60946] = 32'b00000000000000001100011010101111;
assign LUT_4[60947] = 32'b00000000000000000101100110100111;
assign LUT_4[60948] = 32'b00000000000000001010000000100111;
assign LUT_4[60949] = 32'b00000000000000000011001100011111;
assign LUT_4[60950] = 32'b00000000000000001001011011001011;
assign LUT_4[60951] = 32'b00000000000000000010100111000011;
assign LUT_4[60952] = 32'b00000000000000000110001100100000;
assign LUT_4[60953] = 32'b11111111111111111111011000011000;
assign LUT_4[60954] = 32'b00000000000000000101100111000100;
assign LUT_4[60955] = 32'b11111111111111111110110010111100;
assign LUT_4[60956] = 32'b00000000000000000011001100111100;
assign LUT_4[60957] = 32'b11111111111111111100011000110100;
assign LUT_4[60958] = 32'b00000000000000000010100111100000;
assign LUT_4[60959] = 32'b11111111111111111011110011011000;
assign LUT_4[60960] = 32'b00000000000000001101101001100100;
assign LUT_4[60961] = 32'b00000000000000000110110101011100;
assign LUT_4[60962] = 32'b00000000000000001101000100001000;
assign LUT_4[60963] = 32'b00000000000000000110010000000000;
assign LUT_4[60964] = 32'b00000000000000001010101010000000;
assign LUT_4[60965] = 32'b00000000000000000011110101111000;
assign LUT_4[60966] = 32'b00000000000000001010000100100100;
assign LUT_4[60967] = 32'b00000000000000000011010000011100;
assign LUT_4[60968] = 32'b00000000000000000110110101111001;
assign LUT_4[60969] = 32'b00000000000000000000000001110001;
assign LUT_4[60970] = 32'b00000000000000000110010000011101;
assign LUT_4[60971] = 32'b11111111111111111111011100010101;
assign LUT_4[60972] = 32'b00000000000000000011110110010101;
assign LUT_4[60973] = 32'b11111111111111111101000010001101;
assign LUT_4[60974] = 32'b00000000000000000011010000111001;
assign LUT_4[60975] = 32'b11111111111111111100011100110001;
assign LUT_4[60976] = 32'b00000000000000001011011011010010;
assign LUT_4[60977] = 32'b00000000000000000100100111001010;
assign LUT_4[60978] = 32'b00000000000000001010110101110110;
assign LUT_4[60979] = 32'b00000000000000000100000001101110;
assign LUT_4[60980] = 32'b00000000000000001000011011101110;
assign LUT_4[60981] = 32'b00000000000000000001100111100110;
assign LUT_4[60982] = 32'b00000000000000000111110110010010;
assign LUT_4[60983] = 32'b00000000000000000001000010001010;
assign LUT_4[60984] = 32'b00000000000000000100100111100111;
assign LUT_4[60985] = 32'b11111111111111111101110011011111;
assign LUT_4[60986] = 32'b00000000000000000100000010001011;
assign LUT_4[60987] = 32'b11111111111111111101001110000011;
assign LUT_4[60988] = 32'b00000000000000000001101000000011;
assign LUT_4[60989] = 32'b11111111111111111010110011111011;
assign LUT_4[60990] = 32'b00000000000000000001000010100111;
assign LUT_4[60991] = 32'b11111111111111111010001110011111;
assign LUT_4[60992] = 32'b00000000000000010000100101110001;
assign LUT_4[60993] = 32'b00000000000000001001110001101001;
assign LUT_4[60994] = 32'b00000000000000010000000000010101;
assign LUT_4[60995] = 32'b00000000000000001001001100001101;
assign LUT_4[60996] = 32'b00000000000000001101100110001101;
assign LUT_4[60997] = 32'b00000000000000000110110010000101;
assign LUT_4[60998] = 32'b00000000000000001101000000110001;
assign LUT_4[60999] = 32'b00000000000000000110001100101001;
assign LUT_4[61000] = 32'b00000000000000001001110010000110;
assign LUT_4[61001] = 32'b00000000000000000010111101111110;
assign LUT_4[61002] = 32'b00000000000000001001001100101010;
assign LUT_4[61003] = 32'b00000000000000000010011000100010;
assign LUT_4[61004] = 32'b00000000000000000110110010100010;
assign LUT_4[61005] = 32'b11111111111111111111111110011010;
assign LUT_4[61006] = 32'b00000000000000000110001101000110;
assign LUT_4[61007] = 32'b11111111111111111111011000111110;
assign LUT_4[61008] = 32'b00000000000000001110010111011111;
assign LUT_4[61009] = 32'b00000000000000000111100011010111;
assign LUT_4[61010] = 32'b00000000000000001101110010000011;
assign LUT_4[61011] = 32'b00000000000000000110111101111011;
assign LUT_4[61012] = 32'b00000000000000001011010111111011;
assign LUT_4[61013] = 32'b00000000000000000100100011110011;
assign LUT_4[61014] = 32'b00000000000000001010110010011111;
assign LUT_4[61015] = 32'b00000000000000000011111110010111;
assign LUT_4[61016] = 32'b00000000000000000111100011110100;
assign LUT_4[61017] = 32'b00000000000000000000101111101100;
assign LUT_4[61018] = 32'b00000000000000000110111110011000;
assign LUT_4[61019] = 32'b00000000000000000000001010010000;
assign LUT_4[61020] = 32'b00000000000000000100100100010000;
assign LUT_4[61021] = 32'b11111111111111111101110000001000;
assign LUT_4[61022] = 32'b00000000000000000011111110110100;
assign LUT_4[61023] = 32'b11111111111111111101001010101100;
assign LUT_4[61024] = 32'b00000000000000001111000000111000;
assign LUT_4[61025] = 32'b00000000000000001000001100110000;
assign LUT_4[61026] = 32'b00000000000000001110011011011100;
assign LUT_4[61027] = 32'b00000000000000000111100111010100;
assign LUT_4[61028] = 32'b00000000000000001100000001010100;
assign LUT_4[61029] = 32'b00000000000000000101001101001100;
assign LUT_4[61030] = 32'b00000000000000001011011011111000;
assign LUT_4[61031] = 32'b00000000000000000100100111110000;
assign LUT_4[61032] = 32'b00000000000000001000001101001101;
assign LUT_4[61033] = 32'b00000000000000000001011001000101;
assign LUT_4[61034] = 32'b00000000000000000111100111110001;
assign LUT_4[61035] = 32'b00000000000000000000110011101001;
assign LUT_4[61036] = 32'b00000000000000000101001101101001;
assign LUT_4[61037] = 32'b11111111111111111110011001100001;
assign LUT_4[61038] = 32'b00000000000000000100101000001101;
assign LUT_4[61039] = 32'b11111111111111111101110100000101;
assign LUT_4[61040] = 32'b00000000000000001100110010100110;
assign LUT_4[61041] = 32'b00000000000000000101111110011110;
assign LUT_4[61042] = 32'b00000000000000001100001101001010;
assign LUT_4[61043] = 32'b00000000000000000101011001000010;
assign LUT_4[61044] = 32'b00000000000000001001110011000010;
assign LUT_4[61045] = 32'b00000000000000000010111110111010;
assign LUT_4[61046] = 32'b00000000000000001001001101100110;
assign LUT_4[61047] = 32'b00000000000000000010011001011110;
assign LUT_4[61048] = 32'b00000000000000000101111110111011;
assign LUT_4[61049] = 32'b11111111111111111111001010110011;
assign LUT_4[61050] = 32'b00000000000000000101011001011111;
assign LUT_4[61051] = 32'b11111111111111111110100101010111;
assign LUT_4[61052] = 32'b00000000000000000010111111010111;
assign LUT_4[61053] = 32'b11111111111111111100001011001111;
assign LUT_4[61054] = 32'b00000000000000000010011001111011;
assign LUT_4[61055] = 32'b11111111111111111011100101110011;
assign LUT_4[61056] = 32'b00000000000000010001110100100101;
assign LUT_4[61057] = 32'b00000000000000001011000000011101;
assign LUT_4[61058] = 32'b00000000000000010001001111001001;
assign LUT_4[61059] = 32'b00000000000000001010011011000001;
assign LUT_4[61060] = 32'b00000000000000001110110101000001;
assign LUT_4[61061] = 32'b00000000000000001000000000111001;
assign LUT_4[61062] = 32'b00000000000000001110001111100101;
assign LUT_4[61063] = 32'b00000000000000000111011011011101;
assign LUT_4[61064] = 32'b00000000000000001011000000111010;
assign LUT_4[61065] = 32'b00000000000000000100001100110010;
assign LUT_4[61066] = 32'b00000000000000001010011011011110;
assign LUT_4[61067] = 32'b00000000000000000011100111010110;
assign LUT_4[61068] = 32'b00000000000000001000000001010110;
assign LUT_4[61069] = 32'b00000000000000000001001101001110;
assign LUT_4[61070] = 32'b00000000000000000111011011111010;
assign LUT_4[61071] = 32'b00000000000000000000100111110010;
assign LUT_4[61072] = 32'b00000000000000001111100110010011;
assign LUT_4[61073] = 32'b00000000000000001000110010001011;
assign LUT_4[61074] = 32'b00000000000000001111000000110111;
assign LUT_4[61075] = 32'b00000000000000001000001100101111;
assign LUT_4[61076] = 32'b00000000000000001100100110101111;
assign LUT_4[61077] = 32'b00000000000000000101110010100111;
assign LUT_4[61078] = 32'b00000000000000001100000001010011;
assign LUT_4[61079] = 32'b00000000000000000101001101001011;
assign LUT_4[61080] = 32'b00000000000000001000110010101000;
assign LUT_4[61081] = 32'b00000000000000000001111110100000;
assign LUT_4[61082] = 32'b00000000000000001000001101001100;
assign LUT_4[61083] = 32'b00000000000000000001011001000100;
assign LUT_4[61084] = 32'b00000000000000000101110011000100;
assign LUT_4[61085] = 32'b11111111111111111110111110111100;
assign LUT_4[61086] = 32'b00000000000000000101001101101000;
assign LUT_4[61087] = 32'b11111111111111111110011001100000;
assign LUT_4[61088] = 32'b00000000000000010000001111101100;
assign LUT_4[61089] = 32'b00000000000000001001011011100100;
assign LUT_4[61090] = 32'b00000000000000001111101010010000;
assign LUT_4[61091] = 32'b00000000000000001000110110001000;
assign LUT_4[61092] = 32'b00000000000000001101010000001000;
assign LUT_4[61093] = 32'b00000000000000000110011100000000;
assign LUT_4[61094] = 32'b00000000000000001100101010101100;
assign LUT_4[61095] = 32'b00000000000000000101110110100100;
assign LUT_4[61096] = 32'b00000000000000001001011100000001;
assign LUT_4[61097] = 32'b00000000000000000010100111111001;
assign LUT_4[61098] = 32'b00000000000000001000110110100101;
assign LUT_4[61099] = 32'b00000000000000000010000010011101;
assign LUT_4[61100] = 32'b00000000000000000110011100011101;
assign LUT_4[61101] = 32'b11111111111111111111101000010101;
assign LUT_4[61102] = 32'b00000000000000000101110111000001;
assign LUT_4[61103] = 32'b11111111111111111111000010111001;
assign LUT_4[61104] = 32'b00000000000000001110000001011010;
assign LUT_4[61105] = 32'b00000000000000000111001101010010;
assign LUT_4[61106] = 32'b00000000000000001101011011111110;
assign LUT_4[61107] = 32'b00000000000000000110100111110110;
assign LUT_4[61108] = 32'b00000000000000001011000001110110;
assign LUT_4[61109] = 32'b00000000000000000100001101101110;
assign LUT_4[61110] = 32'b00000000000000001010011100011010;
assign LUT_4[61111] = 32'b00000000000000000011101000010010;
assign LUT_4[61112] = 32'b00000000000000000111001101101111;
assign LUT_4[61113] = 32'b00000000000000000000011001100111;
assign LUT_4[61114] = 32'b00000000000000000110101000010011;
assign LUT_4[61115] = 32'b11111111111111111111110100001011;
assign LUT_4[61116] = 32'b00000000000000000100001110001011;
assign LUT_4[61117] = 32'b11111111111111111101011010000011;
assign LUT_4[61118] = 32'b00000000000000000011101000101111;
assign LUT_4[61119] = 32'b11111111111111111100110100100111;
assign LUT_4[61120] = 32'b00000000000000010011001011111001;
assign LUT_4[61121] = 32'b00000000000000001100010111110001;
assign LUT_4[61122] = 32'b00000000000000010010100110011101;
assign LUT_4[61123] = 32'b00000000000000001011110010010101;
assign LUT_4[61124] = 32'b00000000000000010000001100010101;
assign LUT_4[61125] = 32'b00000000000000001001011000001101;
assign LUT_4[61126] = 32'b00000000000000001111100110111001;
assign LUT_4[61127] = 32'b00000000000000001000110010110001;
assign LUT_4[61128] = 32'b00000000000000001100011000001110;
assign LUT_4[61129] = 32'b00000000000000000101100100000110;
assign LUT_4[61130] = 32'b00000000000000001011110010110010;
assign LUT_4[61131] = 32'b00000000000000000100111110101010;
assign LUT_4[61132] = 32'b00000000000000001001011000101010;
assign LUT_4[61133] = 32'b00000000000000000010100100100010;
assign LUT_4[61134] = 32'b00000000000000001000110011001110;
assign LUT_4[61135] = 32'b00000000000000000001111111000110;
assign LUT_4[61136] = 32'b00000000000000010000111101100111;
assign LUT_4[61137] = 32'b00000000000000001010001001011111;
assign LUT_4[61138] = 32'b00000000000000010000011000001011;
assign LUT_4[61139] = 32'b00000000000000001001100100000011;
assign LUT_4[61140] = 32'b00000000000000001101111110000011;
assign LUT_4[61141] = 32'b00000000000000000111001001111011;
assign LUT_4[61142] = 32'b00000000000000001101011000100111;
assign LUT_4[61143] = 32'b00000000000000000110100100011111;
assign LUT_4[61144] = 32'b00000000000000001010001001111100;
assign LUT_4[61145] = 32'b00000000000000000011010101110100;
assign LUT_4[61146] = 32'b00000000000000001001100100100000;
assign LUT_4[61147] = 32'b00000000000000000010110000011000;
assign LUT_4[61148] = 32'b00000000000000000111001010011000;
assign LUT_4[61149] = 32'b00000000000000000000010110010000;
assign LUT_4[61150] = 32'b00000000000000000110100100111100;
assign LUT_4[61151] = 32'b11111111111111111111110000110100;
assign LUT_4[61152] = 32'b00000000000000010001100111000000;
assign LUT_4[61153] = 32'b00000000000000001010110010111000;
assign LUT_4[61154] = 32'b00000000000000010001000001100100;
assign LUT_4[61155] = 32'b00000000000000001010001101011100;
assign LUT_4[61156] = 32'b00000000000000001110100111011100;
assign LUT_4[61157] = 32'b00000000000000000111110011010100;
assign LUT_4[61158] = 32'b00000000000000001110000010000000;
assign LUT_4[61159] = 32'b00000000000000000111001101111000;
assign LUT_4[61160] = 32'b00000000000000001010110011010101;
assign LUT_4[61161] = 32'b00000000000000000011111111001101;
assign LUT_4[61162] = 32'b00000000000000001010001101111001;
assign LUT_4[61163] = 32'b00000000000000000011011001110001;
assign LUT_4[61164] = 32'b00000000000000000111110011110001;
assign LUT_4[61165] = 32'b00000000000000000000111111101001;
assign LUT_4[61166] = 32'b00000000000000000111001110010101;
assign LUT_4[61167] = 32'b00000000000000000000011010001101;
assign LUT_4[61168] = 32'b00000000000000001111011000101110;
assign LUT_4[61169] = 32'b00000000000000001000100100100110;
assign LUT_4[61170] = 32'b00000000000000001110110011010010;
assign LUT_4[61171] = 32'b00000000000000000111111111001010;
assign LUT_4[61172] = 32'b00000000000000001100011001001010;
assign LUT_4[61173] = 32'b00000000000000000101100101000010;
assign LUT_4[61174] = 32'b00000000000000001011110011101110;
assign LUT_4[61175] = 32'b00000000000000000100111111100110;
assign LUT_4[61176] = 32'b00000000000000001000100101000011;
assign LUT_4[61177] = 32'b00000000000000000001110000111011;
assign LUT_4[61178] = 32'b00000000000000000111111111100111;
assign LUT_4[61179] = 32'b00000000000000000001001011011111;
assign LUT_4[61180] = 32'b00000000000000000101100101011111;
assign LUT_4[61181] = 32'b11111111111111111110110001010111;
assign LUT_4[61182] = 32'b00000000000000000101000000000011;
assign LUT_4[61183] = 32'b11111111111111111110001011111011;
assign LUT_4[61184] = 32'b00000000000000010100001010000000;
assign LUT_4[61185] = 32'b00000000000000001101010101111000;
assign LUT_4[61186] = 32'b00000000000000010011100100100100;
assign LUT_4[61187] = 32'b00000000000000001100110000011100;
assign LUT_4[61188] = 32'b00000000000000010001001010011100;
assign LUT_4[61189] = 32'b00000000000000001010010110010100;
assign LUT_4[61190] = 32'b00000000000000010000100101000000;
assign LUT_4[61191] = 32'b00000000000000001001110000111000;
assign LUT_4[61192] = 32'b00000000000000001101010110010101;
assign LUT_4[61193] = 32'b00000000000000000110100010001101;
assign LUT_4[61194] = 32'b00000000000000001100110000111001;
assign LUT_4[61195] = 32'b00000000000000000101111100110001;
assign LUT_4[61196] = 32'b00000000000000001010010110110001;
assign LUT_4[61197] = 32'b00000000000000000011100010101001;
assign LUT_4[61198] = 32'b00000000000000001001110001010101;
assign LUT_4[61199] = 32'b00000000000000000010111101001101;
assign LUT_4[61200] = 32'b00000000000000010001111011101110;
assign LUT_4[61201] = 32'b00000000000000001011000111100110;
assign LUT_4[61202] = 32'b00000000000000010001010110010010;
assign LUT_4[61203] = 32'b00000000000000001010100010001010;
assign LUT_4[61204] = 32'b00000000000000001110111100001010;
assign LUT_4[61205] = 32'b00000000000000001000001000000010;
assign LUT_4[61206] = 32'b00000000000000001110010110101110;
assign LUT_4[61207] = 32'b00000000000000000111100010100110;
assign LUT_4[61208] = 32'b00000000000000001011001000000011;
assign LUT_4[61209] = 32'b00000000000000000100010011111011;
assign LUT_4[61210] = 32'b00000000000000001010100010100111;
assign LUT_4[61211] = 32'b00000000000000000011101110011111;
assign LUT_4[61212] = 32'b00000000000000001000001000011111;
assign LUT_4[61213] = 32'b00000000000000000001010100010111;
assign LUT_4[61214] = 32'b00000000000000000111100011000011;
assign LUT_4[61215] = 32'b00000000000000000000101110111011;
assign LUT_4[61216] = 32'b00000000000000010010100101000111;
assign LUT_4[61217] = 32'b00000000000000001011110000111111;
assign LUT_4[61218] = 32'b00000000000000010001111111101011;
assign LUT_4[61219] = 32'b00000000000000001011001011100011;
assign LUT_4[61220] = 32'b00000000000000001111100101100011;
assign LUT_4[61221] = 32'b00000000000000001000110001011011;
assign LUT_4[61222] = 32'b00000000000000001111000000000111;
assign LUT_4[61223] = 32'b00000000000000001000001011111111;
assign LUT_4[61224] = 32'b00000000000000001011110001011100;
assign LUT_4[61225] = 32'b00000000000000000100111101010100;
assign LUT_4[61226] = 32'b00000000000000001011001100000000;
assign LUT_4[61227] = 32'b00000000000000000100010111111000;
assign LUT_4[61228] = 32'b00000000000000001000110001111000;
assign LUT_4[61229] = 32'b00000000000000000001111101110000;
assign LUT_4[61230] = 32'b00000000000000001000001100011100;
assign LUT_4[61231] = 32'b00000000000000000001011000010100;
assign LUT_4[61232] = 32'b00000000000000010000010110110101;
assign LUT_4[61233] = 32'b00000000000000001001100010101101;
assign LUT_4[61234] = 32'b00000000000000001111110001011001;
assign LUT_4[61235] = 32'b00000000000000001000111101010001;
assign LUT_4[61236] = 32'b00000000000000001101010111010001;
assign LUT_4[61237] = 32'b00000000000000000110100011001001;
assign LUT_4[61238] = 32'b00000000000000001100110001110101;
assign LUT_4[61239] = 32'b00000000000000000101111101101101;
assign LUT_4[61240] = 32'b00000000000000001001100011001010;
assign LUT_4[61241] = 32'b00000000000000000010101111000010;
assign LUT_4[61242] = 32'b00000000000000001000111101101110;
assign LUT_4[61243] = 32'b00000000000000000010001001100110;
assign LUT_4[61244] = 32'b00000000000000000110100011100110;
assign LUT_4[61245] = 32'b11111111111111111111101111011110;
assign LUT_4[61246] = 32'b00000000000000000101111110001010;
assign LUT_4[61247] = 32'b11111111111111111111001010000010;
assign LUT_4[61248] = 32'b00000000000000010101100001010100;
assign LUT_4[61249] = 32'b00000000000000001110101101001100;
assign LUT_4[61250] = 32'b00000000000000010100111011111000;
assign LUT_4[61251] = 32'b00000000000000001110000111110000;
assign LUT_4[61252] = 32'b00000000000000010010100001110000;
assign LUT_4[61253] = 32'b00000000000000001011101101101000;
assign LUT_4[61254] = 32'b00000000000000010001111100010100;
assign LUT_4[61255] = 32'b00000000000000001011001000001100;
assign LUT_4[61256] = 32'b00000000000000001110101101101001;
assign LUT_4[61257] = 32'b00000000000000000111111001100001;
assign LUT_4[61258] = 32'b00000000000000001110001000001101;
assign LUT_4[61259] = 32'b00000000000000000111010100000101;
assign LUT_4[61260] = 32'b00000000000000001011101110000101;
assign LUT_4[61261] = 32'b00000000000000000100111001111101;
assign LUT_4[61262] = 32'b00000000000000001011001000101001;
assign LUT_4[61263] = 32'b00000000000000000100010100100001;
assign LUT_4[61264] = 32'b00000000000000010011010011000010;
assign LUT_4[61265] = 32'b00000000000000001100011110111010;
assign LUT_4[61266] = 32'b00000000000000010010101101100110;
assign LUT_4[61267] = 32'b00000000000000001011111001011110;
assign LUT_4[61268] = 32'b00000000000000010000010011011110;
assign LUT_4[61269] = 32'b00000000000000001001011111010110;
assign LUT_4[61270] = 32'b00000000000000001111101110000010;
assign LUT_4[61271] = 32'b00000000000000001000111001111010;
assign LUT_4[61272] = 32'b00000000000000001100011111010111;
assign LUT_4[61273] = 32'b00000000000000000101101011001111;
assign LUT_4[61274] = 32'b00000000000000001011111001111011;
assign LUT_4[61275] = 32'b00000000000000000101000101110011;
assign LUT_4[61276] = 32'b00000000000000001001011111110011;
assign LUT_4[61277] = 32'b00000000000000000010101011101011;
assign LUT_4[61278] = 32'b00000000000000001000111010010111;
assign LUT_4[61279] = 32'b00000000000000000010000110001111;
assign LUT_4[61280] = 32'b00000000000000010011111100011011;
assign LUT_4[61281] = 32'b00000000000000001101001000010011;
assign LUT_4[61282] = 32'b00000000000000010011010110111111;
assign LUT_4[61283] = 32'b00000000000000001100100010110111;
assign LUT_4[61284] = 32'b00000000000000010000111100110111;
assign LUT_4[61285] = 32'b00000000000000001010001000101111;
assign LUT_4[61286] = 32'b00000000000000010000010111011011;
assign LUT_4[61287] = 32'b00000000000000001001100011010011;
assign LUT_4[61288] = 32'b00000000000000001101001000110000;
assign LUT_4[61289] = 32'b00000000000000000110010100101000;
assign LUT_4[61290] = 32'b00000000000000001100100011010100;
assign LUT_4[61291] = 32'b00000000000000000101101111001100;
assign LUT_4[61292] = 32'b00000000000000001010001001001100;
assign LUT_4[61293] = 32'b00000000000000000011010101000100;
assign LUT_4[61294] = 32'b00000000000000001001100011110000;
assign LUT_4[61295] = 32'b00000000000000000010101111101000;
assign LUT_4[61296] = 32'b00000000000000010001101110001001;
assign LUT_4[61297] = 32'b00000000000000001010111010000001;
assign LUT_4[61298] = 32'b00000000000000010001001000101101;
assign LUT_4[61299] = 32'b00000000000000001010010100100101;
assign LUT_4[61300] = 32'b00000000000000001110101110100101;
assign LUT_4[61301] = 32'b00000000000000000111111010011101;
assign LUT_4[61302] = 32'b00000000000000001110001001001001;
assign LUT_4[61303] = 32'b00000000000000000111010101000001;
assign LUT_4[61304] = 32'b00000000000000001010111010011110;
assign LUT_4[61305] = 32'b00000000000000000100000110010110;
assign LUT_4[61306] = 32'b00000000000000001010010101000010;
assign LUT_4[61307] = 32'b00000000000000000011100000111010;
assign LUT_4[61308] = 32'b00000000000000000111111010111010;
assign LUT_4[61309] = 32'b00000000000000000001000110110010;
assign LUT_4[61310] = 32'b00000000000000000111010101011110;
assign LUT_4[61311] = 32'b00000000000000000000100001010110;
assign LUT_4[61312] = 32'b00000000000000010110110000001000;
assign LUT_4[61313] = 32'b00000000000000001111111100000000;
assign LUT_4[61314] = 32'b00000000000000010110001010101100;
assign LUT_4[61315] = 32'b00000000000000001111010110100100;
assign LUT_4[61316] = 32'b00000000000000010011110000100100;
assign LUT_4[61317] = 32'b00000000000000001100111100011100;
assign LUT_4[61318] = 32'b00000000000000010011001011001000;
assign LUT_4[61319] = 32'b00000000000000001100010111000000;
assign LUT_4[61320] = 32'b00000000000000001111111100011101;
assign LUT_4[61321] = 32'b00000000000000001001001000010101;
assign LUT_4[61322] = 32'b00000000000000001111010111000001;
assign LUT_4[61323] = 32'b00000000000000001000100010111001;
assign LUT_4[61324] = 32'b00000000000000001100111100111001;
assign LUT_4[61325] = 32'b00000000000000000110001000110001;
assign LUT_4[61326] = 32'b00000000000000001100010111011101;
assign LUT_4[61327] = 32'b00000000000000000101100011010101;
assign LUT_4[61328] = 32'b00000000000000010100100001110110;
assign LUT_4[61329] = 32'b00000000000000001101101101101110;
assign LUT_4[61330] = 32'b00000000000000010011111100011010;
assign LUT_4[61331] = 32'b00000000000000001101001000010010;
assign LUT_4[61332] = 32'b00000000000000010001100010010010;
assign LUT_4[61333] = 32'b00000000000000001010101110001010;
assign LUT_4[61334] = 32'b00000000000000010000111100110110;
assign LUT_4[61335] = 32'b00000000000000001010001000101110;
assign LUT_4[61336] = 32'b00000000000000001101101110001011;
assign LUT_4[61337] = 32'b00000000000000000110111010000011;
assign LUT_4[61338] = 32'b00000000000000001101001000101111;
assign LUT_4[61339] = 32'b00000000000000000110010100100111;
assign LUT_4[61340] = 32'b00000000000000001010101110100111;
assign LUT_4[61341] = 32'b00000000000000000011111010011111;
assign LUT_4[61342] = 32'b00000000000000001010001001001011;
assign LUT_4[61343] = 32'b00000000000000000011010101000011;
assign LUT_4[61344] = 32'b00000000000000010101001011001111;
assign LUT_4[61345] = 32'b00000000000000001110010111000111;
assign LUT_4[61346] = 32'b00000000000000010100100101110011;
assign LUT_4[61347] = 32'b00000000000000001101110001101011;
assign LUT_4[61348] = 32'b00000000000000010010001011101011;
assign LUT_4[61349] = 32'b00000000000000001011010111100011;
assign LUT_4[61350] = 32'b00000000000000010001100110001111;
assign LUT_4[61351] = 32'b00000000000000001010110010000111;
assign LUT_4[61352] = 32'b00000000000000001110010111100100;
assign LUT_4[61353] = 32'b00000000000000000111100011011100;
assign LUT_4[61354] = 32'b00000000000000001101110010001000;
assign LUT_4[61355] = 32'b00000000000000000110111110000000;
assign LUT_4[61356] = 32'b00000000000000001011011000000000;
assign LUT_4[61357] = 32'b00000000000000000100100011111000;
assign LUT_4[61358] = 32'b00000000000000001010110010100100;
assign LUT_4[61359] = 32'b00000000000000000011111110011100;
assign LUT_4[61360] = 32'b00000000000000010010111100111101;
assign LUT_4[61361] = 32'b00000000000000001100001000110101;
assign LUT_4[61362] = 32'b00000000000000010010010111100001;
assign LUT_4[61363] = 32'b00000000000000001011100011011001;
assign LUT_4[61364] = 32'b00000000000000001111111101011001;
assign LUT_4[61365] = 32'b00000000000000001001001001010001;
assign LUT_4[61366] = 32'b00000000000000001111010111111101;
assign LUT_4[61367] = 32'b00000000000000001000100011110101;
assign LUT_4[61368] = 32'b00000000000000001100001001010010;
assign LUT_4[61369] = 32'b00000000000000000101010101001010;
assign LUT_4[61370] = 32'b00000000000000001011100011110110;
assign LUT_4[61371] = 32'b00000000000000000100101111101110;
assign LUT_4[61372] = 32'b00000000000000001001001001101110;
assign LUT_4[61373] = 32'b00000000000000000010010101100110;
assign LUT_4[61374] = 32'b00000000000000001000100100010010;
assign LUT_4[61375] = 32'b00000000000000000001110000001010;
assign LUT_4[61376] = 32'b00000000000000011000000111011100;
assign LUT_4[61377] = 32'b00000000000000010001010011010100;
assign LUT_4[61378] = 32'b00000000000000010111100010000000;
assign LUT_4[61379] = 32'b00000000000000010000101101111000;
assign LUT_4[61380] = 32'b00000000000000010101000111111000;
assign LUT_4[61381] = 32'b00000000000000001110010011110000;
assign LUT_4[61382] = 32'b00000000000000010100100010011100;
assign LUT_4[61383] = 32'b00000000000000001101101110010100;
assign LUT_4[61384] = 32'b00000000000000010001010011110001;
assign LUT_4[61385] = 32'b00000000000000001010011111101001;
assign LUT_4[61386] = 32'b00000000000000010000101110010101;
assign LUT_4[61387] = 32'b00000000000000001001111010001101;
assign LUT_4[61388] = 32'b00000000000000001110010100001101;
assign LUT_4[61389] = 32'b00000000000000000111100000000101;
assign LUT_4[61390] = 32'b00000000000000001101101110110001;
assign LUT_4[61391] = 32'b00000000000000000110111010101001;
assign LUT_4[61392] = 32'b00000000000000010101111001001010;
assign LUT_4[61393] = 32'b00000000000000001111000101000010;
assign LUT_4[61394] = 32'b00000000000000010101010011101110;
assign LUT_4[61395] = 32'b00000000000000001110011111100110;
assign LUT_4[61396] = 32'b00000000000000010010111001100110;
assign LUT_4[61397] = 32'b00000000000000001100000101011110;
assign LUT_4[61398] = 32'b00000000000000010010010100001010;
assign LUT_4[61399] = 32'b00000000000000001011100000000010;
assign LUT_4[61400] = 32'b00000000000000001111000101011111;
assign LUT_4[61401] = 32'b00000000000000001000010001010111;
assign LUT_4[61402] = 32'b00000000000000001110100000000011;
assign LUT_4[61403] = 32'b00000000000000000111101011111011;
assign LUT_4[61404] = 32'b00000000000000001100000101111011;
assign LUT_4[61405] = 32'b00000000000000000101010001110011;
assign LUT_4[61406] = 32'b00000000000000001011100000011111;
assign LUT_4[61407] = 32'b00000000000000000100101100010111;
assign LUT_4[61408] = 32'b00000000000000010110100010100011;
assign LUT_4[61409] = 32'b00000000000000001111101110011011;
assign LUT_4[61410] = 32'b00000000000000010101111101000111;
assign LUT_4[61411] = 32'b00000000000000001111001000111111;
assign LUT_4[61412] = 32'b00000000000000010011100010111111;
assign LUT_4[61413] = 32'b00000000000000001100101110110111;
assign LUT_4[61414] = 32'b00000000000000010010111101100011;
assign LUT_4[61415] = 32'b00000000000000001100001001011011;
assign LUT_4[61416] = 32'b00000000000000001111101110111000;
assign LUT_4[61417] = 32'b00000000000000001000111010110000;
assign LUT_4[61418] = 32'b00000000000000001111001001011100;
assign LUT_4[61419] = 32'b00000000000000001000010101010100;
assign LUT_4[61420] = 32'b00000000000000001100101111010100;
assign LUT_4[61421] = 32'b00000000000000000101111011001100;
assign LUT_4[61422] = 32'b00000000000000001100001001111000;
assign LUT_4[61423] = 32'b00000000000000000101010101110000;
assign LUT_4[61424] = 32'b00000000000000010100010100010001;
assign LUT_4[61425] = 32'b00000000000000001101100000001001;
assign LUT_4[61426] = 32'b00000000000000010011101110110101;
assign LUT_4[61427] = 32'b00000000000000001100111010101101;
assign LUT_4[61428] = 32'b00000000000000010001010100101101;
assign LUT_4[61429] = 32'b00000000000000001010100000100101;
assign LUT_4[61430] = 32'b00000000000000010000101111010001;
assign LUT_4[61431] = 32'b00000000000000001001111011001001;
assign LUT_4[61432] = 32'b00000000000000001101100000100110;
assign LUT_4[61433] = 32'b00000000000000000110101100011110;
assign LUT_4[61434] = 32'b00000000000000001100111011001010;
assign LUT_4[61435] = 32'b00000000000000000110000111000010;
assign LUT_4[61436] = 32'b00000000000000001010100001000010;
assign LUT_4[61437] = 32'b00000000000000000011101100111010;
assign LUT_4[61438] = 32'b00000000000000001001111011100110;
assign LUT_4[61439] = 32'b00000000000000000011000111011110;
assign LUT_4[61440] = 32'b00000000000000001111010000011101;
assign LUT_4[61441] = 32'b00000000000000001000011100010101;
assign LUT_4[61442] = 32'b00000000000000001110101011000001;
assign LUT_4[61443] = 32'b00000000000000000111110110111001;
assign LUT_4[61444] = 32'b00000000000000001100010000111001;
assign LUT_4[61445] = 32'b00000000000000000101011100110001;
assign LUT_4[61446] = 32'b00000000000000001011101011011101;
assign LUT_4[61447] = 32'b00000000000000000100110111010101;
assign LUT_4[61448] = 32'b00000000000000001000011100110010;
assign LUT_4[61449] = 32'b00000000000000000001101000101010;
assign LUT_4[61450] = 32'b00000000000000000111110111010110;
assign LUT_4[61451] = 32'b00000000000000000001000011001110;
assign LUT_4[61452] = 32'b00000000000000000101011101001110;
assign LUT_4[61453] = 32'b11111111111111111110101001000110;
assign LUT_4[61454] = 32'b00000000000000000100110111110010;
assign LUT_4[61455] = 32'b11111111111111111110000011101010;
assign LUT_4[61456] = 32'b00000000000000001101000010001011;
assign LUT_4[61457] = 32'b00000000000000000110001110000011;
assign LUT_4[61458] = 32'b00000000000000001100011100101111;
assign LUT_4[61459] = 32'b00000000000000000101101000100111;
assign LUT_4[61460] = 32'b00000000000000001010000010100111;
assign LUT_4[61461] = 32'b00000000000000000011001110011111;
assign LUT_4[61462] = 32'b00000000000000001001011101001011;
assign LUT_4[61463] = 32'b00000000000000000010101001000011;
assign LUT_4[61464] = 32'b00000000000000000110001110100000;
assign LUT_4[61465] = 32'b11111111111111111111011010011000;
assign LUT_4[61466] = 32'b00000000000000000101101001000100;
assign LUT_4[61467] = 32'b11111111111111111110110100111100;
assign LUT_4[61468] = 32'b00000000000000000011001110111100;
assign LUT_4[61469] = 32'b11111111111111111100011010110100;
assign LUT_4[61470] = 32'b00000000000000000010101001100000;
assign LUT_4[61471] = 32'b11111111111111111011110101011000;
assign LUT_4[61472] = 32'b00000000000000001101101011100100;
assign LUT_4[61473] = 32'b00000000000000000110110111011100;
assign LUT_4[61474] = 32'b00000000000000001101000110001000;
assign LUT_4[61475] = 32'b00000000000000000110010010000000;
assign LUT_4[61476] = 32'b00000000000000001010101100000000;
assign LUT_4[61477] = 32'b00000000000000000011110111111000;
assign LUT_4[61478] = 32'b00000000000000001010000110100100;
assign LUT_4[61479] = 32'b00000000000000000011010010011100;
assign LUT_4[61480] = 32'b00000000000000000110110111111001;
assign LUT_4[61481] = 32'b00000000000000000000000011110001;
assign LUT_4[61482] = 32'b00000000000000000110010010011101;
assign LUT_4[61483] = 32'b11111111111111111111011110010101;
assign LUT_4[61484] = 32'b00000000000000000011111000010101;
assign LUT_4[61485] = 32'b11111111111111111101000100001101;
assign LUT_4[61486] = 32'b00000000000000000011010010111001;
assign LUT_4[61487] = 32'b11111111111111111100011110110001;
assign LUT_4[61488] = 32'b00000000000000001011011101010010;
assign LUT_4[61489] = 32'b00000000000000000100101001001010;
assign LUT_4[61490] = 32'b00000000000000001010110111110110;
assign LUT_4[61491] = 32'b00000000000000000100000011101110;
assign LUT_4[61492] = 32'b00000000000000001000011101101110;
assign LUT_4[61493] = 32'b00000000000000000001101001100110;
assign LUT_4[61494] = 32'b00000000000000000111111000010010;
assign LUT_4[61495] = 32'b00000000000000000001000100001010;
assign LUT_4[61496] = 32'b00000000000000000100101001100111;
assign LUT_4[61497] = 32'b11111111111111111101110101011111;
assign LUT_4[61498] = 32'b00000000000000000100000100001011;
assign LUT_4[61499] = 32'b11111111111111111101010000000011;
assign LUT_4[61500] = 32'b00000000000000000001101010000011;
assign LUT_4[61501] = 32'b11111111111111111010110101111011;
assign LUT_4[61502] = 32'b00000000000000000001000100100111;
assign LUT_4[61503] = 32'b11111111111111111010010000011111;
assign LUT_4[61504] = 32'b00000000000000010000100111110001;
assign LUT_4[61505] = 32'b00000000000000001001110011101001;
assign LUT_4[61506] = 32'b00000000000000010000000010010101;
assign LUT_4[61507] = 32'b00000000000000001001001110001101;
assign LUT_4[61508] = 32'b00000000000000001101101000001101;
assign LUT_4[61509] = 32'b00000000000000000110110100000101;
assign LUT_4[61510] = 32'b00000000000000001101000010110001;
assign LUT_4[61511] = 32'b00000000000000000110001110101001;
assign LUT_4[61512] = 32'b00000000000000001001110100000110;
assign LUT_4[61513] = 32'b00000000000000000010111111111110;
assign LUT_4[61514] = 32'b00000000000000001001001110101010;
assign LUT_4[61515] = 32'b00000000000000000010011010100010;
assign LUT_4[61516] = 32'b00000000000000000110110100100010;
assign LUT_4[61517] = 32'b00000000000000000000000000011010;
assign LUT_4[61518] = 32'b00000000000000000110001111000110;
assign LUT_4[61519] = 32'b11111111111111111111011010111110;
assign LUT_4[61520] = 32'b00000000000000001110011001011111;
assign LUT_4[61521] = 32'b00000000000000000111100101010111;
assign LUT_4[61522] = 32'b00000000000000001101110100000011;
assign LUT_4[61523] = 32'b00000000000000000110111111111011;
assign LUT_4[61524] = 32'b00000000000000001011011001111011;
assign LUT_4[61525] = 32'b00000000000000000100100101110011;
assign LUT_4[61526] = 32'b00000000000000001010110100011111;
assign LUT_4[61527] = 32'b00000000000000000100000000010111;
assign LUT_4[61528] = 32'b00000000000000000111100101110100;
assign LUT_4[61529] = 32'b00000000000000000000110001101100;
assign LUT_4[61530] = 32'b00000000000000000111000000011000;
assign LUT_4[61531] = 32'b00000000000000000000001100010000;
assign LUT_4[61532] = 32'b00000000000000000100100110010000;
assign LUT_4[61533] = 32'b11111111111111111101110010001000;
assign LUT_4[61534] = 32'b00000000000000000100000000110100;
assign LUT_4[61535] = 32'b11111111111111111101001100101100;
assign LUT_4[61536] = 32'b00000000000000001111000010111000;
assign LUT_4[61537] = 32'b00000000000000001000001110110000;
assign LUT_4[61538] = 32'b00000000000000001110011101011100;
assign LUT_4[61539] = 32'b00000000000000000111101001010100;
assign LUT_4[61540] = 32'b00000000000000001100000011010100;
assign LUT_4[61541] = 32'b00000000000000000101001111001100;
assign LUT_4[61542] = 32'b00000000000000001011011101111000;
assign LUT_4[61543] = 32'b00000000000000000100101001110000;
assign LUT_4[61544] = 32'b00000000000000001000001111001101;
assign LUT_4[61545] = 32'b00000000000000000001011011000101;
assign LUT_4[61546] = 32'b00000000000000000111101001110001;
assign LUT_4[61547] = 32'b00000000000000000000110101101001;
assign LUT_4[61548] = 32'b00000000000000000101001111101001;
assign LUT_4[61549] = 32'b11111111111111111110011011100001;
assign LUT_4[61550] = 32'b00000000000000000100101010001101;
assign LUT_4[61551] = 32'b11111111111111111101110110000101;
assign LUT_4[61552] = 32'b00000000000000001100110100100110;
assign LUT_4[61553] = 32'b00000000000000000110000000011110;
assign LUT_4[61554] = 32'b00000000000000001100001111001010;
assign LUT_4[61555] = 32'b00000000000000000101011011000010;
assign LUT_4[61556] = 32'b00000000000000001001110101000010;
assign LUT_4[61557] = 32'b00000000000000000011000000111010;
assign LUT_4[61558] = 32'b00000000000000001001001111100110;
assign LUT_4[61559] = 32'b00000000000000000010011011011110;
assign LUT_4[61560] = 32'b00000000000000000110000000111011;
assign LUT_4[61561] = 32'b11111111111111111111001100110011;
assign LUT_4[61562] = 32'b00000000000000000101011011011111;
assign LUT_4[61563] = 32'b11111111111111111110100111010111;
assign LUT_4[61564] = 32'b00000000000000000011000001010111;
assign LUT_4[61565] = 32'b11111111111111111100001101001111;
assign LUT_4[61566] = 32'b00000000000000000010011011111011;
assign LUT_4[61567] = 32'b11111111111111111011100111110011;
assign LUT_4[61568] = 32'b00000000000000010001110110100101;
assign LUT_4[61569] = 32'b00000000000000001011000010011101;
assign LUT_4[61570] = 32'b00000000000000010001010001001001;
assign LUT_4[61571] = 32'b00000000000000001010011101000001;
assign LUT_4[61572] = 32'b00000000000000001110110111000001;
assign LUT_4[61573] = 32'b00000000000000001000000010111001;
assign LUT_4[61574] = 32'b00000000000000001110010001100101;
assign LUT_4[61575] = 32'b00000000000000000111011101011101;
assign LUT_4[61576] = 32'b00000000000000001011000010111010;
assign LUT_4[61577] = 32'b00000000000000000100001110110010;
assign LUT_4[61578] = 32'b00000000000000001010011101011110;
assign LUT_4[61579] = 32'b00000000000000000011101001010110;
assign LUT_4[61580] = 32'b00000000000000001000000011010110;
assign LUT_4[61581] = 32'b00000000000000000001001111001110;
assign LUT_4[61582] = 32'b00000000000000000111011101111010;
assign LUT_4[61583] = 32'b00000000000000000000101001110010;
assign LUT_4[61584] = 32'b00000000000000001111101000010011;
assign LUT_4[61585] = 32'b00000000000000001000110100001011;
assign LUT_4[61586] = 32'b00000000000000001111000010110111;
assign LUT_4[61587] = 32'b00000000000000001000001110101111;
assign LUT_4[61588] = 32'b00000000000000001100101000101111;
assign LUT_4[61589] = 32'b00000000000000000101110100100111;
assign LUT_4[61590] = 32'b00000000000000001100000011010011;
assign LUT_4[61591] = 32'b00000000000000000101001111001011;
assign LUT_4[61592] = 32'b00000000000000001000110100101000;
assign LUT_4[61593] = 32'b00000000000000000010000000100000;
assign LUT_4[61594] = 32'b00000000000000001000001111001100;
assign LUT_4[61595] = 32'b00000000000000000001011011000100;
assign LUT_4[61596] = 32'b00000000000000000101110101000100;
assign LUT_4[61597] = 32'b11111111111111111111000000111100;
assign LUT_4[61598] = 32'b00000000000000000101001111101000;
assign LUT_4[61599] = 32'b11111111111111111110011011100000;
assign LUT_4[61600] = 32'b00000000000000010000010001101100;
assign LUT_4[61601] = 32'b00000000000000001001011101100100;
assign LUT_4[61602] = 32'b00000000000000001111101100010000;
assign LUT_4[61603] = 32'b00000000000000001000111000001000;
assign LUT_4[61604] = 32'b00000000000000001101010010001000;
assign LUT_4[61605] = 32'b00000000000000000110011110000000;
assign LUT_4[61606] = 32'b00000000000000001100101100101100;
assign LUT_4[61607] = 32'b00000000000000000101111000100100;
assign LUT_4[61608] = 32'b00000000000000001001011110000001;
assign LUT_4[61609] = 32'b00000000000000000010101001111001;
assign LUT_4[61610] = 32'b00000000000000001000111000100101;
assign LUT_4[61611] = 32'b00000000000000000010000100011101;
assign LUT_4[61612] = 32'b00000000000000000110011110011101;
assign LUT_4[61613] = 32'b11111111111111111111101010010101;
assign LUT_4[61614] = 32'b00000000000000000101111001000001;
assign LUT_4[61615] = 32'b11111111111111111111000100111001;
assign LUT_4[61616] = 32'b00000000000000001110000011011010;
assign LUT_4[61617] = 32'b00000000000000000111001111010010;
assign LUT_4[61618] = 32'b00000000000000001101011101111110;
assign LUT_4[61619] = 32'b00000000000000000110101001110110;
assign LUT_4[61620] = 32'b00000000000000001011000011110110;
assign LUT_4[61621] = 32'b00000000000000000100001111101110;
assign LUT_4[61622] = 32'b00000000000000001010011110011010;
assign LUT_4[61623] = 32'b00000000000000000011101010010010;
assign LUT_4[61624] = 32'b00000000000000000111001111101111;
assign LUT_4[61625] = 32'b00000000000000000000011011100111;
assign LUT_4[61626] = 32'b00000000000000000110101010010011;
assign LUT_4[61627] = 32'b11111111111111111111110110001011;
assign LUT_4[61628] = 32'b00000000000000000100010000001011;
assign LUT_4[61629] = 32'b11111111111111111101011100000011;
assign LUT_4[61630] = 32'b00000000000000000011101010101111;
assign LUT_4[61631] = 32'b11111111111111111100110110100111;
assign LUT_4[61632] = 32'b00000000000000010011001101111001;
assign LUT_4[61633] = 32'b00000000000000001100011001110001;
assign LUT_4[61634] = 32'b00000000000000010010101000011101;
assign LUT_4[61635] = 32'b00000000000000001011110100010101;
assign LUT_4[61636] = 32'b00000000000000010000001110010101;
assign LUT_4[61637] = 32'b00000000000000001001011010001101;
assign LUT_4[61638] = 32'b00000000000000001111101000111001;
assign LUT_4[61639] = 32'b00000000000000001000110100110001;
assign LUT_4[61640] = 32'b00000000000000001100011010001110;
assign LUT_4[61641] = 32'b00000000000000000101100110000110;
assign LUT_4[61642] = 32'b00000000000000001011110100110010;
assign LUT_4[61643] = 32'b00000000000000000101000000101010;
assign LUT_4[61644] = 32'b00000000000000001001011010101010;
assign LUT_4[61645] = 32'b00000000000000000010100110100010;
assign LUT_4[61646] = 32'b00000000000000001000110101001110;
assign LUT_4[61647] = 32'b00000000000000000010000001000110;
assign LUT_4[61648] = 32'b00000000000000010000111111100111;
assign LUT_4[61649] = 32'b00000000000000001010001011011111;
assign LUT_4[61650] = 32'b00000000000000010000011010001011;
assign LUT_4[61651] = 32'b00000000000000001001100110000011;
assign LUT_4[61652] = 32'b00000000000000001110000000000011;
assign LUT_4[61653] = 32'b00000000000000000111001011111011;
assign LUT_4[61654] = 32'b00000000000000001101011010100111;
assign LUT_4[61655] = 32'b00000000000000000110100110011111;
assign LUT_4[61656] = 32'b00000000000000001010001011111100;
assign LUT_4[61657] = 32'b00000000000000000011010111110100;
assign LUT_4[61658] = 32'b00000000000000001001100110100000;
assign LUT_4[61659] = 32'b00000000000000000010110010011000;
assign LUT_4[61660] = 32'b00000000000000000111001100011000;
assign LUT_4[61661] = 32'b00000000000000000000011000010000;
assign LUT_4[61662] = 32'b00000000000000000110100110111100;
assign LUT_4[61663] = 32'b11111111111111111111110010110100;
assign LUT_4[61664] = 32'b00000000000000010001101001000000;
assign LUT_4[61665] = 32'b00000000000000001010110100111000;
assign LUT_4[61666] = 32'b00000000000000010001000011100100;
assign LUT_4[61667] = 32'b00000000000000001010001111011100;
assign LUT_4[61668] = 32'b00000000000000001110101001011100;
assign LUT_4[61669] = 32'b00000000000000000111110101010100;
assign LUT_4[61670] = 32'b00000000000000001110000100000000;
assign LUT_4[61671] = 32'b00000000000000000111001111111000;
assign LUT_4[61672] = 32'b00000000000000001010110101010101;
assign LUT_4[61673] = 32'b00000000000000000100000001001101;
assign LUT_4[61674] = 32'b00000000000000001010001111111001;
assign LUT_4[61675] = 32'b00000000000000000011011011110001;
assign LUT_4[61676] = 32'b00000000000000000111110101110001;
assign LUT_4[61677] = 32'b00000000000000000001000001101001;
assign LUT_4[61678] = 32'b00000000000000000111010000010101;
assign LUT_4[61679] = 32'b00000000000000000000011100001101;
assign LUT_4[61680] = 32'b00000000000000001111011010101110;
assign LUT_4[61681] = 32'b00000000000000001000100110100110;
assign LUT_4[61682] = 32'b00000000000000001110110101010010;
assign LUT_4[61683] = 32'b00000000000000001000000001001010;
assign LUT_4[61684] = 32'b00000000000000001100011011001010;
assign LUT_4[61685] = 32'b00000000000000000101100111000010;
assign LUT_4[61686] = 32'b00000000000000001011110101101110;
assign LUT_4[61687] = 32'b00000000000000000101000001100110;
assign LUT_4[61688] = 32'b00000000000000001000100111000011;
assign LUT_4[61689] = 32'b00000000000000000001110010111011;
assign LUT_4[61690] = 32'b00000000000000001000000001100111;
assign LUT_4[61691] = 32'b00000000000000000001001101011111;
assign LUT_4[61692] = 32'b00000000000000000101100111011111;
assign LUT_4[61693] = 32'b11111111111111111110110011010111;
assign LUT_4[61694] = 32'b00000000000000000101000010000011;
assign LUT_4[61695] = 32'b11111111111111111110001101111011;
assign LUT_4[61696] = 32'b00000000000000010100001100000000;
assign LUT_4[61697] = 32'b00000000000000001101010111111000;
assign LUT_4[61698] = 32'b00000000000000010011100110100100;
assign LUT_4[61699] = 32'b00000000000000001100110010011100;
assign LUT_4[61700] = 32'b00000000000000010001001100011100;
assign LUT_4[61701] = 32'b00000000000000001010011000010100;
assign LUT_4[61702] = 32'b00000000000000010000100111000000;
assign LUT_4[61703] = 32'b00000000000000001001110010111000;
assign LUT_4[61704] = 32'b00000000000000001101011000010101;
assign LUT_4[61705] = 32'b00000000000000000110100100001101;
assign LUT_4[61706] = 32'b00000000000000001100110010111001;
assign LUT_4[61707] = 32'b00000000000000000101111110110001;
assign LUT_4[61708] = 32'b00000000000000001010011000110001;
assign LUT_4[61709] = 32'b00000000000000000011100100101001;
assign LUT_4[61710] = 32'b00000000000000001001110011010101;
assign LUT_4[61711] = 32'b00000000000000000010111111001101;
assign LUT_4[61712] = 32'b00000000000000010001111101101110;
assign LUT_4[61713] = 32'b00000000000000001011001001100110;
assign LUT_4[61714] = 32'b00000000000000010001011000010010;
assign LUT_4[61715] = 32'b00000000000000001010100100001010;
assign LUT_4[61716] = 32'b00000000000000001110111110001010;
assign LUT_4[61717] = 32'b00000000000000001000001010000010;
assign LUT_4[61718] = 32'b00000000000000001110011000101110;
assign LUT_4[61719] = 32'b00000000000000000111100100100110;
assign LUT_4[61720] = 32'b00000000000000001011001010000011;
assign LUT_4[61721] = 32'b00000000000000000100010101111011;
assign LUT_4[61722] = 32'b00000000000000001010100100100111;
assign LUT_4[61723] = 32'b00000000000000000011110000011111;
assign LUT_4[61724] = 32'b00000000000000001000001010011111;
assign LUT_4[61725] = 32'b00000000000000000001010110010111;
assign LUT_4[61726] = 32'b00000000000000000111100101000011;
assign LUT_4[61727] = 32'b00000000000000000000110000111011;
assign LUT_4[61728] = 32'b00000000000000010010100111000111;
assign LUT_4[61729] = 32'b00000000000000001011110010111111;
assign LUT_4[61730] = 32'b00000000000000010010000001101011;
assign LUT_4[61731] = 32'b00000000000000001011001101100011;
assign LUT_4[61732] = 32'b00000000000000001111100111100011;
assign LUT_4[61733] = 32'b00000000000000001000110011011011;
assign LUT_4[61734] = 32'b00000000000000001111000010000111;
assign LUT_4[61735] = 32'b00000000000000001000001101111111;
assign LUT_4[61736] = 32'b00000000000000001011110011011100;
assign LUT_4[61737] = 32'b00000000000000000100111111010100;
assign LUT_4[61738] = 32'b00000000000000001011001110000000;
assign LUT_4[61739] = 32'b00000000000000000100011001111000;
assign LUT_4[61740] = 32'b00000000000000001000110011111000;
assign LUT_4[61741] = 32'b00000000000000000001111111110000;
assign LUT_4[61742] = 32'b00000000000000001000001110011100;
assign LUT_4[61743] = 32'b00000000000000000001011010010100;
assign LUT_4[61744] = 32'b00000000000000010000011000110101;
assign LUT_4[61745] = 32'b00000000000000001001100100101101;
assign LUT_4[61746] = 32'b00000000000000001111110011011001;
assign LUT_4[61747] = 32'b00000000000000001000111111010001;
assign LUT_4[61748] = 32'b00000000000000001101011001010001;
assign LUT_4[61749] = 32'b00000000000000000110100101001001;
assign LUT_4[61750] = 32'b00000000000000001100110011110101;
assign LUT_4[61751] = 32'b00000000000000000101111111101101;
assign LUT_4[61752] = 32'b00000000000000001001100101001010;
assign LUT_4[61753] = 32'b00000000000000000010110001000010;
assign LUT_4[61754] = 32'b00000000000000001000111111101110;
assign LUT_4[61755] = 32'b00000000000000000010001011100110;
assign LUT_4[61756] = 32'b00000000000000000110100101100110;
assign LUT_4[61757] = 32'b11111111111111111111110001011110;
assign LUT_4[61758] = 32'b00000000000000000110000000001010;
assign LUT_4[61759] = 32'b11111111111111111111001100000010;
assign LUT_4[61760] = 32'b00000000000000010101100011010100;
assign LUT_4[61761] = 32'b00000000000000001110101111001100;
assign LUT_4[61762] = 32'b00000000000000010100111101111000;
assign LUT_4[61763] = 32'b00000000000000001110001001110000;
assign LUT_4[61764] = 32'b00000000000000010010100011110000;
assign LUT_4[61765] = 32'b00000000000000001011101111101000;
assign LUT_4[61766] = 32'b00000000000000010001111110010100;
assign LUT_4[61767] = 32'b00000000000000001011001010001100;
assign LUT_4[61768] = 32'b00000000000000001110101111101001;
assign LUT_4[61769] = 32'b00000000000000000111111011100001;
assign LUT_4[61770] = 32'b00000000000000001110001010001101;
assign LUT_4[61771] = 32'b00000000000000000111010110000101;
assign LUT_4[61772] = 32'b00000000000000001011110000000101;
assign LUT_4[61773] = 32'b00000000000000000100111011111101;
assign LUT_4[61774] = 32'b00000000000000001011001010101001;
assign LUT_4[61775] = 32'b00000000000000000100010110100001;
assign LUT_4[61776] = 32'b00000000000000010011010101000010;
assign LUT_4[61777] = 32'b00000000000000001100100000111010;
assign LUT_4[61778] = 32'b00000000000000010010101111100110;
assign LUT_4[61779] = 32'b00000000000000001011111011011110;
assign LUT_4[61780] = 32'b00000000000000010000010101011110;
assign LUT_4[61781] = 32'b00000000000000001001100001010110;
assign LUT_4[61782] = 32'b00000000000000001111110000000010;
assign LUT_4[61783] = 32'b00000000000000001000111011111010;
assign LUT_4[61784] = 32'b00000000000000001100100001010111;
assign LUT_4[61785] = 32'b00000000000000000101101101001111;
assign LUT_4[61786] = 32'b00000000000000001011111011111011;
assign LUT_4[61787] = 32'b00000000000000000101000111110011;
assign LUT_4[61788] = 32'b00000000000000001001100001110011;
assign LUT_4[61789] = 32'b00000000000000000010101101101011;
assign LUT_4[61790] = 32'b00000000000000001000111100010111;
assign LUT_4[61791] = 32'b00000000000000000010001000001111;
assign LUT_4[61792] = 32'b00000000000000010011111110011011;
assign LUT_4[61793] = 32'b00000000000000001101001010010011;
assign LUT_4[61794] = 32'b00000000000000010011011000111111;
assign LUT_4[61795] = 32'b00000000000000001100100100110111;
assign LUT_4[61796] = 32'b00000000000000010000111110110111;
assign LUT_4[61797] = 32'b00000000000000001010001010101111;
assign LUT_4[61798] = 32'b00000000000000010000011001011011;
assign LUT_4[61799] = 32'b00000000000000001001100101010011;
assign LUT_4[61800] = 32'b00000000000000001101001010110000;
assign LUT_4[61801] = 32'b00000000000000000110010110101000;
assign LUT_4[61802] = 32'b00000000000000001100100101010100;
assign LUT_4[61803] = 32'b00000000000000000101110001001100;
assign LUT_4[61804] = 32'b00000000000000001010001011001100;
assign LUT_4[61805] = 32'b00000000000000000011010111000100;
assign LUT_4[61806] = 32'b00000000000000001001100101110000;
assign LUT_4[61807] = 32'b00000000000000000010110001101000;
assign LUT_4[61808] = 32'b00000000000000010001110000001001;
assign LUT_4[61809] = 32'b00000000000000001010111100000001;
assign LUT_4[61810] = 32'b00000000000000010001001010101101;
assign LUT_4[61811] = 32'b00000000000000001010010110100101;
assign LUT_4[61812] = 32'b00000000000000001110110000100101;
assign LUT_4[61813] = 32'b00000000000000000111111100011101;
assign LUT_4[61814] = 32'b00000000000000001110001011001001;
assign LUT_4[61815] = 32'b00000000000000000111010111000001;
assign LUT_4[61816] = 32'b00000000000000001010111100011110;
assign LUT_4[61817] = 32'b00000000000000000100001000010110;
assign LUT_4[61818] = 32'b00000000000000001010010111000010;
assign LUT_4[61819] = 32'b00000000000000000011100010111010;
assign LUT_4[61820] = 32'b00000000000000000111111100111010;
assign LUT_4[61821] = 32'b00000000000000000001001000110010;
assign LUT_4[61822] = 32'b00000000000000000111010111011110;
assign LUT_4[61823] = 32'b00000000000000000000100011010110;
assign LUT_4[61824] = 32'b00000000000000010110110010001000;
assign LUT_4[61825] = 32'b00000000000000001111111110000000;
assign LUT_4[61826] = 32'b00000000000000010110001100101100;
assign LUT_4[61827] = 32'b00000000000000001111011000100100;
assign LUT_4[61828] = 32'b00000000000000010011110010100100;
assign LUT_4[61829] = 32'b00000000000000001100111110011100;
assign LUT_4[61830] = 32'b00000000000000010011001101001000;
assign LUT_4[61831] = 32'b00000000000000001100011001000000;
assign LUT_4[61832] = 32'b00000000000000001111111110011101;
assign LUT_4[61833] = 32'b00000000000000001001001010010101;
assign LUT_4[61834] = 32'b00000000000000001111011001000001;
assign LUT_4[61835] = 32'b00000000000000001000100100111001;
assign LUT_4[61836] = 32'b00000000000000001100111110111001;
assign LUT_4[61837] = 32'b00000000000000000110001010110001;
assign LUT_4[61838] = 32'b00000000000000001100011001011101;
assign LUT_4[61839] = 32'b00000000000000000101100101010101;
assign LUT_4[61840] = 32'b00000000000000010100100011110110;
assign LUT_4[61841] = 32'b00000000000000001101101111101110;
assign LUT_4[61842] = 32'b00000000000000010011111110011010;
assign LUT_4[61843] = 32'b00000000000000001101001010010010;
assign LUT_4[61844] = 32'b00000000000000010001100100010010;
assign LUT_4[61845] = 32'b00000000000000001010110000001010;
assign LUT_4[61846] = 32'b00000000000000010000111110110110;
assign LUT_4[61847] = 32'b00000000000000001010001010101110;
assign LUT_4[61848] = 32'b00000000000000001101110000001011;
assign LUT_4[61849] = 32'b00000000000000000110111100000011;
assign LUT_4[61850] = 32'b00000000000000001101001010101111;
assign LUT_4[61851] = 32'b00000000000000000110010110100111;
assign LUT_4[61852] = 32'b00000000000000001010110000100111;
assign LUT_4[61853] = 32'b00000000000000000011111100011111;
assign LUT_4[61854] = 32'b00000000000000001010001011001011;
assign LUT_4[61855] = 32'b00000000000000000011010111000011;
assign LUT_4[61856] = 32'b00000000000000010101001101001111;
assign LUT_4[61857] = 32'b00000000000000001110011001000111;
assign LUT_4[61858] = 32'b00000000000000010100100111110011;
assign LUT_4[61859] = 32'b00000000000000001101110011101011;
assign LUT_4[61860] = 32'b00000000000000010010001101101011;
assign LUT_4[61861] = 32'b00000000000000001011011001100011;
assign LUT_4[61862] = 32'b00000000000000010001101000001111;
assign LUT_4[61863] = 32'b00000000000000001010110100000111;
assign LUT_4[61864] = 32'b00000000000000001110011001100100;
assign LUT_4[61865] = 32'b00000000000000000111100101011100;
assign LUT_4[61866] = 32'b00000000000000001101110100001000;
assign LUT_4[61867] = 32'b00000000000000000111000000000000;
assign LUT_4[61868] = 32'b00000000000000001011011010000000;
assign LUT_4[61869] = 32'b00000000000000000100100101111000;
assign LUT_4[61870] = 32'b00000000000000001010110100100100;
assign LUT_4[61871] = 32'b00000000000000000100000000011100;
assign LUT_4[61872] = 32'b00000000000000010010111110111101;
assign LUT_4[61873] = 32'b00000000000000001100001010110101;
assign LUT_4[61874] = 32'b00000000000000010010011001100001;
assign LUT_4[61875] = 32'b00000000000000001011100101011001;
assign LUT_4[61876] = 32'b00000000000000001111111111011001;
assign LUT_4[61877] = 32'b00000000000000001001001011010001;
assign LUT_4[61878] = 32'b00000000000000001111011001111101;
assign LUT_4[61879] = 32'b00000000000000001000100101110101;
assign LUT_4[61880] = 32'b00000000000000001100001011010010;
assign LUT_4[61881] = 32'b00000000000000000101010111001010;
assign LUT_4[61882] = 32'b00000000000000001011100101110110;
assign LUT_4[61883] = 32'b00000000000000000100110001101110;
assign LUT_4[61884] = 32'b00000000000000001001001011101110;
assign LUT_4[61885] = 32'b00000000000000000010010111100110;
assign LUT_4[61886] = 32'b00000000000000001000100110010010;
assign LUT_4[61887] = 32'b00000000000000000001110010001010;
assign LUT_4[61888] = 32'b00000000000000011000001001011100;
assign LUT_4[61889] = 32'b00000000000000010001010101010100;
assign LUT_4[61890] = 32'b00000000000000010111100100000000;
assign LUT_4[61891] = 32'b00000000000000010000101111111000;
assign LUT_4[61892] = 32'b00000000000000010101001001111000;
assign LUT_4[61893] = 32'b00000000000000001110010101110000;
assign LUT_4[61894] = 32'b00000000000000010100100100011100;
assign LUT_4[61895] = 32'b00000000000000001101110000010100;
assign LUT_4[61896] = 32'b00000000000000010001010101110001;
assign LUT_4[61897] = 32'b00000000000000001010100001101001;
assign LUT_4[61898] = 32'b00000000000000010000110000010101;
assign LUT_4[61899] = 32'b00000000000000001001111100001101;
assign LUT_4[61900] = 32'b00000000000000001110010110001101;
assign LUT_4[61901] = 32'b00000000000000000111100010000101;
assign LUT_4[61902] = 32'b00000000000000001101110000110001;
assign LUT_4[61903] = 32'b00000000000000000110111100101001;
assign LUT_4[61904] = 32'b00000000000000010101111011001010;
assign LUT_4[61905] = 32'b00000000000000001111000111000010;
assign LUT_4[61906] = 32'b00000000000000010101010101101110;
assign LUT_4[61907] = 32'b00000000000000001110100001100110;
assign LUT_4[61908] = 32'b00000000000000010010111011100110;
assign LUT_4[61909] = 32'b00000000000000001100000111011110;
assign LUT_4[61910] = 32'b00000000000000010010010110001010;
assign LUT_4[61911] = 32'b00000000000000001011100010000010;
assign LUT_4[61912] = 32'b00000000000000001111000111011111;
assign LUT_4[61913] = 32'b00000000000000001000010011010111;
assign LUT_4[61914] = 32'b00000000000000001110100010000011;
assign LUT_4[61915] = 32'b00000000000000000111101101111011;
assign LUT_4[61916] = 32'b00000000000000001100000111111011;
assign LUT_4[61917] = 32'b00000000000000000101010011110011;
assign LUT_4[61918] = 32'b00000000000000001011100010011111;
assign LUT_4[61919] = 32'b00000000000000000100101110010111;
assign LUT_4[61920] = 32'b00000000000000010110100100100011;
assign LUT_4[61921] = 32'b00000000000000001111110000011011;
assign LUT_4[61922] = 32'b00000000000000010101111111000111;
assign LUT_4[61923] = 32'b00000000000000001111001010111111;
assign LUT_4[61924] = 32'b00000000000000010011100100111111;
assign LUT_4[61925] = 32'b00000000000000001100110000110111;
assign LUT_4[61926] = 32'b00000000000000010010111111100011;
assign LUT_4[61927] = 32'b00000000000000001100001011011011;
assign LUT_4[61928] = 32'b00000000000000001111110000111000;
assign LUT_4[61929] = 32'b00000000000000001000111100110000;
assign LUT_4[61930] = 32'b00000000000000001111001011011100;
assign LUT_4[61931] = 32'b00000000000000001000010111010100;
assign LUT_4[61932] = 32'b00000000000000001100110001010100;
assign LUT_4[61933] = 32'b00000000000000000101111101001100;
assign LUT_4[61934] = 32'b00000000000000001100001011111000;
assign LUT_4[61935] = 32'b00000000000000000101010111110000;
assign LUT_4[61936] = 32'b00000000000000010100010110010001;
assign LUT_4[61937] = 32'b00000000000000001101100010001001;
assign LUT_4[61938] = 32'b00000000000000010011110000110101;
assign LUT_4[61939] = 32'b00000000000000001100111100101101;
assign LUT_4[61940] = 32'b00000000000000010001010110101101;
assign LUT_4[61941] = 32'b00000000000000001010100010100101;
assign LUT_4[61942] = 32'b00000000000000010000110001010001;
assign LUT_4[61943] = 32'b00000000000000001001111101001001;
assign LUT_4[61944] = 32'b00000000000000001101100010100110;
assign LUT_4[61945] = 32'b00000000000000000110101110011110;
assign LUT_4[61946] = 32'b00000000000000001100111101001010;
assign LUT_4[61947] = 32'b00000000000000000110001001000010;
assign LUT_4[61948] = 32'b00000000000000001010100011000010;
assign LUT_4[61949] = 32'b00000000000000000011101110111010;
assign LUT_4[61950] = 32'b00000000000000001001111101100110;
assign LUT_4[61951] = 32'b00000000000000000011001001011110;
assign LUT_4[61952] = 32'b00000000000000001110010100100101;
assign LUT_4[61953] = 32'b00000000000000000111100000011101;
assign LUT_4[61954] = 32'b00000000000000001101101111001001;
assign LUT_4[61955] = 32'b00000000000000000110111011000001;
assign LUT_4[61956] = 32'b00000000000000001011010101000001;
assign LUT_4[61957] = 32'b00000000000000000100100000111001;
assign LUT_4[61958] = 32'b00000000000000001010101111100101;
assign LUT_4[61959] = 32'b00000000000000000011111011011101;
assign LUT_4[61960] = 32'b00000000000000000111100000111010;
assign LUT_4[61961] = 32'b00000000000000000000101100110010;
assign LUT_4[61962] = 32'b00000000000000000110111011011110;
assign LUT_4[61963] = 32'b00000000000000000000000111010110;
assign LUT_4[61964] = 32'b00000000000000000100100001010110;
assign LUT_4[61965] = 32'b11111111111111111101101101001110;
assign LUT_4[61966] = 32'b00000000000000000011111011111010;
assign LUT_4[61967] = 32'b11111111111111111101000111110010;
assign LUT_4[61968] = 32'b00000000000000001100000110010011;
assign LUT_4[61969] = 32'b00000000000000000101010010001011;
assign LUT_4[61970] = 32'b00000000000000001011100000110111;
assign LUT_4[61971] = 32'b00000000000000000100101100101111;
assign LUT_4[61972] = 32'b00000000000000001001000110101111;
assign LUT_4[61973] = 32'b00000000000000000010010010100111;
assign LUT_4[61974] = 32'b00000000000000001000100001010011;
assign LUT_4[61975] = 32'b00000000000000000001101101001011;
assign LUT_4[61976] = 32'b00000000000000000101010010101000;
assign LUT_4[61977] = 32'b11111111111111111110011110100000;
assign LUT_4[61978] = 32'b00000000000000000100101101001100;
assign LUT_4[61979] = 32'b11111111111111111101111001000100;
assign LUT_4[61980] = 32'b00000000000000000010010011000100;
assign LUT_4[61981] = 32'b11111111111111111011011110111100;
assign LUT_4[61982] = 32'b00000000000000000001101101101000;
assign LUT_4[61983] = 32'b11111111111111111010111001100000;
assign LUT_4[61984] = 32'b00000000000000001100101111101100;
assign LUT_4[61985] = 32'b00000000000000000101111011100100;
assign LUT_4[61986] = 32'b00000000000000001100001010010000;
assign LUT_4[61987] = 32'b00000000000000000101010110001000;
assign LUT_4[61988] = 32'b00000000000000001001110000001000;
assign LUT_4[61989] = 32'b00000000000000000010111100000000;
assign LUT_4[61990] = 32'b00000000000000001001001010101100;
assign LUT_4[61991] = 32'b00000000000000000010010110100100;
assign LUT_4[61992] = 32'b00000000000000000101111100000001;
assign LUT_4[61993] = 32'b11111111111111111111000111111001;
assign LUT_4[61994] = 32'b00000000000000000101010110100101;
assign LUT_4[61995] = 32'b11111111111111111110100010011101;
assign LUT_4[61996] = 32'b00000000000000000010111100011101;
assign LUT_4[61997] = 32'b11111111111111111100001000010101;
assign LUT_4[61998] = 32'b00000000000000000010010111000001;
assign LUT_4[61999] = 32'b11111111111111111011100010111001;
assign LUT_4[62000] = 32'b00000000000000001010100001011010;
assign LUT_4[62001] = 32'b00000000000000000011101101010010;
assign LUT_4[62002] = 32'b00000000000000001001111011111110;
assign LUT_4[62003] = 32'b00000000000000000011000111110110;
assign LUT_4[62004] = 32'b00000000000000000111100001110110;
assign LUT_4[62005] = 32'b00000000000000000000101101101110;
assign LUT_4[62006] = 32'b00000000000000000110111100011010;
assign LUT_4[62007] = 32'b00000000000000000000001000010010;
assign LUT_4[62008] = 32'b00000000000000000011101101101111;
assign LUT_4[62009] = 32'b11111111111111111100111001100111;
assign LUT_4[62010] = 32'b00000000000000000011001000010011;
assign LUT_4[62011] = 32'b11111111111111111100010100001011;
assign LUT_4[62012] = 32'b00000000000000000000101110001011;
assign LUT_4[62013] = 32'b11111111111111111001111010000011;
assign LUT_4[62014] = 32'b00000000000000000000001000101111;
assign LUT_4[62015] = 32'b11111111111111111001010100100111;
assign LUT_4[62016] = 32'b00000000000000001111101011111001;
assign LUT_4[62017] = 32'b00000000000000001000110111110001;
assign LUT_4[62018] = 32'b00000000000000001111000110011101;
assign LUT_4[62019] = 32'b00000000000000001000010010010101;
assign LUT_4[62020] = 32'b00000000000000001100101100010101;
assign LUT_4[62021] = 32'b00000000000000000101111000001101;
assign LUT_4[62022] = 32'b00000000000000001100000110111001;
assign LUT_4[62023] = 32'b00000000000000000101010010110001;
assign LUT_4[62024] = 32'b00000000000000001000111000001110;
assign LUT_4[62025] = 32'b00000000000000000010000100000110;
assign LUT_4[62026] = 32'b00000000000000001000010010110010;
assign LUT_4[62027] = 32'b00000000000000000001011110101010;
assign LUT_4[62028] = 32'b00000000000000000101111000101010;
assign LUT_4[62029] = 32'b11111111111111111111000100100010;
assign LUT_4[62030] = 32'b00000000000000000101010011001110;
assign LUT_4[62031] = 32'b11111111111111111110011111000110;
assign LUT_4[62032] = 32'b00000000000000001101011101100111;
assign LUT_4[62033] = 32'b00000000000000000110101001011111;
assign LUT_4[62034] = 32'b00000000000000001100111000001011;
assign LUT_4[62035] = 32'b00000000000000000110000100000011;
assign LUT_4[62036] = 32'b00000000000000001010011110000011;
assign LUT_4[62037] = 32'b00000000000000000011101001111011;
assign LUT_4[62038] = 32'b00000000000000001001111000100111;
assign LUT_4[62039] = 32'b00000000000000000011000100011111;
assign LUT_4[62040] = 32'b00000000000000000110101001111100;
assign LUT_4[62041] = 32'b11111111111111111111110101110100;
assign LUT_4[62042] = 32'b00000000000000000110000100100000;
assign LUT_4[62043] = 32'b11111111111111111111010000011000;
assign LUT_4[62044] = 32'b00000000000000000011101010011000;
assign LUT_4[62045] = 32'b11111111111111111100110110010000;
assign LUT_4[62046] = 32'b00000000000000000011000100111100;
assign LUT_4[62047] = 32'b11111111111111111100010000110100;
assign LUT_4[62048] = 32'b00000000000000001110000111000000;
assign LUT_4[62049] = 32'b00000000000000000111010010111000;
assign LUT_4[62050] = 32'b00000000000000001101100001100100;
assign LUT_4[62051] = 32'b00000000000000000110101101011100;
assign LUT_4[62052] = 32'b00000000000000001011000111011100;
assign LUT_4[62053] = 32'b00000000000000000100010011010100;
assign LUT_4[62054] = 32'b00000000000000001010100010000000;
assign LUT_4[62055] = 32'b00000000000000000011101101111000;
assign LUT_4[62056] = 32'b00000000000000000111010011010101;
assign LUT_4[62057] = 32'b00000000000000000000011111001101;
assign LUT_4[62058] = 32'b00000000000000000110101101111001;
assign LUT_4[62059] = 32'b11111111111111111111111001110001;
assign LUT_4[62060] = 32'b00000000000000000100010011110001;
assign LUT_4[62061] = 32'b11111111111111111101011111101001;
assign LUT_4[62062] = 32'b00000000000000000011101110010101;
assign LUT_4[62063] = 32'b11111111111111111100111010001101;
assign LUT_4[62064] = 32'b00000000000000001011111000101110;
assign LUT_4[62065] = 32'b00000000000000000101000100100110;
assign LUT_4[62066] = 32'b00000000000000001011010011010010;
assign LUT_4[62067] = 32'b00000000000000000100011111001010;
assign LUT_4[62068] = 32'b00000000000000001000111001001010;
assign LUT_4[62069] = 32'b00000000000000000010000101000010;
assign LUT_4[62070] = 32'b00000000000000001000010011101110;
assign LUT_4[62071] = 32'b00000000000000000001011111100110;
assign LUT_4[62072] = 32'b00000000000000000101000101000011;
assign LUT_4[62073] = 32'b11111111111111111110010000111011;
assign LUT_4[62074] = 32'b00000000000000000100011111100111;
assign LUT_4[62075] = 32'b11111111111111111101101011011111;
assign LUT_4[62076] = 32'b00000000000000000010000101011111;
assign LUT_4[62077] = 32'b11111111111111111011010001010111;
assign LUT_4[62078] = 32'b00000000000000000001100000000011;
assign LUT_4[62079] = 32'b11111111111111111010101011111011;
assign LUT_4[62080] = 32'b00000000000000010000111010101101;
assign LUT_4[62081] = 32'b00000000000000001010000110100101;
assign LUT_4[62082] = 32'b00000000000000010000010101010001;
assign LUT_4[62083] = 32'b00000000000000001001100001001001;
assign LUT_4[62084] = 32'b00000000000000001101111011001001;
assign LUT_4[62085] = 32'b00000000000000000111000111000001;
assign LUT_4[62086] = 32'b00000000000000001101010101101101;
assign LUT_4[62087] = 32'b00000000000000000110100001100101;
assign LUT_4[62088] = 32'b00000000000000001010000111000010;
assign LUT_4[62089] = 32'b00000000000000000011010010111010;
assign LUT_4[62090] = 32'b00000000000000001001100001100110;
assign LUT_4[62091] = 32'b00000000000000000010101101011110;
assign LUT_4[62092] = 32'b00000000000000000111000111011110;
assign LUT_4[62093] = 32'b00000000000000000000010011010110;
assign LUT_4[62094] = 32'b00000000000000000110100010000010;
assign LUT_4[62095] = 32'b11111111111111111111101101111010;
assign LUT_4[62096] = 32'b00000000000000001110101100011011;
assign LUT_4[62097] = 32'b00000000000000000111111000010011;
assign LUT_4[62098] = 32'b00000000000000001110000110111111;
assign LUT_4[62099] = 32'b00000000000000000111010010110111;
assign LUT_4[62100] = 32'b00000000000000001011101100110111;
assign LUT_4[62101] = 32'b00000000000000000100111000101111;
assign LUT_4[62102] = 32'b00000000000000001011000111011011;
assign LUT_4[62103] = 32'b00000000000000000100010011010011;
assign LUT_4[62104] = 32'b00000000000000000111111000110000;
assign LUT_4[62105] = 32'b00000000000000000001000100101000;
assign LUT_4[62106] = 32'b00000000000000000111010011010100;
assign LUT_4[62107] = 32'b00000000000000000000011111001100;
assign LUT_4[62108] = 32'b00000000000000000100111001001100;
assign LUT_4[62109] = 32'b11111111111111111110000101000100;
assign LUT_4[62110] = 32'b00000000000000000100010011110000;
assign LUT_4[62111] = 32'b11111111111111111101011111101000;
assign LUT_4[62112] = 32'b00000000000000001111010101110100;
assign LUT_4[62113] = 32'b00000000000000001000100001101100;
assign LUT_4[62114] = 32'b00000000000000001110110000011000;
assign LUT_4[62115] = 32'b00000000000000000111111100010000;
assign LUT_4[62116] = 32'b00000000000000001100010110010000;
assign LUT_4[62117] = 32'b00000000000000000101100010001000;
assign LUT_4[62118] = 32'b00000000000000001011110000110100;
assign LUT_4[62119] = 32'b00000000000000000100111100101100;
assign LUT_4[62120] = 32'b00000000000000001000100010001001;
assign LUT_4[62121] = 32'b00000000000000000001101110000001;
assign LUT_4[62122] = 32'b00000000000000000111111100101101;
assign LUT_4[62123] = 32'b00000000000000000001001000100101;
assign LUT_4[62124] = 32'b00000000000000000101100010100101;
assign LUT_4[62125] = 32'b11111111111111111110101110011101;
assign LUT_4[62126] = 32'b00000000000000000100111101001001;
assign LUT_4[62127] = 32'b11111111111111111110001001000001;
assign LUT_4[62128] = 32'b00000000000000001101000111100010;
assign LUT_4[62129] = 32'b00000000000000000110010011011010;
assign LUT_4[62130] = 32'b00000000000000001100100010000110;
assign LUT_4[62131] = 32'b00000000000000000101101101111110;
assign LUT_4[62132] = 32'b00000000000000001010000111111110;
assign LUT_4[62133] = 32'b00000000000000000011010011110110;
assign LUT_4[62134] = 32'b00000000000000001001100010100010;
assign LUT_4[62135] = 32'b00000000000000000010101110011010;
assign LUT_4[62136] = 32'b00000000000000000110010011110111;
assign LUT_4[62137] = 32'b11111111111111111111011111101111;
assign LUT_4[62138] = 32'b00000000000000000101101110011011;
assign LUT_4[62139] = 32'b11111111111111111110111010010011;
assign LUT_4[62140] = 32'b00000000000000000011010100010011;
assign LUT_4[62141] = 32'b11111111111111111100100000001011;
assign LUT_4[62142] = 32'b00000000000000000010101110110111;
assign LUT_4[62143] = 32'b11111111111111111011111010101111;
assign LUT_4[62144] = 32'b00000000000000010010010010000001;
assign LUT_4[62145] = 32'b00000000000000001011011101111001;
assign LUT_4[62146] = 32'b00000000000000010001101100100101;
assign LUT_4[62147] = 32'b00000000000000001010111000011101;
assign LUT_4[62148] = 32'b00000000000000001111010010011101;
assign LUT_4[62149] = 32'b00000000000000001000011110010101;
assign LUT_4[62150] = 32'b00000000000000001110101101000001;
assign LUT_4[62151] = 32'b00000000000000000111111000111001;
assign LUT_4[62152] = 32'b00000000000000001011011110010110;
assign LUT_4[62153] = 32'b00000000000000000100101010001110;
assign LUT_4[62154] = 32'b00000000000000001010111000111010;
assign LUT_4[62155] = 32'b00000000000000000100000100110010;
assign LUT_4[62156] = 32'b00000000000000001000011110110010;
assign LUT_4[62157] = 32'b00000000000000000001101010101010;
assign LUT_4[62158] = 32'b00000000000000000111111001010110;
assign LUT_4[62159] = 32'b00000000000000000001000101001110;
assign LUT_4[62160] = 32'b00000000000000010000000011101111;
assign LUT_4[62161] = 32'b00000000000000001001001111100111;
assign LUT_4[62162] = 32'b00000000000000001111011110010011;
assign LUT_4[62163] = 32'b00000000000000001000101010001011;
assign LUT_4[62164] = 32'b00000000000000001101000100001011;
assign LUT_4[62165] = 32'b00000000000000000110010000000011;
assign LUT_4[62166] = 32'b00000000000000001100011110101111;
assign LUT_4[62167] = 32'b00000000000000000101101010100111;
assign LUT_4[62168] = 32'b00000000000000001001010000000100;
assign LUT_4[62169] = 32'b00000000000000000010011011111100;
assign LUT_4[62170] = 32'b00000000000000001000101010101000;
assign LUT_4[62171] = 32'b00000000000000000001110110100000;
assign LUT_4[62172] = 32'b00000000000000000110010000100000;
assign LUT_4[62173] = 32'b11111111111111111111011100011000;
assign LUT_4[62174] = 32'b00000000000000000101101011000100;
assign LUT_4[62175] = 32'b11111111111111111110110110111100;
assign LUT_4[62176] = 32'b00000000000000010000101101001000;
assign LUT_4[62177] = 32'b00000000000000001001111001000000;
assign LUT_4[62178] = 32'b00000000000000010000000111101100;
assign LUT_4[62179] = 32'b00000000000000001001010011100100;
assign LUT_4[62180] = 32'b00000000000000001101101101100100;
assign LUT_4[62181] = 32'b00000000000000000110111001011100;
assign LUT_4[62182] = 32'b00000000000000001101001000001000;
assign LUT_4[62183] = 32'b00000000000000000110010100000000;
assign LUT_4[62184] = 32'b00000000000000001001111001011101;
assign LUT_4[62185] = 32'b00000000000000000011000101010101;
assign LUT_4[62186] = 32'b00000000000000001001010100000001;
assign LUT_4[62187] = 32'b00000000000000000010011111111001;
assign LUT_4[62188] = 32'b00000000000000000110111001111001;
assign LUT_4[62189] = 32'b00000000000000000000000101110001;
assign LUT_4[62190] = 32'b00000000000000000110010100011101;
assign LUT_4[62191] = 32'b11111111111111111111100000010101;
assign LUT_4[62192] = 32'b00000000000000001110011110110110;
assign LUT_4[62193] = 32'b00000000000000000111101010101110;
assign LUT_4[62194] = 32'b00000000000000001101111001011010;
assign LUT_4[62195] = 32'b00000000000000000111000101010010;
assign LUT_4[62196] = 32'b00000000000000001011011111010010;
assign LUT_4[62197] = 32'b00000000000000000100101011001010;
assign LUT_4[62198] = 32'b00000000000000001010111001110110;
assign LUT_4[62199] = 32'b00000000000000000100000101101110;
assign LUT_4[62200] = 32'b00000000000000000111101011001011;
assign LUT_4[62201] = 32'b00000000000000000000110111000011;
assign LUT_4[62202] = 32'b00000000000000000111000101101111;
assign LUT_4[62203] = 32'b00000000000000000000010001100111;
assign LUT_4[62204] = 32'b00000000000000000100101011100111;
assign LUT_4[62205] = 32'b11111111111111111101110111011111;
assign LUT_4[62206] = 32'b00000000000000000100000110001011;
assign LUT_4[62207] = 32'b11111111111111111101010010000011;
assign LUT_4[62208] = 32'b00000000000000010011010000001000;
assign LUT_4[62209] = 32'b00000000000000001100011100000000;
assign LUT_4[62210] = 32'b00000000000000010010101010101100;
assign LUT_4[62211] = 32'b00000000000000001011110110100100;
assign LUT_4[62212] = 32'b00000000000000010000010000100100;
assign LUT_4[62213] = 32'b00000000000000001001011100011100;
assign LUT_4[62214] = 32'b00000000000000001111101011001000;
assign LUT_4[62215] = 32'b00000000000000001000110111000000;
assign LUT_4[62216] = 32'b00000000000000001100011100011101;
assign LUT_4[62217] = 32'b00000000000000000101101000010101;
assign LUT_4[62218] = 32'b00000000000000001011110111000001;
assign LUT_4[62219] = 32'b00000000000000000101000010111001;
assign LUT_4[62220] = 32'b00000000000000001001011100111001;
assign LUT_4[62221] = 32'b00000000000000000010101000110001;
assign LUT_4[62222] = 32'b00000000000000001000110111011101;
assign LUT_4[62223] = 32'b00000000000000000010000011010101;
assign LUT_4[62224] = 32'b00000000000000010001000001110110;
assign LUT_4[62225] = 32'b00000000000000001010001101101110;
assign LUT_4[62226] = 32'b00000000000000010000011100011010;
assign LUT_4[62227] = 32'b00000000000000001001101000010010;
assign LUT_4[62228] = 32'b00000000000000001110000010010010;
assign LUT_4[62229] = 32'b00000000000000000111001110001010;
assign LUT_4[62230] = 32'b00000000000000001101011100110110;
assign LUT_4[62231] = 32'b00000000000000000110101000101110;
assign LUT_4[62232] = 32'b00000000000000001010001110001011;
assign LUT_4[62233] = 32'b00000000000000000011011010000011;
assign LUT_4[62234] = 32'b00000000000000001001101000101111;
assign LUT_4[62235] = 32'b00000000000000000010110100100111;
assign LUT_4[62236] = 32'b00000000000000000111001110100111;
assign LUT_4[62237] = 32'b00000000000000000000011010011111;
assign LUT_4[62238] = 32'b00000000000000000110101001001011;
assign LUT_4[62239] = 32'b11111111111111111111110101000011;
assign LUT_4[62240] = 32'b00000000000000010001101011001111;
assign LUT_4[62241] = 32'b00000000000000001010110111000111;
assign LUT_4[62242] = 32'b00000000000000010001000101110011;
assign LUT_4[62243] = 32'b00000000000000001010010001101011;
assign LUT_4[62244] = 32'b00000000000000001110101011101011;
assign LUT_4[62245] = 32'b00000000000000000111110111100011;
assign LUT_4[62246] = 32'b00000000000000001110000110001111;
assign LUT_4[62247] = 32'b00000000000000000111010010000111;
assign LUT_4[62248] = 32'b00000000000000001010110111100100;
assign LUT_4[62249] = 32'b00000000000000000100000011011100;
assign LUT_4[62250] = 32'b00000000000000001010010010001000;
assign LUT_4[62251] = 32'b00000000000000000011011110000000;
assign LUT_4[62252] = 32'b00000000000000000111111000000000;
assign LUT_4[62253] = 32'b00000000000000000001000011111000;
assign LUT_4[62254] = 32'b00000000000000000111010010100100;
assign LUT_4[62255] = 32'b00000000000000000000011110011100;
assign LUT_4[62256] = 32'b00000000000000001111011100111101;
assign LUT_4[62257] = 32'b00000000000000001000101000110101;
assign LUT_4[62258] = 32'b00000000000000001110110111100001;
assign LUT_4[62259] = 32'b00000000000000001000000011011001;
assign LUT_4[62260] = 32'b00000000000000001100011101011001;
assign LUT_4[62261] = 32'b00000000000000000101101001010001;
assign LUT_4[62262] = 32'b00000000000000001011110111111101;
assign LUT_4[62263] = 32'b00000000000000000101000011110101;
assign LUT_4[62264] = 32'b00000000000000001000101001010010;
assign LUT_4[62265] = 32'b00000000000000000001110101001010;
assign LUT_4[62266] = 32'b00000000000000001000000011110110;
assign LUT_4[62267] = 32'b00000000000000000001001111101110;
assign LUT_4[62268] = 32'b00000000000000000101101001101110;
assign LUT_4[62269] = 32'b11111111111111111110110101100110;
assign LUT_4[62270] = 32'b00000000000000000101000100010010;
assign LUT_4[62271] = 32'b11111111111111111110010000001010;
assign LUT_4[62272] = 32'b00000000000000010100100111011100;
assign LUT_4[62273] = 32'b00000000000000001101110011010100;
assign LUT_4[62274] = 32'b00000000000000010100000010000000;
assign LUT_4[62275] = 32'b00000000000000001101001101111000;
assign LUT_4[62276] = 32'b00000000000000010001100111111000;
assign LUT_4[62277] = 32'b00000000000000001010110011110000;
assign LUT_4[62278] = 32'b00000000000000010001000010011100;
assign LUT_4[62279] = 32'b00000000000000001010001110010100;
assign LUT_4[62280] = 32'b00000000000000001101110011110001;
assign LUT_4[62281] = 32'b00000000000000000110111111101001;
assign LUT_4[62282] = 32'b00000000000000001101001110010101;
assign LUT_4[62283] = 32'b00000000000000000110011010001101;
assign LUT_4[62284] = 32'b00000000000000001010110100001101;
assign LUT_4[62285] = 32'b00000000000000000100000000000101;
assign LUT_4[62286] = 32'b00000000000000001010001110110001;
assign LUT_4[62287] = 32'b00000000000000000011011010101001;
assign LUT_4[62288] = 32'b00000000000000010010011001001010;
assign LUT_4[62289] = 32'b00000000000000001011100101000010;
assign LUT_4[62290] = 32'b00000000000000010001110011101110;
assign LUT_4[62291] = 32'b00000000000000001010111111100110;
assign LUT_4[62292] = 32'b00000000000000001111011001100110;
assign LUT_4[62293] = 32'b00000000000000001000100101011110;
assign LUT_4[62294] = 32'b00000000000000001110110100001010;
assign LUT_4[62295] = 32'b00000000000000001000000000000010;
assign LUT_4[62296] = 32'b00000000000000001011100101011111;
assign LUT_4[62297] = 32'b00000000000000000100110001010111;
assign LUT_4[62298] = 32'b00000000000000001011000000000011;
assign LUT_4[62299] = 32'b00000000000000000100001011111011;
assign LUT_4[62300] = 32'b00000000000000001000100101111011;
assign LUT_4[62301] = 32'b00000000000000000001110001110011;
assign LUT_4[62302] = 32'b00000000000000001000000000011111;
assign LUT_4[62303] = 32'b00000000000000000001001100010111;
assign LUT_4[62304] = 32'b00000000000000010011000010100011;
assign LUT_4[62305] = 32'b00000000000000001100001110011011;
assign LUT_4[62306] = 32'b00000000000000010010011101000111;
assign LUT_4[62307] = 32'b00000000000000001011101000111111;
assign LUT_4[62308] = 32'b00000000000000010000000010111111;
assign LUT_4[62309] = 32'b00000000000000001001001110110111;
assign LUT_4[62310] = 32'b00000000000000001111011101100011;
assign LUT_4[62311] = 32'b00000000000000001000101001011011;
assign LUT_4[62312] = 32'b00000000000000001100001110111000;
assign LUT_4[62313] = 32'b00000000000000000101011010110000;
assign LUT_4[62314] = 32'b00000000000000001011101001011100;
assign LUT_4[62315] = 32'b00000000000000000100110101010100;
assign LUT_4[62316] = 32'b00000000000000001001001111010100;
assign LUT_4[62317] = 32'b00000000000000000010011011001100;
assign LUT_4[62318] = 32'b00000000000000001000101001111000;
assign LUT_4[62319] = 32'b00000000000000000001110101110000;
assign LUT_4[62320] = 32'b00000000000000010000110100010001;
assign LUT_4[62321] = 32'b00000000000000001010000000001001;
assign LUT_4[62322] = 32'b00000000000000010000001110110101;
assign LUT_4[62323] = 32'b00000000000000001001011010101101;
assign LUT_4[62324] = 32'b00000000000000001101110100101101;
assign LUT_4[62325] = 32'b00000000000000000111000000100101;
assign LUT_4[62326] = 32'b00000000000000001101001111010001;
assign LUT_4[62327] = 32'b00000000000000000110011011001001;
assign LUT_4[62328] = 32'b00000000000000001010000000100110;
assign LUT_4[62329] = 32'b00000000000000000011001100011110;
assign LUT_4[62330] = 32'b00000000000000001001011011001010;
assign LUT_4[62331] = 32'b00000000000000000010100111000010;
assign LUT_4[62332] = 32'b00000000000000000111000001000010;
assign LUT_4[62333] = 32'b00000000000000000000001100111010;
assign LUT_4[62334] = 32'b00000000000000000110011011100110;
assign LUT_4[62335] = 32'b11111111111111111111100111011110;
assign LUT_4[62336] = 32'b00000000000000010101110110010000;
assign LUT_4[62337] = 32'b00000000000000001111000010001000;
assign LUT_4[62338] = 32'b00000000000000010101010000110100;
assign LUT_4[62339] = 32'b00000000000000001110011100101100;
assign LUT_4[62340] = 32'b00000000000000010010110110101100;
assign LUT_4[62341] = 32'b00000000000000001100000010100100;
assign LUT_4[62342] = 32'b00000000000000010010010001010000;
assign LUT_4[62343] = 32'b00000000000000001011011101001000;
assign LUT_4[62344] = 32'b00000000000000001111000010100101;
assign LUT_4[62345] = 32'b00000000000000001000001110011101;
assign LUT_4[62346] = 32'b00000000000000001110011101001001;
assign LUT_4[62347] = 32'b00000000000000000111101001000001;
assign LUT_4[62348] = 32'b00000000000000001100000011000001;
assign LUT_4[62349] = 32'b00000000000000000101001110111001;
assign LUT_4[62350] = 32'b00000000000000001011011101100101;
assign LUT_4[62351] = 32'b00000000000000000100101001011101;
assign LUT_4[62352] = 32'b00000000000000010011100111111110;
assign LUT_4[62353] = 32'b00000000000000001100110011110110;
assign LUT_4[62354] = 32'b00000000000000010011000010100010;
assign LUT_4[62355] = 32'b00000000000000001100001110011010;
assign LUT_4[62356] = 32'b00000000000000010000101000011010;
assign LUT_4[62357] = 32'b00000000000000001001110100010010;
assign LUT_4[62358] = 32'b00000000000000010000000010111110;
assign LUT_4[62359] = 32'b00000000000000001001001110110110;
assign LUT_4[62360] = 32'b00000000000000001100110100010011;
assign LUT_4[62361] = 32'b00000000000000000110000000001011;
assign LUT_4[62362] = 32'b00000000000000001100001110110111;
assign LUT_4[62363] = 32'b00000000000000000101011010101111;
assign LUT_4[62364] = 32'b00000000000000001001110100101111;
assign LUT_4[62365] = 32'b00000000000000000011000000100111;
assign LUT_4[62366] = 32'b00000000000000001001001111010011;
assign LUT_4[62367] = 32'b00000000000000000010011011001011;
assign LUT_4[62368] = 32'b00000000000000010100010001010111;
assign LUT_4[62369] = 32'b00000000000000001101011101001111;
assign LUT_4[62370] = 32'b00000000000000010011101011111011;
assign LUT_4[62371] = 32'b00000000000000001100110111110011;
assign LUT_4[62372] = 32'b00000000000000010001010001110011;
assign LUT_4[62373] = 32'b00000000000000001010011101101011;
assign LUT_4[62374] = 32'b00000000000000010000101100010111;
assign LUT_4[62375] = 32'b00000000000000001001111000001111;
assign LUT_4[62376] = 32'b00000000000000001101011101101100;
assign LUT_4[62377] = 32'b00000000000000000110101001100100;
assign LUT_4[62378] = 32'b00000000000000001100111000010000;
assign LUT_4[62379] = 32'b00000000000000000110000100001000;
assign LUT_4[62380] = 32'b00000000000000001010011110001000;
assign LUT_4[62381] = 32'b00000000000000000011101010000000;
assign LUT_4[62382] = 32'b00000000000000001001111000101100;
assign LUT_4[62383] = 32'b00000000000000000011000100100100;
assign LUT_4[62384] = 32'b00000000000000010010000011000101;
assign LUT_4[62385] = 32'b00000000000000001011001110111101;
assign LUT_4[62386] = 32'b00000000000000010001011101101001;
assign LUT_4[62387] = 32'b00000000000000001010101001100001;
assign LUT_4[62388] = 32'b00000000000000001111000011100001;
assign LUT_4[62389] = 32'b00000000000000001000001111011001;
assign LUT_4[62390] = 32'b00000000000000001110011110000101;
assign LUT_4[62391] = 32'b00000000000000000111101001111101;
assign LUT_4[62392] = 32'b00000000000000001011001111011010;
assign LUT_4[62393] = 32'b00000000000000000100011011010010;
assign LUT_4[62394] = 32'b00000000000000001010101001111110;
assign LUT_4[62395] = 32'b00000000000000000011110101110110;
assign LUT_4[62396] = 32'b00000000000000001000001111110110;
assign LUT_4[62397] = 32'b00000000000000000001011011101110;
assign LUT_4[62398] = 32'b00000000000000000111101010011010;
assign LUT_4[62399] = 32'b00000000000000000000110110010010;
assign LUT_4[62400] = 32'b00000000000000010111001101100100;
assign LUT_4[62401] = 32'b00000000000000010000011001011100;
assign LUT_4[62402] = 32'b00000000000000010110101000001000;
assign LUT_4[62403] = 32'b00000000000000001111110100000000;
assign LUT_4[62404] = 32'b00000000000000010100001110000000;
assign LUT_4[62405] = 32'b00000000000000001101011001111000;
assign LUT_4[62406] = 32'b00000000000000010011101000100100;
assign LUT_4[62407] = 32'b00000000000000001100110100011100;
assign LUT_4[62408] = 32'b00000000000000010000011001111001;
assign LUT_4[62409] = 32'b00000000000000001001100101110001;
assign LUT_4[62410] = 32'b00000000000000001111110100011101;
assign LUT_4[62411] = 32'b00000000000000001001000000010101;
assign LUT_4[62412] = 32'b00000000000000001101011010010101;
assign LUT_4[62413] = 32'b00000000000000000110100110001101;
assign LUT_4[62414] = 32'b00000000000000001100110100111001;
assign LUT_4[62415] = 32'b00000000000000000110000000110001;
assign LUT_4[62416] = 32'b00000000000000010100111111010010;
assign LUT_4[62417] = 32'b00000000000000001110001011001010;
assign LUT_4[62418] = 32'b00000000000000010100011001110110;
assign LUT_4[62419] = 32'b00000000000000001101100101101110;
assign LUT_4[62420] = 32'b00000000000000010001111111101110;
assign LUT_4[62421] = 32'b00000000000000001011001011100110;
assign LUT_4[62422] = 32'b00000000000000010001011010010010;
assign LUT_4[62423] = 32'b00000000000000001010100110001010;
assign LUT_4[62424] = 32'b00000000000000001110001011100111;
assign LUT_4[62425] = 32'b00000000000000000111010111011111;
assign LUT_4[62426] = 32'b00000000000000001101100110001011;
assign LUT_4[62427] = 32'b00000000000000000110110010000011;
assign LUT_4[62428] = 32'b00000000000000001011001100000011;
assign LUT_4[62429] = 32'b00000000000000000100010111111011;
assign LUT_4[62430] = 32'b00000000000000001010100110100111;
assign LUT_4[62431] = 32'b00000000000000000011110010011111;
assign LUT_4[62432] = 32'b00000000000000010101101000101011;
assign LUT_4[62433] = 32'b00000000000000001110110100100011;
assign LUT_4[62434] = 32'b00000000000000010101000011001111;
assign LUT_4[62435] = 32'b00000000000000001110001111000111;
assign LUT_4[62436] = 32'b00000000000000010010101001000111;
assign LUT_4[62437] = 32'b00000000000000001011110100111111;
assign LUT_4[62438] = 32'b00000000000000010010000011101011;
assign LUT_4[62439] = 32'b00000000000000001011001111100011;
assign LUT_4[62440] = 32'b00000000000000001110110101000000;
assign LUT_4[62441] = 32'b00000000000000001000000000111000;
assign LUT_4[62442] = 32'b00000000000000001110001111100100;
assign LUT_4[62443] = 32'b00000000000000000111011011011100;
assign LUT_4[62444] = 32'b00000000000000001011110101011100;
assign LUT_4[62445] = 32'b00000000000000000101000001010100;
assign LUT_4[62446] = 32'b00000000000000001011010000000000;
assign LUT_4[62447] = 32'b00000000000000000100011011111000;
assign LUT_4[62448] = 32'b00000000000000010011011010011001;
assign LUT_4[62449] = 32'b00000000000000001100100110010001;
assign LUT_4[62450] = 32'b00000000000000010010110100111101;
assign LUT_4[62451] = 32'b00000000000000001100000000110101;
assign LUT_4[62452] = 32'b00000000000000010000011010110101;
assign LUT_4[62453] = 32'b00000000000000001001100110101101;
assign LUT_4[62454] = 32'b00000000000000001111110101011001;
assign LUT_4[62455] = 32'b00000000000000001001000001010001;
assign LUT_4[62456] = 32'b00000000000000001100100110101110;
assign LUT_4[62457] = 32'b00000000000000000101110010100110;
assign LUT_4[62458] = 32'b00000000000000001100000001010010;
assign LUT_4[62459] = 32'b00000000000000000101001101001010;
assign LUT_4[62460] = 32'b00000000000000001001100111001010;
assign LUT_4[62461] = 32'b00000000000000000010110011000010;
assign LUT_4[62462] = 32'b00000000000000001001000001101110;
assign LUT_4[62463] = 32'b00000000000000000010001101100110;
assign LUT_4[62464] = 32'b00000000000000010000111010111100;
assign LUT_4[62465] = 32'b00000000000000001010000110110100;
assign LUT_4[62466] = 32'b00000000000000010000010101100000;
assign LUT_4[62467] = 32'b00000000000000001001100001011000;
assign LUT_4[62468] = 32'b00000000000000001101111011011000;
assign LUT_4[62469] = 32'b00000000000000000111000111010000;
assign LUT_4[62470] = 32'b00000000000000001101010101111100;
assign LUT_4[62471] = 32'b00000000000000000110100001110100;
assign LUT_4[62472] = 32'b00000000000000001010000111010001;
assign LUT_4[62473] = 32'b00000000000000000011010011001001;
assign LUT_4[62474] = 32'b00000000000000001001100001110101;
assign LUT_4[62475] = 32'b00000000000000000010101101101101;
assign LUT_4[62476] = 32'b00000000000000000111000111101101;
assign LUT_4[62477] = 32'b00000000000000000000010011100101;
assign LUT_4[62478] = 32'b00000000000000000110100010010001;
assign LUT_4[62479] = 32'b11111111111111111111101110001001;
assign LUT_4[62480] = 32'b00000000000000001110101100101010;
assign LUT_4[62481] = 32'b00000000000000000111111000100010;
assign LUT_4[62482] = 32'b00000000000000001110000111001110;
assign LUT_4[62483] = 32'b00000000000000000111010011000110;
assign LUT_4[62484] = 32'b00000000000000001011101101000110;
assign LUT_4[62485] = 32'b00000000000000000100111000111110;
assign LUT_4[62486] = 32'b00000000000000001011000111101010;
assign LUT_4[62487] = 32'b00000000000000000100010011100010;
assign LUT_4[62488] = 32'b00000000000000000111111000111111;
assign LUT_4[62489] = 32'b00000000000000000001000100110111;
assign LUT_4[62490] = 32'b00000000000000000111010011100011;
assign LUT_4[62491] = 32'b00000000000000000000011111011011;
assign LUT_4[62492] = 32'b00000000000000000100111001011011;
assign LUT_4[62493] = 32'b11111111111111111110000101010011;
assign LUT_4[62494] = 32'b00000000000000000100010011111111;
assign LUT_4[62495] = 32'b11111111111111111101011111110111;
assign LUT_4[62496] = 32'b00000000000000001111010110000011;
assign LUT_4[62497] = 32'b00000000000000001000100001111011;
assign LUT_4[62498] = 32'b00000000000000001110110000100111;
assign LUT_4[62499] = 32'b00000000000000000111111100011111;
assign LUT_4[62500] = 32'b00000000000000001100010110011111;
assign LUT_4[62501] = 32'b00000000000000000101100010010111;
assign LUT_4[62502] = 32'b00000000000000001011110001000011;
assign LUT_4[62503] = 32'b00000000000000000100111100111011;
assign LUT_4[62504] = 32'b00000000000000001000100010011000;
assign LUT_4[62505] = 32'b00000000000000000001101110010000;
assign LUT_4[62506] = 32'b00000000000000000111111100111100;
assign LUT_4[62507] = 32'b00000000000000000001001000110100;
assign LUT_4[62508] = 32'b00000000000000000101100010110100;
assign LUT_4[62509] = 32'b11111111111111111110101110101100;
assign LUT_4[62510] = 32'b00000000000000000100111101011000;
assign LUT_4[62511] = 32'b11111111111111111110001001010000;
assign LUT_4[62512] = 32'b00000000000000001101000111110001;
assign LUT_4[62513] = 32'b00000000000000000110010011101001;
assign LUT_4[62514] = 32'b00000000000000001100100010010101;
assign LUT_4[62515] = 32'b00000000000000000101101110001101;
assign LUT_4[62516] = 32'b00000000000000001010001000001101;
assign LUT_4[62517] = 32'b00000000000000000011010100000101;
assign LUT_4[62518] = 32'b00000000000000001001100010110001;
assign LUT_4[62519] = 32'b00000000000000000010101110101001;
assign LUT_4[62520] = 32'b00000000000000000110010100000110;
assign LUT_4[62521] = 32'b11111111111111111111011111111110;
assign LUT_4[62522] = 32'b00000000000000000101101110101010;
assign LUT_4[62523] = 32'b11111111111111111110111010100010;
assign LUT_4[62524] = 32'b00000000000000000011010100100010;
assign LUT_4[62525] = 32'b11111111111111111100100000011010;
assign LUT_4[62526] = 32'b00000000000000000010101111000110;
assign LUT_4[62527] = 32'b11111111111111111011111010111110;
assign LUT_4[62528] = 32'b00000000000000010010010010010000;
assign LUT_4[62529] = 32'b00000000000000001011011110001000;
assign LUT_4[62530] = 32'b00000000000000010001101100110100;
assign LUT_4[62531] = 32'b00000000000000001010111000101100;
assign LUT_4[62532] = 32'b00000000000000001111010010101100;
assign LUT_4[62533] = 32'b00000000000000001000011110100100;
assign LUT_4[62534] = 32'b00000000000000001110101101010000;
assign LUT_4[62535] = 32'b00000000000000000111111001001000;
assign LUT_4[62536] = 32'b00000000000000001011011110100101;
assign LUT_4[62537] = 32'b00000000000000000100101010011101;
assign LUT_4[62538] = 32'b00000000000000001010111001001001;
assign LUT_4[62539] = 32'b00000000000000000100000101000001;
assign LUT_4[62540] = 32'b00000000000000001000011111000001;
assign LUT_4[62541] = 32'b00000000000000000001101010111001;
assign LUT_4[62542] = 32'b00000000000000000111111001100101;
assign LUT_4[62543] = 32'b00000000000000000001000101011101;
assign LUT_4[62544] = 32'b00000000000000010000000011111110;
assign LUT_4[62545] = 32'b00000000000000001001001111110110;
assign LUT_4[62546] = 32'b00000000000000001111011110100010;
assign LUT_4[62547] = 32'b00000000000000001000101010011010;
assign LUT_4[62548] = 32'b00000000000000001101000100011010;
assign LUT_4[62549] = 32'b00000000000000000110010000010010;
assign LUT_4[62550] = 32'b00000000000000001100011110111110;
assign LUT_4[62551] = 32'b00000000000000000101101010110110;
assign LUT_4[62552] = 32'b00000000000000001001010000010011;
assign LUT_4[62553] = 32'b00000000000000000010011100001011;
assign LUT_4[62554] = 32'b00000000000000001000101010110111;
assign LUT_4[62555] = 32'b00000000000000000001110110101111;
assign LUT_4[62556] = 32'b00000000000000000110010000101111;
assign LUT_4[62557] = 32'b11111111111111111111011100100111;
assign LUT_4[62558] = 32'b00000000000000000101101011010011;
assign LUT_4[62559] = 32'b11111111111111111110110111001011;
assign LUT_4[62560] = 32'b00000000000000010000101101010111;
assign LUT_4[62561] = 32'b00000000000000001001111001001111;
assign LUT_4[62562] = 32'b00000000000000010000000111111011;
assign LUT_4[62563] = 32'b00000000000000001001010011110011;
assign LUT_4[62564] = 32'b00000000000000001101101101110011;
assign LUT_4[62565] = 32'b00000000000000000110111001101011;
assign LUT_4[62566] = 32'b00000000000000001101001000010111;
assign LUT_4[62567] = 32'b00000000000000000110010100001111;
assign LUT_4[62568] = 32'b00000000000000001001111001101100;
assign LUT_4[62569] = 32'b00000000000000000011000101100100;
assign LUT_4[62570] = 32'b00000000000000001001010100010000;
assign LUT_4[62571] = 32'b00000000000000000010100000001000;
assign LUT_4[62572] = 32'b00000000000000000110111010001000;
assign LUT_4[62573] = 32'b00000000000000000000000110000000;
assign LUT_4[62574] = 32'b00000000000000000110010100101100;
assign LUT_4[62575] = 32'b11111111111111111111100000100100;
assign LUT_4[62576] = 32'b00000000000000001110011111000101;
assign LUT_4[62577] = 32'b00000000000000000111101010111101;
assign LUT_4[62578] = 32'b00000000000000001101111001101001;
assign LUT_4[62579] = 32'b00000000000000000111000101100001;
assign LUT_4[62580] = 32'b00000000000000001011011111100001;
assign LUT_4[62581] = 32'b00000000000000000100101011011001;
assign LUT_4[62582] = 32'b00000000000000001010111010000101;
assign LUT_4[62583] = 32'b00000000000000000100000101111101;
assign LUT_4[62584] = 32'b00000000000000000111101011011010;
assign LUT_4[62585] = 32'b00000000000000000000110111010010;
assign LUT_4[62586] = 32'b00000000000000000111000101111110;
assign LUT_4[62587] = 32'b00000000000000000000010001110110;
assign LUT_4[62588] = 32'b00000000000000000100101011110110;
assign LUT_4[62589] = 32'b11111111111111111101110111101110;
assign LUT_4[62590] = 32'b00000000000000000100000110011010;
assign LUT_4[62591] = 32'b11111111111111111101010010010010;
assign LUT_4[62592] = 32'b00000000000000010011100001000100;
assign LUT_4[62593] = 32'b00000000000000001100101100111100;
assign LUT_4[62594] = 32'b00000000000000010010111011101000;
assign LUT_4[62595] = 32'b00000000000000001100000111100000;
assign LUT_4[62596] = 32'b00000000000000010000100001100000;
assign LUT_4[62597] = 32'b00000000000000001001101101011000;
assign LUT_4[62598] = 32'b00000000000000001111111100000100;
assign LUT_4[62599] = 32'b00000000000000001001000111111100;
assign LUT_4[62600] = 32'b00000000000000001100101101011001;
assign LUT_4[62601] = 32'b00000000000000000101111001010001;
assign LUT_4[62602] = 32'b00000000000000001100000111111101;
assign LUT_4[62603] = 32'b00000000000000000101010011110101;
assign LUT_4[62604] = 32'b00000000000000001001101101110101;
assign LUT_4[62605] = 32'b00000000000000000010111001101101;
assign LUT_4[62606] = 32'b00000000000000001001001000011001;
assign LUT_4[62607] = 32'b00000000000000000010010100010001;
assign LUT_4[62608] = 32'b00000000000000010001010010110010;
assign LUT_4[62609] = 32'b00000000000000001010011110101010;
assign LUT_4[62610] = 32'b00000000000000010000101101010110;
assign LUT_4[62611] = 32'b00000000000000001001111001001110;
assign LUT_4[62612] = 32'b00000000000000001110010011001110;
assign LUT_4[62613] = 32'b00000000000000000111011111000110;
assign LUT_4[62614] = 32'b00000000000000001101101101110010;
assign LUT_4[62615] = 32'b00000000000000000110111001101010;
assign LUT_4[62616] = 32'b00000000000000001010011111000111;
assign LUT_4[62617] = 32'b00000000000000000011101010111111;
assign LUT_4[62618] = 32'b00000000000000001001111001101011;
assign LUT_4[62619] = 32'b00000000000000000011000101100011;
assign LUT_4[62620] = 32'b00000000000000000111011111100011;
assign LUT_4[62621] = 32'b00000000000000000000101011011011;
assign LUT_4[62622] = 32'b00000000000000000110111010000111;
assign LUT_4[62623] = 32'b00000000000000000000000101111111;
assign LUT_4[62624] = 32'b00000000000000010001111100001011;
assign LUT_4[62625] = 32'b00000000000000001011001000000011;
assign LUT_4[62626] = 32'b00000000000000010001010110101111;
assign LUT_4[62627] = 32'b00000000000000001010100010100111;
assign LUT_4[62628] = 32'b00000000000000001110111100100111;
assign LUT_4[62629] = 32'b00000000000000001000001000011111;
assign LUT_4[62630] = 32'b00000000000000001110010111001011;
assign LUT_4[62631] = 32'b00000000000000000111100011000011;
assign LUT_4[62632] = 32'b00000000000000001011001000100000;
assign LUT_4[62633] = 32'b00000000000000000100010100011000;
assign LUT_4[62634] = 32'b00000000000000001010100011000100;
assign LUT_4[62635] = 32'b00000000000000000011101110111100;
assign LUT_4[62636] = 32'b00000000000000001000001000111100;
assign LUT_4[62637] = 32'b00000000000000000001010100110100;
assign LUT_4[62638] = 32'b00000000000000000111100011100000;
assign LUT_4[62639] = 32'b00000000000000000000101111011000;
assign LUT_4[62640] = 32'b00000000000000001111101101111001;
assign LUT_4[62641] = 32'b00000000000000001000111001110001;
assign LUT_4[62642] = 32'b00000000000000001111001000011101;
assign LUT_4[62643] = 32'b00000000000000001000010100010101;
assign LUT_4[62644] = 32'b00000000000000001100101110010101;
assign LUT_4[62645] = 32'b00000000000000000101111010001101;
assign LUT_4[62646] = 32'b00000000000000001100001000111001;
assign LUT_4[62647] = 32'b00000000000000000101010100110001;
assign LUT_4[62648] = 32'b00000000000000001000111010001110;
assign LUT_4[62649] = 32'b00000000000000000010000110000110;
assign LUT_4[62650] = 32'b00000000000000001000010100110010;
assign LUT_4[62651] = 32'b00000000000000000001100000101010;
assign LUT_4[62652] = 32'b00000000000000000101111010101010;
assign LUT_4[62653] = 32'b11111111111111111111000110100010;
assign LUT_4[62654] = 32'b00000000000000000101010101001110;
assign LUT_4[62655] = 32'b11111111111111111110100001000110;
assign LUT_4[62656] = 32'b00000000000000010100111000011000;
assign LUT_4[62657] = 32'b00000000000000001110000100010000;
assign LUT_4[62658] = 32'b00000000000000010100010010111100;
assign LUT_4[62659] = 32'b00000000000000001101011110110100;
assign LUT_4[62660] = 32'b00000000000000010001111000110100;
assign LUT_4[62661] = 32'b00000000000000001011000100101100;
assign LUT_4[62662] = 32'b00000000000000010001010011011000;
assign LUT_4[62663] = 32'b00000000000000001010011111010000;
assign LUT_4[62664] = 32'b00000000000000001110000100101101;
assign LUT_4[62665] = 32'b00000000000000000111010000100101;
assign LUT_4[62666] = 32'b00000000000000001101011111010001;
assign LUT_4[62667] = 32'b00000000000000000110101011001001;
assign LUT_4[62668] = 32'b00000000000000001011000101001001;
assign LUT_4[62669] = 32'b00000000000000000100010001000001;
assign LUT_4[62670] = 32'b00000000000000001010011111101101;
assign LUT_4[62671] = 32'b00000000000000000011101011100101;
assign LUT_4[62672] = 32'b00000000000000010010101010000110;
assign LUT_4[62673] = 32'b00000000000000001011110101111110;
assign LUT_4[62674] = 32'b00000000000000010010000100101010;
assign LUT_4[62675] = 32'b00000000000000001011010000100010;
assign LUT_4[62676] = 32'b00000000000000001111101010100010;
assign LUT_4[62677] = 32'b00000000000000001000110110011010;
assign LUT_4[62678] = 32'b00000000000000001111000101000110;
assign LUT_4[62679] = 32'b00000000000000001000010000111110;
assign LUT_4[62680] = 32'b00000000000000001011110110011011;
assign LUT_4[62681] = 32'b00000000000000000101000010010011;
assign LUT_4[62682] = 32'b00000000000000001011010000111111;
assign LUT_4[62683] = 32'b00000000000000000100011100110111;
assign LUT_4[62684] = 32'b00000000000000001000110110110111;
assign LUT_4[62685] = 32'b00000000000000000010000010101111;
assign LUT_4[62686] = 32'b00000000000000001000010001011011;
assign LUT_4[62687] = 32'b00000000000000000001011101010011;
assign LUT_4[62688] = 32'b00000000000000010011010011011111;
assign LUT_4[62689] = 32'b00000000000000001100011111010111;
assign LUT_4[62690] = 32'b00000000000000010010101110000011;
assign LUT_4[62691] = 32'b00000000000000001011111001111011;
assign LUT_4[62692] = 32'b00000000000000010000010011111011;
assign LUT_4[62693] = 32'b00000000000000001001011111110011;
assign LUT_4[62694] = 32'b00000000000000001111101110011111;
assign LUT_4[62695] = 32'b00000000000000001000111010010111;
assign LUT_4[62696] = 32'b00000000000000001100011111110100;
assign LUT_4[62697] = 32'b00000000000000000101101011101100;
assign LUT_4[62698] = 32'b00000000000000001011111010011000;
assign LUT_4[62699] = 32'b00000000000000000101000110010000;
assign LUT_4[62700] = 32'b00000000000000001001100000010000;
assign LUT_4[62701] = 32'b00000000000000000010101100001000;
assign LUT_4[62702] = 32'b00000000000000001000111010110100;
assign LUT_4[62703] = 32'b00000000000000000010000110101100;
assign LUT_4[62704] = 32'b00000000000000010001000101001101;
assign LUT_4[62705] = 32'b00000000000000001010010001000101;
assign LUT_4[62706] = 32'b00000000000000010000011111110001;
assign LUT_4[62707] = 32'b00000000000000001001101011101001;
assign LUT_4[62708] = 32'b00000000000000001110000101101001;
assign LUT_4[62709] = 32'b00000000000000000111010001100001;
assign LUT_4[62710] = 32'b00000000000000001101100000001101;
assign LUT_4[62711] = 32'b00000000000000000110101100000101;
assign LUT_4[62712] = 32'b00000000000000001010010001100010;
assign LUT_4[62713] = 32'b00000000000000000011011101011010;
assign LUT_4[62714] = 32'b00000000000000001001101100000110;
assign LUT_4[62715] = 32'b00000000000000000010110111111110;
assign LUT_4[62716] = 32'b00000000000000000111010001111110;
assign LUT_4[62717] = 32'b00000000000000000000011101110110;
assign LUT_4[62718] = 32'b00000000000000000110101100100010;
assign LUT_4[62719] = 32'b11111111111111111111111000011010;
assign LUT_4[62720] = 32'b00000000000000010101110110011111;
assign LUT_4[62721] = 32'b00000000000000001111000010010111;
assign LUT_4[62722] = 32'b00000000000000010101010001000011;
assign LUT_4[62723] = 32'b00000000000000001110011100111011;
assign LUT_4[62724] = 32'b00000000000000010010110110111011;
assign LUT_4[62725] = 32'b00000000000000001100000010110011;
assign LUT_4[62726] = 32'b00000000000000010010010001011111;
assign LUT_4[62727] = 32'b00000000000000001011011101010111;
assign LUT_4[62728] = 32'b00000000000000001111000010110100;
assign LUT_4[62729] = 32'b00000000000000001000001110101100;
assign LUT_4[62730] = 32'b00000000000000001110011101011000;
assign LUT_4[62731] = 32'b00000000000000000111101001010000;
assign LUT_4[62732] = 32'b00000000000000001100000011010000;
assign LUT_4[62733] = 32'b00000000000000000101001111001000;
assign LUT_4[62734] = 32'b00000000000000001011011101110100;
assign LUT_4[62735] = 32'b00000000000000000100101001101100;
assign LUT_4[62736] = 32'b00000000000000010011101000001101;
assign LUT_4[62737] = 32'b00000000000000001100110100000101;
assign LUT_4[62738] = 32'b00000000000000010011000010110001;
assign LUT_4[62739] = 32'b00000000000000001100001110101001;
assign LUT_4[62740] = 32'b00000000000000010000101000101001;
assign LUT_4[62741] = 32'b00000000000000001001110100100001;
assign LUT_4[62742] = 32'b00000000000000010000000011001101;
assign LUT_4[62743] = 32'b00000000000000001001001111000101;
assign LUT_4[62744] = 32'b00000000000000001100110100100010;
assign LUT_4[62745] = 32'b00000000000000000110000000011010;
assign LUT_4[62746] = 32'b00000000000000001100001111000110;
assign LUT_4[62747] = 32'b00000000000000000101011010111110;
assign LUT_4[62748] = 32'b00000000000000001001110100111110;
assign LUT_4[62749] = 32'b00000000000000000011000000110110;
assign LUT_4[62750] = 32'b00000000000000001001001111100010;
assign LUT_4[62751] = 32'b00000000000000000010011011011010;
assign LUT_4[62752] = 32'b00000000000000010100010001100110;
assign LUT_4[62753] = 32'b00000000000000001101011101011110;
assign LUT_4[62754] = 32'b00000000000000010011101100001010;
assign LUT_4[62755] = 32'b00000000000000001100111000000010;
assign LUT_4[62756] = 32'b00000000000000010001010010000010;
assign LUT_4[62757] = 32'b00000000000000001010011101111010;
assign LUT_4[62758] = 32'b00000000000000010000101100100110;
assign LUT_4[62759] = 32'b00000000000000001001111000011110;
assign LUT_4[62760] = 32'b00000000000000001101011101111011;
assign LUT_4[62761] = 32'b00000000000000000110101001110011;
assign LUT_4[62762] = 32'b00000000000000001100111000011111;
assign LUT_4[62763] = 32'b00000000000000000110000100010111;
assign LUT_4[62764] = 32'b00000000000000001010011110010111;
assign LUT_4[62765] = 32'b00000000000000000011101010001111;
assign LUT_4[62766] = 32'b00000000000000001001111000111011;
assign LUT_4[62767] = 32'b00000000000000000011000100110011;
assign LUT_4[62768] = 32'b00000000000000010010000011010100;
assign LUT_4[62769] = 32'b00000000000000001011001111001100;
assign LUT_4[62770] = 32'b00000000000000010001011101111000;
assign LUT_4[62771] = 32'b00000000000000001010101001110000;
assign LUT_4[62772] = 32'b00000000000000001111000011110000;
assign LUT_4[62773] = 32'b00000000000000001000001111101000;
assign LUT_4[62774] = 32'b00000000000000001110011110010100;
assign LUT_4[62775] = 32'b00000000000000000111101010001100;
assign LUT_4[62776] = 32'b00000000000000001011001111101001;
assign LUT_4[62777] = 32'b00000000000000000100011011100001;
assign LUT_4[62778] = 32'b00000000000000001010101010001101;
assign LUT_4[62779] = 32'b00000000000000000011110110000101;
assign LUT_4[62780] = 32'b00000000000000001000010000000101;
assign LUT_4[62781] = 32'b00000000000000000001011011111101;
assign LUT_4[62782] = 32'b00000000000000000111101010101001;
assign LUT_4[62783] = 32'b00000000000000000000110110100001;
assign LUT_4[62784] = 32'b00000000000000010111001101110011;
assign LUT_4[62785] = 32'b00000000000000010000011001101011;
assign LUT_4[62786] = 32'b00000000000000010110101000010111;
assign LUT_4[62787] = 32'b00000000000000001111110100001111;
assign LUT_4[62788] = 32'b00000000000000010100001110001111;
assign LUT_4[62789] = 32'b00000000000000001101011010000111;
assign LUT_4[62790] = 32'b00000000000000010011101000110011;
assign LUT_4[62791] = 32'b00000000000000001100110100101011;
assign LUT_4[62792] = 32'b00000000000000010000011010001000;
assign LUT_4[62793] = 32'b00000000000000001001100110000000;
assign LUT_4[62794] = 32'b00000000000000001111110100101100;
assign LUT_4[62795] = 32'b00000000000000001001000000100100;
assign LUT_4[62796] = 32'b00000000000000001101011010100100;
assign LUT_4[62797] = 32'b00000000000000000110100110011100;
assign LUT_4[62798] = 32'b00000000000000001100110101001000;
assign LUT_4[62799] = 32'b00000000000000000110000001000000;
assign LUT_4[62800] = 32'b00000000000000010100111111100001;
assign LUT_4[62801] = 32'b00000000000000001110001011011001;
assign LUT_4[62802] = 32'b00000000000000010100011010000101;
assign LUT_4[62803] = 32'b00000000000000001101100101111101;
assign LUT_4[62804] = 32'b00000000000000010001111111111101;
assign LUT_4[62805] = 32'b00000000000000001011001011110101;
assign LUT_4[62806] = 32'b00000000000000010001011010100001;
assign LUT_4[62807] = 32'b00000000000000001010100110011001;
assign LUT_4[62808] = 32'b00000000000000001110001011110110;
assign LUT_4[62809] = 32'b00000000000000000111010111101110;
assign LUT_4[62810] = 32'b00000000000000001101100110011010;
assign LUT_4[62811] = 32'b00000000000000000110110010010010;
assign LUT_4[62812] = 32'b00000000000000001011001100010010;
assign LUT_4[62813] = 32'b00000000000000000100011000001010;
assign LUT_4[62814] = 32'b00000000000000001010100110110110;
assign LUT_4[62815] = 32'b00000000000000000011110010101110;
assign LUT_4[62816] = 32'b00000000000000010101101000111010;
assign LUT_4[62817] = 32'b00000000000000001110110100110010;
assign LUT_4[62818] = 32'b00000000000000010101000011011110;
assign LUT_4[62819] = 32'b00000000000000001110001111010110;
assign LUT_4[62820] = 32'b00000000000000010010101001010110;
assign LUT_4[62821] = 32'b00000000000000001011110101001110;
assign LUT_4[62822] = 32'b00000000000000010010000011111010;
assign LUT_4[62823] = 32'b00000000000000001011001111110010;
assign LUT_4[62824] = 32'b00000000000000001110110101001111;
assign LUT_4[62825] = 32'b00000000000000001000000001000111;
assign LUT_4[62826] = 32'b00000000000000001110001111110011;
assign LUT_4[62827] = 32'b00000000000000000111011011101011;
assign LUT_4[62828] = 32'b00000000000000001011110101101011;
assign LUT_4[62829] = 32'b00000000000000000101000001100011;
assign LUT_4[62830] = 32'b00000000000000001011010000001111;
assign LUT_4[62831] = 32'b00000000000000000100011100000111;
assign LUT_4[62832] = 32'b00000000000000010011011010101000;
assign LUT_4[62833] = 32'b00000000000000001100100110100000;
assign LUT_4[62834] = 32'b00000000000000010010110101001100;
assign LUT_4[62835] = 32'b00000000000000001100000001000100;
assign LUT_4[62836] = 32'b00000000000000010000011011000100;
assign LUT_4[62837] = 32'b00000000000000001001100110111100;
assign LUT_4[62838] = 32'b00000000000000001111110101101000;
assign LUT_4[62839] = 32'b00000000000000001001000001100000;
assign LUT_4[62840] = 32'b00000000000000001100100110111101;
assign LUT_4[62841] = 32'b00000000000000000101110010110101;
assign LUT_4[62842] = 32'b00000000000000001100000001100001;
assign LUT_4[62843] = 32'b00000000000000000101001101011001;
assign LUT_4[62844] = 32'b00000000000000001001100111011001;
assign LUT_4[62845] = 32'b00000000000000000010110011010001;
assign LUT_4[62846] = 32'b00000000000000001001000001111101;
assign LUT_4[62847] = 32'b00000000000000000010001101110101;
assign LUT_4[62848] = 32'b00000000000000011000011100100111;
assign LUT_4[62849] = 32'b00000000000000010001101000011111;
assign LUT_4[62850] = 32'b00000000000000010111110111001011;
assign LUT_4[62851] = 32'b00000000000000010001000011000011;
assign LUT_4[62852] = 32'b00000000000000010101011101000011;
assign LUT_4[62853] = 32'b00000000000000001110101000111011;
assign LUT_4[62854] = 32'b00000000000000010100110111100111;
assign LUT_4[62855] = 32'b00000000000000001110000011011111;
assign LUT_4[62856] = 32'b00000000000000010001101000111100;
assign LUT_4[62857] = 32'b00000000000000001010110100110100;
assign LUT_4[62858] = 32'b00000000000000010001000011100000;
assign LUT_4[62859] = 32'b00000000000000001010001111011000;
assign LUT_4[62860] = 32'b00000000000000001110101001011000;
assign LUT_4[62861] = 32'b00000000000000000111110101010000;
assign LUT_4[62862] = 32'b00000000000000001110000011111100;
assign LUT_4[62863] = 32'b00000000000000000111001111110100;
assign LUT_4[62864] = 32'b00000000000000010110001110010101;
assign LUT_4[62865] = 32'b00000000000000001111011010001101;
assign LUT_4[62866] = 32'b00000000000000010101101000111001;
assign LUT_4[62867] = 32'b00000000000000001110110100110001;
assign LUT_4[62868] = 32'b00000000000000010011001110110001;
assign LUT_4[62869] = 32'b00000000000000001100011010101001;
assign LUT_4[62870] = 32'b00000000000000010010101001010101;
assign LUT_4[62871] = 32'b00000000000000001011110101001101;
assign LUT_4[62872] = 32'b00000000000000001111011010101010;
assign LUT_4[62873] = 32'b00000000000000001000100110100010;
assign LUT_4[62874] = 32'b00000000000000001110110101001110;
assign LUT_4[62875] = 32'b00000000000000001000000001000110;
assign LUT_4[62876] = 32'b00000000000000001100011011000110;
assign LUT_4[62877] = 32'b00000000000000000101100110111110;
assign LUT_4[62878] = 32'b00000000000000001011110101101010;
assign LUT_4[62879] = 32'b00000000000000000101000001100010;
assign LUT_4[62880] = 32'b00000000000000010110110111101110;
assign LUT_4[62881] = 32'b00000000000000010000000011100110;
assign LUT_4[62882] = 32'b00000000000000010110010010010010;
assign LUT_4[62883] = 32'b00000000000000001111011110001010;
assign LUT_4[62884] = 32'b00000000000000010011111000001010;
assign LUT_4[62885] = 32'b00000000000000001101000100000010;
assign LUT_4[62886] = 32'b00000000000000010011010010101110;
assign LUT_4[62887] = 32'b00000000000000001100011110100110;
assign LUT_4[62888] = 32'b00000000000000010000000100000011;
assign LUT_4[62889] = 32'b00000000000000001001001111111011;
assign LUT_4[62890] = 32'b00000000000000001111011110100111;
assign LUT_4[62891] = 32'b00000000000000001000101010011111;
assign LUT_4[62892] = 32'b00000000000000001101000100011111;
assign LUT_4[62893] = 32'b00000000000000000110010000010111;
assign LUT_4[62894] = 32'b00000000000000001100011111000011;
assign LUT_4[62895] = 32'b00000000000000000101101010111011;
assign LUT_4[62896] = 32'b00000000000000010100101001011100;
assign LUT_4[62897] = 32'b00000000000000001101110101010100;
assign LUT_4[62898] = 32'b00000000000000010100000100000000;
assign LUT_4[62899] = 32'b00000000000000001101001111111000;
assign LUT_4[62900] = 32'b00000000000000010001101001111000;
assign LUT_4[62901] = 32'b00000000000000001010110101110000;
assign LUT_4[62902] = 32'b00000000000000010001000100011100;
assign LUT_4[62903] = 32'b00000000000000001010010000010100;
assign LUT_4[62904] = 32'b00000000000000001101110101110001;
assign LUT_4[62905] = 32'b00000000000000000111000001101001;
assign LUT_4[62906] = 32'b00000000000000001101010000010101;
assign LUT_4[62907] = 32'b00000000000000000110011100001101;
assign LUT_4[62908] = 32'b00000000000000001010110110001101;
assign LUT_4[62909] = 32'b00000000000000000100000010000101;
assign LUT_4[62910] = 32'b00000000000000001010010000110001;
assign LUT_4[62911] = 32'b00000000000000000011011100101001;
assign LUT_4[62912] = 32'b00000000000000011001110011111011;
assign LUT_4[62913] = 32'b00000000000000010010111111110011;
assign LUT_4[62914] = 32'b00000000000000011001001110011111;
assign LUT_4[62915] = 32'b00000000000000010010011010010111;
assign LUT_4[62916] = 32'b00000000000000010110110100010111;
assign LUT_4[62917] = 32'b00000000000000010000000000001111;
assign LUT_4[62918] = 32'b00000000000000010110001110111011;
assign LUT_4[62919] = 32'b00000000000000001111011010110011;
assign LUT_4[62920] = 32'b00000000000000010011000000010000;
assign LUT_4[62921] = 32'b00000000000000001100001100001000;
assign LUT_4[62922] = 32'b00000000000000010010011010110100;
assign LUT_4[62923] = 32'b00000000000000001011100110101100;
assign LUT_4[62924] = 32'b00000000000000010000000000101100;
assign LUT_4[62925] = 32'b00000000000000001001001100100100;
assign LUT_4[62926] = 32'b00000000000000001111011011010000;
assign LUT_4[62927] = 32'b00000000000000001000100111001000;
assign LUT_4[62928] = 32'b00000000000000010111100101101001;
assign LUT_4[62929] = 32'b00000000000000010000110001100001;
assign LUT_4[62930] = 32'b00000000000000010111000000001101;
assign LUT_4[62931] = 32'b00000000000000010000001100000101;
assign LUT_4[62932] = 32'b00000000000000010100100110000101;
assign LUT_4[62933] = 32'b00000000000000001101110001111101;
assign LUT_4[62934] = 32'b00000000000000010100000000101001;
assign LUT_4[62935] = 32'b00000000000000001101001100100001;
assign LUT_4[62936] = 32'b00000000000000010000110001111110;
assign LUT_4[62937] = 32'b00000000000000001001111101110110;
assign LUT_4[62938] = 32'b00000000000000010000001100100010;
assign LUT_4[62939] = 32'b00000000000000001001011000011010;
assign LUT_4[62940] = 32'b00000000000000001101110010011010;
assign LUT_4[62941] = 32'b00000000000000000110111110010010;
assign LUT_4[62942] = 32'b00000000000000001101001100111110;
assign LUT_4[62943] = 32'b00000000000000000110011000110110;
assign LUT_4[62944] = 32'b00000000000000011000001111000010;
assign LUT_4[62945] = 32'b00000000000000010001011010111010;
assign LUT_4[62946] = 32'b00000000000000010111101001100110;
assign LUT_4[62947] = 32'b00000000000000010000110101011110;
assign LUT_4[62948] = 32'b00000000000000010101001111011110;
assign LUT_4[62949] = 32'b00000000000000001110011011010110;
assign LUT_4[62950] = 32'b00000000000000010100101010000010;
assign LUT_4[62951] = 32'b00000000000000001101110101111010;
assign LUT_4[62952] = 32'b00000000000000010001011011010111;
assign LUT_4[62953] = 32'b00000000000000001010100111001111;
assign LUT_4[62954] = 32'b00000000000000010000110101111011;
assign LUT_4[62955] = 32'b00000000000000001010000001110011;
assign LUT_4[62956] = 32'b00000000000000001110011011110011;
assign LUT_4[62957] = 32'b00000000000000000111100111101011;
assign LUT_4[62958] = 32'b00000000000000001101110110010111;
assign LUT_4[62959] = 32'b00000000000000000111000010001111;
assign LUT_4[62960] = 32'b00000000000000010110000000110000;
assign LUT_4[62961] = 32'b00000000000000001111001100101000;
assign LUT_4[62962] = 32'b00000000000000010101011011010100;
assign LUT_4[62963] = 32'b00000000000000001110100111001100;
assign LUT_4[62964] = 32'b00000000000000010011000001001100;
assign LUT_4[62965] = 32'b00000000000000001100001101000100;
assign LUT_4[62966] = 32'b00000000000000010010011011110000;
assign LUT_4[62967] = 32'b00000000000000001011100111101000;
assign LUT_4[62968] = 32'b00000000000000001111001101000101;
assign LUT_4[62969] = 32'b00000000000000001000011000111101;
assign LUT_4[62970] = 32'b00000000000000001110100111101001;
assign LUT_4[62971] = 32'b00000000000000000111110011100001;
assign LUT_4[62972] = 32'b00000000000000001100001101100001;
assign LUT_4[62973] = 32'b00000000000000000101011001011001;
assign LUT_4[62974] = 32'b00000000000000001011101000000101;
assign LUT_4[62975] = 32'b00000000000000000100110011111101;
assign LUT_4[62976] = 32'b00000000000000001111111111000100;
assign LUT_4[62977] = 32'b00000000000000001001001010111100;
assign LUT_4[62978] = 32'b00000000000000001111011001101000;
assign LUT_4[62979] = 32'b00000000000000001000100101100000;
assign LUT_4[62980] = 32'b00000000000000001100111111100000;
assign LUT_4[62981] = 32'b00000000000000000110001011011000;
assign LUT_4[62982] = 32'b00000000000000001100011010000100;
assign LUT_4[62983] = 32'b00000000000000000101100101111100;
assign LUT_4[62984] = 32'b00000000000000001001001011011001;
assign LUT_4[62985] = 32'b00000000000000000010010111010001;
assign LUT_4[62986] = 32'b00000000000000001000100101111101;
assign LUT_4[62987] = 32'b00000000000000000001110001110101;
assign LUT_4[62988] = 32'b00000000000000000110001011110101;
assign LUT_4[62989] = 32'b11111111111111111111010111101101;
assign LUT_4[62990] = 32'b00000000000000000101100110011001;
assign LUT_4[62991] = 32'b11111111111111111110110010010001;
assign LUT_4[62992] = 32'b00000000000000001101110000110010;
assign LUT_4[62993] = 32'b00000000000000000110111100101010;
assign LUT_4[62994] = 32'b00000000000000001101001011010110;
assign LUT_4[62995] = 32'b00000000000000000110010111001110;
assign LUT_4[62996] = 32'b00000000000000001010110001001110;
assign LUT_4[62997] = 32'b00000000000000000011111101000110;
assign LUT_4[62998] = 32'b00000000000000001010001011110010;
assign LUT_4[62999] = 32'b00000000000000000011010111101010;
assign LUT_4[63000] = 32'b00000000000000000110111101000111;
assign LUT_4[63001] = 32'b00000000000000000000001000111111;
assign LUT_4[63002] = 32'b00000000000000000110010111101011;
assign LUT_4[63003] = 32'b11111111111111111111100011100011;
assign LUT_4[63004] = 32'b00000000000000000011111101100011;
assign LUT_4[63005] = 32'b11111111111111111101001001011011;
assign LUT_4[63006] = 32'b00000000000000000011011000000111;
assign LUT_4[63007] = 32'b11111111111111111100100011111111;
assign LUT_4[63008] = 32'b00000000000000001110011010001011;
assign LUT_4[63009] = 32'b00000000000000000111100110000011;
assign LUT_4[63010] = 32'b00000000000000001101110100101111;
assign LUT_4[63011] = 32'b00000000000000000111000000100111;
assign LUT_4[63012] = 32'b00000000000000001011011010100111;
assign LUT_4[63013] = 32'b00000000000000000100100110011111;
assign LUT_4[63014] = 32'b00000000000000001010110101001011;
assign LUT_4[63015] = 32'b00000000000000000100000001000011;
assign LUT_4[63016] = 32'b00000000000000000111100110100000;
assign LUT_4[63017] = 32'b00000000000000000000110010011000;
assign LUT_4[63018] = 32'b00000000000000000111000001000100;
assign LUT_4[63019] = 32'b00000000000000000000001100111100;
assign LUT_4[63020] = 32'b00000000000000000100100110111100;
assign LUT_4[63021] = 32'b11111111111111111101110010110100;
assign LUT_4[63022] = 32'b00000000000000000100000001100000;
assign LUT_4[63023] = 32'b11111111111111111101001101011000;
assign LUT_4[63024] = 32'b00000000000000001100001011111001;
assign LUT_4[63025] = 32'b00000000000000000101010111110001;
assign LUT_4[63026] = 32'b00000000000000001011100110011101;
assign LUT_4[63027] = 32'b00000000000000000100110010010101;
assign LUT_4[63028] = 32'b00000000000000001001001100010101;
assign LUT_4[63029] = 32'b00000000000000000010011000001101;
assign LUT_4[63030] = 32'b00000000000000001000100110111001;
assign LUT_4[63031] = 32'b00000000000000000001110010110001;
assign LUT_4[63032] = 32'b00000000000000000101011000001110;
assign LUT_4[63033] = 32'b11111111111111111110100100000110;
assign LUT_4[63034] = 32'b00000000000000000100110010110010;
assign LUT_4[63035] = 32'b11111111111111111101111110101010;
assign LUT_4[63036] = 32'b00000000000000000010011000101010;
assign LUT_4[63037] = 32'b11111111111111111011100100100010;
assign LUT_4[63038] = 32'b00000000000000000001110011001110;
assign LUT_4[63039] = 32'b11111111111111111010111111000110;
assign LUT_4[63040] = 32'b00000000000000010001010110011000;
assign LUT_4[63041] = 32'b00000000000000001010100010010000;
assign LUT_4[63042] = 32'b00000000000000010000110000111100;
assign LUT_4[63043] = 32'b00000000000000001001111100110100;
assign LUT_4[63044] = 32'b00000000000000001110010110110100;
assign LUT_4[63045] = 32'b00000000000000000111100010101100;
assign LUT_4[63046] = 32'b00000000000000001101110001011000;
assign LUT_4[63047] = 32'b00000000000000000110111101010000;
assign LUT_4[63048] = 32'b00000000000000001010100010101101;
assign LUT_4[63049] = 32'b00000000000000000011101110100101;
assign LUT_4[63050] = 32'b00000000000000001001111101010001;
assign LUT_4[63051] = 32'b00000000000000000011001001001001;
assign LUT_4[63052] = 32'b00000000000000000111100011001001;
assign LUT_4[63053] = 32'b00000000000000000000101111000001;
assign LUT_4[63054] = 32'b00000000000000000110111101101101;
assign LUT_4[63055] = 32'b00000000000000000000001001100101;
assign LUT_4[63056] = 32'b00000000000000001111001000000110;
assign LUT_4[63057] = 32'b00000000000000001000010011111110;
assign LUT_4[63058] = 32'b00000000000000001110100010101010;
assign LUT_4[63059] = 32'b00000000000000000111101110100010;
assign LUT_4[63060] = 32'b00000000000000001100001000100010;
assign LUT_4[63061] = 32'b00000000000000000101010100011010;
assign LUT_4[63062] = 32'b00000000000000001011100011000110;
assign LUT_4[63063] = 32'b00000000000000000100101110111110;
assign LUT_4[63064] = 32'b00000000000000001000010100011011;
assign LUT_4[63065] = 32'b00000000000000000001100000010011;
assign LUT_4[63066] = 32'b00000000000000000111101110111111;
assign LUT_4[63067] = 32'b00000000000000000000111010110111;
assign LUT_4[63068] = 32'b00000000000000000101010100110111;
assign LUT_4[63069] = 32'b11111111111111111110100000101111;
assign LUT_4[63070] = 32'b00000000000000000100101111011011;
assign LUT_4[63071] = 32'b11111111111111111101111011010011;
assign LUT_4[63072] = 32'b00000000000000001111110001011111;
assign LUT_4[63073] = 32'b00000000000000001000111101010111;
assign LUT_4[63074] = 32'b00000000000000001111001100000011;
assign LUT_4[63075] = 32'b00000000000000001000010111111011;
assign LUT_4[63076] = 32'b00000000000000001100110001111011;
assign LUT_4[63077] = 32'b00000000000000000101111101110011;
assign LUT_4[63078] = 32'b00000000000000001100001100011111;
assign LUT_4[63079] = 32'b00000000000000000101011000010111;
assign LUT_4[63080] = 32'b00000000000000001000111101110100;
assign LUT_4[63081] = 32'b00000000000000000010001001101100;
assign LUT_4[63082] = 32'b00000000000000001000011000011000;
assign LUT_4[63083] = 32'b00000000000000000001100100010000;
assign LUT_4[63084] = 32'b00000000000000000101111110010000;
assign LUT_4[63085] = 32'b11111111111111111111001010001000;
assign LUT_4[63086] = 32'b00000000000000000101011000110100;
assign LUT_4[63087] = 32'b11111111111111111110100100101100;
assign LUT_4[63088] = 32'b00000000000000001101100011001101;
assign LUT_4[63089] = 32'b00000000000000000110101111000101;
assign LUT_4[63090] = 32'b00000000000000001100111101110001;
assign LUT_4[63091] = 32'b00000000000000000110001001101001;
assign LUT_4[63092] = 32'b00000000000000001010100011101001;
assign LUT_4[63093] = 32'b00000000000000000011101111100001;
assign LUT_4[63094] = 32'b00000000000000001001111110001101;
assign LUT_4[63095] = 32'b00000000000000000011001010000101;
assign LUT_4[63096] = 32'b00000000000000000110101111100010;
assign LUT_4[63097] = 32'b11111111111111111111111011011010;
assign LUT_4[63098] = 32'b00000000000000000110001010000110;
assign LUT_4[63099] = 32'b11111111111111111111010101111110;
assign LUT_4[63100] = 32'b00000000000000000011101111111110;
assign LUT_4[63101] = 32'b11111111111111111100111011110110;
assign LUT_4[63102] = 32'b00000000000000000011001010100010;
assign LUT_4[63103] = 32'b11111111111111111100010110011010;
assign LUT_4[63104] = 32'b00000000000000010010100101001100;
assign LUT_4[63105] = 32'b00000000000000001011110001000100;
assign LUT_4[63106] = 32'b00000000000000010001111111110000;
assign LUT_4[63107] = 32'b00000000000000001011001011101000;
assign LUT_4[63108] = 32'b00000000000000001111100101101000;
assign LUT_4[63109] = 32'b00000000000000001000110001100000;
assign LUT_4[63110] = 32'b00000000000000001111000000001100;
assign LUT_4[63111] = 32'b00000000000000001000001100000100;
assign LUT_4[63112] = 32'b00000000000000001011110001100001;
assign LUT_4[63113] = 32'b00000000000000000100111101011001;
assign LUT_4[63114] = 32'b00000000000000001011001100000101;
assign LUT_4[63115] = 32'b00000000000000000100010111111101;
assign LUT_4[63116] = 32'b00000000000000001000110001111101;
assign LUT_4[63117] = 32'b00000000000000000001111101110101;
assign LUT_4[63118] = 32'b00000000000000001000001100100001;
assign LUT_4[63119] = 32'b00000000000000000001011000011001;
assign LUT_4[63120] = 32'b00000000000000010000010110111010;
assign LUT_4[63121] = 32'b00000000000000001001100010110010;
assign LUT_4[63122] = 32'b00000000000000001111110001011110;
assign LUT_4[63123] = 32'b00000000000000001000111101010110;
assign LUT_4[63124] = 32'b00000000000000001101010111010110;
assign LUT_4[63125] = 32'b00000000000000000110100011001110;
assign LUT_4[63126] = 32'b00000000000000001100110001111010;
assign LUT_4[63127] = 32'b00000000000000000101111101110010;
assign LUT_4[63128] = 32'b00000000000000001001100011001111;
assign LUT_4[63129] = 32'b00000000000000000010101111000111;
assign LUT_4[63130] = 32'b00000000000000001000111101110011;
assign LUT_4[63131] = 32'b00000000000000000010001001101011;
assign LUT_4[63132] = 32'b00000000000000000110100011101011;
assign LUT_4[63133] = 32'b11111111111111111111101111100011;
assign LUT_4[63134] = 32'b00000000000000000101111110001111;
assign LUT_4[63135] = 32'b11111111111111111111001010000111;
assign LUT_4[63136] = 32'b00000000000000010001000000010011;
assign LUT_4[63137] = 32'b00000000000000001010001100001011;
assign LUT_4[63138] = 32'b00000000000000010000011010110111;
assign LUT_4[63139] = 32'b00000000000000001001100110101111;
assign LUT_4[63140] = 32'b00000000000000001110000000101111;
assign LUT_4[63141] = 32'b00000000000000000111001100100111;
assign LUT_4[63142] = 32'b00000000000000001101011011010011;
assign LUT_4[63143] = 32'b00000000000000000110100111001011;
assign LUT_4[63144] = 32'b00000000000000001010001100101000;
assign LUT_4[63145] = 32'b00000000000000000011011000100000;
assign LUT_4[63146] = 32'b00000000000000001001100111001100;
assign LUT_4[63147] = 32'b00000000000000000010110011000100;
assign LUT_4[63148] = 32'b00000000000000000111001101000100;
assign LUT_4[63149] = 32'b00000000000000000000011000111100;
assign LUT_4[63150] = 32'b00000000000000000110100111101000;
assign LUT_4[63151] = 32'b11111111111111111111110011100000;
assign LUT_4[63152] = 32'b00000000000000001110110010000001;
assign LUT_4[63153] = 32'b00000000000000000111111101111001;
assign LUT_4[63154] = 32'b00000000000000001110001100100101;
assign LUT_4[63155] = 32'b00000000000000000111011000011101;
assign LUT_4[63156] = 32'b00000000000000001011110010011101;
assign LUT_4[63157] = 32'b00000000000000000100111110010101;
assign LUT_4[63158] = 32'b00000000000000001011001101000001;
assign LUT_4[63159] = 32'b00000000000000000100011000111001;
assign LUT_4[63160] = 32'b00000000000000000111111110010110;
assign LUT_4[63161] = 32'b00000000000000000001001010001110;
assign LUT_4[63162] = 32'b00000000000000000111011000111010;
assign LUT_4[63163] = 32'b00000000000000000000100100110010;
assign LUT_4[63164] = 32'b00000000000000000100111110110010;
assign LUT_4[63165] = 32'b11111111111111111110001010101010;
assign LUT_4[63166] = 32'b00000000000000000100011001010110;
assign LUT_4[63167] = 32'b11111111111111111101100101001110;
assign LUT_4[63168] = 32'b00000000000000010011111100100000;
assign LUT_4[63169] = 32'b00000000000000001101001000011000;
assign LUT_4[63170] = 32'b00000000000000010011010111000100;
assign LUT_4[63171] = 32'b00000000000000001100100010111100;
assign LUT_4[63172] = 32'b00000000000000010000111100111100;
assign LUT_4[63173] = 32'b00000000000000001010001000110100;
assign LUT_4[63174] = 32'b00000000000000010000010111100000;
assign LUT_4[63175] = 32'b00000000000000001001100011011000;
assign LUT_4[63176] = 32'b00000000000000001101001000110101;
assign LUT_4[63177] = 32'b00000000000000000110010100101101;
assign LUT_4[63178] = 32'b00000000000000001100100011011001;
assign LUT_4[63179] = 32'b00000000000000000101101111010001;
assign LUT_4[63180] = 32'b00000000000000001010001001010001;
assign LUT_4[63181] = 32'b00000000000000000011010101001001;
assign LUT_4[63182] = 32'b00000000000000001001100011110101;
assign LUT_4[63183] = 32'b00000000000000000010101111101101;
assign LUT_4[63184] = 32'b00000000000000010001101110001110;
assign LUT_4[63185] = 32'b00000000000000001010111010000110;
assign LUT_4[63186] = 32'b00000000000000010001001000110010;
assign LUT_4[63187] = 32'b00000000000000001010010100101010;
assign LUT_4[63188] = 32'b00000000000000001110101110101010;
assign LUT_4[63189] = 32'b00000000000000000111111010100010;
assign LUT_4[63190] = 32'b00000000000000001110001001001110;
assign LUT_4[63191] = 32'b00000000000000000111010101000110;
assign LUT_4[63192] = 32'b00000000000000001010111010100011;
assign LUT_4[63193] = 32'b00000000000000000100000110011011;
assign LUT_4[63194] = 32'b00000000000000001010010101000111;
assign LUT_4[63195] = 32'b00000000000000000011100000111111;
assign LUT_4[63196] = 32'b00000000000000000111111010111111;
assign LUT_4[63197] = 32'b00000000000000000001000110110111;
assign LUT_4[63198] = 32'b00000000000000000111010101100011;
assign LUT_4[63199] = 32'b00000000000000000000100001011011;
assign LUT_4[63200] = 32'b00000000000000010010010111100111;
assign LUT_4[63201] = 32'b00000000000000001011100011011111;
assign LUT_4[63202] = 32'b00000000000000010001110010001011;
assign LUT_4[63203] = 32'b00000000000000001010111110000011;
assign LUT_4[63204] = 32'b00000000000000001111011000000011;
assign LUT_4[63205] = 32'b00000000000000001000100011111011;
assign LUT_4[63206] = 32'b00000000000000001110110010100111;
assign LUT_4[63207] = 32'b00000000000000000111111110011111;
assign LUT_4[63208] = 32'b00000000000000001011100011111100;
assign LUT_4[63209] = 32'b00000000000000000100101111110100;
assign LUT_4[63210] = 32'b00000000000000001010111110100000;
assign LUT_4[63211] = 32'b00000000000000000100001010011000;
assign LUT_4[63212] = 32'b00000000000000001000100100011000;
assign LUT_4[63213] = 32'b00000000000000000001110000010000;
assign LUT_4[63214] = 32'b00000000000000000111111110111100;
assign LUT_4[63215] = 32'b00000000000000000001001010110100;
assign LUT_4[63216] = 32'b00000000000000010000001001010101;
assign LUT_4[63217] = 32'b00000000000000001001010101001101;
assign LUT_4[63218] = 32'b00000000000000001111100011111001;
assign LUT_4[63219] = 32'b00000000000000001000101111110001;
assign LUT_4[63220] = 32'b00000000000000001101001001110001;
assign LUT_4[63221] = 32'b00000000000000000110010101101001;
assign LUT_4[63222] = 32'b00000000000000001100100100010101;
assign LUT_4[63223] = 32'b00000000000000000101110000001101;
assign LUT_4[63224] = 32'b00000000000000001001010101101010;
assign LUT_4[63225] = 32'b00000000000000000010100001100010;
assign LUT_4[63226] = 32'b00000000000000001000110000001110;
assign LUT_4[63227] = 32'b00000000000000000001111100000110;
assign LUT_4[63228] = 32'b00000000000000000110010110000110;
assign LUT_4[63229] = 32'b11111111111111111111100001111110;
assign LUT_4[63230] = 32'b00000000000000000101110000101010;
assign LUT_4[63231] = 32'b11111111111111111110111100100010;
assign LUT_4[63232] = 32'b00000000000000010100111010100111;
assign LUT_4[63233] = 32'b00000000000000001110000110011111;
assign LUT_4[63234] = 32'b00000000000000010100010101001011;
assign LUT_4[63235] = 32'b00000000000000001101100001000011;
assign LUT_4[63236] = 32'b00000000000000010001111011000011;
assign LUT_4[63237] = 32'b00000000000000001011000110111011;
assign LUT_4[63238] = 32'b00000000000000010001010101100111;
assign LUT_4[63239] = 32'b00000000000000001010100001011111;
assign LUT_4[63240] = 32'b00000000000000001110000110111100;
assign LUT_4[63241] = 32'b00000000000000000111010010110100;
assign LUT_4[63242] = 32'b00000000000000001101100001100000;
assign LUT_4[63243] = 32'b00000000000000000110101101011000;
assign LUT_4[63244] = 32'b00000000000000001011000111011000;
assign LUT_4[63245] = 32'b00000000000000000100010011010000;
assign LUT_4[63246] = 32'b00000000000000001010100001111100;
assign LUT_4[63247] = 32'b00000000000000000011101101110100;
assign LUT_4[63248] = 32'b00000000000000010010101100010101;
assign LUT_4[63249] = 32'b00000000000000001011111000001101;
assign LUT_4[63250] = 32'b00000000000000010010000110111001;
assign LUT_4[63251] = 32'b00000000000000001011010010110001;
assign LUT_4[63252] = 32'b00000000000000001111101100110001;
assign LUT_4[63253] = 32'b00000000000000001000111000101001;
assign LUT_4[63254] = 32'b00000000000000001111000111010101;
assign LUT_4[63255] = 32'b00000000000000001000010011001101;
assign LUT_4[63256] = 32'b00000000000000001011111000101010;
assign LUT_4[63257] = 32'b00000000000000000101000100100010;
assign LUT_4[63258] = 32'b00000000000000001011010011001110;
assign LUT_4[63259] = 32'b00000000000000000100011111000110;
assign LUT_4[63260] = 32'b00000000000000001000111001000110;
assign LUT_4[63261] = 32'b00000000000000000010000100111110;
assign LUT_4[63262] = 32'b00000000000000001000010011101010;
assign LUT_4[63263] = 32'b00000000000000000001011111100010;
assign LUT_4[63264] = 32'b00000000000000010011010101101110;
assign LUT_4[63265] = 32'b00000000000000001100100001100110;
assign LUT_4[63266] = 32'b00000000000000010010110000010010;
assign LUT_4[63267] = 32'b00000000000000001011111100001010;
assign LUT_4[63268] = 32'b00000000000000010000010110001010;
assign LUT_4[63269] = 32'b00000000000000001001100010000010;
assign LUT_4[63270] = 32'b00000000000000001111110000101110;
assign LUT_4[63271] = 32'b00000000000000001000111100100110;
assign LUT_4[63272] = 32'b00000000000000001100100010000011;
assign LUT_4[63273] = 32'b00000000000000000101101101111011;
assign LUT_4[63274] = 32'b00000000000000001011111100100111;
assign LUT_4[63275] = 32'b00000000000000000101001000011111;
assign LUT_4[63276] = 32'b00000000000000001001100010011111;
assign LUT_4[63277] = 32'b00000000000000000010101110010111;
assign LUT_4[63278] = 32'b00000000000000001000111101000011;
assign LUT_4[63279] = 32'b00000000000000000010001000111011;
assign LUT_4[63280] = 32'b00000000000000010001000111011100;
assign LUT_4[63281] = 32'b00000000000000001010010011010100;
assign LUT_4[63282] = 32'b00000000000000010000100010000000;
assign LUT_4[63283] = 32'b00000000000000001001101101111000;
assign LUT_4[63284] = 32'b00000000000000001110000111111000;
assign LUT_4[63285] = 32'b00000000000000000111010011110000;
assign LUT_4[63286] = 32'b00000000000000001101100010011100;
assign LUT_4[63287] = 32'b00000000000000000110101110010100;
assign LUT_4[63288] = 32'b00000000000000001010010011110001;
assign LUT_4[63289] = 32'b00000000000000000011011111101001;
assign LUT_4[63290] = 32'b00000000000000001001101110010101;
assign LUT_4[63291] = 32'b00000000000000000010111010001101;
assign LUT_4[63292] = 32'b00000000000000000111010100001101;
assign LUT_4[63293] = 32'b00000000000000000000100000000101;
assign LUT_4[63294] = 32'b00000000000000000110101110110001;
assign LUT_4[63295] = 32'b11111111111111111111111010101001;
assign LUT_4[63296] = 32'b00000000000000010110010001111011;
assign LUT_4[63297] = 32'b00000000000000001111011101110011;
assign LUT_4[63298] = 32'b00000000000000010101101100011111;
assign LUT_4[63299] = 32'b00000000000000001110111000010111;
assign LUT_4[63300] = 32'b00000000000000010011010010010111;
assign LUT_4[63301] = 32'b00000000000000001100011110001111;
assign LUT_4[63302] = 32'b00000000000000010010101100111011;
assign LUT_4[63303] = 32'b00000000000000001011111000110011;
assign LUT_4[63304] = 32'b00000000000000001111011110010000;
assign LUT_4[63305] = 32'b00000000000000001000101010001000;
assign LUT_4[63306] = 32'b00000000000000001110111000110100;
assign LUT_4[63307] = 32'b00000000000000001000000100101100;
assign LUT_4[63308] = 32'b00000000000000001100011110101100;
assign LUT_4[63309] = 32'b00000000000000000101101010100100;
assign LUT_4[63310] = 32'b00000000000000001011111001010000;
assign LUT_4[63311] = 32'b00000000000000000101000101001000;
assign LUT_4[63312] = 32'b00000000000000010100000011101001;
assign LUT_4[63313] = 32'b00000000000000001101001111100001;
assign LUT_4[63314] = 32'b00000000000000010011011110001101;
assign LUT_4[63315] = 32'b00000000000000001100101010000101;
assign LUT_4[63316] = 32'b00000000000000010001000100000101;
assign LUT_4[63317] = 32'b00000000000000001010001111111101;
assign LUT_4[63318] = 32'b00000000000000010000011110101001;
assign LUT_4[63319] = 32'b00000000000000001001101010100001;
assign LUT_4[63320] = 32'b00000000000000001101001111111110;
assign LUT_4[63321] = 32'b00000000000000000110011011110110;
assign LUT_4[63322] = 32'b00000000000000001100101010100010;
assign LUT_4[63323] = 32'b00000000000000000101110110011010;
assign LUT_4[63324] = 32'b00000000000000001010010000011010;
assign LUT_4[63325] = 32'b00000000000000000011011100010010;
assign LUT_4[63326] = 32'b00000000000000001001101010111110;
assign LUT_4[63327] = 32'b00000000000000000010110110110110;
assign LUT_4[63328] = 32'b00000000000000010100101101000010;
assign LUT_4[63329] = 32'b00000000000000001101111000111010;
assign LUT_4[63330] = 32'b00000000000000010100000111100110;
assign LUT_4[63331] = 32'b00000000000000001101010011011110;
assign LUT_4[63332] = 32'b00000000000000010001101101011110;
assign LUT_4[63333] = 32'b00000000000000001010111001010110;
assign LUT_4[63334] = 32'b00000000000000010001001000000010;
assign LUT_4[63335] = 32'b00000000000000001010010011111010;
assign LUT_4[63336] = 32'b00000000000000001101111001010111;
assign LUT_4[63337] = 32'b00000000000000000111000101001111;
assign LUT_4[63338] = 32'b00000000000000001101010011111011;
assign LUT_4[63339] = 32'b00000000000000000110011111110011;
assign LUT_4[63340] = 32'b00000000000000001010111001110011;
assign LUT_4[63341] = 32'b00000000000000000100000101101011;
assign LUT_4[63342] = 32'b00000000000000001010010100010111;
assign LUT_4[63343] = 32'b00000000000000000011100000001111;
assign LUT_4[63344] = 32'b00000000000000010010011110110000;
assign LUT_4[63345] = 32'b00000000000000001011101010101000;
assign LUT_4[63346] = 32'b00000000000000010001111001010100;
assign LUT_4[63347] = 32'b00000000000000001011000101001100;
assign LUT_4[63348] = 32'b00000000000000001111011111001100;
assign LUT_4[63349] = 32'b00000000000000001000101011000100;
assign LUT_4[63350] = 32'b00000000000000001110111001110000;
assign LUT_4[63351] = 32'b00000000000000001000000101101000;
assign LUT_4[63352] = 32'b00000000000000001011101011000101;
assign LUT_4[63353] = 32'b00000000000000000100110110111101;
assign LUT_4[63354] = 32'b00000000000000001011000101101001;
assign LUT_4[63355] = 32'b00000000000000000100010001100001;
assign LUT_4[63356] = 32'b00000000000000001000101011100001;
assign LUT_4[63357] = 32'b00000000000000000001110111011001;
assign LUT_4[63358] = 32'b00000000000000001000000110000101;
assign LUT_4[63359] = 32'b00000000000000000001010001111101;
assign LUT_4[63360] = 32'b00000000000000010111100000101111;
assign LUT_4[63361] = 32'b00000000000000010000101100100111;
assign LUT_4[63362] = 32'b00000000000000010110111011010011;
assign LUT_4[63363] = 32'b00000000000000010000000111001011;
assign LUT_4[63364] = 32'b00000000000000010100100001001011;
assign LUT_4[63365] = 32'b00000000000000001101101101000011;
assign LUT_4[63366] = 32'b00000000000000010011111011101111;
assign LUT_4[63367] = 32'b00000000000000001101000111100111;
assign LUT_4[63368] = 32'b00000000000000010000101101000100;
assign LUT_4[63369] = 32'b00000000000000001001111000111100;
assign LUT_4[63370] = 32'b00000000000000010000000111101000;
assign LUT_4[63371] = 32'b00000000000000001001010011100000;
assign LUT_4[63372] = 32'b00000000000000001101101101100000;
assign LUT_4[63373] = 32'b00000000000000000110111001011000;
assign LUT_4[63374] = 32'b00000000000000001101001000000100;
assign LUT_4[63375] = 32'b00000000000000000110010011111100;
assign LUT_4[63376] = 32'b00000000000000010101010010011101;
assign LUT_4[63377] = 32'b00000000000000001110011110010101;
assign LUT_4[63378] = 32'b00000000000000010100101101000001;
assign LUT_4[63379] = 32'b00000000000000001101111000111001;
assign LUT_4[63380] = 32'b00000000000000010010010010111001;
assign LUT_4[63381] = 32'b00000000000000001011011110110001;
assign LUT_4[63382] = 32'b00000000000000010001101101011101;
assign LUT_4[63383] = 32'b00000000000000001010111001010101;
assign LUT_4[63384] = 32'b00000000000000001110011110110010;
assign LUT_4[63385] = 32'b00000000000000000111101010101010;
assign LUT_4[63386] = 32'b00000000000000001101111001010110;
assign LUT_4[63387] = 32'b00000000000000000111000101001110;
assign LUT_4[63388] = 32'b00000000000000001011011111001110;
assign LUT_4[63389] = 32'b00000000000000000100101011000110;
assign LUT_4[63390] = 32'b00000000000000001010111001110010;
assign LUT_4[63391] = 32'b00000000000000000100000101101010;
assign LUT_4[63392] = 32'b00000000000000010101111011110110;
assign LUT_4[63393] = 32'b00000000000000001111000111101110;
assign LUT_4[63394] = 32'b00000000000000010101010110011010;
assign LUT_4[63395] = 32'b00000000000000001110100010010010;
assign LUT_4[63396] = 32'b00000000000000010010111100010010;
assign LUT_4[63397] = 32'b00000000000000001100001000001010;
assign LUT_4[63398] = 32'b00000000000000010010010110110110;
assign LUT_4[63399] = 32'b00000000000000001011100010101110;
assign LUT_4[63400] = 32'b00000000000000001111001000001011;
assign LUT_4[63401] = 32'b00000000000000001000010100000011;
assign LUT_4[63402] = 32'b00000000000000001110100010101111;
assign LUT_4[63403] = 32'b00000000000000000111101110100111;
assign LUT_4[63404] = 32'b00000000000000001100001000100111;
assign LUT_4[63405] = 32'b00000000000000000101010100011111;
assign LUT_4[63406] = 32'b00000000000000001011100011001011;
assign LUT_4[63407] = 32'b00000000000000000100101111000011;
assign LUT_4[63408] = 32'b00000000000000010011101101100100;
assign LUT_4[63409] = 32'b00000000000000001100111001011100;
assign LUT_4[63410] = 32'b00000000000000010011001000001000;
assign LUT_4[63411] = 32'b00000000000000001100010100000000;
assign LUT_4[63412] = 32'b00000000000000010000101110000000;
assign LUT_4[63413] = 32'b00000000000000001001111001111000;
assign LUT_4[63414] = 32'b00000000000000010000001000100100;
assign LUT_4[63415] = 32'b00000000000000001001010100011100;
assign LUT_4[63416] = 32'b00000000000000001100111001111001;
assign LUT_4[63417] = 32'b00000000000000000110000101110001;
assign LUT_4[63418] = 32'b00000000000000001100010100011101;
assign LUT_4[63419] = 32'b00000000000000000101100000010101;
assign LUT_4[63420] = 32'b00000000000000001001111010010101;
assign LUT_4[63421] = 32'b00000000000000000011000110001101;
assign LUT_4[63422] = 32'b00000000000000001001010100111001;
assign LUT_4[63423] = 32'b00000000000000000010100000110001;
assign LUT_4[63424] = 32'b00000000000000011000111000000011;
assign LUT_4[63425] = 32'b00000000000000010010000011111011;
assign LUT_4[63426] = 32'b00000000000000011000010010100111;
assign LUT_4[63427] = 32'b00000000000000010001011110011111;
assign LUT_4[63428] = 32'b00000000000000010101111000011111;
assign LUT_4[63429] = 32'b00000000000000001111000100010111;
assign LUT_4[63430] = 32'b00000000000000010101010011000011;
assign LUT_4[63431] = 32'b00000000000000001110011110111011;
assign LUT_4[63432] = 32'b00000000000000010010000100011000;
assign LUT_4[63433] = 32'b00000000000000001011010000010000;
assign LUT_4[63434] = 32'b00000000000000010001011110111100;
assign LUT_4[63435] = 32'b00000000000000001010101010110100;
assign LUT_4[63436] = 32'b00000000000000001111000100110100;
assign LUT_4[63437] = 32'b00000000000000001000010000101100;
assign LUT_4[63438] = 32'b00000000000000001110011111011000;
assign LUT_4[63439] = 32'b00000000000000000111101011010000;
assign LUT_4[63440] = 32'b00000000000000010110101001110001;
assign LUT_4[63441] = 32'b00000000000000001111110101101001;
assign LUT_4[63442] = 32'b00000000000000010110000100010101;
assign LUT_4[63443] = 32'b00000000000000001111010000001101;
assign LUT_4[63444] = 32'b00000000000000010011101010001101;
assign LUT_4[63445] = 32'b00000000000000001100110110000101;
assign LUT_4[63446] = 32'b00000000000000010011000100110001;
assign LUT_4[63447] = 32'b00000000000000001100010000101001;
assign LUT_4[63448] = 32'b00000000000000001111110110000110;
assign LUT_4[63449] = 32'b00000000000000001001000001111110;
assign LUT_4[63450] = 32'b00000000000000001111010000101010;
assign LUT_4[63451] = 32'b00000000000000001000011100100010;
assign LUT_4[63452] = 32'b00000000000000001100110110100010;
assign LUT_4[63453] = 32'b00000000000000000110000010011010;
assign LUT_4[63454] = 32'b00000000000000001100010001000110;
assign LUT_4[63455] = 32'b00000000000000000101011100111110;
assign LUT_4[63456] = 32'b00000000000000010111010011001010;
assign LUT_4[63457] = 32'b00000000000000010000011111000010;
assign LUT_4[63458] = 32'b00000000000000010110101101101110;
assign LUT_4[63459] = 32'b00000000000000001111111001100110;
assign LUT_4[63460] = 32'b00000000000000010100010011100110;
assign LUT_4[63461] = 32'b00000000000000001101011111011110;
assign LUT_4[63462] = 32'b00000000000000010011101110001010;
assign LUT_4[63463] = 32'b00000000000000001100111010000010;
assign LUT_4[63464] = 32'b00000000000000010000011111011111;
assign LUT_4[63465] = 32'b00000000000000001001101011010111;
assign LUT_4[63466] = 32'b00000000000000001111111010000011;
assign LUT_4[63467] = 32'b00000000000000001001000101111011;
assign LUT_4[63468] = 32'b00000000000000001101011111111011;
assign LUT_4[63469] = 32'b00000000000000000110101011110011;
assign LUT_4[63470] = 32'b00000000000000001100111010011111;
assign LUT_4[63471] = 32'b00000000000000000110000110010111;
assign LUT_4[63472] = 32'b00000000000000010101000100111000;
assign LUT_4[63473] = 32'b00000000000000001110010000110000;
assign LUT_4[63474] = 32'b00000000000000010100011111011100;
assign LUT_4[63475] = 32'b00000000000000001101101011010100;
assign LUT_4[63476] = 32'b00000000000000010010000101010100;
assign LUT_4[63477] = 32'b00000000000000001011010001001100;
assign LUT_4[63478] = 32'b00000000000000010001011111111000;
assign LUT_4[63479] = 32'b00000000000000001010101011110000;
assign LUT_4[63480] = 32'b00000000000000001110010001001101;
assign LUT_4[63481] = 32'b00000000000000000111011101000101;
assign LUT_4[63482] = 32'b00000000000000001101101011110001;
assign LUT_4[63483] = 32'b00000000000000000110110111101001;
assign LUT_4[63484] = 32'b00000000000000001011010001101001;
assign LUT_4[63485] = 32'b00000000000000000100011101100001;
assign LUT_4[63486] = 32'b00000000000000001010101100001101;
assign LUT_4[63487] = 32'b00000000000000000011111000000101;
assign LUT_4[63488] = 32'b00000000000000001010101111100111;
assign LUT_4[63489] = 32'b00000000000000000011111011011111;
assign LUT_4[63490] = 32'b00000000000000001010001010001011;
assign LUT_4[63491] = 32'b00000000000000000011010110000011;
assign LUT_4[63492] = 32'b00000000000000000111110000000011;
assign LUT_4[63493] = 32'b00000000000000000000111011111011;
assign LUT_4[63494] = 32'b00000000000000000111001010100111;
assign LUT_4[63495] = 32'b00000000000000000000010110011111;
assign LUT_4[63496] = 32'b00000000000000000011111011111100;
assign LUT_4[63497] = 32'b11111111111111111101000111110100;
assign LUT_4[63498] = 32'b00000000000000000011010110100000;
assign LUT_4[63499] = 32'b11111111111111111100100010011000;
assign LUT_4[63500] = 32'b00000000000000000000111100011000;
assign LUT_4[63501] = 32'b11111111111111111010001000010000;
assign LUT_4[63502] = 32'b00000000000000000000010110111100;
assign LUT_4[63503] = 32'b11111111111111111001100010110100;
assign LUT_4[63504] = 32'b00000000000000001000100001010101;
assign LUT_4[63505] = 32'b00000000000000000001101101001101;
assign LUT_4[63506] = 32'b00000000000000000111111011111001;
assign LUT_4[63507] = 32'b00000000000000000001000111110001;
assign LUT_4[63508] = 32'b00000000000000000101100001110001;
assign LUT_4[63509] = 32'b11111111111111111110101101101001;
assign LUT_4[63510] = 32'b00000000000000000100111100010101;
assign LUT_4[63511] = 32'b11111111111111111110001000001101;
assign LUT_4[63512] = 32'b00000000000000000001101101101010;
assign LUT_4[63513] = 32'b11111111111111111010111001100010;
assign LUT_4[63514] = 32'b00000000000000000001001000001110;
assign LUT_4[63515] = 32'b11111111111111111010010100000110;
assign LUT_4[63516] = 32'b11111111111111111110101110000110;
assign LUT_4[63517] = 32'b11111111111111110111111001111110;
assign LUT_4[63518] = 32'b11111111111111111110001000101010;
assign LUT_4[63519] = 32'b11111111111111110111010100100010;
assign LUT_4[63520] = 32'b00000000000000001001001010101110;
assign LUT_4[63521] = 32'b00000000000000000010010110100110;
assign LUT_4[63522] = 32'b00000000000000001000100101010010;
assign LUT_4[63523] = 32'b00000000000000000001110001001010;
assign LUT_4[63524] = 32'b00000000000000000110001011001010;
assign LUT_4[63525] = 32'b11111111111111111111010111000010;
assign LUT_4[63526] = 32'b00000000000000000101100101101110;
assign LUT_4[63527] = 32'b11111111111111111110110001100110;
assign LUT_4[63528] = 32'b00000000000000000010010111000011;
assign LUT_4[63529] = 32'b11111111111111111011100010111011;
assign LUT_4[63530] = 32'b00000000000000000001110001100111;
assign LUT_4[63531] = 32'b11111111111111111010111101011111;
assign LUT_4[63532] = 32'b11111111111111111111010111011111;
assign LUT_4[63533] = 32'b11111111111111111000100011010111;
assign LUT_4[63534] = 32'b11111111111111111110110010000011;
assign LUT_4[63535] = 32'b11111111111111110111111101111011;
assign LUT_4[63536] = 32'b00000000000000000110111100011100;
assign LUT_4[63537] = 32'b00000000000000000000001000010100;
assign LUT_4[63538] = 32'b00000000000000000110010111000000;
assign LUT_4[63539] = 32'b11111111111111111111100010111000;
assign LUT_4[63540] = 32'b00000000000000000011111100111000;
assign LUT_4[63541] = 32'b11111111111111111101001000110000;
assign LUT_4[63542] = 32'b00000000000000000011010111011100;
assign LUT_4[63543] = 32'b11111111111111111100100011010100;
assign LUT_4[63544] = 32'b00000000000000000000001000110001;
assign LUT_4[63545] = 32'b11111111111111111001010100101001;
assign LUT_4[63546] = 32'b11111111111111111111100011010101;
assign LUT_4[63547] = 32'b11111111111111111000101111001101;
assign LUT_4[63548] = 32'b11111111111111111101001001001101;
assign LUT_4[63549] = 32'b11111111111111110110010101000101;
assign LUT_4[63550] = 32'b11111111111111111100100011110001;
assign LUT_4[63551] = 32'b11111111111111110101101111101001;
assign LUT_4[63552] = 32'b00000000000000001100000110111011;
assign LUT_4[63553] = 32'b00000000000000000101010010110011;
assign LUT_4[63554] = 32'b00000000000000001011100001011111;
assign LUT_4[63555] = 32'b00000000000000000100101101010111;
assign LUT_4[63556] = 32'b00000000000000001001000111010111;
assign LUT_4[63557] = 32'b00000000000000000010010011001111;
assign LUT_4[63558] = 32'b00000000000000001000100001111011;
assign LUT_4[63559] = 32'b00000000000000000001101101110011;
assign LUT_4[63560] = 32'b00000000000000000101010011010000;
assign LUT_4[63561] = 32'b11111111111111111110011111001000;
assign LUT_4[63562] = 32'b00000000000000000100101101110100;
assign LUT_4[63563] = 32'b11111111111111111101111001101100;
assign LUT_4[63564] = 32'b00000000000000000010010011101100;
assign LUT_4[63565] = 32'b11111111111111111011011111100100;
assign LUT_4[63566] = 32'b00000000000000000001101110010000;
assign LUT_4[63567] = 32'b11111111111111111010111010001000;
assign LUT_4[63568] = 32'b00000000000000001001111000101001;
assign LUT_4[63569] = 32'b00000000000000000011000100100001;
assign LUT_4[63570] = 32'b00000000000000001001010011001101;
assign LUT_4[63571] = 32'b00000000000000000010011111000101;
assign LUT_4[63572] = 32'b00000000000000000110111001000101;
assign LUT_4[63573] = 32'b00000000000000000000000100111101;
assign LUT_4[63574] = 32'b00000000000000000110010011101001;
assign LUT_4[63575] = 32'b11111111111111111111011111100001;
assign LUT_4[63576] = 32'b00000000000000000011000100111110;
assign LUT_4[63577] = 32'b11111111111111111100010000110110;
assign LUT_4[63578] = 32'b00000000000000000010011111100010;
assign LUT_4[63579] = 32'b11111111111111111011101011011010;
assign LUT_4[63580] = 32'b00000000000000000000000101011010;
assign LUT_4[63581] = 32'b11111111111111111001010001010010;
assign LUT_4[63582] = 32'b11111111111111111111011111111110;
assign LUT_4[63583] = 32'b11111111111111111000101011110110;
assign LUT_4[63584] = 32'b00000000000000001010100010000010;
assign LUT_4[63585] = 32'b00000000000000000011101101111010;
assign LUT_4[63586] = 32'b00000000000000001001111100100110;
assign LUT_4[63587] = 32'b00000000000000000011001000011110;
assign LUT_4[63588] = 32'b00000000000000000111100010011110;
assign LUT_4[63589] = 32'b00000000000000000000101110010110;
assign LUT_4[63590] = 32'b00000000000000000110111101000010;
assign LUT_4[63591] = 32'b00000000000000000000001000111010;
assign LUT_4[63592] = 32'b00000000000000000011101110010111;
assign LUT_4[63593] = 32'b11111111111111111100111010001111;
assign LUT_4[63594] = 32'b00000000000000000011001000111011;
assign LUT_4[63595] = 32'b11111111111111111100010100110011;
assign LUT_4[63596] = 32'b00000000000000000000101110110011;
assign LUT_4[63597] = 32'b11111111111111111001111010101011;
assign LUT_4[63598] = 32'b00000000000000000000001001010111;
assign LUT_4[63599] = 32'b11111111111111111001010101001111;
assign LUT_4[63600] = 32'b00000000000000001000010011110000;
assign LUT_4[63601] = 32'b00000000000000000001011111101000;
assign LUT_4[63602] = 32'b00000000000000000111101110010100;
assign LUT_4[63603] = 32'b00000000000000000000111010001100;
assign LUT_4[63604] = 32'b00000000000000000101010100001100;
assign LUT_4[63605] = 32'b11111111111111111110100000000100;
assign LUT_4[63606] = 32'b00000000000000000100101110110000;
assign LUT_4[63607] = 32'b11111111111111111101111010101000;
assign LUT_4[63608] = 32'b00000000000000000001100000000101;
assign LUT_4[63609] = 32'b11111111111111111010101011111101;
assign LUT_4[63610] = 32'b00000000000000000000111010101001;
assign LUT_4[63611] = 32'b11111111111111111010000110100001;
assign LUT_4[63612] = 32'b11111111111111111110100000100001;
assign LUT_4[63613] = 32'b11111111111111110111101100011001;
assign LUT_4[63614] = 32'b11111111111111111101111011000101;
assign LUT_4[63615] = 32'b11111111111111110111000110111101;
assign LUT_4[63616] = 32'b00000000000000001101010101101111;
assign LUT_4[63617] = 32'b00000000000000000110100001100111;
assign LUT_4[63618] = 32'b00000000000000001100110000010011;
assign LUT_4[63619] = 32'b00000000000000000101111100001011;
assign LUT_4[63620] = 32'b00000000000000001010010110001011;
assign LUT_4[63621] = 32'b00000000000000000011100010000011;
assign LUT_4[63622] = 32'b00000000000000001001110000101111;
assign LUT_4[63623] = 32'b00000000000000000010111100100111;
assign LUT_4[63624] = 32'b00000000000000000110100010000100;
assign LUT_4[63625] = 32'b11111111111111111111101101111100;
assign LUT_4[63626] = 32'b00000000000000000101111100101000;
assign LUT_4[63627] = 32'b11111111111111111111001000100000;
assign LUT_4[63628] = 32'b00000000000000000011100010100000;
assign LUT_4[63629] = 32'b11111111111111111100101110011000;
assign LUT_4[63630] = 32'b00000000000000000010111101000100;
assign LUT_4[63631] = 32'b11111111111111111100001000111100;
assign LUT_4[63632] = 32'b00000000000000001011000111011101;
assign LUT_4[63633] = 32'b00000000000000000100010011010101;
assign LUT_4[63634] = 32'b00000000000000001010100010000001;
assign LUT_4[63635] = 32'b00000000000000000011101101111001;
assign LUT_4[63636] = 32'b00000000000000001000000111111001;
assign LUT_4[63637] = 32'b00000000000000000001010011110001;
assign LUT_4[63638] = 32'b00000000000000000111100010011101;
assign LUT_4[63639] = 32'b00000000000000000000101110010101;
assign LUT_4[63640] = 32'b00000000000000000100010011110010;
assign LUT_4[63641] = 32'b11111111111111111101011111101010;
assign LUT_4[63642] = 32'b00000000000000000011101110010110;
assign LUT_4[63643] = 32'b11111111111111111100111010001110;
assign LUT_4[63644] = 32'b00000000000000000001010100001110;
assign LUT_4[63645] = 32'b11111111111111111010100000000110;
assign LUT_4[63646] = 32'b00000000000000000000101110110010;
assign LUT_4[63647] = 32'b11111111111111111001111010101010;
assign LUT_4[63648] = 32'b00000000000000001011110000110110;
assign LUT_4[63649] = 32'b00000000000000000100111100101110;
assign LUT_4[63650] = 32'b00000000000000001011001011011010;
assign LUT_4[63651] = 32'b00000000000000000100010111010010;
assign LUT_4[63652] = 32'b00000000000000001000110001010010;
assign LUT_4[63653] = 32'b00000000000000000001111101001010;
assign LUT_4[63654] = 32'b00000000000000001000001011110110;
assign LUT_4[63655] = 32'b00000000000000000001010111101110;
assign LUT_4[63656] = 32'b00000000000000000100111101001011;
assign LUT_4[63657] = 32'b11111111111111111110001001000011;
assign LUT_4[63658] = 32'b00000000000000000100010111101111;
assign LUT_4[63659] = 32'b11111111111111111101100011100111;
assign LUT_4[63660] = 32'b00000000000000000001111101100111;
assign LUT_4[63661] = 32'b11111111111111111011001001011111;
assign LUT_4[63662] = 32'b00000000000000000001011000001011;
assign LUT_4[63663] = 32'b11111111111111111010100100000011;
assign LUT_4[63664] = 32'b00000000000000001001100010100100;
assign LUT_4[63665] = 32'b00000000000000000010101110011100;
assign LUT_4[63666] = 32'b00000000000000001000111101001000;
assign LUT_4[63667] = 32'b00000000000000000010001001000000;
assign LUT_4[63668] = 32'b00000000000000000110100011000000;
assign LUT_4[63669] = 32'b11111111111111111111101110111000;
assign LUT_4[63670] = 32'b00000000000000000101111101100100;
assign LUT_4[63671] = 32'b11111111111111111111001001011100;
assign LUT_4[63672] = 32'b00000000000000000010101110111001;
assign LUT_4[63673] = 32'b11111111111111111011111010110001;
assign LUT_4[63674] = 32'b00000000000000000010001001011101;
assign LUT_4[63675] = 32'b11111111111111111011010101010101;
assign LUT_4[63676] = 32'b11111111111111111111101111010101;
assign LUT_4[63677] = 32'b11111111111111111000111011001101;
assign LUT_4[63678] = 32'b11111111111111111111001001111001;
assign LUT_4[63679] = 32'b11111111111111111000010101110001;
assign LUT_4[63680] = 32'b00000000000000001110101101000011;
assign LUT_4[63681] = 32'b00000000000000000111111000111011;
assign LUT_4[63682] = 32'b00000000000000001110000111100111;
assign LUT_4[63683] = 32'b00000000000000000111010011011111;
assign LUT_4[63684] = 32'b00000000000000001011101101011111;
assign LUT_4[63685] = 32'b00000000000000000100111001010111;
assign LUT_4[63686] = 32'b00000000000000001011001000000011;
assign LUT_4[63687] = 32'b00000000000000000100010011111011;
assign LUT_4[63688] = 32'b00000000000000000111111001011000;
assign LUT_4[63689] = 32'b00000000000000000001000101010000;
assign LUT_4[63690] = 32'b00000000000000000111010011111100;
assign LUT_4[63691] = 32'b00000000000000000000011111110100;
assign LUT_4[63692] = 32'b00000000000000000100111001110100;
assign LUT_4[63693] = 32'b11111111111111111110000101101100;
assign LUT_4[63694] = 32'b00000000000000000100010100011000;
assign LUT_4[63695] = 32'b11111111111111111101100000010000;
assign LUT_4[63696] = 32'b00000000000000001100011110110001;
assign LUT_4[63697] = 32'b00000000000000000101101010101001;
assign LUT_4[63698] = 32'b00000000000000001011111001010101;
assign LUT_4[63699] = 32'b00000000000000000101000101001101;
assign LUT_4[63700] = 32'b00000000000000001001011111001101;
assign LUT_4[63701] = 32'b00000000000000000010101011000101;
assign LUT_4[63702] = 32'b00000000000000001000111001110001;
assign LUT_4[63703] = 32'b00000000000000000010000101101001;
assign LUT_4[63704] = 32'b00000000000000000101101011000110;
assign LUT_4[63705] = 32'b11111111111111111110110110111110;
assign LUT_4[63706] = 32'b00000000000000000101000101101010;
assign LUT_4[63707] = 32'b11111111111111111110010001100010;
assign LUT_4[63708] = 32'b00000000000000000010101011100010;
assign LUT_4[63709] = 32'b11111111111111111011110111011010;
assign LUT_4[63710] = 32'b00000000000000000010000110000110;
assign LUT_4[63711] = 32'b11111111111111111011010001111110;
assign LUT_4[63712] = 32'b00000000000000001101001000001010;
assign LUT_4[63713] = 32'b00000000000000000110010100000010;
assign LUT_4[63714] = 32'b00000000000000001100100010101110;
assign LUT_4[63715] = 32'b00000000000000000101101110100110;
assign LUT_4[63716] = 32'b00000000000000001010001000100110;
assign LUT_4[63717] = 32'b00000000000000000011010100011110;
assign LUT_4[63718] = 32'b00000000000000001001100011001010;
assign LUT_4[63719] = 32'b00000000000000000010101111000010;
assign LUT_4[63720] = 32'b00000000000000000110010100011111;
assign LUT_4[63721] = 32'b11111111111111111111100000010111;
assign LUT_4[63722] = 32'b00000000000000000101101111000011;
assign LUT_4[63723] = 32'b11111111111111111110111010111011;
assign LUT_4[63724] = 32'b00000000000000000011010100111011;
assign LUT_4[63725] = 32'b11111111111111111100100000110011;
assign LUT_4[63726] = 32'b00000000000000000010101111011111;
assign LUT_4[63727] = 32'b11111111111111111011111011010111;
assign LUT_4[63728] = 32'b00000000000000001010111001111000;
assign LUT_4[63729] = 32'b00000000000000000100000101110000;
assign LUT_4[63730] = 32'b00000000000000001010010100011100;
assign LUT_4[63731] = 32'b00000000000000000011100000010100;
assign LUT_4[63732] = 32'b00000000000000000111111010010100;
assign LUT_4[63733] = 32'b00000000000000000001000110001100;
assign LUT_4[63734] = 32'b00000000000000000111010100111000;
assign LUT_4[63735] = 32'b00000000000000000000100000110000;
assign LUT_4[63736] = 32'b00000000000000000100000110001101;
assign LUT_4[63737] = 32'b11111111111111111101010010000101;
assign LUT_4[63738] = 32'b00000000000000000011100000110001;
assign LUT_4[63739] = 32'b11111111111111111100101100101001;
assign LUT_4[63740] = 32'b00000000000000000001000110101001;
assign LUT_4[63741] = 32'b11111111111111111010010010100001;
assign LUT_4[63742] = 32'b00000000000000000000100001001101;
assign LUT_4[63743] = 32'b11111111111111111001101101000101;
assign LUT_4[63744] = 32'b00000000000000001111101011001010;
assign LUT_4[63745] = 32'b00000000000000001000110111000010;
assign LUT_4[63746] = 32'b00000000000000001111000101101110;
assign LUT_4[63747] = 32'b00000000000000001000010001100110;
assign LUT_4[63748] = 32'b00000000000000001100101011100110;
assign LUT_4[63749] = 32'b00000000000000000101110111011110;
assign LUT_4[63750] = 32'b00000000000000001100000110001010;
assign LUT_4[63751] = 32'b00000000000000000101010010000010;
assign LUT_4[63752] = 32'b00000000000000001000110111011111;
assign LUT_4[63753] = 32'b00000000000000000010000011010111;
assign LUT_4[63754] = 32'b00000000000000001000010010000011;
assign LUT_4[63755] = 32'b00000000000000000001011101111011;
assign LUT_4[63756] = 32'b00000000000000000101110111111011;
assign LUT_4[63757] = 32'b11111111111111111111000011110011;
assign LUT_4[63758] = 32'b00000000000000000101010010011111;
assign LUT_4[63759] = 32'b11111111111111111110011110010111;
assign LUT_4[63760] = 32'b00000000000000001101011100111000;
assign LUT_4[63761] = 32'b00000000000000000110101000110000;
assign LUT_4[63762] = 32'b00000000000000001100110111011100;
assign LUT_4[63763] = 32'b00000000000000000110000011010100;
assign LUT_4[63764] = 32'b00000000000000001010011101010100;
assign LUT_4[63765] = 32'b00000000000000000011101001001100;
assign LUT_4[63766] = 32'b00000000000000001001110111111000;
assign LUT_4[63767] = 32'b00000000000000000011000011110000;
assign LUT_4[63768] = 32'b00000000000000000110101001001101;
assign LUT_4[63769] = 32'b11111111111111111111110101000101;
assign LUT_4[63770] = 32'b00000000000000000110000011110001;
assign LUT_4[63771] = 32'b11111111111111111111001111101001;
assign LUT_4[63772] = 32'b00000000000000000011101001101001;
assign LUT_4[63773] = 32'b11111111111111111100110101100001;
assign LUT_4[63774] = 32'b00000000000000000011000100001101;
assign LUT_4[63775] = 32'b11111111111111111100010000000101;
assign LUT_4[63776] = 32'b00000000000000001110000110010001;
assign LUT_4[63777] = 32'b00000000000000000111010010001001;
assign LUT_4[63778] = 32'b00000000000000001101100000110101;
assign LUT_4[63779] = 32'b00000000000000000110101100101101;
assign LUT_4[63780] = 32'b00000000000000001011000110101101;
assign LUT_4[63781] = 32'b00000000000000000100010010100101;
assign LUT_4[63782] = 32'b00000000000000001010100001010001;
assign LUT_4[63783] = 32'b00000000000000000011101101001001;
assign LUT_4[63784] = 32'b00000000000000000111010010100110;
assign LUT_4[63785] = 32'b00000000000000000000011110011110;
assign LUT_4[63786] = 32'b00000000000000000110101101001010;
assign LUT_4[63787] = 32'b11111111111111111111111001000010;
assign LUT_4[63788] = 32'b00000000000000000100010011000010;
assign LUT_4[63789] = 32'b11111111111111111101011110111010;
assign LUT_4[63790] = 32'b00000000000000000011101101100110;
assign LUT_4[63791] = 32'b11111111111111111100111001011110;
assign LUT_4[63792] = 32'b00000000000000001011110111111111;
assign LUT_4[63793] = 32'b00000000000000000101000011110111;
assign LUT_4[63794] = 32'b00000000000000001011010010100011;
assign LUT_4[63795] = 32'b00000000000000000100011110011011;
assign LUT_4[63796] = 32'b00000000000000001000111000011011;
assign LUT_4[63797] = 32'b00000000000000000010000100010011;
assign LUT_4[63798] = 32'b00000000000000001000010010111111;
assign LUT_4[63799] = 32'b00000000000000000001011110110111;
assign LUT_4[63800] = 32'b00000000000000000101000100010100;
assign LUT_4[63801] = 32'b11111111111111111110010000001100;
assign LUT_4[63802] = 32'b00000000000000000100011110111000;
assign LUT_4[63803] = 32'b11111111111111111101101010110000;
assign LUT_4[63804] = 32'b00000000000000000010000100110000;
assign LUT_4[63805] = 32'b11111111111111111011010000101000;
assign LUT_4[63806] = 32'b00000000000000000001011111010100;
assign LUT_4[63807] = 32'b11111111111111111010101011001100;
assign LUT_4[63808] = 32'b00000000000000010001000010011110;
assign LUT_4[63809] = 32'b00000000000000001010001110010110;
assign LUT_4[63810] = 32'b00000000000000010000011101000010;
assign LUT_4[63811] = 32'b00000000000000001001101000111010;
assign LUT_4[63812] = 32'b00000000000000001110000010111010;
assign LUT_4[63813] = 32'b00000000000000000111001110110010;
assign LUT_4[63814] = 32'b00000000000000001101011101011110;
assign LUT_4[63815] = 32'b00000000000000000110101001010110;
assign LUT_4[63816] = 32'b00000000000000001010001110110011;
assign LUT_4[63817] = 32'b00000000000000000011011010101011;
assign LUT_4[63818] = 32'b00000000000000001001101001010111;
assign LUT_4[63819] = 32'b00000000000000000010110101001111;
assign LUT_4[63820] = 32'b00000000000000000111001111001111;
assign LUT_4[63821] = 32'b00000000000000000000011011000111;
assign LUT_4[63822] = 32'b00000000000000000110101001110011;
assign LUT_4[63823] = 32'b11111111111111111111110101101011;
assign LUT_4[63824] = 32'b00000000000000001110110100001100;
assign LUT_4[63825] = 32'b00000000000000001000000000000100;
assign LUT_4[63826] = 32'b00000000000000001110001110110000;
assign LUT_4[63827] = 32'b00000000000000000111011010101000;
assign LUT_4[63828] = 32'b00000000000000001011110100101000;
assign LUT_4[63829] = 32'b00000000000000000101000000100000;
assign LUT_4[63830] = 32'b00000000000000001011001111001100;
assign LUT_4[63831] = 32'b00000000000000000100011011000100;
assign LUT_4[63832] = 32'b00000000000000001000000000100001;
assign LUT_4[63833] = 32'b00000000000000000001001100011001;
assign LUT_4[63834] = 32'b00000000000000000111011011000101;
assign LUT_4[63835] = 32'b00000000000000000000100110111101;
assign LUT_4[63836] = 32'b00000000000000000101000000111101;
assign LUT_4[63837] = 32'b11111111111111111110001100110101;
assign LUT_4[63838] = 32'b00000000000000000100011011100001;
assign LUT_4[63839] = 32'b11111111111111111101100111011001;
assign LUT_4[63840] = 32'b00000000000000001111011101100101;
assign LUT_4[63841] = 32'b00000000000000001000101001011101;
assign LUT_4[63842] = 32'b00000000000000001110111000001001;
assign LUT_4[63843] = 32'b00000000000000001000000100000001;
assign LUT_4[63844] = 32'b00000000000000001100011110000001;
assign LUT_4[63845] = 32'b00000000000000000101101001111001;
assign LUT_4[63846] = 32'b00000000000000001011111000100101;
assign LUT_4[63847] = 32'b00000000000000000101000100011101;
assign LUT_4[63848] = 32'b00000000000000001000101001111010;
assign LUT_4[63849] = 32'b00000000000000000001110101110010;
assign LUT_4[63850] = 32'b00000000000000001000000100011110;
assign LUT_4[63851] = 32'b00000000000000000001010000010110;
assign LUT_4[63852] = 32'b00000000000000000101101010010110;
assign LUT_4[63853] = 32'b11111111111111111110110110001110;
assign LUT_4[63854] = 32'b00000000000000000101000100111010;
assign LUT_4[63855] = 32'b11111111111111111110010000110010;
assign LUT_4[63856] = 32'b00000000000000001101001111010011;
assign LUT_4[63857] = 32'b00000000000000000110011011001011;
assign LUT_4[63858] = 32'b00000000000000001100101001110111;
assign LUT_4[63859] = 32'b00000000000000000101110101101111;
assign LUT_4[63860] = 32'b00000000000000001010001111101111;
assign LUT_4[63861] = 32'b00000000000000000011011011100111;
assign LUT_4[63862] = 32'b00000000000000001001101010010011;
assign LUT_4[63863] = 32'b00000000000000000010110110001011;
assign LUT_4[63864] = 32'b00000000000000000110011011101000;
assign LUT_4[63865] = 32'b11111111111111111111100111100000;
assign LUT_4[63866] = 32'b00000000000000000101110110001100;
assign LUT_4[63867] = 32'b11111111111111111111000010000100;
assign LUT_4[63868] = 32'b00000000000000000011011100000100;
assign LUT_4[63869] = 32'b11111111111111111100100111111100;
assign LUT_4[63870] = 32'b00000000000000000010110110101000;
assign LUT_4[63871] = 32'b11111111111111111100000010100000;
assign LUT_4[63872] = 32'b00000000000000010010010001010010;
assign LUT_4[63873] = 32'b00000000000000001011011101001010;
assign LUT_4[63874] = 32'b00000000000000010001101011110110;
assign LUT_4[63875] = 32'b00000000000000001010110111101110;
assign LUT_4[63876] = 32'b00000000000000001111010001101110;
assign LUT_4[63877] = 32'b00000000000000001000011101100110;
assign LUT_4[63878] = 32'b00000000000000001110101100010010;
assign LUT_4[63879] = 32'b00000000000000000111111000001010;
assign LUT_4[63880] = 32'b00000000000000001011011101100111;
assign LUT_4[63881] = 32'b00000000000000000100101001011111;
assign LUT_4[63882] = 32'b00000000000000001010111000001011;
assign LUT_4[63883] = 32'b00000000000000000100000100000011;
assign LUT_4[63884] = 32'b00000000000000001000011110000011;
assign LUT_4[63885] = 32'b00000000000000000001101001111011;
assign LUT_4[63886] = 32'b00000000000000000111111000100111;
assign LUT_4[63887] = 32'b00000000000000000001000100011111;
assign LUT_4[63888] = 32'b00000000000000010000000011000000;
assign LUT_4[63889] = 32'b00000000000000001001001110111000;
assign LUT_4[63890] = 32'b00000000000000001111011101100100;
assign LUT_4[63891] = 32'b00000000000000001000101001011100;
assign LUT_4[63892] = 32'b00000000000000001101000011011100;
assign LUT_4[63893] = 32'b00000000000000000110001111010100;
assign LUT_4[63894] = 32'b00000000000000001100011110000000;
assign LUT_4[63895] = 32'b00000000000000000101101001111000;
assign LUT_4[63896] = 32'b00000000000000001001001111010101;
assign LUT_4[63897] = 32'b00000000000000000010011011001101;
assign LUT_4[63898] = 32'b00000000000000001000101001111001;
assign LUT_4[63899] = 32'b00000000000000000001110101110001;
assign LUT_4[63900] = 32'b00000000000000000110001111110001;
assign LUT_4[63901] = 32'b11111111111111111111011011101001;
assign LUT_4[63902] = 32'b00000000000000000101101010010101;
assign LUT_4[63903] = 32'b11111111111111111110110110001101;
assign LUT_4[63904] = 32'b00000000000000010000101100011001;
assign LUT_4[63905] = 32'b00000000000000001001111000010001;
assign LUT_4[63906] = 32'b00000000000000010000000110111101;
assign LUT_4[63907] = 32'b00000000000000001001010010110101;
assign LUT_4[63908] = 32'b00000000000000001101101100110101;
assign LUT_4[63909] = 32'b00000000000000000110111000101101;
assign LUT_4[63910] = 32'b00000000000000001101000111011001;
assign LUT_4[63911] = 32'b00000000000000000110010011010001;
assign LUT_4[63912] = 32'b00000000000000001001111000101110;
assign LUT_4[63913] = 32'b00000000000000000011000100100110;
assign LUT_4[63914] = 32'b00000000000000001001010011010010;
assign LUT_4[63915] = 32'b00000000000000000010011111001010;
assign LUT_4[63916] = 32'b00000000000000000110111001001010;
assign LUT_4[63917] = 32'b00000000000000000000000101000010;
assign LUT_4[63918] = 32'b00000000000000000110010011101110;
assign LUT_4[63919] = 32'b11111111111111111111011111100110;
assign LUT_4[63920] = 32'b00000000000000001110011110000111;
assign LUT_4[63921] = 32'b00000000000000000111101001111111;
assign LUT_4[63922] = 32'b00000000000000001101111000101011;
assign LUT_4[63923] = 32'b00000000000000000111000100100011;
assign LUT_4[63924] = 32'b00000000000000001011011110100011;
assign LUT_4[63925] = 32'b00000000000000000100101010011011;
assign LUT_4[63926] = 32'b00000000000000001010111001000111;
assign LUT_4[63927] = 32'b00000000000000000100000100111111;
assign LUT_4[63928] = 32'b00000000000000000111101010011100;
assign LUT_4[63929] = 32'b00000000000000000000110110010100;
assign LUT_4[63930] = 32'b00000000000000000111000101000000;
assign LUT_4[63931] = 32'b00000000000000000000010000111000;
assign LUT_4[63932] = 32'b00000000000000000100101010111000;
assign LUT_4[63933] = 32'b11111111111111111101110110110000;
assign LUT_4[63934] = 32'b00000000000000000100000101011100;
assign LUT_4[63935] = 32'b11111111111111111101010001010100;
assign LUT_4[63936] = 32'b00000000000000010011101000100110;
assign LUT_4[63937] = 32'b00000000000000001100110100011110;
assign LUT_4[63938] = 32'b00000000000000010011000011001010;
assign LUT_4[63939] = 32'b00000000000000001100001111000010;
assign LUT_4[63940] = 32'b00000000000000010000101001000010;
assign LUT_4[63941] = 32'b00000000000000001001110100111010;
assign LUT_4[63942] = 32'b00000000000000010000000011100110;
assign LUT_4[63943] = 32'b00000000000000001001001111011110;
assign LUT_4[63944] = 32'b00000000000000001100110100111011;
assign LUT_4[63945] = 32'b00000000000000000110000000110011;
assign LUT_4[63946] = 32'b00000000000000001100001111011111;
assign LUT_4[63947] = 32'b00000000000000000101011011010111;
assign LUT_4[63948] = 32'b00000000000000001001110101010111;
assign LUT_4[63949] = 32'b00000000000000000011000001001111;
assign LUT_4[63950] = 32'b00000000000000001001001111111011;
assign LUT_4[63951] = 32'b00000000000000000010011011110011;
assign LUT_4[63952] = 32'b00000000000000010001011010010100;
assign LUT_4[63953] = 32'b00000000000000001010100110001100;
assign LUT_4[63954] = 32'b00000000000000010000110100111000;
assign LUT_4[63955] = 32'b00000000000000001010000000110000;
assign LUT_4[63956] = 32'b00000000000000001110011010110000;
assign LUT_4[63957] = 32'b00000000000000000111100110101000;
assign LUT_4[63958] = 32'b00000000000000001101110101010100;
assign LUT_4[63959] = 32'b00000000000000000111000001001100;
assign LUT_4[63960] = 32'b00000000000000001010100110101001;
assign LUT_4[63961] = 32'b00000000000000000011110010100001;
assign LUT_4[63962] = 32'b00000000000000001010000001001101;
assign LUT_4[63963] = 32'b00000000000000000011001101000101;
assign LUT_4[63964] = 32'b00000000000000000111100111000101;
assign LUT_4[63965] = 32'b00000000000000000000110010111101;
assign LUT_4[63966] = 32'b00000000000000000111000001101001;
assign LUT_4[63967] = 32'b00000000000000000000001101100001;
assign LUT_4[63968] = 32'b00000000000000010010000011101101;
assign LUT_4[63969] = 32'b00000000000000001011001111100101;
assign LUT_4[63970] = 32'b00000000000000010001011110010001;
assign LUT_4[63971] = 32'b00000000000000001010101010001001;
assign LUT_4[63972] = 32'b00000000000000001111000100001001;
assign LUT_4[63973] = 32'b00000000000000001000010000000001;
assign LUT_4[63974] = 32'b00000000000000001110011110101101;
assign LUT_4[63975] = 32'b00000000000000000111101010100101;
assign LUT_4[63976] = 32'b00000000000000001011010000000010;
assign LUT_4[63977] = 32'b00000000000000000100011011111010;
assign LUT_4[63978] = 32'b00000000000000001010101010100110;
assign LUT_4[63979] = 32'b00000000000000000011110110011110;
assign LUT_4[63980] = 32'b00000000000000001000010000011110;
assign LUT_4[63981] = 32'b00000000000000000001011100010110;
assign LUT_4[63982] = 32'b00000000000000000111101011000010;
assign LUT_4[63983] = 32'b00000000000000000000110110111010;
assign LUT_4[63984] = 32'b00000000000000001111110101011011;
assign LUT_4[63985] = 32'b00000000000000001001000001010011;
assign LUT_4[63986] = 32'b00000000000000001111001111111111;
assign LUT_4[63987] = 32'b00000000000000001000011011110111;
assign LUT_4[63988] = 32'b00000000000000001100110101110111;
assign LUT_4[63989] = 32'b00000000000000000110000001101111;
assign LUT_4[63990] = 32'b00000000000000001100010000011011;
assign LUT_4[63991] = 32'b00000000000000000101011100010011;
assign LUT_4[63992] = 32'b00000000000000001001000001110000;
assign LUT_4[63993] = 32'b00000000000000000010001101101000;
assign LUT_4[63994] = 32'b00000000000000001000011100010100;
assign LUT_4[63995] = 32'b00000000000000000001101000001100;
assign LUT_4[63996] = 32'b00000000000000000110000010001100;
assign LUT_4[63997] = 32'b11111111111111111111001110000100;
assign LUT_4[63998] = 32'b00000000000000000101011100110000;
assign LUT_4[63999] = 32'b11111111111111111110101000101000;
assign LUT_4[64000] = 32'b00000000000000001001110011101111;
assign LUT_4[64001] = 32'b00000000000000000010111111100111;
assign LUT_4[64002] = 32'b00000000000000001001001110010011;
assign LUT_4[64003] = 32'b00000000000000000010011010001011;
assign LUT_4[64004] = 32'b00000000000000000110110100001011;
assign LUT_4[64005] = 32'b00000000000000000000000000000011;
assign LUT_4[64006] = 32'b00000000000000000110001110101111;
assign LUT_4[64007] = 32'b11111111111111111111011010100111;
assign LUT_4[64008] = 32'b00000000000000000011000000000100;
assign LUT_4[64009] = 32'b11111111111111111100001011111100;
assign LUT_4[64010] = 32'b00000000000000000010011010101000;
assign LUT_4[64011] = 32'b11111111111111111011100110100000;
assign LUT_4[64012] = 32'b00000000000000000000000000100000;
assign LUT_4[64013] = 32'b11111111111111111001001100011000;
assign LUT_4[64014] = 32'b11111111111111111111011011000100;
assign LUT_4[64015] = 32'b11111111111111111000100110111100;
assign LUT_4[64016] = 32'b00000000000000000111100101011101;
assign LUT_4[64017] = 32'b00000000000000000000110001010101;
assign LUT_4[64018] = 32'b00000000000000000111000000000001;
assign LUT_4[64019] = 32'b00000000000000000000001011111001;
assign LUT_4[64020] = 32'b00000000000000000100100101111001;
assign LUT_4[64021] = 32'b11111111111111111101110001110001;
assign LUT_4[64022] = 32'b00000000000000000100000000011101;
assign LUT_4[64023] = 32'b11111111111111111101001100010101;
assign LUT_4[64024] = 32'b00000000000000000000110001110010;
assign LUT_4[64025] = 32'b11111111111111111001111101101010;
assign LUT_4[64026] = 32'b00000000000000000000001100010110;
assign LUT_4[64027] = 32'b11111111111111111001011000001110;
assign LUT_4[64028] = 32'b11111111111111111101110010001110;
assign LUT_4[64029] = 32'b11111111111111110110111110000110;
assign LUT_4[64030] = 32'b11111111111111111101001100110010;
assign LUT_4[64031] = 32'b11111111111111110110011000101010;
assign LUT_4[64032] = 32'b00000000000000001000001110110110;
assign LUT_4[64033] = 32'b00000000000000000001011010101110;
assign LUT_4[64034] = 32'b00000000000000000111101001011010;
assign LUT_4[64035] = 32'b00000000000000000000110101010010;
assign LUT_4[64036] = 32'b00000000000000000101001111010010;
assign LUT_4[64037] = 32'b11111111111111111110011011001010;
assign LUT_4[64038] = 32'b00000000000000000100101001110110;
assign LUT_4[64039] = 32'b11111111111111111101110101101110;
assign LUT_4[64040] = 32'b00000000000000000001011011001011;
assign LUT_4[64041] = 32'b11111111111111111010100111000011;
assign LUT_4[64042] = 32'b00000000000000000000110101101111;
assign LUT_4[64043] = 32'b11111111111111111010000001100111;
assign LUT_4[64044] = 32'b11111111111111111110011011100111;
assign LUT_4[64045] = 32'b11111111111111110111100111011111;
assign LUT_4[64046] = 32'b11111111111111111101110110001011;
assign LUT_4[64047] = 32'b11111111111111110111000010000011;
assign LUT_4[64048] = 32'b00000000000000000110000000100100;
assign LUT_4[64049] = 32'b11111111111111111111001100011100;
assign LUT_4[64050] = 32'b00000000000000000101011011001000;
assign LUT_4[64051] = 32'b11111111111111111110100111000000;
assign LUT_4[64052] = 32'b00000000000000000011000001000000;
assign LUT_4[64053] = 32'b11111111111111111100001100111000;
assign LUT_4[64054] = 32'b00000000000000000010011011100100;
assign LUT_4[64055] = 32'b11111111111111111011100111011100;
assign LUT_4[64056] = 32'b11111111111111111111001100111001;
assign LUT_4[64057] = 32'b11111111111111111000011000110001;
assign LUT_4[64058] = 32'b11111111111111111110100111011101;
assign LUT_4[64059] = 32'b11111111111111110111110011010101;
assign LUT_4[64060] = 32'b11111111111111111100001101010101;
assign LUT_4[64061] = 32'b11111111111111110101011001001101;
assign LUT_4[64062] = 32'b11111111111111111011100111111001;
assign LUT_4[64063] = 32'b11111111111111110100110011110001;
assign LUT_4[64064] = 32'b00000000000000001011001011000011;
assign LUT_4[64065] = 32'b00000000000000000100010110111011;
assign LUT_4[64066] = 32'b00000000000000001010100101100111;
assign LUT_4[64067] = 32'b00000000000000000011110001011111;
assign LUT_4[64068] = 32'b00000000000000001000001011011111;
assign LUT_4[64069] = 32'b00000000000000000001010111010111;
assign LUT_4[64070] = 32'b00000000000000000111100110000011;
assign LUT_4[64071] = 32'b00000000000000000000110001111011;
assign LUT_4[64072] = 32'b00000000000000000100010111011000;
assign LUT_4[64073] = 32'b11111111111111111101100011010000;
assign LUT_4[64074] = 32'b00000000000000000011110001111100;
assign LUT_4[64075] = 32'b11111111111111111100111101110100;
assign LUT_4[64076] = 32'b00000000000000000001010111110100;
assign LUT_4[64077] = 32'b11111111111111111010100011101100;
assign LUT_4[64078] = 32'b00000000000000000000110010011000;
assign LUT_4[64079] = 32'b11111111111111111001111110010000;
assign LUT_4[64080] = 32'b00000000000000001000111100110001;
assign LUT_4[64081] = 32'b00000000000000000010001000101001;
assign LUT_4[64082] = 32'b00000000000000001000010111010101;
assign LUT_4[64083] = 32'b00000000000000000001100011001101;
assign LUT_4[64084] = 32'b00000000000000000101111101001101;
assign LUT_4[64085] = 32'b11111111111111111111001001000101;
assign LUT_4[64086] = 32'b00000000000000000101010111110001;
assign LUT_4[64087] = 32'b11111111111111111110100011101001;
assign LUT_4[64088] = 32'b00000000000000000010001001000110;
assign LUT_4[64089] = 32'b11111111111111111011010100111110;
assign LUT_4[64090] = 32'b00000000000000000001100011101010;
assign LUT_4[64091] = 32'b11111111111111111010101111100010;
assign LUT_4[64092] = 32'b11111111111111111111001001100010;
assign LUT_4[64093] = 32'b11111111111111111000010101011010;
assign LUT_4[64094] = 32'b11111111111111111110100100000110;
assign LUT_4[64095] = 32'b11111111111111110111101111111110;
assign LUT_4[64096] = 32'b00000000000000001001100110001010;
assign LUT_4[64097] = 32'b00000000000000000010110010000010;
assign LUT_4[64098] = 32'b00000000000000001001000000101110;
assign LUT_4[64099] = 32'b00000000000000000010001100100110;
assign LUT_4[64100] = 32'b00000000000000000110100110100110;
assign LUT_4[64101] = 32'b11111111111111111111110010011110;
assign LUT_4[64102] = 32'b00000000000000000110000001001010;
assign LUT_4[64103] = 32'b11111111111111111111001101000010;
assign LUT_4[64104] = 32'b00000000000000000010110010011111;
assign LUT_4[64105] = 32'b11111111111111111011111110010111;
assign LUT_4[64106] = 32'b00000000000000000010001101000011;
assign LUT_4[64107] = 32'b11111111111111111011011000111011;
assign LUT_4[64108] = 32'b11111111111111111111110010111011;
assign LUT_4[64109] = 32'b11111111111111111000111110110011;
assign LUT_4[64110] = 32'b11111111111111111111001101011111;
assign LUT_4[64111] = 32'b11111111111111111000011001010111;
assign LUT_4[64112] = 32'b00000000000000000111010111111000;
assign LUT_4[64113] = 32'b00000000000000000000100011110000;
assign LUT_4[64114] = 32'b00000000000000000110110010011100;
assign LUT_4[64115] = 32'b11111111111111111111111110010100;
assign LUT_4[64116] = 32'b00000000000000000100011000010100;
assign LUT_4[64117] = 32'b11111111111111111101100100001100;
assign LUT_4[64118] = 32'b00000000000000000011110010111000;
assign LUT_4[64119] = 32'b11111111111111111100111110110000;
assign LUT_4[64120] = 32'b00000000000000000000100100001101;
assign LUT_4[64121] = 32'b11111111111111111001110000000101;
assign LUT_4[64122] = 32'b11111111111111111111111110110001;
assign LUT_4[64123] = 32'b11111111111111111001001010101001;
assign LUT_4[64124] = 32'b11111111111111111101100100101001;
assign LUT_4[64125] = 32'b11111111111111110110110000100001;
assign LUT_4[64126] = 32'b11111111111111111100111111001101;
assign LUT_4[64127] = 32'b11111111111111110110001011000101;
assign LUT_4[64128] = 32'b00000000000000001100011001110111;
assign LUT_4[64129] = 32'b00000000000000000101100101101111;
assign LUT_4[64130] = 32'b00000000000000001011110100011011;
assign LUT_4[64131] = 32'b00000000000000000101000000010011;
assign LUT_4[64132] = 32'b00000000000000001001011010010011;
assign LUT_4[64133] = 32'b00000000000000000010100110001011;
assign LUT_4[64134] = 32'b00000000000000001000110100110111;
assign LUT_4[64135] = 32'b00000000000000000010000000101111;
assign LUT_4[64136] = 32'b00000000000000000101100110001100;
assign LUT_4[64137] = 32'b11111111111111111110110010000100;
assign LUT_4[64138] = 32'b00000000000000000101000000110000;
assign LUT_4[64139] = 32'b11111111111111111110001100101000;
assign LUT_4[64140] = 32'b00000000000000000010100110101000;
assign LUT_4[64141] = 32'b11111111111111111011110010100000;
assign LUT_4[64142] = 32'b00000000000000000010000001001100;
assign LUT_4[64143] = 32'b11111111111111111011001101000100;
assign LUT_4[64144] = 32'b00000000000000001010001011100101;
assign LUT_4[64145] = 32'b00000000000000000011010111011101;
assign LUT_4[64146] = 32'b00000000000000001001100110001001;
assign LUT_4[64147] = 32'b00000000000000000010110010000001;
assign LUT_4[64148] = 32'b00000000000000000111001100000001;
assign LUT_4[64149] = 32'b00000000000000000000010111111001;
assign LUT_4[64150] = 32'b00000000000000000110100110100101;
assign LUT_4[64151] = 32'b11111111111111111111110010011101;
assign LUT_4[64152] = 32'b00000000000000000011010111111010;
assign LUT_4[64153] = 32'b11111111111111111100100011110010;
assign LUT_4[64154] = 32'b00000000000000000010110010011110;
assign LUT_4[64155] = 32'b11111111111111111011111110010110;
assign LUT_4[64156] = 32'b00000000000000000000011000010110;
assign LUT_4[64157] = 32'b11111111111111111001100100001110;
assign LUT_4[64158] = 32'b11111111111111111111110010111010;
assign LUT_4[64159] = 32'b11111111111111111000111110110010;
assign LUT_4[64160] = 32'b00000000000000001010110100111110;
assign LUT_4[64161] = 32'b00000000000000000100000000110110;
assign LUT_4[64162] = 32'b00000000000000001010001111100010;
assign LUT_4[64163] = 32'b00000000000000000011011011011010;
assign LUT_4[64164] = 32'b00000000000000000111110101011010;
assign LUT_4[64165] = 32'b00000000000000000001000001010010;
assign LUT_4[64166] = 32'b00000000000000000111001111111110;
assign LUT_4[64167] = 32'b00000000000000000000011011110110;
assign LUT_4[64168] = 32'b00000000000000000100000001010011;
assign LUT_4[64169] = 32'b11111111111111111101001101001011;
assign LUT_4[64170] = 32'b00000000000000000011011011110111;
assign LUT_4[64171] = 32'b11111111111111111100100111101111;
assign LUT_4[64172] = 32'b00000000000000000001000001101111;
assign LUT_4[64173] = 32'b11111111111111111010001101100111;
assign LUT_4[64174] = 32'b00000000000000000000011100010011;
assign LUT_4[64175] = 32'b11111111111111111001101000001011;
assign LUT_4[64176] = 32'b00000000000000001000100110101100;
assign LUT_4[64177] = 32'b00000000000000000001110010100100;
assign LUT_4[64178] = 32'b00000000000000001000000001010000;
assign LUT_4[64179] = 32'b00000000000000000001001101001000;
assign LUT_4[64180] = 32'b00000000000000000101100111001000;
assign LUT_4[64181] = 32'b11111111111111111110110011000000;
assign LUT_4[64182] = 32'b00000000000000000101000001101100;
assign LUT_4[64183] = 32'b11111111111111111110001101100100;
assign LUT_4[64184] = 32'b00000000000000000001110011000001;
assign LUT_4[64185] = 32'b11111111111111111010111110111001;
assign LUT_4[64186] = 32'b00000000000000000001001101100101;
assign LUT_4[64187] = 32'b11111111111111111010011001011101;
assign LUT_4[64188] = 32'b11111111111111111110110011011101;
assign LUT_4[64189] = 32'b11111111111111110111111111010101;
assign LUT_4[64190] = 32'b11111111111111111110001110000001;
assign LUT_4[64191] = 32'b11111111111111110111011001111001;
assign LUT_4[64192] = 32'b00000000000000001101110001001011;
assign LUT_4[64193] = 32'b00000000000000000110111101000011;
assign LUT_4[64194] = 32'b00000000000000001101001011101111;
assign LUT_4[64195] = 32'b00000000000000000110010111100111;
assign LUT_4[64196] = 32'b00000000000000001010110001100111;
assign LUT_4[64197] = 32'b00000000000000000011111101011111;
assign LUT_4[64198] = 32'b00000000000000001010001100001011;
assign LUT_4[64199] = 32'b00000000000000000011011000000011;
assign LUT_4[64200] = 32'b00000000000000000110111101100000;
assign LUT_4[64201] = 32'b00000000000000000000001001011000;
assign LUT_4[64202] = 32'b00000000000000000110011000000100;
assign LUT_4[64203] = 32'b11111111111111111111100011111100;
assign LUT_4[64204] = 32'b00000000000000000011111101111100;
assign LUT_4[64205] = 32'b11111111111111111101001001110100;
assign LUT_4[64206] = 32'b00000000000000000011011000100000;
assign LUT_4[64207] = 32'b11111111111111111100100100011000;
assign LUT_4[64208] = 32'b00000000000000001011100010111001;
assign LUT_4[64209] = 32'b00000000000000000100101110110001;
assign LUT_4[64210] = 32'b00000000000000001010111101011101;
assign LUT_4[64211] = 32'b00000000000000000100001001010101;
assign LUT_4[64212] = 32'b00000000000000001000100011010101;
assign LUT_4[64213] = 32'b00000000000000000001101111001101;
assign LUT_4[64214] = 32'b00000000000000000111111101111001;
assign LUT_4[64215] = 32'b00000000000000000001001001110001;
assign LUT_4[64216] = 32'b00000000000000000100101111001110;
assign LUT_4[64217] = 32'b11111111111111111101111011000110;
assign LUT_4[64218] = 32'b00000000000000000100001001110010;
assign LUT_4[64219] = 32'b11111111111111111101010101101010;
assign LUT_4[64220] = 32'b00000000000000000001101111101010;
assign LUT_4[64221] = 32'b11111111111111111010111011100010;
assign LUT_4[64222] = 32'b00000000000000000001001010001110;
assign LUT_4[64223] = 32'b11111111111111111010010110000110;
assign LUT_4[64224] = 32'b00000000000000001100001100010010;
assign LUT_4[64225] = 32'b00000000000000000101011000001010;
assign LUT_4[64226] = 32'b00000000000000001011100110110110;
assign LUT_4[64227] = 32'b00000000000000000100110010101110;
assign LUT_4[64228] = 32'b00000000000000001001001100101110;
assign LUT_4[64229] = 32'b00000000000000000010011000100110;
assign LUT_4[64230] = 32'b00000000000000001000100111010010;
assign LUT_4[64231] = 32'b00000000000000000001110011001010;
assign LUT_4[64232] = 32'b00000000000000000101011000100111;
assign LUT_4[64233] = 32'b11111111111111111110100100011111;
assign LUT_4[64234] = 32'b00000000000000000100110011001011;
assign LUT_4[64235] = 32'b11111111111111111101111111000011;
assign LUT_4[64236] = 32'b00000000000000000010011001000011;
assign LUT_4[64237] = 32'b11111111111111111011100100111011;
assign LUT_4[64238] = 32'b00000000000000000001110011100111;
assign LUT_4[64239] = 32'b11111111111111111010111111011111;
assign LUT_4[64240] = 32'b00000000000000001001111110000000;
assign LUT_4[64241] = 32'b00000000000000000011001001111000;
assign LUT_4[64242] = 32'b00000000000000001001011000100100;
assign LUT_4[64243] = 32'b00000000000000000010100100011100;
assign LUT_4[64244] = 32'b00000000000000000110111110011100;
assign LUT_4[64245] = 32'b00000000000000000000001010010100;
assign LUT_4[64246] = 32'b00000000000000000110011001000000;
assign LUT_4[64247] = 32'b11111111111111111111100100111000;
assign LUT_4[64248] = 32'b00000000000000000011001010010101;
assign LUT_4[64249] = 32'b11111111111111111100010110001101;
assign LUT_4[64250] = 32'b00000000000000000010100100111001;
assign LUT_4[64251] = 32'b11111111111111111011110000110001;
assign LUT_4[64252] = 32'b00000000000000000000001010110001;
assign LUT_4[64253] = 32'b11111111111111111001010110101001;
assign LUT_4[64254] = 32'b11111111111111111111100101010101;
assign LUT_4[64255] = 32'b11111111111111111000110001001101;
assign LUT_4[64256] = 32'b00000000000000001110101111010010;
assign LUT_4[64257] = 32'b00000000000000000111111011001010;
assign LUT_4[64258] = 32'b00000000000000001110001001110110;
assign LUT_4[64259] = 32'b00000000000000000111010101101110;
assign LUT_4[64260] = 32'b00000000000000001011101111101110;
assign LUT_4[64261] = 32'b00000000000000000100111011100110;
assign LUT_4[64262] = 32'b00000000000000001011001010010010;
assign LUT_4[64263] = 32'b00000000000000000100010110001010;
assign LUT_4[64264] = 32'b00000000000000000111111011100111;
assign LUT_4[64265] = 32'b00000000000000000001000111011111;
assign LUT_4[64266] = 32'b00000000000000000111010110001011;
assign LUT_4[64267] = 32'b00000000000000000000100010000011;
assign LUT_4[64268] = 32'b00000000000000000100111100000011;
assign LUT_4[64269] = 32'b11111111111111111110000111111011;
assign LUT_4[64270] = 32'b00000000000000000100010110100111;
assign LUT_4[64271] = 32'b11111111111111111101100010011111;
assign LUT_4[64272] = 32'b00000000000000001100100001000000;
assign LUT_4[64273] = 32'b00000000000000000101101100111000;
assign LUT_4[64274] = 32'b00000000000000001011111011100100;
assign LUT_4[64275] = 32'b00000000000000000101000111011100;
assign LUT_4[64276] = 32'b00000000000000001001100001011100;
assign LUT_4[64277] = 32'b00000000000000000010101101010100;
assign LUT_4[64278] = 32'b00000000000000001000111100000000;
assign LUT_4[64279] = 32'b00000000000000000010000111111000;
assign LUT_4[64280] = 32'b00000000000000000101101101010101;
assign LUT_4[64281] = 32'b11111111111111111110111001001101;
assign LUT_4[64282] = 32'b00000000000000000101000111111001;
assign LUT_4[64283] = 32'b11111111111111111110010011110001;
assign LUT_4[64284] = 32'b00000000000000000010101101110001;
assign LUT_4[64285] = 32'b11111111111111111011111001101001;
assign LUT_4[64286] = 32'b00000000000000000010001000010101;
assign LUT_4[64287] = 32'b11111111111111111011010100001101;
assign LUT_4[64288] = 32'b00000000000000001101001010011001;
assign LUT_4[64289] = 32'b00000000000000000110010110010001;
assign LUT_4[64290] = 32'b00000000000000001100100100111101;
assign LUT_4[64291] = 32'b00000000000000000101110000110101;
assign LUT_4[64292] = 32'b00000000000000001010001010110101;
assign LUT_4[64293] = 32'b00000000000000000011010110101101;
assign LUT_4[64294] = 32'b00000000000000001001100101011001;
assign LUT_4[64295] = 32'b00000000000000000010110001010001;
assign LUT_4[64296] = 32'b00000000000000000110010110101110;
assign LUT_4[64297] = 32'b11111111111111111111100010100110;
assign LUT_4[64298] = 32'b00000000000000000101110001010010;
assign LUT_4[64299] = 32'b11111111111111111110111101001010;
assign LUT_4[64300] = 32'b00000000000000000011010111001010;
assign LUT_4[64301] = 32'b11111111111111111100100011000010;
assign LUT_4[64302] = 32'b00000000000000000010110001101110;
assign LUT_4[64303] = 32'b11111111111111111011111101100110;
assign LUT_4[64304] = 32'b00000000000000001010111100000111;
assign LUT_4[64305] = 32'b00000000000000000100000111111111;
assign LUT_4[64306] = 32'b00000000000000001010010110101011;
assign LUT_4[64307] = 32'b00000000000000000011100010100011;
assign LUT_4[64308] = 32'b00000000000000000111111100100011;
assign LUT_4[64309] = 32'b00000000000000000001001000011011;
assign LUT_4[64310] = 32'b00000000000000000111010111000111;
assign LUT_4[64311] = 32'b00000000000000000000100010111111;
assign LUT_4[64312] = 32'b00000000000000000100001000011100;
assign LUT_4[64313] = 32'b11111111111111111101010100010100;
assign LUT_4[64314] = 32'b00000000000000000011100011000000;
assign LUT_4[64315] = 32'b11111111111111111100101110111000;
assign LUT_4[64316] = 32'b00000000000000000001001000111000;
assign LUT_4[64317] = 32'b11111111111111111010010100110000;
assign LUT_4[64318] = 32'b00000000000000000000100011011100;
assign LUT_4[64319] = 32'b11111111111111111001101111010100;
assign LUT_4[64320] = 32'b00000000000000010000000110100110;
assign LUT_4[64321] = 32'b00000000000000001001010010011110;
assign LUT_4[64322] = 32'b00000000000000001111100001001010;
assign LUT_4[64323] = 32'b00000000000000001000101101000010;
assign LUT_4[64324] = 32'b00000000000000001101000111000010;
assign LUT_4[64325] = 32'b00000000000000000110010010111010;
assign LUT_4[64326] = 32'b00000000000000001100100001100110;
assign LUT_4[64327] = 32'b00000000000000000101101101011110;
assign LUT_4[64328] = 32'b00000000000000001001010010111011;
assign LUT_4[64329] = 32'b00000000000000000010011110110011;
assign LUT_4[64330] = 32'b00000000000000001000101101011111;
assign LUT_4[64331] = 32'b00000000000000000001111001010111;
assign LUT_4[64332] = 32'b00000000000000000110010011010111;
assign LUT_4[64333] = 32'b11111111111111111111011111001111;
assign LUT_4[64334] = 32'b00000000000000000101101101111011;
assign LUT_4[64335] = 32'b11111111111111111110111001110011;
assign LUT_4[64336] = 32'b00000000000000001101111000010100;
assign LUT_4[64337] = 32'b00000000000000000111000100001100;
assign LUT_4[64338] = 32'b00000000000000001101010010111000;
assign LUT_4[64339] = 32'b00000000000000000110011110110000;
assign LUT_4[64340] = 32'b00000000000000001010111000110000;
assign LUT_4[64341] = 32'b00000000000000000100000100101000;
assign LUT_4[64342] = 32'b00000000000000001010010011010100;
assign LUT_4[64343] = 32'b00000000000000000011011111001100;
assign LUT_4[64344] = 32'b00000000000000000111000100101001;
assign LUT_4[64345] = 32'b00000000000000000000010000100001;
assign LUT_4[64346] = 32'b00000000000000000110011111001101;
assign LUT_4[64347] = 32'b11111111111111111111101011000101;
assign LUT_4[64348] = 32'b00000000000000000100000101000101;
assign LUT_4[64349] = 32'b11111111111111111101010000111101;
assign LUT_4[64350] = 32'b00000000000000000011011111101001;
assign LUT_4[64351] = 32'b11111111111111111100101011100001;
assign LUT_4[64352] = 32'b00000000000000001110100001101101;
assign LUT_4[64353] = 32'b00000000000000000111101101100101;
assign LUT_4[64354] = 32'b00000000000000001101111100010001;
assign LUT_4[64355] = 32'b00000000000000000111001000001001;
assign LUT_4[64356] = 32'b00000000000000001011100010001001;
assign LUT_4[64357] = 32'b00000000000000000100101110000001;
assign LUT_4[64358] = 32'b00000000000000001010111100101101;
assign LUT_4[64359] = 32'b00000000000000000100001000100101;
assign LUT_4[64360] = 32'b00000000000000000111101110000010;
assign LUT_4[64361] = 32'b00000000000000000000111001111010;
assign LUT_4[64362] = 32'b00000000000000000111001000100110;
assign LUT_4[64363] = 32'b00000000000000000000010100011110;
assign LUT_4[64364] = 32'b00000000000000000100101110011110;
assign LUT_4[64365] = 32'b11111111111111111101111010010110;
assign LUT_4[64366] = 32'b00000000000000000100001001000010;
assign LUT_4[64367] = 32'b11111111111111111101010100111010;
assign LUT_4[64368] = 32'b00000000000000001100010011011011;
assign LUT_4[64369] = 32'b00000000000000000101011111010011;
assign LUT_4[64370] = 32'b00000000000000001011101101111111;
assign LUT_4[64371] = 32'b00000000000000000100111001110111;
assign LUT_4[64372] = 32'b00000000000000001001010011110111;
assign LUT_4[64373] = 32'b00000000000000000010011111101111;
assign LUT_4[64374] = 32'b00000000000000001000101110011011;
assign LUT_4[64375] = 32'b00000000000000000001111010010011;
assign LUT_4[64376] = 32'b00000000000000000101011111110000;
assign LUT_4[64377] = 32'b11111111111111111110101011101000;
assign LUT_4[64378] = 32'b00000000000000000100111010010100;
assign LUT_4[64379] = 32'b11111111111111111110000110001100;
assign LUT_4[64380] = 32'b00000000000000000010100000001100;
assign LUT_4[64381] = 32'b11111111111111111011101100000100;
assign LUT_4[64382] = 32'b00000000000000000001111010110000;
assign LUT_4[64383] = 32'b11111111111111111011000110101000;
assign LUT_4[64384] = 32'b00000000000000010001010101011010;
assign LUT_4[64385] = 32'b00000000000000001010100001010010;
assign LUT_4[64386] = 32'b00000000000000010000101111111110;
assign LUT_4[64387] = 32'b00000000000000001001111011110110;
assign LUT_4[64388] = 32'b00000000000000001110010101110110;
assign LUT_4[64389] = 32'b00000000000000000111100001101110;
assign LUT_4[64390] = 32'b00000000000000001101110000011010;
assign LUT_4[64391] = 32'b00000000000000000110111100010010;
assign LUT_4[64392] = 32'b00000000000000001010100001101111;
assign LUT_4[64393] = 32'b00000000000000000011101101100111;
assign LUT_4[64394] = 32'b00000000000000001001111100010011;
assign LUT_4[64395] = 32'b00000000000000000011001000001011;
assign LUT_4[64396] = 32'b00000000000000000111100010001011;
assign LUT_4[64397] = 32'b00000000000000000000101110000011;
assign LUT_4[64398] = 32'b00000000000000000110111100101111;
assign LUT_4[64399] = 32'b00000000000000000000001000100111;
assign LUT_4[64400] = 32'b00000000000000001111000111001000;
assign LUT_4[64401] = 32'b00000000000000001000010011000000;
assign LUT_4[64402] = 32'b00000000000000001110100001101100;
assign LUT_4[64403] = 32'b00000000000000000111101101100100;
assign LUT_4[64404] = 32'b00000000000000001100000111100100;
assign LUT_4[64405] = 32'b00000000000000000101010011011100;
assign LUT_4[64406] = 32'b00000000000000001011100010001000;
assign LUT_4[64407] = 32'b00000000000000000100101110000000;
assign LUT_4[64408] = 32'b00000000000000001000010011011101;
assign LUT_4[64409] = 32'b00000000000000000001011111010101;
assign LUT_4[64410] = 32'b00000000000000000111101110000001;
assign LUT_4[64411] = 32'b00000000000000000000111001111001;
assign LUT_4[64412] = 32'b00000000000000000101010011111001;
assign LUT_4[64413] = 32'b11111111111111111110011111110001;
assign LUT_4[64414] = 32'b00000000000000000100101110011101;
assign LUT_4[64415] = 32'b11111111111111111101111010010101;
assign LUT_4[64416] = 32'b00000000000000001111110000100001;
assign LUT_4[64417] = 32'b00000000000000001000111100011001;
assign LUT_4[64418] = 32'b00000000000000001111001011000101;
assign LUT_4[64419] = 32'b00000000000000001000010110111101;
assign LUT_4[64420] = 32'b00000000000000001100110000111101;
assign LUT_4[64421] = 32'b00000000000000000101111100110101;
assign LUT_4[64422] = 32'b00000000000000001100001011100001;
assign LUT_4[64423] = 32'b00000000000000000101010111011001;
assign LUT_4[64424] = 32'b00000000000000001000111100110110;
assign LUT_4[64425] = 32'b00000000000000000010001000101110;
assign LUT_4[64426] = 32'b00000000000000001000010111011010;
assign LUT_4[64427] = 32'b00000000000000000001100011010010;
assign LUT_4[64428] = 32'b00000000000000000101111101010010;
assign LUT_4[64429] = 32'b11111111111111111111001001001010;
assign LUT_4[64430] = 32'b00000000000000000101010111110110;
assign LUT_4[64431] = 32'b11111111111111111110100011101110;
assign LUT_4[64432] = 32'b00000000000000001101100010001111;
assign LUT_4[64433] = 32'b00000000000000000110101110000111;
assign LUT_4[64434] = 32'b00000000000000001100111100110011;
assign LUT_4[64435] = 32'b00000000000000000110001000101011;
assign LUT_4[64436] = 32'b00000000000000001010100010101011;
assign LUT_4[64437] = 32'b00000000000000000011101110100011;
assign LUT_4[64438] = 32'b00000000000000001001111101001111;
assign LUT_4[64439] = 32'b00000000000000000011001001000111;
assign LUT_4[64440] = 32'b00000000000000000110101110100100;
assign LUT_4[64441] = 32'b11111111111111111111111010011100;
assign LUT_4[64442] = 32'b00000000000000000110001001001000;
assign LUT_4[64443] = 32'b11111111111111111111010101000000;
assign LUT_4[64444] = 32'b00000000000000000011101111000000;
assign LUT_4[64445] = 32'b11111111111111111100111010111000;
assign LUT_4[64446] = 32'b00000000000000000011001001100100;
assign LUT_4[64447] = 32'b11111111111111111100010101011100;
assign LUT_4[64448] = 32'b00000000000000010010101100101110;
assign LUT_4[64449] = 32'b00000000000000001011111000100110;
assign LUT_4[64450] = 32'b00000000000000010010000111010010;
assign LUT_4[64451] = 32'b00000000000000001011010011001010;
assign LUT_4[64452] = 32'b00000000000000001111101101001010;
assign LUT_4[64453] = 32'b00000000000000001000111001000010;
assign LUT_4[64454] = 32'b00000000000000001111000111101110;
assign LUT_4[64455] = 32'b00000000000000001000010011100110;
assign LUT_4[64456] = 32'b00000000000000001011111001000011;
assign LUT_4[64457] = 32'b00000000000000000101000100111011;
assign LUT_4[64458] = 32'b00000000000000001011010011100111;
assign LUT_4[64459] = 32'b00000000000000000100011111011111;
assign LUT_4[64460] = 32'b00000000000000001000111001011111;
assign LUT_4[64461] = 32'b00000000000000000010000101010111;
assign LUT_4[64462] = 32'b00000000000000001000010100000011;
assign LUT_4[64463] = 32'b00000000000000000001011111111011;
assign LUT_4[64464] = 32'b00000000000000010000011110011100;
assign LUT_4[64465] = 32'b00000000000000001001101010010100;
assign LUT_4[64466] = 32'b00000000000000001111111001000000;
assign LUT_4[64467] = 32'b00000000000000001001000100111000;
assign LUT_4[64468] = 32'b00000000000000001101011110111000;
assign LUT_4[64469] = 32'b00000000000000000110101010110000;
assign LUT_4[64470] = 32'b00000000000000001100111001011100;
assign LUT_4[64471] = 32'b00000000000000000110000101010100;
assign LUT_4[64472] = 32'b00000000000000001001101010110001;
assign LUT_4[64473] = 32'b00000000000000000010110110101001;
assign LUT_4[64474] = 32'b00000000000000001001000101010101;
assign LUT_4[64475] = 32'b00000000000000000010010001001101;
assign LUT_4[64476] = 32'b00000000000000000110101011001101;
assign LUT_4[64477] = 32'b11111111111111111111110111000101;
assign LUT_4[64478] = 32'b00000000000000000110000101110001;
assign LUT_4[64479] = 32'b11111111111111111111010001101001;
assign LUT_4[64480] = 32'b00000000000000010001000111110101;
assign LUT_4[64481] = 32'b00000000000000001010010011101101;
assign LUT_4[64482] = 32'b00000000000000010000100010011001;
assign LUT_4[64483] = 32'b00000000000000001001101110010001;
assign LUT_4[64484] = 32'b00000000000000001110001000010001;
assign LUT_4[64485] = 32'b00000000000000000111010100001001;
assign LUT_4[64486] = 32'b00000000000000001101100010110101;
assign LUT_4[64487] = 32'b00000000000000000110101110101101;
assign LUT_4[64488] = 32'b00000000000000001010010100001010;
assign LUT_4[64489] = 32'b00000000000000000011100000000010;
assign LUT_4[64490] = 32'b00000000000000001001101110101110;
assign LUT_4[64491] = 32'b00000000000000000010111010100110;
assign LUT_4[64492] = 32'b00000000000000000111010100100110;
assign LUT_4[64493] = 32'b00000000000000000000100000011110;
assign LUT_4[64494] = 32'b00000000000000000110101111001010;
assign LUT_4[64495] = 32'b11111111111111111111111011000010;
assign LUT_4[64496] = 32'b00000000000000001110111001100011;
assign LUT_4[64497] = 32'b00000000000000001000000101011011;
assign LUT_4[64498] = 32'b00000000000000001110010100000111;
assign LUT_4[64499] = 32'b00000000000000000111011111111111;
assign LUT_4[64500] = 32'b00000000000000001011111001111111;
assign LUT_4[64501] = 32'b00000000000000000101000101110111;
assign LUT_4[64502] = 32'b00000000000000001011010100100011;
assign LUT_4[64503] = 32'b00000000000000000100100000011011;
assign LUT_4[64504] = 32'b00000000000000001000000101111000;
assign LUT_4[64505] = 32'b00000000000000000001010001110000;
assign LUT_4[64506] = 32'b00000000000000000111100000011100;
assign LUT_4[64507] = 32'b00000000000000000000101100010100;
assign LUT_4[64508] = 32'b00000000000000000101000110010100;
assign LUT_4[64509] = 32'b11111111111111111110010010001100;
assign LUT_4[64510] = 32'b00000000000000000100100000111000;
assign LUT_4[64511] = 32'b11111111111111111101101100110000;
assign LUT_4[64512] = 32'b00000000000000001100011010000110;
assign LUT_4[64513] = 32'b00000000000000000101100101111110;
assign LUT_4[64514] = 32'b00000000000000001011110100101010;
assign LUT_4[64515] = 32'b00000000000000000101000000100010;
assign LUT_4[64516] = 32'b00000000000000001001011010100010;
assign LUT_4[64517] = 32'b00000000000000000010100110011010;
assign LUT_4[64518] = 32'b00000000000000001000110101000110;
assign LUT_4[64519] = 32'b00000000000000000010000000111110;
assign LUT_4[64520] = 32'b00000000000000000101100110011011;
assign LUT_4[64521] = 32'b11111111111111111110110010010011;
assign LUT_4[64522] = 32'b00000000000000000101000000111111;
assign LUT_4[64523] = 32'b11111111111111111110001100110111;
assign LUT_4[64524] = 32'b00000000000000000010100110110111;
assign LUT_4[64525] = 32'b11111111111111111011110010101111;
assign LUT_4[64526] = 32'b00000000000000000010000001011011;
assign LUT_4[64527] = 32'b11111111111111111011001101010011;
assign LUT_4[64528] = 32'b00000000000000001010001011110100;
assign LUT_4[64529] = 32'b00000000000000000011010111101100;
assign LUT_4[64530] = 32'b00000000000000001001100110011000;
assign LUT_4[64531] = 32'b00000000000000000010110010010000;
assign LUT_4[64532] = 32'b00000000000000000111001100010000;
assign LUT_4[64533] = 32'b00000000000000000000011000001000;
assign LUT_4[64534] = 32'b00000000000000000110100110110100;
assign LUT_4[64535] = 32'b11111111111111111111110010101100;
assign LUT_4[64536] = 32'b00000000000000000011011000001001;
assign LUT_4[64537] = 32'b11111111111111111100100100000001;
assign LUT_4[64538] = 32'b00000000000000000010110010101101;
assign LUT_4[64539] = 32'b11111111111111111011111110100101;
assign LUT_4[64540] = 32'b00000000000000000000011000100101;
assign LUT_4[64541] = 32'b11111111111111111001100100011101;
assign LUT_4[64542] = 32'b11111111111111111111110011001001;
assign LUT_4[64543] = 32'b11111111111111111000111111000001;
assign LUT_4[64544] = 32'b00000000000000001010110101001101;
assign LUT_4[64545] = 32'b00000000000000000100000001000101;
assign LUT_4[64546] = 32'b00000000000000001010001111110001;
assign LUT_4[64547] = 32'b00000000000000000011011011101001;
assign LUT_4[64548] = 32'b00000000000000000111110101101001;
assign LUT_4[64549] = 32'b00000000000000000001000001100001;
assign LUT_4[64550] = 32'b00000000000000000111010000001101;
assign LUT_4[64551] = 32'b00000000000000000000011100000101;
assign LUT_4[64552] = 32'b00000000000000000100000001100010;
assign LUT_4[64553] = 32'b11111111111111111101001101011010;
assign LUT_4[64554] = 32'b00000000000000000011011100000110;
assign LUT_4[64555] = 32'b11111111111111111100100111111110;
assign LUT_4[64556] = 32'b00000000000000000001000001111110;
assign LUT_4[64557] = 32'b11111111111111111010001101110110;
assign LUT_4[64558] = 32'b00000000000000000000011100100010;
assign LUT_4[64559] = 32'b11111111111111111001101000011010;
assign LUT_4[64560] = 32'b00000000000000001000100110111011;
assign LUT_4[64561] = 32'b00000000000000000001110010110011;
assign LUT_4[64562] = 32'b00000000000000001000000001011111;
assign LUT_4[64563] = 32'b00000000000000000001001101010111;
assign LUT_4[64564] = 32'b00000000000000000101100111010111;
assign LUT_4[64565] = 32'b11111111111111111110110011001111;
assign LUT_4[64566] = 32'b00000000000000000101000001111011;
assign LUT_4[64567] = 32'b11111111111111111110001101110011;
assign LUT_4[64568] = 32'b00000000000000000001110011010000;
assign LUT_4[64569] = 32'b11111111111111111010111111001000;
assign LUT_4[64570] = 32'b00000000000000000001001101110100;
assign LUT_4[64571] = 32'b11111111111111111010011001101100;
assign LUT_4[64572] = 32'b11111111111111111110110011101100;
assign LUT_4[64573] = 32'b11111111111111110111111111100100;
assign LUT_4[64574] = 32'b11111111111111111110001110010000;
assign LUT_4[64575] = 32'b11111111111111110111011010001000;
assign LUT_4[64576] = 32'b00000000000000001101110001011010;
assign LUT_4[64577] = 32'b00000000000000000110111101010010;
assign LUT_4[64578] = 32'b00000000000000001101001011111110;
assign LUT_4[64579] = 32'b00000000000000000110010111110110;
assign LUT_4[64580] = 32'b00000000000000001010110001110110;
assign LUT_4[64581] = 32'b00000000000000000011111101101110;
assign LUT_4[64582] = 32'b00000000000000001010001100011010;
assign LUT_4[64583] = 32'b00000000000000000011011000010010;
assign LUT_4[64584] = 32'b00000000000000000110111101101111;
assign LUT_4[64585] = 32'b00000000000000000000001001100111;
assign LUT_4[64586] = 32'b00000000000000000110011000010011;
assign LUT_4[64587] = 32'b11111111111111111111100100001011;
assign LUT_4[64588] = 32'b00000000000000000011111110001011;
assign LUT_4[64589] = 32'b11111111111111111101001010000011;
assign LUT_4[64590] = 32'b00000000000000000011011000101111;
assign LUT_4[64591] = 32'b11111111111111111100100100100111;
assign LUT_4[64592] = 32'b00000000000000001011100011001000;
assign LUT_4[64593] = 32'b00000000000000000100101111000000;
assign LUT_4[64594] = 32'b00000000000000001010111101101100;
assign LUT_4[64595] = 32'b00000000000000000100001001100100;
assign LUT_4[64596] = 32'b00000000000000001000100011100100;
assign LUT_4[64597] = 32'b00000000000000000001101111011100;
assign LUT_4[64598] = 32'b00000000000000000111111110001000;
assign LUT_4[64599] = 32'b00000000000000000001001010000000;
assign LUT_4[64600] = 32'b00000000000000000100101111011101;
assign LUT_4[64601] = 32'b11111111111111111101111011010101;
assign LUT_4[64602] = 32'b00000000000000000100001010000001;
assign LUT_4[64603] = 32'b11111111111111111101010101111001;
assign LUT_4[64604] = 32'b00000000000000000001101111111001;
assign LUT_4[64605] = 32'b11111111111111111010111011110001;
assign LUT_4[64606] = 32'b00000000000000000001001010011101;
assign LUT_4[64607] = 32'b11111111111111111010010110010101;
assign LUT_4[64608] = 32'b00000000000000001100001100100001;
assign LUT_4[64609] = 32'b00000000000000000101011000011001;
assign LUT_4[64610] = 32'b00000000000000001011100111000101;
assign LUT_4[64611] = 32'b00000000000000000100110010111101;
assign LUT_4[64612] = 32'b00000000000000001001001100111101;
assign LUT_4[64613] = 32'b00000000000000000010011000110101;
assign LUT_4[64614] = 32'b00000000000000001000100111100001;
assign LUT_4[64615] = 32'b00000000000000000001110011011001;
assign LUT_4[64616] = 32'b00000000000000000101011000110110;
assign LUT_4[64617] = 32'b11111111111111111110100100101110;
assign LUT_4[64618] = 32'b00000000000000000100110011011010;
assign LUT_4[64619] = 32'b11111111111111111101111111010010;
assign LUT_4[64620] = 32'b00000000000000000010011001010010;
assign LUT_4[64621] = 32'b11111111111111111011100101001010;
assign LUT_4[64622] = 32'b00000000000000000001110011110110;
assign LUT_4[64623] = 32'b11111111111111111010111111101110;
assign LUT_4[64624] = 32'b00000000000000001001111110001111;
assign LUT_4[64625] = 32'b00000000000000000011001010000111;
assign LUT_4[64626] = 32'b00000000000000001001011000110011;
assign LUT_4[64627] = 32'b00000000000000000010100100101011;
assign LUT_4[64628] = 32'b00000000000000000110111110101011;
assign LUT_4[64629] = 32'b00000000000000000000001010100011;
assign LUT_4[64630] = 32'b00000000000000000110011001001111;
assign LUT_4[64631] = 32'b11111111111111111111100101000111;
assign LUT_4[64632] = 32'b00000000000000000011001010100100;
assign LUT_4[64633] = 32'b11111111111111111100010110011100;
assign LUT_4[64634] = 32'b00000000000000000010100101001000;
assign LUT_4[64635] = 32'b11111111111111111011110001000000;
assign LUT_4[64636] = 32'b00000000000000000000001011000000;
assign LUT_4[64637] = 32'b11111111111111111001010110111000;
assign LUT_4[64638] = 32'b11111111111111111111100101100100;
assign LUT_4[64639] = 32'b11111111111111111000110001011100;
assign LUT_4[64640] = 32'b00000000000000001111000000001110;
assign LUT_4[64641] = 32'b00000000000000001000001100000110;
assign LUT_4[64642] = 32'b00000000000000001110011010110010;
assign LUT_4[64643] = 32'b00000000000000000111100110101010;
assign LUT_4[64644] = 32'b00000000000000001100000000101010;
assign LUT_4[64645] = 32'b00000000000000000101001100100010;
assign LUT_4[64646] = 32'b00000000000000001011011011001110;
assign LUT_4[64647] = 32'b00000000000000000100100111000110;
assign LUT_4[64648] = 32'b00000000000000001000001100100011;
assign LUT_4[64649] = 32'b00000000000000000001011000011011;
assign LUT_4[64650] = 32'b00000000000000000111100111000111;
assign LUT_4[64651] = 32'b00000000000000000000110010111111;
assign LUT_4[64652] = 32'b00000000000000000101001100111111;
assign LUT_4[64653] = 32'b11111111111111111110011000110111;
assign LUT_4[64654] = 32'b00000000000000000100100111100011;
assign LUT_4[64655] = 32'b11111111111111111101110011011011;
assign LUT_4[64656] = 32'b00000000000000001100110001111100;
assign LUT_4[64657] = 32'b00000000000000000101111101110100;
assign LUT_4[64658] = 32'b00000000000000001100001100100000;
assign LUT_4[64659] = 32'b00000000000000000101011000011000;
assign LUT_4[64660] = 32'b00000000000000001001110010011000;
assign LUT_4[64661] = 32'b00000000000000000010111110010000;
assign LUT_4[64662] = 32'b00000000000000001001001100111100;
assign LUT_4[64663] = 32'b00000000000000000010011000110100;
assign LUT_4[64664] = 32'b00000000000000000101111110010001;
assign LUT_4[64665] = 32'b11111111111111111111001010001001;
assign LUT_4[64666] = 32'b00000000000000000101011000110101;
assign LUT_4[64667] = 32'b11111111111111111110100100101101;
assign LUT_4[64668] = 32'b00000000000000000010111110101101;
assign LUT_4[64669] = 32'b11111111111111111100001010100101;
assign LUT_4[64670] = 32'b00000000000000000010011001010001;
assign LUT_4[64671] = 32'b11111111111111111011100101001001;
assign LUT_4[64672] = 32'b00000000000000001101011011010101;
assign LUT_4[64673] = 32'b00000000000000000110100111001101;
assign LUT_4[64674] = 32'b00000000000000001100110101111001;
assign LUT_4[64675] = 32'b00000000000000000110000001110001;
assign LUT_4[64676] = 32'b00000000000000001010011011110001;
assign LUT_4[64677] = 32'b00000000000000000011100111101001;
assign LUT_4[64678] = 32'b00000000000000001001110110010101;
assign LUT_4[64679] = 32'b00000000000000000011000010001101;
assign LUT_4[64680] = 32'b00000000000000000110100111101010;
assign LUT_4[64681] = 32'b11111111111111111111110011100010;
assign LUT_4[64682] = 32'b00000000000000000110000010001110;
assign LUT_4[64683] = 32'b11111111111111111111001110000110;
assign LUT_4[64684] = 32'b00000000000000000011101000000110;
assign LUT_4[64685] = 32'b11111111111111111100110011111110;
assign LUT_4[64686] = 32'b00000000000000000011000010101010;
assign LUT_4[64687] = 32'b11111111111111111100001110100010;
assign LUT_4[64688] = 32'b00000000000000001011001101000011;
assign LUT_4[64689] = 32'b00000000000000000100011000111011;
assign LUT_4[64690] = 32'b00000000000000001010100111100111;
assign LUT_4[64691] = 32'b00000000000000000011110011011111;
assign LUT_4[64692] = 32'b00000000000000001000001101011111;
assign LUT_4[64693] = 32'b00000000000000000001011001010111;
assign LUT_4[64694] = 32'b00000000000000000111101000000011;
assign LUT_4[64695] = 32'b00000000000000000000110011111011;
assign LUT_4[64696] = 32'b00000000000000000100011001011000;
assign LUT_4[64697] = 32'b11111111111111111101100101010000;
assign LUT_4[64698] = 32'b00000000000000000011110011111100;
assign LUT_4[64699] = 32'b11111111111111111100111111110100;
assign LUT_4[64700] = 32'b00000000000000000001011001110100;
assign LUT_4[64701] = 32'b11111111111111111010100101101100;
assign LUT_4[64702] = 32'b00000000000000000000110100011000;
assign LUT_4[64703] = 32'b11111111111111111010000000010000;
assign LUT_4[64704] = 32'b00000000000000010000010111100010;
assign LUT_4[64705] = 32'b00000000000000001001100011011010;
assign LUT_4[64706] = 32'b00000000000000001111110010000110;
assign LUT_4[64707] = 32'b00000000000000001000111101111110;
assign LUT_4[64708] = 32'b00000000000000001101010111111110;
assign LUT_4[64709] = 32'b00000000000000000110100011110110;
assign LUT_4[64710] = 32'b00000000000000001100110010100010;
assign LUT_4[64711] = 32'b00000000000000000101111110011010;
assign LUT_4[64712] = 32'b00000000000000001001100011110111;
assign LUT_4[64713] = 32'b00000000000000000010101111101111;
assign LUT_4[64714] = 32'b00000000000000001000111110011011;
assign LUT_4[64715] = 32'b00000000000000000010001010010011;
assign LUT_4[64716] = 32'b00000000000000000110100100010011;
assign LUT_4[64717] = 32'b11111111111111111111110000001011;
assign LUT_4[64718] = 32'b00000000000000000101111110110111;
assign LUT_4[64719] = 32'b11111111111111111111001010101111;
assign LUT_4[64720] = 32'b00000000000000001110001001010000;
assign LUT_4[64721] = 32'b00000000000000000111010101001000;
assign LUT_4[64722] = 32'b00000000000000001101100011110100;
assign LUT_4[64723] = 32'b00000000000000000110101111101100;
assign LUT_4[64724] = 32'b00000000000000001011001001101100;
assign LUT_4[64725] = 32'b00000000000000000100010101100100;
assign LUT_4[64726] = 32'b00000000000000001010100100010000;
assign LUT_4[64727] = 32'b00000000000000000011110000001000;
assign LUT_4[64728] = 32'b00000000000000000111010101100101;
assign LUT_4[64729] = 32'b00000000000000000000100001011101;
assign LUT_4[64730] = 32'b00000000000000000110110000001001;
assign LUT_4[64731] = 32'b11111111111111111111111100000001;
assign LUT_4[64732] = 32'b00000000000000000100010110000001;
assign LUT_4[64733] = 32'b11111111111111111101100001111001;
assign LUT_4[64734] = 32'b00000000000000000011110000100101;
assign LUT_4[64735] = 32'b11111111111111111100111100011101;
assign LUT_4[64736] = 32'b00000000000000001110110010101001;
assign LUT_4[64737] = 32'b00000000000000000111111110100001;
assign LUT_4[64738] = 32'b00000000000000001110001101001101;
assign LUT_4[64739] = 32'b00000000000000000111011001000101;
assign LUT_4[64740] = 32'b00000000000000001011110011000101;
assign LUT_4[64741] = 32'b00000000000000000100111110111101;
assign LUT_4[64742] = 32'b00000000000000001011001101101001;
assign LUT_4[64743] = 32'b00000000000000000100011001100001;
assign LUT_4[64744] = 32'b00000000000000000111111110111110;
assign LUT_4[64745] = 32'b00000000000000000001001010110110;
assign LUT_4[64746] = 32'b00000000000000000111011001100010;
assign LUT_4[64747] = 32'b00000000000000000000100101011010;
assign LUT_4[64748] = 32'b00000000000000000100111111011010;
assign LUT_4[64749] = 32'b11111111111111111110001011010010;
assign LUT_4[64750] = 32'b00000000000000000100011001111110;
assign LUT_4[64751] = 32'b11111111111111111101100101110110;
assign LUT_4[64752] = 32'b00000000000000001100100100010111;
assign LUT_4[64753] = 32'b00000000000000000101110000001111;
assign LUT_4[64754] = 32'b00000000000000001011111110111011;
assign LUT_4[64755] = 32'b00000000000000000101001010110011;
assign LUT_4[64756] = 32'b00000000000000001001100100110011;
assign LUT_4[64757] = 32'b00000000000000000010110000101011;
assign LUT_4[64758] = 32'b00000000000000001000111111010111;
assign LUT_4[64759] = 32'b00000000000000000010001011001111;
assign LUT_4[64760] = 32'b00000000000000000101110000101100;
assign LUT_4[64761] = 32'b11111111111111111110111100100100;
assign LUT_4[64762] = 32'b00000000000000000101001011010000;
assign LUT_4[64763] = 32'b11111111111111111110010111001000;
assign LUT_4[64764] = 32'b00000000000000000010110001001000;
assign LUT_4[64765] = 32'b11111111111111111011111101000000;
assign LUT_4[64766] = 32'b00000000000000000010001011101100;
assign LUT_4[64767] = 32'b11111111111111111011010111100100;
assign LUT_4[64768] = 32'b00000000000000010001010101101001;
assign LUT_4[64769] = 32'b00000000000000001010100001100001;
assign LUT_4[64770] = 32'b00000000000000010000110000001101;
assign LUT_4[64771] = 32'b00000000000000001001111100000101;
assign LUT_4[64772] = 32'b00000000000000001110010110000101;
assign LUT_4[64773] = 32'b00000000000000000111100001111101;
assign LUT_4[64774] = 32'b00000000000000001101110000101001;
assign LUT_4[64775] = 32'b00000000000000000110111100100001;
assign LUT_4[64776] = 32'b00000000000000001010100001111110;
assign LUT_4[64777] = 32'b00000000000000000011101101110110;
assign LUT_4[64778] = 32'b00000000000000001001111100100010;
assign LUT_4[64779] = 32'b00000000000000000011001000011010;
assign LUT_4[64780] = 32'b00000000000000000111100010011010;
assign LUT_4[64781] = 32'b00000000000000000000101110010010;
assign LUT_4[64782] = 32'b00000000000000000110111100111110;
assign LUT_4[64783] = 32'b00000000000000000000001000110110;
assign LUT_4[64784] = 32'b00000000000000001111000111010111;
assign LUT_4[64785] = 32'b00000000000000001000010011001111;
assign LUT_4[64786] = 32'b00000000000000001110100001111011;
assign LUT_4[64787] = 32'b00000000000000000111101101110011;
assign LUT_4[64788] = 32'b00000000000000001100000111110011;
assign LUT_4[64789] = 32'b00000000000000000101010011101011;
assign LUT_4[64790] = 32'b00000000000000001011100010010111;
assign LUT_4[64791] = 32'b00000000000000000100101110001111;
assign LUT_4[64792] = 32'b00000000000000001000010011101100;
assign LUT_4[64793] = 32'b00000000000000000001011111100100;
assign LUT_4[64794] = 32'b00000000000000000111101110010000;
assign LUT_4[64795] = 32'b00000000000000000000111010001000;
assign LUT_4[64796] = 32'b00000000000000000101010100001000;
assign LUT_4[64797] = 32'b11111111111111111110100000000000;
assign LUT_4[64798] = 32'b00000000000000000100101110101100;
assign LUT_4[64799] = 32'b11111111111111111101111010100100;
assign LUT_4[64800] = 32'b00000000000000001111110000110000;
assign LUT_4[64801] = 32'b00000000000000001000111100101000;
assign LUT_4[64802] = 32'b00000000000000001111001011010100;
assign LUT_4[64803] = 32'b00000000000000001000010111001100;
assign LUT_4[64804] = 32'b00000000000000001100110001001100;
assign LUT_4[64805] = 32'b00000000000000000101111101000100;
assign LUT_4[64806] = 32'b00000000000000001100001011110000;
assign LUT_4[64807] = 32'b00000000000000000101010111101000;
assign LUT_4[64808] = 32'b00000000000000001000111101000101;
assign LUT_4[64809] = 32'b00000000000000000010001000111101;
assign LUT_4[64810] = 32'b00000000000000001000010111101001;
assign LUT_4[64811] = 32'b00000000000000000001100011100001;
assign LUT_4[64812] = 32'b00000000000000000101111101100001;
assign LUT_4[64813] = 32'b11111111111111111111001001011001;
assign LUT_4[64814] = 32'b00000000000000000101011000000101;
assign LUT_4[64815] = 32'b11111111111111111110100011111101;
assign LUT_4[64816] = 32'b00000000000000001101100010011110;
assign LUT_4[64817] = 32'b00000000000000000110101110010110;
assign LUT_4[64818] = 32'b00000000000000001100111101000010;
assign LUT_4[64819] = 32'b00000000000000000110001000111010;
assign LUT_4[64820] = 32'b00000000000000001010100010111010;
assign LUT_4[64821] = 32'b00000000000000000011101110110010;
assign LUT_4[64822] = 32'b00000000000000001001111101011110;
assign LUT_4[64823] = 32'b00000000000000000011001001010110;
assign LUT_4[64824] = 32'b00000000000000000110101110110011;
assign LUT_4[64825] = 32'b11111111111111111111111010101011;
assign LUT_4[64826] = 32'b00000000000000000110001001010111;
assign LUT_4[64827] = 32'b11111111111111111111010101001111;
assign LUT_4[64828] = 32'b00000000000000000011101111001111;
assign LUT_4[64829] = 32'b11111111111111111100111011000111;
assign LUT_4[64830] = 32'b00000000000000000011001001110011;
assign LUT_4[64831] = 32'b11111111111111111100010101101011;
assign LUT_4[64832] = 32'b00000000000000010010101100111101;
assign LUT_4[64833] = 32'b00000000000000001011111000110101;
assign LUT_4[64834] = 32'b00000000000000010010000111100001;
assign LUT_4[64835] = 32'b00000000000000001011010011011001;
assign LUT_4[64836] = 32'b00000000000000001111101101011001;
assign LUT_4[64837] = 32'b00000000000000001000111001010001;
assign LUT_4[64838] = 32'b00000000000000001111000111111101;
assign LUT_4[64839] = 32'b00000000000000001000010011110101;
assign LUT_4[64840] = 32'b00000000000000001011111001010010;
assign LUT_4[64841] = 32'b00000000000000000101000101001010;
assign LUT_4[64842] = 32'b00000000000000001011010011110110;
assign LUT_4[64843] = 32'b00000000000000000100011111101110;
assign LUT_4[64844] = 32'b00000000000000001000111001101110;
assign LUT_4[64845] = 32'b00000000000000000010000101100110;
assign LUT_4[64846] = 32'b00000000000000001000010100010010;
assign LUT_4[64847] = 32'b00000000000000000001100000001010;
assign LUT_4[64848] = 32'b00000000000000010000011110101011;
assign LUT_4[64849] = 32'b00000000000000001001101010100011;
assign LUT_4[64850] = 32'b00000000000000001111111001001111;
assign LUT_4[64851] = 32'b00000000000000001001000101000111;
assign LUT_4[64852] = 32'b00000000000000001101011111000111;
assign LUT_4[64853] = 32'b00000000000000000110101010111111;
assign LUT_4[64854] = 32'b00000000000000001100111001101011;
assign LUT_4[64855] = 32'b00000000000000000110000101100011;
assign LUT_4[64856] = 32'b00000000000000001001101011000000;
assign LUT_4[64857] = 32'b00000000000000000010110110111000;
assign LUT_4[64858] = 32'b00000000000000001001000101100100;
assign LUT_4[64859] = 32'b00000000000000000010010001011100;
assign LUT_4[64860] = 32'b00000000000000000110101011011100;
assign LUT_4[64861] = 32'b11111111111111111111110111010100;
assign LUT_4[64862] = 32'b00000000000000000110000110000000;
assign LUT_4[64863] = 32'b11111111111111111111010001111000;
assign LUT_4[64864] = 32'b00000000000000010001001000000100;
assign LUT_4[64865] = 32'b00000000000000001010010011111100;
assign LUT_4[64866] = 32'b00000000000000010000100010101000;
assign LUT_4[64867] = 32'b00000000000000001001101110100000;
assign LUT_4[64868] = 32'b00000000000000001110001000100000;
assign LUT_4[64869] = 32'b00000000000000000111010100011000;
assign LUT_4[64870] = 32'b00000000000000001101100011000100;
assign LUT_4[64871] = 32'b00000000000000000110101110111100;
assign LUT_4[64872] = 32'b00000000000000001010010100011001;
assign LUT_4[64873] = 32'b00000000000000000011100000010001;
assign LUT_4[64874] = 32'b00000000000000001001101110111101;
assign LUT_4[64875] = 32'b00000000000000000010111010110101;
assign LUT_4[64876] = 32'b00000000000000000111010100110101;
assign LUT_4[64877] = 32'b00000000000000000000100000101101;
assign LUT_4[64878] = 32'b00000000000000000110101111011001;
assign LUT_4[64879] = 32'b11111111111111111111111011010001;
assign LUT_4[64880] = 32'b00000000000000001110111001110010;
assign LUT_4[64881] = 32'b00000000000000001000000101101010;
assign LUT_4[64882] = 32'b00000000000000001110010100010110;
assign LUT_4[64883] = 32'b00000000000000000111100000001110;
assign LUT_4[64884] = 32'b00000000000000001011111010001110;
assign LUT_4[64885] = 32'b00000000000000000101000110000110;
assign LUT_4[64886] = 32'b00000000000000001011010100110010;
assign LUT_4[64887] = 32'b00000000000000000100100000101010;
assign LUT_4[64888] = 32'b00000000000000001000000110000111;
assign LUT_4[64889] = 32'b00000000000000000001010001111111;
assign LUT_4[64890] = 32'b00000000000000000111100000101011;
assign LUT_4[64891] = 32'b00000000000000000000101100100011;
assign LUT_4[64892] = 32'b00000000000000000101000110100011;
assign LUT_4[64893] = 32'b11111111111111111110010010011011;
assign LUT_4[64894] = 32'b00000000000000000100100001000111;
assign LUT_4[64895] = 32'b11111111111111111101101100111111;
assign LUT_4[64896] = 32'b00000000000000010011111011110001;
assign LUT_4[64897] = 32'b00000000000000001101000111101001;
assign LUT_4[64898] = 32'b00000000000000010011010110010101;
assign LUT_4[64899] = 32'b00000000000000001100100010001101;
assign LUT_4[64900] = 32'b00000000000000010000111100001101;
assign LUT_4[64901] = 32'b00000000000000001010001000000101;
assign LUT_4[64902] = 32'b00000000000000010000010110110001;
assign LUT_4[64903] = 32'b00000000000000001001100010101001;
assign LUT_4[64904] = 32'b00000000000000001101001000000110;
assign LUT_4[64905] = 32'b00000000000000000110010011111110;
assign LUT_4[64906] = 32'b00000000000000001100100010101010;
assign LUT_4[64907] = 32'b00000000000000000101101110100010;
assign LUT_4[64908] = 32'b00000000000000001010001000100010;
assign LUT_4[64909] = 32'b00000000000000000011010100011010;
assign LUT_4[64910] = 32'b00000000000000001001100011000110;
assign LUT_4[64911] = 32'b00000000000000000010101110111110;
assign LUT_4[64912] = 32'b00000000000000010001101101011111;
assign LUT_4[64913] = 32'b00000000000000001010111001010111;
assign LUT_4[64914] = 32'b00000000000000010001001000000011;
assign LUT_4[64915] = 32'b00000000000000001010010011111011;
assign LUT_4[64916] = 32'b00000000000000001110101101111011;
assign LUT_4[64917] = 32'b00000000000000000111111001110011;
assign LUT_4[64918] = 32'b00000000000000001110001000011111;
assign LUT_4[64919] = 32'b00000000000000000111010100010111;
assign LUT_4[64920] = 32'b00000000000000001010111001110100;
assign LUT_4[64921] = 32'b00000000000000000100000101101100;
assign LUT_4[64922] = 32'b00000000000000001010010100011000;
assign LUT_4[64923] = 32'b00000000000000000011100000010000;
assign LUT_4[64924] = 32'b00000000000000000111111010010000;
assign LUT_4[64925] = 32'b00000000000000000001000110001000;
assign LUT_4[64926] = 32'b00000000000000000111010100110100;
assign LUT_4[64927] = 32'b00000000000000000000100000101100;
assign LUT_4[64928] = 32'b00000000000000010010010110111000;
assign LUT_4[64929] = 32'b00000000000000001011100010110000;
assign LUT_4[64930] = 32'b00000000000000010001110001011100;
assign LUT_4[64931] = 32'b00000000000000001010111101010100;
assign LUT_4[64932] = 32'b00000000000000001111010111010100;
assign LUT_4[64933] = 32'b00000000000000001000100011001100;
assign LUT_4[64934] = 32'b00000000000000001110110001111000;
assign LUT_4[64935] = 32'b00000000000000000111111101110000;
assign LUT_4[64936] = 32'b00000000000000001011100011001101;
assign LUT_4[64937] = 32'b00000000000000000100101111000101;
assign LUT_4[64938] = 32'b00000000000000001010111101110001;
assign LUT_4[64939] = 32'b00000000000000000100001001101001;
assign LUT_4[64940] = 32'b00000000000000001000100011101001;
assign LUT_4[64941] = 32'b00000000000000000001101111100001;
assign LUT_4[64942] = 32'b00000000000000000111111110001101;
assign LUT_4[64943] = 32'b00000000000000000001001010000101;
assign LUT_4[64944] = 32'b00000000000000010000001000100110;
assign LUT_4[64945] = 32'b00000000000000001001010100011110;
assign LUT_4[64946] = 32'b00000000000000001111100011001010;
assign LUT_4[64947] = 32'b00000000000000001000101111000010;
assign LUT_4[64948] = 32'b00000000000000001101001001000010;
assign LUT_4[64949] = 32'b00000000000000000110010100111010;
assign LUT_4[64950] = 32'b00000000000000001100100011100110;
assign LUT_4[64951] = 32'b00000000000000000101101111011110;
assign LUT_4[64952] = 32'b00000000000000001001010100111011;
assign LUT_4[64953] = 32'b00000000000000000010100000110011;
assign LUT_4[64954] = 32'b00000000000000001000101111011111;
assign LUT_4[64955] = 32'b00000000000000000001111011010111;
assign LUT_4[64956] = 32'b00000000000000000110010101010111;
assign LUT_4[64957] = 32'b11111111111111111111100001001111;
assign LUT_4[64958] = 32'b00000000000000000101101111111011;
assign LUT_4[64959] = 32'b11111111111111111110111011110011;
assign LUT_4[64960] = 32'b00000000000000010101010011000101;
assign LUT_4[64961] = 32'b00000000000000001110011110111101;
assign LUT_4[64962] = 32'b00000000000000010100101101101001;
assign LUT_4[64963] = 32'b00000000000000001101111001100001;
assign LUT_4[64964] = 32'b00000000000000010010010011100001;
assign LUT_4[64965] = 32'b00000000000000001011011111011001;
assign LUT_4[64966] = 32'b00000000000000010001101110000101;
assign LUT_4[64967] = 32'b00000000000000001010111001111101;
assign LUT_4[64968] = 32'b00000000000000001110011111011010;
assign LUT_4[64969] = 32'b00000000000000000111101011010010;
assign LUT_4[64970] = 32'b00000000000000001101111001111110;
assign LUT_4[64971] = 32'b00000000000000000111000101110110;
assign LUT_4[64972] = 32'b00000000000000001011011111110110;
assign LUT_4[64973] = 32'b00000000000000000100101011101110;
assign LUT_4[64974] = 32'b00000000000000001010111010011010;
assign LUT_4[64975] = 32'b00000000000000000100000110010010;
assign LUT_4[64976] = 32'b00000000000000010011000100110011;
assign LUT_4[64977] = 32'b00000000000000001100010000101011;
assign LUT_4[64978] = 32'b00000000000000010010011111010111;
assign LUT_4[64979] = 32'b00000000000000001011101011001111;
assign LUT_4[64980] = 32'b00000000000000010000000101001111;
assign LUT_4[64981] = 32'b00000000000000001001010001000111;
assign LUT_4[64982] = 32'b00000000000000001111011111110011;
assign LUT_4[64983] = 32'b00000000000000001000101011101011;
assign LUT_4[64984] = 32'b00000000000000001100010001001000;
assign LUT_4[64985] = 32'b00000000000000000101011101000000;
assign LUT_4[64986] = 32'b00000000000000001011101011101100;
assign LUT_4[64987] = 32'b00000000000000000100110111100100;
assign LUT_4[64988] = 32'b00000000000000001001010001100100;
assign LUT_4[64989] = 32'b00000000000000000010011101011100;
assign LUT_4[64990] = 32'b00000000000000001000101100001000;
assign LUT_4[64991] = 32'b00000000000000000001111000000000;
assign LUT_4[64992] = 32'b00000000000000010011101110001100;
assign LUT_4[64993] = 32'b00000000000000001100111010000100;
assign LUT_4[64994] = 32'b00000000000000010011001000110000;
assign LUT_4[64995] = 32'b00000000000000001100010100101000;
assign LUT_4[64996] = 32'b00000000000000010000101110101000;
assign LUT_4[64997] = 32'b00000000000000001001111010100000;
assign LUT_4[64998] = 32'b00000000000000010000001001001100;
assign LUT_4[64999] = 32'b00000000000000001001010101000100;
assign LUT_4[65000] = 32'b00000000000000001100111010100001;
assign LUT_4[65001] = 32'b00000000000000000110000110011001;
assign LUT_4[65002] = 32'b00000000000000001100010101000101;
assign LUT_4[65003] = 32'b00000000000000000101100000111101;
assign LUT_4[65004] = 32'b00000000000000001001111010111101;
assign LUT_4[65005] = 32'b00000000000000000011000110110101;
assign LUT_4[65006] = 32'b00000000000000001001010101100001;
assign LUT_4[65007] = 32'b00000000000000000010100001011001;
assign LUT_4[65008] = 32'b00000000000000010001011111111010;
assign LUT_4[65009] = 32'b00000000000000001010101011110010;
assign LUT_4[65010] = 32'b00000000000000010000111010011110;
assign LUT_4[65011] = 32'b00000000000000001010000110010110;
assign LUT_4[65012] = 32'b00000000000000001110100000010110;
assign LUT_4[65013] = 32'b00000000000000000111101100001110;
assign LUT_4[65014] = 32'b00000000000000001101111010111010;
assign LUT_4[65015] = 32'b00000000000000000111000110110010;
assign LUT_4[65016] = 32'b00000000000000001010101100001111;
assign LUT_4[65017] = 32'b00000000000000000011111000000111;
assign LUT_4[65018] = 32'b00000000000000001010000110110011;
assign LUT_4[65019] = 32'b00000000000000000011010010101011;
assign LUT_4[65020] = 32'b00000000000000000111101100101011;
assign LUT_4[65021] = 32'b00000000000000000000111000100011;
assign LUT_4[65022] = 32'b00000000000000000111000111001111;
assign LUT_4[65023] = 32'b00000000000000000000010011000111;
assign LUT_4[65024] = 32'b00000000000000001011011110001110;
assign LUT_4[65025] = 32'b00000000000000000100101010000110;
assign LUT_4[65026] = 32'b00000000000000001010111000110010;
assign LUT_4[65027] = 32'b00000000000000000100000100101010;
assign LUT_4[65028] = 32'b00000000000000001000011110101010;
assign LUT_4[65029] = 32'b00000000000000000001101010100010;
assign LUT_4[65030] = 32'b00000000000000000111111001001110;
assign LUT_4[65031] = 32'b00000000000000000001000101000110;
assign LUT_4[65032] = 32'b00000000000000000100101010100011;
assign LUT_4[65033] = 32'b11111111111111111101110110011011;
assign LUT_4[65034] = 32'b00000000000000000100000101000111;
assign LUT_4[65035] = 32'b11111111111111111101010000111111;
assign LUT_4[65036] = 32'b00000000000000000001101010111111;
assign LUT_4[65037] = 32'b11111111111111111010110110110111;
assign LUT_4[65038] = 32'b00000000000000000001000101100011;
assign LUT_4[65039] = 32'b11111111111111111010010001011011;
assign LUT_4[65040] = 32'b00000000000000001001001111111100;
assign LUT_4[65041] = 32'b00000000000000000010011011110100;
assign LUT_4[65042] = 32'b00000000000000001000101010100000;
assign LUT_4[65043] = 32'b00000000000000000001110110011000;
assign LUT_4[65044] = 32'b00000000000000000110010000011000;
assign LUT_4[65045] = 32'b11111111111111111111011100010000;
assign LUT_4[65046] = 32'b00000000000000000101101010111100;
assign LUT_4[65047] = 32'b11111111111111111110110110110100;
assign LUT_4[65048] = 32'b00000000000000000010011100010001;
assign LUT_4[65049] = 32'b11111111111111111011101000001001;
assign LUT_4[65050] = 32'b00000000000000000001110110110101;
assign LUT_4[65051] = 32'b11111111111111111011000010101101;
assign LUT_4[65052] = 32'b11111111111111111111011100101101;
assign LUT_4[65053] = 32'b11111111111111111000101000100101;
assign LUT_4[65054] = 32'b11111111111111111110110111010001;
assign LUT_4[65055] = 32'b11111111111111111000000011001001;
assign LUT_4[65056] = 32'b00000000000000001001111001010101;
assign LUT_4[65057] = 32'b00000000000000000011000101001101;
assign LUT_4[65058] = 32'b00000000000000001001010011111001;
assign LUT_4[65059] = 32'b00000000000000000010011111110001;
assign LUT_4[65060] = 32'b00000000000000000110111001110001;
assign LUT_4[65061] = 32'b00000000000000000000000101101001;
assign LUT_4[65062] = 32'b00000000000000000110010100010101;
assign LUT_4[65063] = 32'b11111111111111111111100000001101;
assign LUT_4[65064] = 32'b00000000000000000011000101101010;
assign LUT_4[65065] = 32'b11111111111111111100010001100010;
assign LUT_4[65066] = 32'b00000000000000000010100000001110;
assign LUT_4[65067] = 32'b11111111111111111011101100000110;
assign LUT_4[65068] = 32'b00000000000000000000000110000110;
assign LUT_4[65069] = 32'b11111111111111111001010001111110;
assign LUT_4[65070] = 32'b11111111111111111111100000101010;
assign LUT_4[65071] = 32'b11111111111111111000101100100010;
assign LUT_4[65072] = 32'b00000000000000000111101011000011;
assign LUT_4[65073] = 32'b00000000000000000000110110111011;
assign LUT_4[65074] = 32'b00000000000000000111000101100111;
assign LUT_4[65075] = 32'b00000000000000000000010001011111;
assign LUT_4[65076] = 32'b00000000000000000100101011011111;
assign LUT_4[65077] = 32'b11111111111111111101110111010111;
assign LUT_4[65078] = 32'b00000000000000000100000110000011;
assign LUT_4[65079] = 32'b11111111111111111101010001111011;
assign LUT_4[65080] = 32'b00000000000000000000110111011000;
assign LUT_4[65081] = 32'b11111111111111111010000011010000;
assign LUT_4[65082] = 32'b00000000000000000000010001111100;
assign LUT_4[65083] = 32'b11111111111111111001011101110100;
assign LUT_4[65084] = 32'b11111111111111111101110111110100;
assign LUT_4[65085] = 32'b11111111111111110111000011101100;
assign LUT_4[65086] = 32'b11111111111111111101010010011000;
assign LUT_4[65087] = 32'b11111111111111110110011110010000;
assign LUT_4[65088] = 32'b00000000000000001100110101100010;
assign LUT_4[65089] = 32'b00000000000000000110000001011010;
assign LUT_4[65090] = 32'b00000000000000001100010000000110;
assign LUT_4[65091] = 32'b00000000000000000101011011111110;
assign LUT_4[65092] = 32'b00000000000000001001110101111110;
assign LUT_4[65093] = 32'b00000000000000000011000001110110;
assign LUT_4[65094] = 32'b00000000000000001001010000100010;
assign LUT_4[65095] = 32'b00000000000000000010011100011010;
assign LUT_4[65096] = 32'b00000000000000000110000001110111;
assign LUT_4[65097] = 32'b11111111111111111111001101101111;
assign LUT_4[65098] = 32'b00000000000000000101011100011011;
assign LUT_4[65099] = 32'b11111111111111111110101000010011;
assign LUT_4[65100] = 32'b00000000000000000011000010010011;
assign LUT_4[65101] = 32'b11111111111111111100001110001011;
assign LUT_4[65102] = 32'b00000000000000000010011100110111;
assign LUT_4[65103] = 32'b11111111111111111011101000101111;
assign LUT_4[65104] = 32'b00000000000000001010100111010000;
assign LUT_4[65105] = 32'b00000000000000000011110011001000;
assign LUT_4[65106] = 32'b00000000000000001010000001110100;
assign LUT_4[65107] = 32'b00000000000000000011001101101100;
assign LUT_4[65108] = 32'b00000000000000000111100111101100;
assign LUT_4[65109] = 32'b00000000000000000000110011100100;
assign LUT_4[65110] = 32'b00000000000000000111000010010000;
assign LUT_4[65111] = 32'b00000000000000000000001110001000;
assign LUT_4[65112] = 32'b00000000000000000011110011100101;
assign LUT_4[65113] = 32'b11111111111111111100111111011101;
assign LUT_4[65114] = 32'b00000000000000000011001110001001;
assign LUT_4[65115] = 32'b11111111111111111100011010000001;
assign LUT_4[65116] = 32'b00000000000000000000110100000001;
assign LUT_4[65117] = 32'b11111111111111111001111111111001;
assign LUT_4[65118] = 32'b00000000000000000000001110100101;
assign LUT_4[65119] = 32'b11111111111111111001011010011101;
assign LUT_4[65120] = 32'b00000000000000001011010000101001;
assign LUT_4[65121] = 32'b00000000000000000100011100100001;
assign LUT_4[65122] = 32'b00000000000000001010101011001101;
assign LUT_4[65123] = 32'b00000000000000000011110111000101;
assign LUT_4[65124] = 32'b00000000000000001000010001000101;
assign LUT_4[65125] = 32'b00000000000000000001011100111101;
assign LUT_4[65126] = 32'b00000000000000000111101011101001;
assign LUT_4[65127] = 32'b00000000000000000000110111100001;
assign LUT_4[65128] = 32'b00000000000000000100011100111110;
assign LUT_4[65129] = 32'b11111111111111111101101000110110;
assign LUT_4[65130] = 32'b00000000000000000011110111100010;
assign LUT_4[65131] = 32'b11111111111111111101000011011010;
assign LUT_4[65132] = 32'b00000000000000000001011101011010;
assign LUT_4[65133] = 32'b11111111111111111010101001010010;
assign LUT_4[65134] = 32'b00000000000000000000110111111110;
assign LUT_4[65135] = 32'b11111111111111111010000011110110;
assign LUT_4[65136] = 32'b00000000000000001001000010010111;
assign LUT_4[65137] = 32'b00000000000000000010001110001111;
assign LUT_4[65138] = 32'b00000000000000001000011100111011;
assign LUT_4[65139] = 32'b00000000000000000001101000110011;
assign LUT_4[65140] = 32'b00000000000000000110000010110011;
assign LUT_4[65141] = 32'b11111111111111111111001110101011;
assign LUT_4[65142] = 32'b00000000000000000101011101010111;
assign LUT_4[65143] = 32'b11111111111111111110101001001111;
assign LUT_4[65144] = 32'b00000000000000000010001110101100;
assign LUT_4[65145] = 32'b11111111111111111011011010100100;
assign LUT_4[65146] = 32'b00000000000000000001101001010000;
assign LUT_4[65147] = 32'b11111111111111111010110101001000;
assign LUT_4[65148] = 32'b11111111111111111111001111001000;
assign LUT_4[65149] = 32'b11111111111111111000011011000000;
assign LUT_4[65150] = 32'b11111111111111111110101001101100;
assign LUT_4[65151] = 32'b11111111111111110111110101100100;
assign LUT_4[65152] = 32'b00000000000000001110000100010110;
assign LUT_4[65153] = 32'b00000000000000000111010000001110;
assign LUT_4[65154] = 32'b00000000000000001101011110111010;
assign LUT_4[65155] = 32'b00000000000000000110101010110010;
assign LUT_4[65156] = 32'b00000000000000001011000100110010;
assign LUT_4[65157] = 32'b00000000000000000100010000101010;
assign LUT_4[65158] = 32'b00000000000000001010011111010110;
assign LUT_4[65159] = 32'b00000000000000000011101011001110;
assign LUT_4[65160] = 32'b00000000000000000111010000101011;
assign LUT_4[65161] = 32'b00000000000000000000011100100011;
assign LUT_4[65162] = 32'b00000000000000000110101011001111;
assign LUT_4[65163] = 32'b11111111111111111111110111000111;
assign LUT_4[65164] = 32'b00000000000000000100010001000111;
assign LUT_4[65165] = 32'b11111111111111111101011100111111;
assign LUT_4[65166] = 32'b00000000000000000011101011101011;
assign LUT_4[65167] = 32'b11111111111111111100110111100011;
assign LUT_4[65168] = 32'b00000000000000001011110110000100;
assign LUT_4[65169] = 32'b00000000000000000101000001111100;
assign LUT_4[65170] = 32'b00000000000000001011010000101000;
assign LUT_4[65171] = 32'b00000000000000000100011100100000;
assign LUT_4[65172] = 32'b00000000000000001000110110100000;
assign LUT_4[65173] = 32'b00000000000000000010000010011000;
assign LUT_4[65174] = 32'b00000000000000001000010001000100;
assign LUT_4[65175] = 32'b00000000000000000001011100111100;
assign LUT_4[65176] = 32'b00000000000000000101000010011001;
assign LUT_4[65177] = 32'b11111111111111111110001110010001;
assign LUT_4[65178] = 32'b00000000000000000100011100111101;
assign LUT_4[65179] = 32'b11111111111111111101101000110101;
assign LUT_4[65180] = 32'b00000000000000000010000010110101;
assign LUT_4[65181] = 32'b11111111111111111011001110101101;
assign LUT_4[65182] = 32'b00000000000000000001011101011001;
assign LUT_4[65183] = 32'b11111111111111111010101001010001;
assign LUT_4[65184] = 32'b00000000000000001100011111011101;
assign LUT_4[65185] = 32'b00000000000000000101101011010101;
assign LUT_4[65186] = 32'b00000000000000001011111010000001;
assign LUT_4[65187] = 32'b00000000000000000101000101111001;
assign LUT_4[65188] = 32'b00000000000000001001011111111001;
assign LUT_4[65189] = 32'b00000000000000000010101011110001;
assign LUT_4[65190] = 32'b00000000000000001000111010011101;
assign LUT_4[65191] = 32'b00000000000000000010000110010101;
assign LUT_4[65192] = 32'b00000000000000000101101011110010;
assign LUT_4[65193] = 32'b11111111111111111110110111101010;
assign LUT_4[65194] = 32'b00000000000000000101000110010110;
assign LUT_4[65195] = 32'b11111111111111111110010010001110;
assign LUT_4[65196] = 32'b00000000000000000010101100001110;
assign LUT_4[65197] = 32'b11111111111111111011111000000110;
assign LUT_4[65198] = 32'b00000000000000000010000110110010;
assign LUT_4[65199] = 32'b11111111111111111011010010101010;
assign LUT_4[65200] = 32'b00000000000000001010010001001011;
assign LUT_4[65201] = 32'b00000000000000000011011101000011;
assign LUT_4[65202] = 32'b00000000000000001001101011101111;
assign LUT_4[65203] = 32'b00000000000000000010110111100111;
assign LUT_4[65204] = 32'b00000000000000000111010001100111;
assign LUT_4[65205] = 32'b00000000000000000000011101011111;
assign LUT_4[65206] = 32'b00000000000000000110101100001011;
assign LUT_4[65207] = 32'b11111111111111111111111000000011;
assign LUT_4[65208] = 32'b00000000000000000011011101100000;
assign LUT_4[65209] = 32'b11111111111111111100101001011000;
assign LUT_4[65210] = 32'b00000000000000000010111000000100;
assign LUT_4[65211] = 32'b11111111111111111100000011111100;
assign LUT_4[65212] = 32'b00000000000000000000011101111100;
assign LUT_4[65213] = 32'b11111111111111111001101001110100;
assign LUT_4[65214] = 32'b11111111111111111111111000100000;
assign LUT_4[65215] = 32'b11111111111111111001000100011000;
assign LUT_4[65216] = 32'b00000000000000001111011011101010;
assign LUT_4[65217] = 32'b00000000000000001000100111100010;
assign LUT_4[65218] = 32'b00000000000000001110110110001110;
assign LUT_4[65219] = 32'b00000000000000001000000010000110;
assign LUT_4[65220] = 32'b00000000000000001100011100000110;
assign LUT_4[65221] = 32'b00000000000000000101100111111110;
assign LUT_4[65222] = 32'b00000000000000001011110110101010;
assign LUT_4[65223] = 32'b00000000000000000101000010100010;
assign LUT_4[65224] = 32'b00000000000000001000100111111111;
assign LUT_4[65225] = 32'b00000000000000000001110011110111;
assign LUT_4[65226] = 32'b00000000000000001000000010100011;
assign LUT_4[65227] = 32'b00000000000000000001001110011011;
assign LUT_4[65228] = 32'b00000000000000000101101000011011;
assign LUT_4[65229] = 32'b11111111111111111110110100010011;
assign LUT_4[65230] = 32'b00000000000000000101000010111111;
assign LUT_4[65231] = 32'b11111111111111111110001110110111;
assign LUT_4[65232] = 32'b00000000000000001101001101011000;
assign LUT_4[65233] = 32'b00000000000000000110011001010000;
assign LUT_4[65234] = 32'b00000000000000001100100111111100;
assign LUT_4[65235] = 32'b00000000000000000101110011110100;
assign LUT_4[65236] = 32'b00000000000000001010001101110100;
assign LUT_4[65237] = 32'b00000000000000000011011001101100;
assign LUT_4[65238] = 32'b00000000000000001001101000011000;
assign LUT_4[65239] = 32'b00000000000000000010110100010000;
assign LUT_4[65240] = 32'b00000000000000000110011001101101;
assign LUT_4[65241] = 32'b11111111111111111111100101100101;
assign LUT_4[65242] = 32'b00000000000000000101110100010001;
assign LUT_4[65243] = 32'b11111111111111111111000000001001;
assign LUT_4[65244] = 32'b00000000000000000011011010001001;
assign LUT_4[65245] = 32'b11111111111111111100100110000001;
assign LUT_4[65246] = 32'b00000000000000000010110100101101;
assign LUT_4[65247] = 32'b11111111111111111100000000100101;
assign LUT_4[65248] = 32'b00000000000000001101110110110001;
assign LUT_4[65249] = 32'b00000000000000000111000010101001;
assign LUT_4[65250] = 32'b00000000000000001101010001010101;
assign LUT_4[65251] = 32'b00000000000000000110011101001101;
assign LUT_4[65252] = 32'b00000000000000001010110111001101;
assign LUT_4[65253] = 32'b00000000000000000100000011000101;
assign LUT_4[65254] = 32'b00000000000000001010010001110001;
assign LUT_4[65255] = 32'b00000000000000000011011101101001;
assign LUT_4[65256] = 32'b00000000000000000111000011000110;
assign LUT_4[65257] = 32'b00000000000000000000001110111110;
assign LUT_4[65258] = 32'b00000000000000000110011101101010;
assign LUT_4[65259] = 32'b11111111111111111111101001100010;
assign LUT_4[65260] = 32'b00000000000000000100000011100010;
assign LUT_4[65261] = 32'b11111111111111111101001111011010;
assign LUT_4[65262] = 32'b00000000000000000011011110000110;
assign LUT_4[65263] = 32'b11111111111111111100101001111110;
assign LUT_4[65264] = 32'b00000000000000001011101000011111;
assign LUT_4[65265] = 32'b00000000000000000100110100010111;
assign LUT_4[65266] = 32'b00000000000000001011000011000011;
assign LUT_4[65267] = 32'b00000000000000000100001110111011;
assign LUT_4[65268] = 32'b00000000000000001000101000111011;
assign LUT_4[65269] = 32'b00000000000000000001110100110011;
assign LUT_4[65270] = 32'b00000000000000001000000011011111;
assign LUT_4[65271] = 32'b00000000000000000001001111010111;
assign LUT_4[65272] = 32'b00000000000000000100110100110100;
assign LUT_4[65273] = 32'b11111111111111111110000000101100;
assign LUT_4[65274] = 32'b00000000000000000100001111011000;
assign LUT_4[65275] = 32'b11111111111111111101011011010000;
assign LUT_4[65276] = 32'b00000000000000000001110101010000;
assign LUT_4[65277] = 32'b11111111111111111011000001001000;
assign LUT_4[65278] = 32'b00000000000000000001001111110100;
assign LUT_4[65279] = 32'b11111111111111111010011011101100;
assign LUT_4[65280] = 32'b00000000000000010000011001110001;
assign LUT_4[65281] = 32'b00000000000000001001100101101001;
assign LUT_4[65282] = 32'b00000000000000001111110100010101;
assign LUT_4[65283] = 32'b00000000000000001001000000001101;
assign LUT_4[65284] = 32'b00000000000000001101011010001101;
assign LUT_4[65285] = 32'b00000000000000000110100110000101;
assign LUT_4[65286] = 32'b00000000000000001100110100110001;
assign LUT_4[65287] = 32'b00000000000000000110000000101001;
assign LUT_4[65288] = 32'b00000000000000001001100110000110;
assign LUT_4[65289] = 32'b00000000000000000010110001111110;
assign LUT_4[65290] = 32'b00000000000000001001000000101010;
assign LUT_4[65291] = 32'b00000000000000000010001100100010;
assign LUT_4[65292] = 32'b00000000000000000110100110100010;
assign LUT_4[65293] = 32'b11111111111111111111110010011010;
assign LUT_4[65294] = 32'b00000000000000000110000001000110;
assign LUT_4[65295] = 32'b11111111111111111111001100111110;
assign LUT_4[65296] = 32'b00000000000000001110001011011111;
assign LUT_4[65297] = 32'b00000000000000000111010111010111;
assign LUT_4[65298] = 32'b00000000000000001101100110000011;
assign LUT_4[65299] = 32'b00000000000000000110110001111011;
assign LUT_4[65300] = 32'b00000000000000001011001011111011;
assign LUT_4[65301] = 32'b00000000000000000100010111110011;
assign LUT_4[65302] = 32'b00000000000000001010100110011111;
assign LUT_4[65303] = 32'b00000000000000000011110010010111;
assign LUT_4[65304] = 32'b00000000000000000111010111110100;
assign LUT_4[65305] = 32'b00000000000000000000100011101100;
assign LUT_4[65306] = 32'b00000000000000000110110010011000;
assign LUT_4[65307] = 32'b11111111111111111111111110010000;
assign LUT_4[65308] = 32'b00000000000000000100011000010000;
assign LUT_4[65309] = 32'b11111111111111111101100100001000;
assign LUT_4[65310] = 32'b00000000000000000011110010110100;
assign LUT_4[65311] = 32'b11111111111111111100111110101100;
assign LUT_4[65312] = 32'b00000000000000001110110100111000;
assign LUT_4[65313] = 32'b00000000000000001000000000110000;
assign LUT_4[65314] = 32'b00000000000000001110001111011100;
assign LUT_4[65315] = 32'b00000000000000000111011011010100;
assign LUT_4[65316] = 32'b00000000000000001011110101010100;
assign LUT_4[65317] = 32'b00000000000000000101000001001100;
assign LUT_4[65318] = 32'b00000000000000001011001111111000;
assign LUT_4[65319] = 32'b00000000000000000100011011110000;
assign LUT_4[65320] = 32'b00000000000000001000000001001101;
assign LUT_4[65321] = 32'b00000000000000000001001101000101;
assign LUT_4[65322] = 32'b00000000000000000111011011110001;
assign LUT_4[65323] = 32'b00000000000000000000100111101001;
assign LUT_4[65324] = 32'b00000000000000000101000001101001;
assign LUT_4[65325] = 32'b11111111111111111110001101100001;
assign LUT_4[65326] = 32'b00000000000000000100011100001101;
assign LUT_4[65327] = 32'b11111111111111111101101000000101;
assign LUT_4[65328] = 32'b00000000000000001100100110100110;
assign LUT_4[65329] = 32'b00000000000000000101110010011110;
assign LUT_4[65330] = 32'b00000000000000001100000001001010;
assign LUT_4[65331] = 32'b00000000000000000101001101000010;
assign LUT_4[65332] = 32'b00000000000000001001100111000010;
assign LUT_4[65333] = 32'b00000000000000000010110010111010;
assign LUT_4[65334] = 32'b00000000000000001001000001100110;
assign LUT_4[65335] = 32'b00000000000000000010001101011110;
assign LUT_4[65336] = 32'b00000000000000000101110010111011;
assign LUT_4[65337] = 32'b11111111111111111110111110110011;
assign LUT_4[65338] = 32'b00000000000000000101001101011111;
assign LUT_4[65339] = 32'b11111111111111111110011001010111;
assign LUT_4[65340] = 32'b00000000000000000010110011010111;
assign LUT_4[65341] = 32'b11111111111111111011111111001111;
assign LUT_4[65342] = 32'b00000000000000000010001101111011;
assign LUT_4[65343] = 32'b11111111111111111011011001110011;
assign LUT_4[65344] = 32'b00000000000000010001110001000101;
assign LUT_4[65345] = 32'b00000000000000001010111100111101;
assign LUT_4[65346] = 32'b00000000000000010001001011101001;
assign LUT_4[65347] = 32'b00000000000000001010010111100001;
assign LUT_4[65348] = 32'b00000000000000001110110001100001;
assign LUT_4[65349] = 32'b00000000000000000111111101011001;
assign LUT_4[65350] = 32'b00000000000000001110001100000101;
assign LUT_4[65351] = 32'b00000000000000000111010111111101;
assign LUT_4[65352] = 32'b00000000000000001010111101011010;
assign LUT_4[65353] = 32'b00000000000000000100001001010010;
assign LUT_4[65354] = 32'b00000000000000001010010111111110;
assign LUT_4[65355] = 32'b00000000000000000011100011110110;
assign LUT_4[65356] = 32'b00000000000000000111111101110110;
assign LUT_4[65357] = 32'b00000000000000000001001001101110;
assign LUT_4[65358] = 32'b00000000000000000111011000011010;
assign LUT_4[65359] = 32'b00000000000000000000100100010010;
assign LUT_4[65360] = 32'b00000000000000001111100010110011;
assign LUT_4[65361] = 32'b00000000000000001000101110101011;
assign LUT_4[65362] = 32'b00000000000000001110111101010111;
assign LUT_4[65363] = 32'b00000000000000001000001001001111;
assign LUT_4[65364] = 32'b00000000000000001100100011001111;
assign LUT_4[65365] = 32'b00000000000000000101101111000111;
assign LUT_4[65366] = 32'b00000000000000001011111101110011;
assign LUT_4[65367] = 32'b00000000000000000101001001101011;
assign LUT_4[65368] = 32'b00000000000000001000101111001000;
assign LUT_4[65369] = 32'b00000000000000000001111011000000;
assign LUT_4[65370] = 32'b00000000000000001000001001101100;
assign LUT_4[65371] = 32'b00000000000000000001010101100100;
assign LUT_4[65372] = 32'b00000000000000000101101111100100;
assign LUT_4[65373] = 32'b11111111111111111110111011011100;
assign LUT_4[65374] = 32'b00000000000000000101001010001000;
assign LUT_4[65375] = 32'b11111111111111111110010110000000;
assign LUT_4[65376] = 32'b00000000000000010000001100001100;
assign LUT_4[65377] = 32'b00000000000000001001011000000100;
assign LUT_4[65378] = 32'b00000000000000001111100110110000;
assign LUT_4[65379] = 32'b00000000000000001000110010101000;
assign LUT_4[65380] = 32'b00000000000000001101001100101000;
assign LUT_4[65381] = 32'b00000000000000000110011000100000;
assign LUT_4[65382] = 32'b00000000000000001100100111001100;
assign LUT_4[65383] = 32'b00000000000000000101110011000100;
assign LUT_4[65384] = 32'b00000000000000001001011000100001;
assign LUT_4[65385] = 32'b00000000000000000010100100011001;
assign LUT_4[65386] = 32'b00000000000000001000110011000101;
assign LUT_4[65387] = 32'b00000000000000000001111110111101;
assign LUT_4[65388] = 32'b00000000000000000110011000111101;
assign LUT_4[65389] = 32'b11111111111111111111100100110101;
assign LUT_4[65390] = 32'b00000000000000000101110011100001;
assign LUT_4[65391] = 32'b11111111111111111110111111011001;
assign LUT_4[65392] = 32'b00000000000000001101111101111010;
assign LUT_4[65393] = 32'b00000000000000000111001001110010;
assign LUT_4[65394] = 32'b00000000000000001101011000011110;
assign LUT_4[65395] = 32'b00000000000000000110100100010110;
assign LUT_4[65396] = 32'b00000000000000001010111110010110;
assign LUT_4[65397] = 32'b00000000000000000100001010001110;
assign LUT_4[65398] = 32'b00000000000000001010011000111010;
assign LUT_4[65399] = 32'b00000000000000000011100100110010;
assign LUT_4[65400] = 32'b00000000000000000111001010001111;
assign LUT_4[65401] = 32'b00000000000000000000010110000111;
assign LUT_4[65402] = 32'b00000000000000000110100100110011;
assign LUT_4[65403] = 32'b11111111111111111111110000101011;
assign LUT_4[65404] = 32'b00000000000000000100001010101011;
assign LUT_4[65405] = 32'b11111111111111111101010110100011;
assign LUT_4[65406] = 32'b00000000000000000011100101001111;
assign LUT_4[65407] = 32'b11111111111111111100110001000111;
assign LUT_4[65408] = 32'b00000000000000010010111111111001;
assign LUT_4[65409] = 32'b00000000000000001100001011110001;
assign LUT_4[65410] = 32'b00000000000000010010011010011101;
assign LUT_4[65411] = 32'b00000000000000001011100110010101;
assign LUT_4[65412] = 32'b00000000000000010000000000010101;
assign LUT_4[65413] = 32'b00000000000000001001001100001101;
assign LUT_4[65414] = 32'b00000000000000001111011010111001;
assign LUT_4[65415] = 32'b00000000000000001000100110110001;
assign LUT_4[65416] = 32'b00000000000000001100001100001110;
assign LUT_4[65417] = 32'b00000000000000000101011000000110;
assign LUT_4[65418] = 32'b00000000000000001011100110110010;
assign LUT_4[65419] = 32'b00000000000000000100110010101010;
assign LUT_4[65420] = 32'b00000000000000001001001100101010;
assign LUT_4[65421] = 32'b00000000000000000010011000100010;
assign LUT_4[65422] = 32'b00000000000000001000100111001110;
assign LUT_4[65423] = 32'b00000000000000000001110011000110;
assign LUT_4[65424] = 32'b00000000000000010000110001100111;
assign LUT_4[65425] = 32'b00000000000000001001111101011111;
assign LUT_4[65426] = 32'b00000000000000010000001100001011;
assign LUT_4[65427] = 32'b00000000000000001001011000000011;
assign LUT_4[65428] = 32'b00000000000000001101110010000011;
assign LUT_4[65429] = 32'b00000000000000000110111101111011;
assign LUT_4[65430] = 32'b00000000000000001101001100100111;
assign LUT_4[65431] = 32'b00000000000000000110011000011111;
assign LUT_4[65432] = 32'b00000000000000001001111101111100;
assign LUT_4[65433] = 32'b00000000000000000011001001110100;
assign LUT_4[65434] = 32'b00000000000000001001011000100000;
assign LUT_4[65435] = 32'b00000000000000000010100100011000;
assign LUT_4[65436] = 32'b00000000000000000110111110011000;
assign LUT_4[65437] = 32'b00000000000000000000001010010000;
assign LUT_4[65438] = 32'b00000000000000000110011000111100;
assign LUT_4[65439] = 32'b11111111111111111111100100110100;
assign LUT_4[65440] = 32'b00000000000000010001011011000000;
assign LUT_4[65441] = 32'b00000000000000001010100110111000;
assign LUT_4[65442] = 32'b00000000000000010000110101100100;
assign LUT_4[65443] = 32'b00000000000000001010000001011100;
assign LUT_4[65444] = 32'b00000000000000001110011011011100;
assign LUT_4[65445] = 32'b00000000000000000111100111010100;
assign LUT_4[65446] = 32'b00000000000000001101110110000000;
assign LUT_4[65447] = 32'b00000000000000000111000001111000;
assign LUT_4[65448] = 32'b00000000000000001010100111010101;
assign LUT_4[65449] = 32'b00000000000000000011110011001101;
assign LUT_4[65450] = 32'b00000000000000001010000001111001;
assign LUT_4[65451] = 32'b00000000000000000011001101110001;
assign LUT_4[65452] = 32'b00000000000000000111100111110001;
assign LUT_4[65453] = 32'b00000000000000000000110011101001;
assign LUT_4[65454] = 32'b00000000000000000111000010010101;
assign LUT_4[65455] = 32'b00000000000000000000001110001101;
assign LUT_4[65456] = 32'b00000000000000001111001100101110;
assign LUT_4[65457] = 32'b00000000000000001000011000100110;
assign LUT_4[65458] = 32'b00000000000000001110100111010010;
assign LUT_4[65459] = 32'b00000000000000000111110011001010;
assign LUT_4[65460] = 32'b00000000000000001100001101001010;
assign LUT_4[65461] = 32'b00000000000000000101011001000010;
assign LUT_4[65462] = 32'b00000000000000001011100111101110;
assign LUT_4[65463] = 32'b00000000000000000100110011100110;
assign LUT_4[65464] = 32'b00000000000000001000011001000011;
assign LUT_4[65465] = 32'b00000000000000000001100100111011;
assign LUT_4[65466] = 32'b00000000000000000111110011100111;
assign LUT_4[65467] = 32'b00000000000000000000111111011111;
assign LUT_4[65468] = 32'b00000000000000000101011001011111;
assign LUT_4[65469] = 32'b11111111111111111110100101010111;
assign LUT_4[65470] = 32'b00000000000000000100110100000011;
assign LUT_4[65471] = 32'b11111111111111111101111111111011;
assign LUT_4[65472] = 32'b00000000000000010100010111001101;
assign LUT_4[65473] = 32'b00000000000000001101100011000101;
assign LUT_4[65474] = 32'b00000000000000010011110001110001;
assign LUT_4[65475] = 32'b00000000000000001100111101101001;
assign LUT_4[65476] = 32'b00000000000000010001010111101001;
assign LUT_4[65477] = 32'b00000000000000001010100011100001;
assign LUT_4[65478] = 32'b00000000000000010000110010001101;
assign LUT_4[65479] = 32'b00000000000000001001111110000101;
assign LUT_4[65480] = 32'b00000000000000001101100011100010;
assign LUT_4[65481] = 32'b00000000000000000110101111011010;
assign LUT_4[65482] = 32'b00000000000000001100111110000110;
assign LUT_4[65483] = 32'b00000000000000000110001001111110;
assign LUT_4[65484] = 32'b00000000000000001010100011111110;
assign LUT_4[65485] = 32'b00000000000000000011101111110110;
assign LUT_4[65486] = 32'b00000000000000001001111110100010;
assign LUT_4[65487] = 32'b00000000000000000011001010011010;
assign LUT_4[65488] = 32'b00000000000000010010001000111011;
assign LUT_4[65489] = 32'b00000000000000001011010100110011;
assign LUT_4[65490] = 32'b00000000000000010001100011011111;
assign LUT_4[65491] = 32'b00000000000000001010101111010111;
assign LUT_4[65492] = 32'b00000000000000001111001001010111;
assign LUT_4[65493] = 32'b00000000000000001000010101001111;
assign LUT_4[65494] = 32'b00000000000000001110100011111011;
assign LUT_4[65495] = 32'b00000000000000000111101111110011;
assign LUT_4[65496] = 32'b00000000000000001011010101010000;
assign LUT_4[65497] = 32'b00000000000000000100100001001000;
assign LUT_4[65498] = 32'b00000000000000001010101111110100;
assign LUT_4[65499] = 32'b00000000000000000011111011101100;
assign LUT_4[65500] = 32'b00000000000000001000010101101100;
assign LUT_4[65501] = 32'b00000000000000000001100001100100;
assign LUT_4[65502] = 32'b00000000000000000111110000010000;
assign LUT_4[65503] = 32'b00000000000000000000111100001000;
assign LUT_4[65504] = 32'b00000000000000010010110010010100;
assign LUT_4[65505] = 32'b00000000000000001011111110001100;
assign LUT_4[65506] = 32'b00000000000000010010001100111000;
assign LUT_4[65507] = 32'b00000000000000001011011000110000;
assign LUT_4[65508] = 32'b00000000000000001111110010110000;
assign LUT_4[65509] = 32'b00000000000000001000111110101000;
assign LUT_4[65510] = 32'b00000000000000001111001101010100;
assign LUT_4[65511] = 32'b00000000000000001000011001001100;
assign LUT_4[65512] = 32'b00000000000000001011111110101001;
assign LUT_4[65513] = 32'b00000000000000000101001010100001;
assign LUT_4[65514] = 32'b00000000000000001011011001001101;
assign LUT_4[65515] = 32'b00000000000000000100100101000101;
assign LUT_4[65516] = 32'b00000000000000001000111111000101;
assign LUT_4[65517] = 32'b00000000000000000010001010111101;
assign LUT_4[65518] = 32'b00000000000000001000011001101001;
assign LUT_4[65519] = 32'b00000000000000000001100101100001;
assign LUT_4[65520] = 32'b00000000000000010000100100000010;
assign LUT_4[65521] = 32'b00000000000000001001101111111010;
assign LUT_4[65522] = 32'b00000000000000001111111110100110;
assign LUT_4[65523] = 32'b00000000000000001001001010011110;
assign LUT_4[65524] = 32'b00000000000000001101100100011110;
assign LUT_4[65525] = 32'b00000000000000000110110000010110;
assign LUT_4[65526] = 32'b00000000000000001100111111000010;
assign LUT_4[65527] = 32'b00000000000000000110001010111010;
assign LUT_4[65528] = 32'b00000000000000001001110000010111;
assign LUT_4[65529] = 32'b00000000000000000010111100001111;
assign LUT_4[65530] = 32'b00000000000000001001001010111011;
assign LUT_4[65531] = 32'b00000000000000000010010110110011;
assign LUT_4[65532] = 32'b00000000000000000110110000110011;
assign LUT_4[65533] = 32'b11111111111111111111111100101011;
assign LUT_4[65534] = 32'b00000000000000000110001011010111;
assign LUT_4[65535] = 32'b11111111111111111111010111001111;
endmodule
